magic
tech sky130A
magscale 1 2
timestamp 1641030212
<< obsli1 >>
rect 1104 2159 99147 197489
<< obsm1 >>
rect 106 1368 99898 197520
<< metal2 >>
rect 386 199200 442 200000
rect 1214 199200 1270 200000
rect 2042 199200 2098 200000
rect 2962 199200 3018 200000
rect 3790 199200 3846 200000
rect 4618 199200 4674 200000
rect 5538 199200 5594 200000
rect 6366 199200 6422 200000
rect 7194 199200 7250 200000
rect 8114 199200 8170 200000
rect 8942 199200 8998 200000
rect 9862 199200 9918 200000
rect 10690 199200 10746 200000
rect 11518 199200 11574 200000
rect 12438 199200 12494 200000
rect 13266 199200 13322 200000
rect 14094 199200 14150 200000
rect 15014 199200 15070 200000
rect 15842 199200 15898 200000
rect 16762 199200 16818 200000
rect 17590 199200 17646 200000
rect 18418 199200 18474 200000
rect 19338 199200 19394 200000
rect 20166 199200 20222 200000
rect 20994 199200 21050 200000
rect 21914 199200 21970 200000
rect 22742 199200 22798 200000
rect 23662 199200 23718 200000
rect 24490 199200 24546 200000
rect 25318 199200 25374 200000
rect 26238 199200 26294 200000
rect 27066 199200 27122 200000
rect 27894 199200 27950 200000
rect 28814 199200 28870 200000
rect 29642 199200 29698 200000
rect 30470 199200 30526 200000
rect 31390 199200 31446 200000
rect 32218 199200 32274 200000
rect 33138 199200 33194 200000
rect 33966 199200 34022 200000
rect 34794 199200 34850 200000
rect 35714 199200 35770 200000
rect 36542 199200 36598 200000
rect 37370 199200 37426 200000
rect 38290 199200 38346 200000
rect 39118 199200 39174 200000
rect 40038 199200 40094 200000
rect 40866 199200 40922 200000
rect 41694 199200 41750 200000
rect 42614 199200 42670 200000
rect 43442 199200 43498 200000
rect 44270 199200 44326 200000
rect 45190 199200 45246 200000
rect 46018 199200 46074 200000
rect 46938 199200 46994 200000
rect 47766 199200 47822 200000
rect 48594 199200 48650 200000
rect 49514 199200 49570 200000
rect 50342 199200 50398 200000
rect 51170 199200 51226 200000
rect 52090 199200 52146 200000
rect 52918 199200 52974 200000
rect 53746 199200 53802 200000
rect 54666 199200 54722 200000
rect 55494 199200 55550 200000
rect 56414 199200 56470 200000
rect 57242 199200 57298 200000
rect 58070 199200 58126 200000
rect 58990 199200 59046 200000
rect 59818 199200 59874 200000
rect 60646 199200 60702 200000
rect 61566 199200 61622 200000
rect 62394 199200 62450 200000
rect 63314 199200 63370 200000
rect 64142 199200 64198 200000
rect 64970 199200 65026 200000
rect 65890 199200 65946 200000
rect 66718 199200 66774 200000
rect 67546 199200 67602 200000
rect 68466 199200 68522 200000
rect 69294 199200 69350 200000
rect 70214 199200 70270 200000
rect 71042 199200 71098 200000
rect 71870 199200 71926 200000
rect 72790 199200 72846 200000
rect 73618 199200 73674 200000
rect 74446 199200 74502 200000
rect 75366 199200 75422 200000
rect 76194 199200 76250 200000
rect 77022 199200 77078 200000
rect 77942 199200 77998 200000
rect 78770 199200 78826 200000
rect 79690 199200 79746 200000
rect 80518 199200 80574 200000
rect 81346 199200 81402 200000
rect 82266 199200 82322 200000
rect 83094 199200 83150 200000
rect 83922 199200 83978 200000
rect 84842 199200 84898 200000
rect 85670 199200 85726 200000
rect 86590 199200 86646 200000
rect 87418 199200 87474 200000
rect 88246 199200 88302 200000
rect 89166 199200 89222 200000
rect 89994 199200 90050 200000
rect 90822 199200 90878 200000
rect 91742 199200 91798 200000
rect 92570 199200 92626 200000
rect 93490 199200 93546 200000
rect 94318 199200 94374 200000
rect 95146 199200 95202 200000
rect 96066 199200 96122 200000
rect 96894 199200 96950 200000
rect 97722 199200 97778 200000
rect 98642 199200 98698 200000
rect 99470 199200 99526 200000
rect 110 0 166 800
rect 294 0 350 800
rect 478 0 534 800
rect 662 0 718 800
rect 846 0 902 800
rect 1030 0 1086 800
rect 1306 0 1362 800
rect 1490 0 1546 800
rect 1674 0 1730 800
rect 1858 0 1914 800
rect 2042 0 2098 800
rect 2318 0 2374 800
rect 2502 0 2558 800
rect 2686 0 2742 800
rect 2870 0 2926 800
rect 3054 0 3110 800
rect 3330 0 3386 800
rect 3514 0 3570 800
rect 3698 0 3754 800
rect 3882 0 3938 800
rect 4066 0 4122 800
rect 4342 0 4398 800
rect 4526 0 4582 800
rect 4710 0 4766 800
rect 4894 0 4950 800
rect 5078 0 5134 800
rect 5262 0 5318 800
rect 5538 0 5594 800
rect 5722 0 5778 800
rect 5906 0 5962 800
rect 6090 0 6146 800
rect 6274 0 6330 800
rect 6550 0 6606 800
rect 6734 0 6790 800
rect 6918 0 6974 800
rect 7102 0 7158 800
rect 7286 0 7342 800
rect 7562 0 7618 800
rect 7746 0 7802 800
rect 7930 0 7986 800
rect 8114 0 8170 800
rect 8298 0 8354 800
rect 8574 0 8630 800
rect 8758 0 8814 800
rect 8942 0 8998 800
rect 9126 0 9182 800
rect 9310 0 9366 800
rect 9586 0 9642 800
rect 9770 0 9826 800
rect 9954 0 10010 800
rect 10138 0 10194 800
rect 10322 0 10378 800
rect 10506 0 10562 800
rect 10782 0 10838 800
rect 10966 0 11022 800
rect 11150 0 11206 800
rect 11334 0 11390 800
rect 11518 0 11574 800
rect 11794 0 11850 800
rect 11978 0 12034 800
rect 12162 0 12218 800
rect 12346 0 12402 800
rect 12530 0 12586 800
rect 12806 0 12862 800
rect 12990 0 13046 800
rect 13174 0 13230 800
rect 13358 0 13414 800
rect 13542 0 13598 800
rect 13818 0 13874 800
rect 14002 0 14058 800
rect 14186 0 14242 800
rect 14370 0 14426 800
rect 14554 0 14610 800
rect 14738 0 14794 800
rect 15014 0 15070 800
rect 15198 0 15254 800
rect 15382 0 15438 800
rect 15566 0 15622 800
rect 15750 0 15806 800
rect 16026 0 16082 800
rect 16210 0 16266 800
rect 16394 0 16450 800
rect 16578 0 16634 800
rect 16762 0 16818 800
rect 17038 0 17094 800
rect 17222 0 17278 800
rect 17406 0 17462 800
rect 17590 0 17646 800
rect 17774 0 17830 800
rect 18050 0 18106 800
rect 18234 0 18290 800
rect 18418 0 18474 800
rect 18602 0 18658 800
rect 18786 0 18842 800
rect 19062 0 19118 800
rect 19246 0 19302 800
rect 19430 0 19486 800
rect 19614 0 19670 800
rect 19798 0 19854 800
rect 19982 0 20038 800
rect 20258 0 20314 800
rect 20442 0 20498 800
rect 20626 0 20682 800
rect 20810 0 20866 800
rect 20994 0 21050 800
rect 21270 0 21326 800
rect 21454 0 21510 800
rect 21638 0 21694 800
rect 21822 0 21878 800
rect 22006 0 22062 800
rect 22282 0 22338 800
rect 22466 0 22522 800
rect 22650 0 22706 800
rect 22834 0 22890 800
rect 23018 0 23074 800
rect 23294 0 23350 800
rect 23478 0 23534 800
rect 23662 0 23718 800
rect 23846 0 23902 800
rect 24030 0 24086 800
rect 24214 0 24270 800
rect 24490 0 24546 800
rect 24674 0 24730 800
rect 24858 0 24914 800
rect 25042 0 25098 800
rect 25226 0 25282 800
rect 25502 0 25558 800
rect 25686 0 25742 800
rect 25870 0 25926 800
rect 26054 0 26110 800
rect 26238 0 26294 800
rect 26514 0 26570 800
rect 26698 0 26754 800
rect 26882 0 26938 800
rect 27066 0 27122 800
rect 27250 0 27306 800
rect 27526 0 27582 800
rect 27710 0 27766 800
rect 27894 0 27950 800
rect 28078 0 28134 800
rect 28262 0 28318 800
rect 28538 0 28594 800
rect 28722 0 28778 800
rect 28906 0 28962 800
rect 29090 0 29146 800
rect 29274 0 29330 800
rect 29458 0 29514 800
rect 29734 0 29790 800
rect 29918 0 29974 800
rect 30102 0 30158 800
rect 30286 0 30342 800
rect 30470 0 30526 800
rect 30746 0 30802 800
rect 30930 0 30986 800
rect 31114 0 31170 800
rect 31298 0 31354 800
rect 31482 0 31538 800
rect 31758 0 31814 800
rect 31942 0 31998 800
rect 32126 0 32182 800
rect 32310 0 32366 800
rect 32494 0 32550 800
rect 32770 0 32826 800
rect 32954 0 33010 800
rect 33138 0 33194 800
rect 33322 0 33378 800
rect 33506 0 33562 800
rect 33690 0 33746 800
rect 33966 0 34022 800
rect 34150 0 34206 800
rect 34334 0 34390 800
rect 34518 0 34574 800
rect 34702 0 34758 800
rect 34978 0 35034 800
rect 35162 0 35218 800
rect 35346 0 35402 800
rect 35530 0 35586 800
rect 35714 0 35770 800
rect 35990 0 36046 800
rect 36174 0 36230 800
rect 36358 0 36414 800
rect 36542 0 36598 800
rect 36726 0 36782 800
rect 37002 0 37058 800
rect 37186 0 37242 800
rect 37370 0 37426 800
rect 37554 0 37610 800
rect 37738 0 37794 800
rect 38014 0 38070 800
rect 38198 0 38254 800
rect 38382 0 38438 800
rect 38566 0 38622 800
rect 38750 0 38806 800
rect 38934 0 38990 800
rect 39210 0 39266 800
rect 39394 0 39450 800
rect 39578 0 39634 800
rect 39762 0 39818 800
rect 39946 0 40002 800
rect 40222 0 40278 800
rect 40406 0 40462 800
rect 40590 0 40646 800
rect 40774 0 40830 800
rect 40958 0 41014 800
rect 41234 0 41290 800
rect 41418 0 41474 800
rect 41602 0 41658 800
rect 41786 0 41842 800
rect 41970 0 42026 800
rect 42246 0 42302 800
rect 42430 0 42486 800
rect 42614 0 42670 800
rect 42798 0 42854 800
rect 42982 0 43038 800
rect 43166 0 43222 800
rect 43442 0 43498 800
rect 43626 0 43682 800
rect 43810 0 43866 800
rect 43994 0 44050 800
rect 44178 0 44234 800
rect 44454 0 44510 800
rect 44638 0 44694 800
rect 44822 0 44878 800
rect 45006 0 45062 800
rect 45190 0 45246 800
rect 45466 0 45522 800
rect 45650 0 45706 800
rect 45834 0 45890 800
rect 46018 0 46074 800
rect 46202 0 46258 800
rect 46478 0 46534 800
rect 46662 0 46718 800
rect 46846 0 46902 800
rect 47030 0 47086 800
rect 47214 0 47270 800
rect 47490 0 47546 800
rect 47674 0 47730 800
rect 47858 0 47914 800
rect 48042 0 48098 800
rect 48226 0 48282 800
rect 48410 0 48466 800
rect 48686 0 48742 800
rect 48870 0 48926 800
rect 49054 0 49110 800
rect 49238 0 49294 800
rect 49422 0 49478 800
rect 49698 0 49754 800
rect 49882 0 49938 800
rect 50066 0 50122 800
rect 50250 0 50306 800
rect 50434 0 50490 800
rect 50710 0 50766 800
rect 50894 0 50950 800
rect 51078 0 51134 800
rect 51262 0 51318 800
rect 51446 0 51502 800
rect 51722 0 51778 800
rect 51906 0 51962 800
rect 52090 0 52146 800
rect 52274 0 52330 800
rect 52458 0 52514 800
rect 52642 0 52698 800
rect 52918 0 52974 800
rect 53102 0 53158 800
rect 53286 0 53342 800
rect 53470 0 53526 800
rect 53654 0 53710 800
rect 53930 0 53986 800
rect 54114 0 54170 800
rect 54298 0 54354 800
rect 54482 0 54538 800
rect 54666 0 54722 800
rect 54942 0 54998 800
rect 55126 0 55182 800
rect 55310 0 55366 800
rect 55494 0 55550 800
rect 55678 0 55734 800
rect 55954 0 56010 800
rect 56138 0 56194 800
rect 56322 0 56378 800
rect 56506 0 56562 800
rect 56690 0 56746 800
rect 56966 0 57022 800
rect 57150 0 57206 800
rect 57334 0 57390 800
rect 57518 0 57574 800
rect 57702 0 57758 800
rect 57886 0 57942 800
rect 58162 0 58218 800
rect 58346 0 58402 800
rect 58530 0 58586 800
rect 58714 0 58770 800
rect 58898 0 58954 800
rect 59174 0 59230 800
rect 59358 0 59414 800
rect 59542 0 59598 800
rect 59726 0 59782 800
rect 59910 0 59966 800
rect 60186 0 60242 800
rect 60370 0 60426 800
rect 60554 0 60610 800
rect 60738 0 60794 800
rect 60922 0 60978 800
rect 61198 0 61254 800
rect 61382 0 61438 800
rect 61566 0 61622 800
rect 61750 0 61806 800
rect 61934 0 61990 800
rect 62118 0 62174 800
rect 62394 0 62450 800
rect 62578 0 62634 800
rect 62762 0 62818 800
rect 62946 0 63002 800
rect 63130 0 63186 800
rect 63406 0 63462 800
rect 63590 0 63646 800
rect 63774 0 63830 800
rect 63958 0 64014 800
rect 64142 0 64198 800
rect 64418 0 64474 800
rect 64602 0 64658 800
rect 64786 0 64842 800
rect 64970 0 65026 800
rect 65154 0 65210 800
rect 65430 0 65486 800
rect 65614 0 65670 800
rect 65798 0 65854 800
rect 65982 0 66038 800
rect 66166 0 66222 800
rect 66442 0 66498 800
rect 66626 0 66682 800
rect 66810 0 66866 800
rect 66994 0 67050 800
rect 67178 0 67234 800
rect 67362 0 67418 800
rect 67638 0 67694 800
rect 67822 0 67878 800
rect 68006 0 68062 800
rect 68190 0 68246 800
rect 68374 0 68430 800
rect 68650 0 68706 800
rect 68834 0 68890 800
rect 69018 0 69074 800
rect 69202 0 69258 800
rect 69386 0 69442 800
rect 69662 0 69718 800
rect 69846 0 69902 800
rect 70030 0 70086 800
rect 70214 0 70270 800
rect 70398 0 70454 800
rect 70674 0 70730 800
rect 70858 0 70914 800
rect 71042 0 71098 800
rect 71226 0 71282 800
rect 71410 0 71466 800
rect 71594 0 71650 800
rect 71870 0 71926 800
rect 72054 0 72110 800
rect 72238 0 72294 800
rect 72422 0 72478 800
rect 72606 0 72662 800
rect 72882 0 72938 800
rect 73066 0 73122 800
rect 73250 0 73306 800
rect 73434 0 73490 800
rect 73618 0 73674 800
rect 73894 0 73950 800
rect 74078 0 74134 800
rect 74262 0 74318 800
rect 74446 0 74502 800
rect 74630 0 74686 800
rect 74906 0 74962 800
rect 75090 0 75146 800
rect 75274 0 75330 800
rect 75458 0 75514 800
rect 75642 0 75698 800
rect 75918 0 75974 800
rect 76102 0 76158 800
rect 76286 0 76342 800
rect 76470 0 76526 800
rect 76654 0 76710 800
rect 76838 0 76894 800
rect 77114 0 77170 800
rect 77298 0 77354 800
rect 77482 0 77538 800
rect 77666 0 77722 800
rect 77850 0 77906 800
rect 78126 0 78182 800
rect 78310 0 78366 800
rect 78494 0 78550 800
rect 78678 0 78734 800
rect 78862 0 78918 800
rect 79138 0 79194 800
rect 79322 0 79378 800
rect 79506 0 79562 800
rect 79690 0 79746 800
rect 79874 0 79930 800
rect 80150 0 80206 800
rect 80334 0 80390 800
rect 80518 0 80574 800
rect 80702 0 80758 800
rect 80886 0 80942 800
rect 81070 0 81126 800
rect 81346 0 81402 800
rect 81530 0 81586 800
rect 81714 0 81770 800
rect 81898 0 81954 800
rect 82082 0 82138 800
rect 82358 0 82414 800
rect 82542 0 82598 800
rect 82726 0 82782 800
rect 82910 0 82966 800
rect 83094 0 83150 800
rect 83370 0 83426 800
rect 83554 0 83610 800
rect 83738 0 83794 800
rect 83922 0 83978 800
rect 84106 0 84162 800
rect 84382 0 84438 800
rect 84566 0 84622 800
rect 84750 0 84806 800
rect 84934 0 84990 800
rect 85118 0 85174 800
rect 85394 0 85450 800
rect 85578 0 85634 800
rect 85762 0 85818 800
rect 85946 0 86002 800
rect 86130 0 86186 800
rect 86314 0 86370 800
rect 86590 0 86646 800
rect 86774 0 86830 800
rect 86958 0 87014 800
rect 87142 0 87198 800
rect 87326 0 87382 800
rect 87602 0 87658 800
rect 87786 0 87842 800
rect 87970 0 88026 800
rect 88154 0 88210 800
rect 88338 0 88394 800
rect 88614 0 88670 800
rect 88798 0 88854 800
rect 88982 0 89038 800
rect 89166 0 89222 800
rect 89350 0 89406 800
rect 89626 0 89682 800
rect 89810 0 89866 800
rect 89994 0 90050 800
rect 90178 0 90234 800
rect 90362 0 90418 800
rect 90546 0 90602 800
rect 90822 0 90878 800
rect 91006 0 91062 800
rect 91190 0 91246 800
rect 91374 0 91430 800
rect 91558 0 91614 800
rect 91834 0 91890 800
rect 92018 0 92074 800
rect 92202 0 92258 800
rect 92386 0 92442 800
rect 92570 0 92626 800
rect 92846 0 92902 800
rect 93030 0 93086 800
rect 93214 0 93270 800
rect 93398 0 93454 800
rect 93582 0 93638 800
rect 93858 0 93914 800
rect 94042 0 94098 800
rect 94226 0 94282 800
rect 94410 0 94466 800
rect 94594 0 94650 800
rect 94870 0 94926 800
rect 95054 0 95110 800
rect 95238 0 95294 800
rect 95422 0 95478 800
rect 95606 0 95662 800
rect 95790 0 95846 800
rect 96066 0 96122 800
rect 96250 0 96306 800
rect 96434 0 96490 800
rect 96618 0 96674 800
rect 96802 0 96858 800
rect 97078 0 97134 800
rect 97262 0 97318 800
rect 97446 0 97502 800
rect 97630 0 97686 800
rect 97814 0 97870 800
rect 98090 0 98146 800
rect 98274 0 98330 800
rect 98458 0 98514 800
rect 98642 0 98698 800
rect 98826 0 98882 800
rect 99102 0 99158 800
rect 99286 0 99342 800
rect 99470 0 99526 800
rect 99654 0 99710 800
rect 99838 0 99894 800
<< obsm2 >>
rect 112 199144 330 199200
rect 498 199144 1158 199200
rect 1326 199144 1986 199200
rect 2154 199144 2906 199200
rect 3074 199144 3734 199200
rect 3902 199144 4562 199200
rect 4730 199144 5482 199200
rect 5650 199144 6310 199200
rect 6478 199144 7138 199200
rect 7306 199144 8058 199200
rect 8226 199144 8886 199200
rect 9054 199144 9806 199200
rect 9974 199144 10634 199200
rect 10802 199144 11462 199200
rect 11630 199144 12382 199200
rect 12550 199144 13210 199200
rect 13378 199144 14038 199200
rect 14206 199144 14958 199200
rect 15126 199144 15786 199200
rect 15954 199144 16706 199200
rect 16874 199144 17534 199200
rect 17702 199144 18362 199200
rect 18530 199144 19282 199200
rect 19450 199144 20110 199200
rect 20278 199144 20938 199200
rect 21106 199144 21858 199200
rect 22026 199144 22686 199200
rect 22854 199144 23606 199200
rect 23774 199144 24434 199200
rect 24602 199144 25262 199200
rect 25430 199144 26182 199200
rect 26350 199144 27010 199200
rect 27178 199144 27838 199200
rect 28006 199144 28758 199200
rect 28926 199144 29586 199200
rect 29754 199144 30414 199200
rect 30582 199144 31334 199200
rect 31502 199144 32162 199200
rect 32330 199144 33082 199200
rect 33250 199144 33910 199200
rect 34078 199144 34738 199200
rect 34906 199144 35658 199200
rect 35826 199144 36486 199200
rect 36654 199144 37314 199200
rect 37482 199144 38234 199200
rect 38402 199144 39062 199200
rect 39230 199144 39982 199200
rect 40150 199144 40810 199200
rect 40978 199144 41638 199200
rect 41806 199144 42558 199200
rect 42726 199144 43386 199200
rect 43554 199144 44214 199200
rect 44382 199144 45134 199200
rect 45302 199144 45962 199200
rect 46130 199144 46882 199200
rect 47050 199144 47710 199200
rect 47878 199144 48538 199200
rect 48706 199144 49458 199200
rect 49626 199144 50286 199200
rect 50454 199144 51114 199200
rect 51282 199144 52034 199200
rect 52202 199144 52862 199200
rect 53030 199144 53690 199200
rect 53858 199144 54610 199200
rect 54778 199144 55438 199200
rect 55606 199144 56358 199200
rect 56526 199144 57186 199200
rect 57354 199144 58014 199200
rect 58182 199144 58934 199200
rect 59102 199144 59762 199200
rect 59930 199144 60590 199200
rect 60758 199144 61510 199200
rect 61678 199144 62338 199200
rect 62506 199144 63258 199200
rect 63426 199144 64086 199200
rect 64254 199144 64914 199200
rect 65082 199144 65834 199200
rect 66002 199144 66662 199200
rect 66830 199144 67490 199200
rect 67658 199144 68410 199200
rect 68578 199144 69238 199200
rect 69406 199144 70158 199200
rect 70326 199144 70986 199200
rect 71154 199144 71814 199200
rect 71982 199144 72734 199200
rect 72902 199144 73562 199200
rect 73730 199144 74390 199200
rect 74558 199144 75310 199200
rect 75478 199144 76138 199200
rect 76306 199144 76966 199200
rect 77134 199144 77886 199200
rect 78054 199144 78714 199200
rect 78882 199144 79634 199200
rect 79802 199144 80462 199200
rect 80630 199144 81290 199200
rect 81458 199144 82210 199200
rect 82378 199144 83038 199200
rect 83206 199144 83866 199200
rect 84034 199144 84786 199200
rect 84954 199144 85614 199200
rect 85782 199144 86534 199200
rect 86702 199144 87362 199200
rect 87530 199144 88190 199200
rect 88358 199144 89110 199200
rect 89278 199144 89938 199200
rect 90106 199144 90766 199200
rect 90934 199144 91686 199200
rect 91854 199144 92514 199200
rect 92682 199144 93434 199200
rect 93602 199144 94262 199200
rect 94430 199144 95090 199200
rect 95258 199144 96010 199200
rect 96178 199144 96838 199200
rect 97006 199144 97666 199200
rect 97834 199144 98586 199200
rect 98754 199144 99414 199200
rect 99582 199144 99892 199200
rect 112 856 99892 199144
rect 222 800 238 856
rect 406 800 422 856
rect 590 800 606 856
rect 774 800 790 856
rect 958 800 974 856
rect 1142 800 1250 856
rect 1418 800 1434 856
rect 1602 800 1618 856
rect 1786 800 1802 856
rect 1970 800 1986 856
rect 2154 800 2262 856
rect 2430 800 2446 856
rect 2614 800 2630 856
rect 2798 800 2814 856
rect 2982 800 2998 856
rect 3166 800 3274 856
rect 3442 800 3458 856
rect 3626 800 3642 856
rect 3810 800 3826 856
rect 3994 800 4010 856
rect 4178 800 4286 856
rect 4454 800 4470 856
rect 4638 800 4654 856
rect 4822 800 4838 856
rect 5006 800 5022 856
rect 5190 800 5206 856
rect 5374 800 5482 856
rect 5650 800 5666 856
rect 5834 800 5850 856
rect 6018 800 6034 856
rect 6202 800 6218 856
rect 6386 800 6494 856
rect 6662 800 6678 856
rect 6846 800 6862 856
rect 7030 800 7046 856
rect 7214 800 7230 856
rect 7398 800 7506 856
rect 7674 800 7690 856
rect 7858 800 7874 856
rect 8042 800 8058 856
rect 8226 800 8242 856
rect 8410 800 8518 856
rect 8686 800 8702 856
rect 8870 800 8886 856
rect 9054 800 9070 856
rect 9238 800 9254 856
rect 9422 800 9530 856
rect 9698 800 9714 856
rect 9882 800 9898 856
rect 10066 800 10082 856
rect 10250 800 10266 856
rect 10434 800 10450 856
rect 10618 800 10726 856
rect 10894 800 10910 856
rect 11078 800 11094 856
rect 11262 800 11278 856
rect 11446 800 11462 856
rect 11630 800 11738 856
rect 11906 800 11922 856
rect 12090 800 12106 856
rect 12274 800 12290 856
rect 12458 800 12474 856
rect 12642 800 12750 856
rect 12918 800 12934 856
rect 13102 800 13118 856
rect 13286 800 13302 856
rect 13470 800 13486 856
rect 13654 800 13762 856
rect 13930 800 13946 856
rect 14114 800 14130 856
rect 14298 800 14314 856
rect 14482 800 14498 856
rect 14666 800 14682 856
rect 14850 800 14958 856
rect 15126 800 15142 856
rect 15310 800 15326 856
rect 15494 800 15510 856
rect 15678 800 15694 856
rect 15862 800 15970 856
rect 16138 800 16154 856
rect 16322 800 16338 856
rect 16506 800 16522 856
rect 16690 800 16706 856
rect 16874 800 16982 856
rect 17150 800 17166 856
rect 17334 800 17350 856
rect 17518 800 17534 856
rect 17702 800 17718 856
rect 17886 800 17994 856
rect 18162 800 18178 856
rect 18346 800 18362 856
rect 18530 800 18546 856
rect 18714 800 18730 856
rect 18898 800 19006 856
rect 19174 800 19190 856
rect 19358 800 19374 856
rect 19542 800 19558 856
rect 19726 800 19742 856
rect 19910 800 19926 856
rect 20094 800 20202 856
rect 20370 800 20386 856
rect 20554 800 20570 856
rect 20738 800 20754 856
rect 20922 800 20938 856
rect 21106 800 21214 856
rect 21382 800 21398 856
rect 21566 800 21582 856
rect 21750 800 21766 856
rect 21934 800 21950 856
rect 22118 800 22226 856
rect 22394 800 22410 856
rect 22578 800 22594 856
rect 22762 800 22778 856
rect 22946 800 22962 856
rect 23130 800 23238 856
rect 23406 800 23422 856
rect 23590 800 23606 856
rect 23774 800 23790 856
rect 23958 800 23974 856
rect 24142 800 24158 856
rect 24326 800 24434 856
rect 24602 800 24618 856
rect 24786 800 24802 856
rect 24970 800 24986 856
rect 25154 800 25170 856
rect 25338 800 25446 856
rect 25614 800 25630 856
rect 25798 800 25814 856
rect 25982 800 25998 856
rect 26166 800 26182 856
rect 26350 800 26458 856
rect 26626 800 26642 856
rect 26810 800 26826 856
rect 26994 800 27010 856
rect 27178 800 27194 856
rect 27362 800 27470 856
rect 27638 800 27654 856
rect 27822 800 27838 856
rect 28006 800 28022 856
rect 28190 800 28206 856
rect 28374 800 28482 856
rect 28650 800 28666 856
rect 28834 800 28850 856
rect 29018 800 29034 856
rect 29202 800 29218 856
rect 29386 800 29402 856
rect 29570 800 29678 856
rect 29846 800 29862 856
rect 30030 800 30046 856
rect 30214 800 30230 856
rect 30398 800 30414 856
rect 30582 800 30690 856
rect 30858 800 30874 856
rect 31042 800 31058 856
rect 31226 800 31242 856
rect 31410 800 31426 856
rect 31594 800 31702 856
rect 31870 800 31886 856
rect 32054 800 32070 856
rect 32238 800 32254 856
rect 32422 800 32438 856
rect 32606 800 32714 856
rect 32882 800 32898 856
rect 33066 800 33082 856
rect 33250 800 33266 856
rect 33434 800 33450 856
rect 33618 800 33634 856
rect 33802 800 33910 856
rect 34078 800 34094 856
rect 34262 800 34278 856
rect 34446 800 34462 856
rect 34630 800 34646 856
rect 34814 800 34922 856
rect 35090 800 35106 856
rect 35274 800 35290 856
rect 35458 800 35474 856
rect 35642 800 35658 856
rect 35826 800 35934 856
rect 36102 800 36118 856
rect 36286 800 36302 856
rect 36470 800 36486 856
rect 36654 800 36670 856
rect 36838 800 36946 856
rect 37114 800 37130 856
rect 37298 800 37314 856
rect 37482 800 37498 856
rect 37666 800 37682 856
rect 37850 800 37958 856
rect 38126 800 38142 856
rect 38310 800 38326 856
rect 38494 800 38510 856
rect 38678 800 38694 856
rect 38862 800 38878 856
rect 39046 800 39154 856
rect 39322 800 39338 856
rect 39506 800 39522 856
rect 39690 800 39706 856
rect 39874 800 39890 856
rect 40058 800 40166 856
rect 40334 800 40350 856
rect 40518 800 40534 856
rect 40702 800 40718 856
rect 40886 800 40902 856
rect 41070 800 41178 856
rect 41346 800 41362 856
rect 41530 800 41546 856
rect 41714 800 41730 856
rect 41898 800 41914 856
rect 42082 800 42190 856
rect 42358 800 42374 856
rect 42542 800 42558 856
rect 42726 800 42742 856
rect 42910 800 42926 856
rect 43094 800 43110 856
rect 43278 800 43386 856
rect 43554 800 43570 856
rect 43738 800 43754 856
rect 43922 800 43938 856
rect 44106 800 44122 856
rect 44290 800 44398 856
rect 44566 800 44582 856
rect 44750 800 44766 856
rect 44934 800 44950 856
rect 45118 800 45134 856
rect 45302 800 45410 856
rect 45578 800 45594 856
rect 45762 800 45778 856
rect 45946 800 45962 856
rect 46130 800 46146 856
rect 46314 800 46422 856
rect 46590 800 46606 856
rect 46774 800 46790 856
rect 46958 800 46974 856
rect 47142 800 47158 856
rect 47326 800 47434 856
rect 47602 800 47618 856
rect 47786 800 47802 856
rect 47970 800 47986 856
rect 48154 800 48170 856
rect 48338 800 48354 856
rect 48522 800 48630 856
rect 48798 800 48814 856
rect 48982 800 48998 856
rect 49166 800 49182 856
rect 49350 800 49366 856
rect 49534 800 49642 856
rect 49810 800 49826 856
rect 49994 800 50010 856
rect 50178 800 50194 856
rect 50362 800 50378 856
rect 50546 800 50654 856
rect 50822 800 50838 856
rect 51006 800 51022 856
rect 51190 800 51206 856
rect 51374 800 51390 856
rect 51558 800 51666 856
rect 51834 800 51850 856
rect 52018 800 52034 856
rect 52202 800 52218 856
rect 52386 800 52402 856
rect 52570 800 52586 856
rect 52754 800 52862 856
rect 53030 800 53046 856
rect 53214 800 53230 856
rect 53398 800 53414 856
rect 53582 800 53598 856
rect 53766 800 53874 856
rect 54042 800 54058 856
rect 54226 800 54242 856
rect 54410 800 54426 856
rect 54594 800 54610 856
rect 54778 800 54886 856
rect 55054 800 55070 856
rect 55238 800 55254 856
rect 55422 800 55438 856
rect 55606 800 55622 856
rect 55790 800 55898 856
rect 56066 800 56082 856
rect 56250 800 56266 856
rect 56434 800 56450 856
rect 56618 800 56634 856
rect 56802 800 56910 856
rect 57078 800 57094 856
rect 57262 800 57278 856
rect 57446 800 57462 856
rect 57630 800 57646 856
rect 57814 800 57830 856
rect 57998 800 58106 856
rect 58274 800 58290 856
rect 58458 800 58474 856
rect 58642 800 58658 856
rect 58826 800 58842 856
rect 59010 800 59118 856
rect 59286 800 59302 856
rect 59470 800 59486 856
rect 59654 800 59670 856
rect 59838 800 59854 856
rect 60022 800 60130 856
rect 60298 800 60314 856
rect 60482 800 60498 856
rect 60666 800 60682 856
rect 60850 800 60866 856
rect 61034 800 61142 856
rect 61310 800 61326 856
rect 61494 800 61510 856
rect 61678 800 61694 856
rect 61862 800 61878 856
rect 62046 800 62062 856
rect 62230 800 62338 856
rect 62506 800 62522 856
rect 62690 800 62706 856
rect 62874 800 62890 856
rect 63058 800 63074 856
rect 63242 800 63350 856
rect 63518 800 63534 856
rect 63702 800 63718 856
rect 63886 800 63902 856
rect 64070 800 64086 856
rect 64254 800 64362 856
rect 64530 800 64546 856
rect 64714 800 64730 856
rect 64898 800 64914 856
rect 65082 800 65098 856
rect 65266 800 65374 856
rect 65542 800 65558 856
rect 65726 800 65742 856
rect 65910 800 65926 856
rect 66094 800 66110 856
rect 66278 800 66386 856
rect 66554 800 66570 856
rect 66738 800 66754 856
rect 66922 800 66938 856
rect 67106 800 67122 856
rect 67290 800 67306 856
rect 67474 800 67582 856
rect 67750 800 67766 856
rect 67934 800 67950 856
rect 68118 800 68134 856
rect 68302 800 68318 856
rect 68486 800 68594 856
rect 68762 800 68778 856
rect 68946 800 68962 856
rect 69130 800 69146 856
rect 69314 800 69330 856
rect 69498 800 69606 856
rect 69774 800 69790 856
rect 69958 800 69974 856
rect 70142 800 70158 856
rect 70326 800 70342 856
rect 70510 800 70618 856
rect 70786 800 70802 856
rect 70970 800 70986 856
rect 71154 800 71170 856
rect 71338 800 71354 856
rect 71522 800 71538 856
rect 71706 800 71814 856
rect 71982 800 71998 856
rect 72166 800 72182 856
rect 72350 800 72366 856
rect 72534 800 72550 856
rect 72718 800 72826 856
rect 72994 800 73010 856
rect 73178 800 73194 856
rect 73362 800 73378 856
rect 73546 800 73562 856
rect 73730 800 73838 856
rect 74006 800 74022 856
rect 74190 800 74206 856
rect 74374 800 74390 856
rect 74558 800 74574 856
rect 74742 800 74850 856
rect 75018 800 75034 856
rect 75202 800 75218 856
rect 75386 800 75402 856
rect 75570 800 75586 856
rect 75754 800 75862 856
rect 76030 800 76046 856
rect 76214 800 76230 856
rect 76398 800 76414 856
rect 76582 800 76598 856
rect 76766 800 76782 856
rect 76950 800 77058 856
rect 77226 800 77242 856
rect 77410 800 77426 856
rect 77594 800 77610 856
rect 77778 800 77794 856
rect 77962 800 78070 856
rect 78238 800 78254 856
rect 78422 800 78438 856
rect 78606 800 78622 856
rect 78790 800 78806 856
rect 78974 800 79082 856
rect 79250 800 79266 856
rect 79434 800 79450 856
rect 79618 800 79634 856
rect 79802 800 79818 856
rect 79986 800 80094 856
rect 80262 800 80278 856
rect 80446 800 80462 856
rect 80630 800 80646 856
rect 80814 800 80830 856
rect 80998 800 81014 856
rect 81182 800 81290 856
rect 81458 800 81474 856
rect 81642 800 81658 856
rect 81826 800 81842 856
rect 82010 800 82026 856
rect 82194 800 82302 856
rect 82470 800 82486 856
rect 82654 800 82670 856
rect 82838 800 82854 856
rect 83022 800 83038 856
rect 83206 800 83314 856
rect 83482 800 83498 856
rect 83666 800 83682 856
rect 83850 800 83866 856
rect 84034 800 84050 856
rect 84218 800 84326 856
rect 84494 800 84510 856
rect 84678 800 84694 856
rect 84862 800 84878 856
rect 85046 800 85062 856
rect 85230 800 85338 856
rect 85506 800 85522 856
rect 85690 800 85706 856
rect 85874 800 85890 856
rect 86058 800 86074 856
rect 86242 800 86258 856
rect 86426 800 86534 856
rect 86702 800 86718 856
rect 86886 800 86902 856
rect 87070 800 87086 856
rect 87254 800 87270 856
rect 87438 800 87546 856
rect 87714 800 87730 856
rect 87898 800 87914 856
rect 88082 800 88098 856
rect 88266 800 88282 856
rect 88450 800 88558 856
rect 88726 800 88742 856
rect 88910 800 88926 856
rect 89094 800 89110 856
rect 89278 800 89294 856
rect 89462 800 89570 856
rect 89738 800 89754 856
rect 89922 800 89938 856
rect 90106 800 90122 856
rect 90290 800 90306 856
rect 90474 800 90490 856
rect 90658 800 90766 856
rect 90934 800 90950 856
rect 91118 800 91134 856
rect 91302 800 91318 856
rect 91486 800 91502 856
rect 91670 800 91778 856
rect 91946 800 91962 856
rect 92130 800 92146 856
rect 92314 800 92330 856
rect 92498 800 92514 856
rect 92682 800 92790 856
rect 92958 800 92974 856
rect 93142 800 93158 856
rect 93326 800 93342 856
rect 93510 800 93526 856
rect 93694 800 93802 856
rect 93970 800 93986 856
rect 94154 800 94170 856
rect 94338 800 94354 856
rect 94522 800 94538 856
rect 94706 800 94814 856
rect 94982 800 94998 856
rect 95166 800 95182 856
rect 95350 800 95366 856
rect 95534 800 95550 856
rect 95718 800 95734 856
rect 95902 800 96010 856
rect 96178 800 96194 856
rect 96362 800 96378 856
rect 96546 800 96562 856
rect 96730 800 96746 856
rect 96914 800 97022 856
rect 97190 800 97206 856
rect 97374 800 97390 856
rect 97558 800 97574 856
rect 97742 800 97758 856
rect 97926 800 98034 856
rect 98202 800 98218 856
rect 98386 800 98402 856
rect 98570 800 98586 856
rect 98754 800 98770 856
rect 98938 800 99046 856
rect 99214 800 99230 856
rect 99398 800 99414 856
rect 99582 800 99598 856
rect 99766 800 99782 856
<< metal3 >>
rect 0 198840 800 198960
rect 99200 198296 100000 198416
rect 0 196664 800 196784
rect 99200 195168 100000 195288
rect 0 194488 800 194608
rect 0 192312 800 192432
rect 99200 191904 100000 192024
rect 0 190136 800 190256
rect 99200 188776 100000 188896
rect 0 187960 800 188080
rect 0 185784 800 185904
rect 99200 185648 100000 185768
rect 0 183608 800 183728
rect 99200 182384 100000 182504
rect 0 181432 800 181552
rect 0 179256 800 179376
rect 99200 179256 100000 179376
rect 0 177080 800 177200
rect 99200 176128 100000 176248
rect 0 174904 800 175024
rect 0 172728 800 172848
rect 99200 172864 100000 172984
rect 0 170552 800 170672
rect 99200 169736 100000 169856
rect 0 168376 800 168496
rect 99200 166608 100000 166728
rect 0 166200 800 166320
rect 0 164024 800 164144
rect 99200 163344 100000 163464
rect 0 161848 800 161968
rect 99200 160216 100000 160336
rect 0 159672 800 159792
rect 0 157496 800 157616
rect 99200 157088 100000 157208
rect 0 155320 800 155440
rect 99200 153824 100000 153944
rect 0 153144 800 153264
rect 0 150968 800 151088
rect 99200 150696 100000 150816
rect 0 148792 800 148912
rect 99200 147568 100000 147688
rect 0 146616 800 146736
rect 0 144440 800 144560
rect 99200 144304 100000 144424
rect 0 142264 800 142384
rect 99200 141176 100000 141296
rect 0 140088 800 140208
rect 0 137912 800 138032
rect 99200 138048 100000 138168
rect 0 135736 800 135856
rect 99200 134784 100000 134904
rect 0 133560 800 133680
rect 99200 131656 100000 131776
rect 0 131384 800 131504
rect 0 129208 800 129328
rect 99200 128392 100000 128512
rect 0 127032 800 127152
rect 99200 125264 100000 125384
rect 0 124856 800 124976
rect 0 122680 800 122800
rect 99200 122136 100000 122256
rect 0 120504 800 120624
rect 99200 118872 100000 118992
rect 0 118328 800 118448
rect 0 116152 800 116272
rect 99200 115744 100000 115864
rect 0 113976 800 114096
rect 99200 112616 100000 112736
rect 0 111800 800 111920
rect 0 109624 800 109744
rect 99200 109352 100000 109472
rect 0 107448 800 107568
rect 99200 106224 100000 106344
rect 0 105272 800 105392
rect 0 103096 800 103216
rect 99200 103096 100000 103216
rect 0 100920 800 101040
rect 99200 99832 100000 99952
rect 0 98744 800 98864
rect 0 96568 800 96688
rect 99200 96704 100000 96824
rect 0 94392 800 94512
rect 99200 93576 100000 93696
rect 0 92216 800 92336
rect 99200 90312 100000 90432
rect 0 90040 800 90160
rect 0 87864 800 87984
rect 99200 87184 100000 87304
rect 0 85688 800 85808
rect 99200 84056 100000 84176
rect 0 83512 800 83632
rect 0 81336 800 81456
rect 99200 80792 100000 80912
rect 0 79160 800 79280
rect 99200 77664 100000 77784
rect 0 76984 800 77104
rect 0 74808 800 74928
rect 99200 74536 100000 74656
rect 0 72632 800 72752
rect 99200 71272 100000 71392
rect 0 70456 800 70576
rect 0 68280 800 68400
rect 99200 68144 100000 68264
rect 0 66104 800 66224
rect 99200 64880 100000 65000
rect 0 63928 800 64048
rect 0 61752 800 61872
rect 99200 61752 100000 61872
rect 0 59576 800 59696
rect 99200 58624 100000 58744
rect 0 57400 800 57520
rect 0 55224 800 55344
rect 99200 55360 100000 55480
rect 0 53048 800 53168
rect 99200 52232 100000 52352
rect 0 50872 800 50992
rect 99200 49104 100000 49224
rect 0 48696 800 48816
rect 0 46520 800 46640
rect 99200 45840 100000 45960
rect 0 44344 800 44464
rect 99200 42712 100000 42832
rect 0 42168 800 42288
rect 0 39992 800 40112
rect 99200 39584 100000 39704
rect 0 37816 800 37936
rect 99200 36320 100000 36440
rect 0 35640 800 35760
rect 0 33464 800 33584
rect 99200 33192 100000 33312
rect 0 31288 800 31408
rect 99200 30064 100000 30184
rect 0 29112 800 29232
rect 0 26936 800 27056
rect 99200 26800 100000 26920
rect 0 24760 800 24880
rect 99200 23672 100000 23792
rect 0 22584 800 22704
rect 0 20408 800 20528
rect 99200 20544 100000 20664
rect 0 18232 800 18352
rect 99200 17280 100000 17400
rect 0 16056 800 16176
rect 99200 14152 100000 14272
rect 0 13880 800 14000
rect 0 11704 800 11824
rect 99200 11024 100000 11144
rect 0 9528 800 9648
rect 99200 7760 100000 7880
rect 0 7352 800 7472
rect 0 5176 800 5296
rect 99200 4632 100000 4752
rect 0 3000 800 3120
rect 99200 1504 100000 1624
rect 0 960 800 1080
<< obsm3 >>
rect 880 198760 99200 198933
rect 800 198496 99200 198760
rect 800 198216 99120 198496
rect 800 196864 99200 198216
rect 880 196584 99200 196864
rect 800 195368 99200 196584
rect 800 195088 99120 195368
rect 800 194688 99200 195088
rect 880 194408 99200 194688
rect 800 192512 99200 194408
rect 880 192232 99200 192512
rect 800 192104 99200 192232
rect 800 191824 99120 192104
rect 800 190336 99200 191824
rect 880 190056 99200 190336
rect 800 188976 99200 190056
rect 800 188696 99120 188976
rect 800 188160 99200 188696
rect 880 187880 99200 188160
rect 800 185984 99200 187880
rect 880 185848 99200 185984
rect 880 185704 99120 185848
rect 800 185568 99120 185704
rect 800 183808 99200 185568
rect 880 183528 99200 183808
rect 800 182584 99200 183528
rect 800 182304 99120 182584
rect 800 181632 99200 182304
rect 880 181352 99200 181632
rect 800 179456 99200 181352
rect 880 179176 99120 179456
rect 800 177280 99200 179176
rect 880 177000 99200 177280
rect 800 176328 99200 177000
rect 800 176048 99120 176328
rect 800 175104 99200 176048
rect 880 174824 99200 175104
rect 800 173064 99200 174824
rect 800 172928 99120 173064
rect 880 172784 99120 172928
rect 880 172648 99200 172784
rect 800 170752 99200 172648
rect 880 170472 99200 170752
rect 800 169936 99200 170472
rect 800 169656 99120 169936
rect 800 168576 99200 169656
rect 880 168296 99200 168576
rect 800 166808 99200 168296
rect 800 166528 99120 166808
rect 800 166400 99200 166528
rect 880 166120 99200 166400
rect 800 164224 99200 166120
rect 880 163944 99200 164224
rect 800 163544 99200 163944
rect 800 163264 99120 163544
rect 800 162048 99200 163264
rect 880 161768 99200 162048
rect 800 160416 99200 161768
rect 800 160136 99120 160416
rect 800 159872 99200 160136
rect 880 159592 99200 159872
rect 800 157696 99200 159592
rect 880 157416 99200 157696
rect 800 157288 99200 157416
rect 800 157008 99120 157288
rect 800 155520 99200 157008
rect 880 155240 99200 155520
rect 800 154024 99200 155240
rect 800 153744 99120 154024
rect 800 153344 99200 153744
rect 880 153064 99200 153344
rect 800 151168 99200 153064
rect 880 150896 99200 151168
rect 880 150888 99120 150896
rect 800 150616 99120 150888
rect 800 148992 99200 150616
rect 880 148712 99200 148992
rect 800 147768 99200 148712
rect 800 147488 99120 147768
rect 800 146816 99200 147488
rect 880 146536 99200 146816
rect 800 144640 99200 146536
rect 880 144504 99200 144640
rect 880 144360 99120 144504
rect 800 144224 99120 144360
rect 800 142464 99200 144224
rect 880 142184 99200 142464
rect 800 141376 99200 142184
rect 800 141096 99120 141376
rect 800 140288 99200 141096
rect 880 140008 99200 140288
rect 800 138248 99200 140008
rect 800 138112 99120 138248
rect 880 137968 99120 138112
rect 880 137832 99200 137968
rect 800 135936 99200 137832
rect 880 135656 99200 135936
rect 800 134984 99200 135656
rect 800 134704 99120 134984
rect 800 133760 99200 134704
rect 880 133480 99200 133760
rect 800 131856 99200 133480
rect 800 131584 99120 131856
rect 880 131576 99120 131584
rect 880 131304 99200 131576
rect 800 129408 99200 131304
rect 880 129128 99200 129408
rect 800 128592 99200 129128
rect 800 128312 99120 128592
rect 800 127232 99200 128312
rect 880 126952 99200 127232
rect 800 125464 99200 126952
rect 800 125184 99120 125464
rect 800 125056 99200 125184
rect 880 124776 99200 125056
rect 800 122880 99200 124776
rect 880 122600 99200 122880
rect 800 122336 99200 122600
rect 800 122056 99120 122336
rect 800 120704 99200 122056
rect 880 120424 99200 120704
rect 800 119072 99200 120424
rect 800 118792 99120 119072
rect 800 118528 99200 118792
rect 880 118248 99200 118528
rect 800 116352 99200 118248
rect 880 116072 99200 116352
rect 800 115944 99200 116072
rect 800 115664 99120 115944
rect 800 114176 99200 115664
rect 880 113896 99200 114176
rect 800 112816 99200 113896
rect 800 112536 99120 112816
rect 800 112000 99200 112536
rect 880 111720 99200 112000
rect 800 109824 99200 111720
rect 880 109552 99200 109824
rect 880 109544 99120 109552
rect 800 109272 99120 109544
rect 800 107648 99200 109272
rect 880 107368 99200 107648
rect 800 106424 99200 107368
rect 800 106144 99120 106424
rect 800 105472 99200 106144
rect 880 105192 99200 105472
rect 800 103296 99200 105192
rect 880 103016 99120 103296
rect 800 101120 99200 103016
rect 880 100840 99200 101120
rect 800 100032 99200 100840
rect 800 99752 99120 100032
rect 800 98944 99200 99752
rect 880 98664 99200 98944
rect 800 96904 99200 98664
rect 800 96768 99120 96904
rect 880 96624 99120 96768
rect 880 96488 99200 96624
rect 800 94592 99200 96488
rect 880 94312 99200 94592
rect 800 93776 99200 94312
rect 800 93496 99120 93776
rect 800 92416 99200 93496
rect 880 92136 99200 92416
rect 800 90512 99200 92136
rect 800 90240 99120 90512
rect 880 90232 99120 90240
rect 880 89960 99200 90232
rect 800 88064 99200 89960
rect 880 87784 99200 88064
rect 800 87384 99200 87784
rect 800 87104 99120 87384
rect 800 85888 99200 87104
rect 880 85608 99200 85888
rect 800 84256 99200 85608
rect 800 83976 99120 84256
rect 800 83712 99200 83976
rect 880 83432 99200 83712
rect 800 81536 99200 83432
rect 880 81256 99200 81536
rect 800 80992 99200 81256
rect 800 80712 99120 80992
rect 800 79360 99200 80712
rect 880 79080 99200 79360
rect 800 77864 99200 79080
rect 800 77584 99120 77864
rect 800 77184 99200 77584
rect 880 76904 99200 77184
rect 800 75008 99200 76904
rect 880 74736 99200 75008
rect 880 74728 99120 74736
rect 800 74456 99120 74728
rect 800 72832 99200 74456
rect 880 72552 99200 72832
rect 800 71472 99200 72552
rect 800 71192 99120 71472
rect 800 70656 99200 71192
rect 880 70376 99200 70656
rect 800 68480 99200 70376
rect 880 68344 99200 68480
rect 880 68200 99120 68344
rect 800 68064 99120 68200
rect 800 66304 99200 68064
rect 880 66024 99200 66304
rect 800 65080 99200 66024
rect 800 64800 99120 65080
rect 800 64128 99200 64800
rect 880 63848 99200 64128
rect 800 61952 99200 63848
rect 880 61672 99120 61952
rect 800 59776 99200 61672
rect 880 59496 99200 59776
rect 800 58824 99200 59496
rect 800 58544 99120 58824
rect 800 57600 99200 58544
rect 880 57320 99200 57600
rect 800 55560 99200 57320
rect 800 55424 99120 55560
rect 880 55280 99120 55424
rect 880 55144 99200 55280
rect 800 53248 99200 55144
rect 880 52968 99200 53248
rect 800 52432 99200 52968
rect 800 52152 99120 52432
rect 800 51072 99200 52152
rect 880 50792 99200 51072
rect 800 49304 99200 50792
rect 800 49024 99120 49304
rect 800 48896 99200 49024
rect 880 48616 99200 48896
rect 800 46720 99200 48616
rect 880 46440 99200 46720
rect 800 46040 99200 46440
rect 800 45760 99120 46040
rect 800 44544 99200 45760
rect 880 44264 99200 44544
rect 800 42912 99200 44264
rect 800 42632 99120 42912
rect 800 42368 99200 42632
rect 880 42088 99200 42368
rect 800 40192 99200 42088
rect 880 39912 99200 40192
rect 800 39784 99200 39912
rect 800 39504 99120 39784
rect 800 38016 99200 39504
rect 880 37736 99200 38016
rect 800 36520 99200 37736
rect 800 36240 99120 36520
rect 800 35840 99200 36240
rect 880 35560 99200 35840
rect 800 33664 99200 35560
rect 880 33392 99200 33664
rect 880 33384 99120 33392
rect 800 33112 99120 33384
rect 800 31488 99200 33112
rect 880 31208 99200 31488
rect 800 30264 99200 31208
rect 800 29984 99120 30264
rect 800 29312 99200 29984
rect 880 29032 99200 29312
rect 800 27136 99200 29032
rect 880 27000 99200 27136
rect 880 26856 99120 27000
rect 800 26720 99120 26856
rect 800 24960 99200 26720
rect 880 24680 99200 24960
rect 800 23872 99200 24680
rect 800 23592 99120 23872
rect 800 22784 99200 23592
rect 880 22504 99200 22784
rect 800 20744 99200 22504
rect 800 20608 99120 20744
rect 880 20464 99120 20608
rect 880 20328 99200 20464
rect 800 18432 99200 20328
rect 880 18152 99200 18432
rect 800 17480 99200 18152
rect 800 17200 99120 17480
rect 800 16256 99200 17200
rect 880 15976 99200 16256
rect 800 14352 99200 15976
rect 800 14080 99120 14352
rect 880 14072 99120 14080
rect 880 13800 99200 14072
rect 800 11904 99200 13800
rect 880 11624 99200 11904
rect 800 11224 99200 11624
rect 800 10944 99120 11224
rect 800 9728 99200 10944
rect 880 9448 99200 9728
rect 800 7960 99200 9448
rect 800 7680 99120 7960
rect 800 7552 99200 7680
rect 880 7272 99200 7552
rect 800 5376 99200 7272
rect 880 5096 99200 5376
rect 800 4832 99200 5096
rect 800 4552 99120 4832
rect 800 3200 99200 4552
rect 880 2920 99200 3200
rect 800 1704 99200 2920
rect 800 1424 99120 1704
rect 800 1160 99200 1424
rect 880 987 99200 1160
<< metal4 >>
rect 4208 2128 4528 197520
rect 19568 2128 19888 197520
rect 34928 2128 35248 197520
rect 50288 2128 50608 197520
rect 65648 2128 65968 197520
rect 81008 2128 81328 197520
rect 96368 2128 96688 197520
<< obsm4 >>
rect 1715 3299 4128 188325
rect 4608 3299 19488 188325
rect 19968 3299 34848 188325
rect 35328 3299 50173 188325
<< labels >>
rlabel metal2 s 386 199200 442 200000 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 26238 199200 26294 200000 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 28814 199200 28870 200000 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 31390 199200 31446 200000 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 33966 199200 34022 200000 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 36542 199200 36598 200000 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 39118 199200 39174 200000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 41694 199200 41750 200000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 44270 199200 44326 200000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 46938 199200 46994 200000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 49514 199200 49570 200000 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 2962 199200 3018 200000 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 52090 199200 52146 200000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 54666 199200 54722 200000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 57242 199200 57298 200000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 59818 199200 59874 200000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 62394 199200 62450 200000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 64970 199200 65026 200000 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 67546 199200 67602 200000 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 70214 199200 70270 200000 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 72790 199200 72846 200000 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 75366 199200 75422 200000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 5538 199200 5594 200000 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 77942 199200 77998 200000 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 80518 199200 80574 200000 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 83094 199200 83150 200000 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 85670 199200 85726 200000 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 88246 199200 88302 200000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 90822 199200 90878 200000 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 93490 199200 93546 200000 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 96066 199200 96122 200000 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 8114 199200 8170 200000 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 10690 199200 10746 200000 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 13266 199200 13322 200000 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 15842 199200 15898 200000 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 18418 199200 18474 200000 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 20994 199200 21050 200000 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 23662 199200 23718 200000 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 1214 199200 1270 200000 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 27066 199200 27122 200000 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 29642 199200 29698 200000 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 32218 199200 32274 200000 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 34794 199200 34850 200000 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 37370 199200 37426 200000 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 40038 199200 40094 200000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 42614 199200 42670 200000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 45190 199200 45246 200000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 47766 199200 47822 200000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 50342 199200 50398 200000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 3790 199200 3846 200000 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 52918 199200 52974 200000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 55494 199200 55550 200000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 58070 199200 58126 200000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 60646 199200 60702 200000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 63314 199200 63370 200000 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 65890 199200 65946 200000 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 68466 199200 68522 200000 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 71042 199200 71098 200000 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 73618 199200 73674 200000 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 76194 199200 76250 200000 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 6366 199200 6422 200000 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 78770 199200 78826 200000 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 81346 199200 81402 200000 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 83922 199200 83978 200000 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 86590 199200 86646 200000 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 89166 199200 89222 200000 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 91742 199200 91798 200000 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 94318 199200 94374 200000 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 96894 199200 96950 200000 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 8942 199200 8998 200000 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 11518 199200 11574 200000 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 14094 199200 14150 200000 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 16762 199200 16818 200000 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 19338 199200 19394 200000 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 21914 199200 21970 200000 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 24490 199200 24546 200000 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 2042 199200 2098 200000 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 27894 199200 27950 200000 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 30470 199200 30526 200000 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 33138 199200 33194 200000 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 35714 199200 35770 200000 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 38290 199200 38346 200000 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 40866 199200 40922 200000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 43442 199200 43498 200000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 46018 199200 46074 200000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 48594 199200 48650 200000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 51170 199200 51226 200000 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 4618 199200 4674 200000 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 53746 199200 53802 200000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 56414 199200 56470 200000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 58990 199200 59046 200000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 61566 199200 61622 200000 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 64142 199200 64198 200000 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 66718 199200 66774 200000 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 69294 199200 69350 200000 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 71870 199200 71926 200000 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 74446 199200 74502 200000 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 77022 199200 77078 200000 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 7194 199200 7250 200000 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 79690 199200 79746 200000 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 82266 199200 82322 200000 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 84842 199200 84898 200000 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 87418 199200 87474 200000 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 89994 199200 90050 200000 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 92570 199200 92626 200000 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 95146 199200 95202 200000 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 97722 199200 97778 200000 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 9862 199200 9918 200000 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 12438 199200 12494 200000 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 15014 199200 15070 200000 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 17590 199200 17646 200000 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 20166 199200 20222 200000 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 22742 199200 22798 200000 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 25318 199200 25374 200000 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 98826 0 98882 800 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 99102 0 99158 800 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 99286 0 99342 800 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 21454 0 21510 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 81898 0 81954 800 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 82542 0 82598 800 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 83094 0 83150 800 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 83738 0 83794 800 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 84382 0 84438 800 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 84934 0 84990 800 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 85578 0 85634 800 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 86130 0 86186 800 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 86774 0 86830 800 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 87326 0 87382 800 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 27526 0 27582 800 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 87970 0 88026 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 88614 0 88670 800 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 89166 0 89222 800 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 89810 0 89866 800 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 90362 0 90418 800 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 91006 0 91062 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 91558 0 91614 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 92202 0 92258 800 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 92846 0 92902 800 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 93398 0 93454 800 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 28078 0 28134 800 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 94042 0 94098 800 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 94594 0 94650 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 95238 0 95294 800 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 95790 0 95846 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 96434 0 96490 800 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 97078 0 97134 800 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 97630 0 97686 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 98274 0 98330 800 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 28722 0 28778 800 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 29274 0 29330 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 29918 0 29974 800 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 30470 0 30526 800 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 31114 0 31170 800 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 31758 0 31814 800 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 32310 0 32366 800 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 32954 0 33010 800 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 22006 0 22062 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 33506 0 33562 800 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 34150 0 34206 800 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 34702 0 34758 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 35346 0 35402 800 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 35990 0 36046 800 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 36542 0 36598 800 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 37186 0 37242 800 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 37738 0 37794 800 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 38382 0 38438 800 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 38934 0 38990 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 22650 0 22706 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 39578 0 39634 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 40222 0 40278 800 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 40774 0 40830 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 41418 0 41474 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 41970 0 42026 800 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 42614 0 42670 800 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 43166 0 43222 800 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 43810 0 43866 800 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 44454 0 44510 800 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 45006 0 45062 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 23294 0 23350 800 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 45650 0 45706 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 46202 0 46258 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 46846 0 46902 800 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 47490 0 47546 800 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 48042 0 48098 800 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 48686 0 48742 800 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 49238 0 49294 800 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 49882 0 49938 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 50434 0 50490 800 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 51078 0 51134 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 23846 0 23902 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 51722 0 51778 800 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 52274 0 52330 800 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 52918 0 52974 800 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 53470 0 53526 800 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 54114 0 54170 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 54666 0 54722 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 55310 0 55366 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 55954 0 56010 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 56506 0 56562 800 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 57150 0 57206 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 24490 0 24546 800 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 57702 0 57758 800 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 58346 0 58402 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 58898 0 58954 800 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 59542 0 59598 800 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 60186 0 60242 800 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 60738 0 60794 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 61382 0 61438 800 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 61934 0 61990 800 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 62578 0 62634 800 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 63130 0 63186 800 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 25042 0 25098 800 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 63774 0 63830 800 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 64418 0 64474 800 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 64970 0 65026 800 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 65614 0 65670 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 66166 0 66222 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 66810 0 66866 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 67362 0 67418 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 68006 0 68062 800 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 68650 0 68706 800 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 69202 0 69258 800 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 25686 0 25742 800 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 69846 0 69902 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 70398 0 70454 800 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 71042 0 71098 800 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 71594 0 71650 800 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 72238 0 72294 800 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 72882 0 72938 800 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 73434 0 73490 800 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 74078 0 74134 800 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 74630 0 74686 800 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 75274 0 75330 800 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 26238 0 26294 800 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 75918 0 75974 800 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 76470 0 76526 800 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 77114 0 77170 800 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 77666 0 77722 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 78310 0 78366 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 78862 0 78918 800 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 79506 0 79562 800 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 80150 0 80206 800 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 80702 0 80758 800 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 81346 0 81402 800 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 26882 0 26938 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 21638 0 21694 800 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 82082 0 82138 800 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 82726 0 82782 800 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 83370 0 83426 800 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 83922 0 83978 800 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 84566 0 84622 800 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 85118 0 85174 800 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 85762 0 85818 800 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 86314 0 86370 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 86958 0 87014 800 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 87602 0 87658 800 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 27710 0 27766 800 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 88154 0 88210 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 88798 0 88854 800 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 89350 0 89406 800 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 89994 0 90050 800 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 90546 0 90602 800 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 91190 0 91246 800 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 91834 0 91890 800 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 92386 0 92442 800 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 93030 0 93086 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 93582 0 93638 800 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 28262 0 28318 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 94226 0 94282 800 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 94870 0 94926 800 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 95422 0 95478 800 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 96066 0 96122 800 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 96618 0 96674 800 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 97262 0 97318 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 97814 0 97870 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 98458 0 98514 800 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 28906 0 28962 800 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 29458 0 29514 800 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 30102 0 30158 800 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 30746 0 30802 800 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 31298 0 31354 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 31942 0 31998 800 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 32494 0 32550 800 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 33138 0 33194 800 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 22282 0 22338 800 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 33690 0 33746 800 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 34334 0 34390 800 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 34978 0 35034 800 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 35530 0 35586 800 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 36174 0 36230 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 36726 0 36782 800 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 37370 0 37426 800 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 38014 0 38070 800 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 38566 0 38622 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 39210 0 39266 800 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 22834 0 22890 800 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 39762 0 39818 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 40406 0 40462 800 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 40958 0 41014 800 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 41602 0 41658 800 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 42246 0 42302 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 42798 0 42854 800 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 43442 0 43498 800 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 43994 0 44050 800 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 44638 0 44694 800 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 45190 0 45246 800 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 23478 0 23534 800 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 45834 0 45890 800 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 46478 0 46534 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 47030 0 47086 800 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 47674 0 47730 800 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 48226 0 48282 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 48870 0 48926 800 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 49422 0 49478 800 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 50066 0 50122 800 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 50710 0 50766 800 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 51262 0 51318 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 24030 0 24086 800 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 51906 0 51962 800 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 52458 0 52514 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 53102 0 53158 800 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 53654 0 53710 800 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 54298 0 54354 800 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 54942 0 54998 800 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 55494 0 55550 800 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 56138 0 56194 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 56690 0 56746 800 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 57334 0 57390 800 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 24674 0 24730 800 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 57886 0 57942 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 58530 0 58586 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 59174 0 59230 800 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 59726 0 59782 800 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 60370 0 60426 800 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 60922 0 60978 800 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 61566 0 61622 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 62118 0 62174 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 62762 0 62818 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 63406 0 63462 800 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 25226 0 25282 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 63958 0 64014 800 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 64602 0 64658 800 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 65154 0 65210 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 65798 0 65854 800 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 66442 0 66498 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 66994 0 67050 800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 67638 0 67694 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 68190 0 68246 800 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 68834 0 68890 800 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 69386 0 69442 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 25870 0 25926 800 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 70030 0 70086 800 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 70674 0 70730 800 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 71226 0 71282 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 71870 0 71926 800 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 72422 0 72478 800 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 73066 0 73122 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 73618 0 73674 800 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 74262 0 74318 800 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 74906 0 74962 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 75458 0 75514 800 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 26514 0 26570 800 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 76102 0 76158 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 76654 0 76710 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 77298 0 77354 800 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 77850 0 77906 800 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 78494 0 78550 800 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 79138 0 79194 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 79690 0 79746 800 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 80334 0 80390 800 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 80886 0 80942 800 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 81530 0 81586 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 27066 0 27122 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 21822 0 21878 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 82358 0 82414 800 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 82910 0 82966 800 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 83554 0 83610 800 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 84106 0 84162 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 84750 0 84806 800 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 85394 0 85450 800 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 85946 0 86002 800 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 86590 0 86646 800 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 87142 0 87198 800 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 87786 0 87842 800 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 27894 0 27950 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 88338 0 88394 800 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 88982 0 89038 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 89626 0 89682 800 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 90178 0 90234 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 90822 0 90878 800 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 91374 0 91430 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 92018 0 92074 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 92570 0 92626 800 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 93214 0 93270 800 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 93858 0 93914 800 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 28538 0 28594 800 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 94410 0 94466 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 95054 0 95110 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 95606 0 95662 800 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 96250 0 96306 800 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 96802 0 96858 800 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 97446 0 97502 800 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 98090 0 98146 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 98642 0 98698 800 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 29090 0 29146 800 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 29734 0 29790 800 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 30286 0 30342 800 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 30930 0 30986 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 31482 0 31538 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 32126 0 32182 800 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 32770 0 32826 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 33322 0 33378 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 22466 0 22522 800 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 33966 0 34022 800 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 34518 0 34574 800 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 35162 0 35218 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 35714 0 35770 800 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 36358 0 36414 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 37002 0 37058 800 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 37554 0 37610 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 38198 0 38254 800 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 38750 0 38806 800 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 39394 0 39450 800 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 23018 0 23074 800 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 39946 0 40002 800 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 40590 0 40646 800 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 41234 0 41290 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 41786 0 41842 800 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 42430 0 42486 800 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 42982 0 43038 800 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 43626 0 43682 800 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 44178 0 44234 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 44822 0 44878 800 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 45466 0 45522 800 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 23662 0 23718 800 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 46018 0 46074 800 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 46662 0 46718 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 47214 0 47270 800 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 47858 0 47914 800 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 48410 0 48466 800 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 49054 0 49110 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 49698 0 49754 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 50250 0 50306 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 50894 0 50950 800 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 51446 0 51502 800 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 24214 0 24270 800 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 52090 0 52146 800 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 52642 0 52698 800 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 53286 0 53342 800 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 53930 0 53986 800 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 54482 0 54538 800 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 55126 0 55182 800 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 55678 0 55734 800 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 56322 0 56378 800 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 56966 0 57022 800 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 57518 0 57574 800 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 24858 0 24914 800 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 58162 0 58218 800 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 58714 0 58770 800 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 59358 0 59414 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 59910 0 59966 800 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 60554 0 60610 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 61198 0 61254 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 61750 0 61806 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 62394 0 62450 800 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 62946 0 63002 800 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 63590 0 63646 800 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 25502 0 25558 800 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 64142 0 64198 800 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 64786 0 64842 800 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 65430 0 65486 800 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 65982 0 66038 800 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 66626 0 66682 800 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 67178 0 67234 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 67822 0 67878 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 68374 0 68430 800 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 69018 0 69074 800 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 69662 0 69718 800 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 26054 0 26110 800 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 70214 0 70270 800 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 70858 0 70914 800 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 71410 0 71466 800 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 72054 0 72110 800 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 72606 0 72662 800 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 73250 0 73306 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 73894 0 73950 800 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 74446 0 74502 800 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 75090 0 75146 800 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 75642 0 75698 800 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 26698 0 26754 800 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 76286 0 76342 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 76838 0 76894 800 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 77482 0 77538 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 78126 0 78182 800 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 78678 0 78734 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 79322 0 79378 800 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 79874 0 79930 800 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 80518 0 80574 800 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 81070 0 81126 800 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 81714 0 81770 800 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 27250 0 27306 800 6 la_oenb[9]
port 501 nsew signal input
rlabel metal2 s 98642 199200 98698 200000 6 ring0_clk
port 502 nsew signal input
rlabel metal3 s 0 122680 800 122800 6 ring0_clkmux[0]
port 503 nsew signal output
rlabel metal3 s 0 124856 800 124976 6 ring0_clkmux[1]
port 504 nsew signal output
rlabel metal3 s 0 127032 800 127152 6 ring0_clkmux[2]
port 505 nsew signal output
rlabel metal3 s 0 129208 800 129328 6 ring0_start
port 506 nsew signal output
rlabel metal3 s 0 960 800 1080 6 ring0_trim_a[0]
port 507 nsew signal output
rlabel metal3 s 0 22584 800 22704 6 ring0_trim_a[10]
port 508 nsew signal output
rlabel metal3 s 0 24760 800 24880 6 ring0_trim_a[11]
port 509 nsew signal output
rlabel metal3 s 0 26936 800 27056 6 ring0_trim_a[12]
port 510 nsew signal output
rlabel metal3 s 0 29112 800 29232 6 ring0_trim_a[13]
port 511 nsew signal output
rlabel metal3 s 0 31288 800 31408 6 ring0_trim_a[14]
port 512 nsew signal output
rlabel metal3 s 0 33464 800 33584 6 ring0_trim_a[15]
port 513 nsew signal output
rlabel metal3 s 0 35640 800 35760 6 ring0_trim_a[16]
port 514 nsew signal output
rlabel metal3 s 0 37816 800 37936 6 ring0_trim_a[17]
port 515 nsew signal output
rlabel metal3 s 0 39992 800 40112 6 ring0_trim_a[18]
port 516 nsew signal output
rlabel metal3 s 0 42168 800 42288 6 ring0_trim_a[19]
port 517 nsew signal output
rlabel metal3 s 0 3000 800 3120 6 ring0_trim_a[1]
port 518 nsew signal output
rlabel metal3 s 0 44344 800 44464 6 ring0_trim_a[20]
port 519 nsew signal output
rlabel metal3 s 0 46520 800 46640 6 ring0_trim_a[21]
port 520 nsew signal output
rlabel metal3 s 0 48696 800 48816 6 ring0_trim_a[22]
port 521 nsew signal output
rlabel metal3 s 0 50872 800 50992 6 ring0_trim_a[23]
port 522 nsew signal output
rlabel metal3 s 0 53048 800 53168 6 ring0_trim_a[24]
port 523 nsew signal output
rlabel metal3 s 0 55224 800 55344 6 ring0_trim_a[25]
port 524 nsew signal output
rlabel metal3 s 0 57400 800 57520 6 ring0_trim_a[26]
port 525 nsew signal output
rlabel metal3 s 0 59576 800 59696 6 ring0_trim_a[27]
port 526 nsew signal output
rlabel metal3 s 0 5176 800 5296 6 ring0_trim_a[2]
port 527 nsew signal output
rlabel metal3 s 0 7352 800 7472 6 ring0_trim_a[3]
port 528 nsew signal output
rlabel metal3 s 0 9528 800 9648 6 ring0_trim_a[4]
port 529 nsew signal output
rlabel metal3 s 0 11704 800 11824 6 ring0_trim_a[5]
port 530 nsew signal output
rlabel metal3 s 0 13880 800 14000 6 ring0_trim_a[6]
port 531 nsew signal output
rlabel metal3 s 0 16056 800 16176 6 ring0_trim_a[7]
port 532 nsew signal output
rlabel metal3 s 0 18232 800 18352 6 ring0_trim_a[8]
port 533 nsew signal output
rlabel metal3 s 0 20408 800 20528 6 ring0_trim_a[9]
port 534 nsew signal output
rlabel metal3 s 0 61752 800 61872 6 ring0_trim_b[0]
port 535 nsew signal output
rlabel metal3 s 0 83512 800 83632 6 ring0_trim_b[10]
port 536 nsew signal output
rlabel metal3 s 0 85688 800 85808 6 ring0_trim_b[11]
port 537 nsew signal output
rlabel metal3 s 0 87864 800 87984 6 ring0_trim_b[12]
port 538 nsew signal output
rlabel metal3 s 0 90040 800 90160 6 ring0_trim_b[13]
port 539 nsew signal output
rlabel metal3 s 0 92216 800 92336 6 ring0_trim_b[14]
port 540 nsew signal output
rlabel metal3 s 0 94392 800 94512 6 ring0_trim_b[15]
port 541 nsew signal output
rlabel metal3 s 0 96568 800 96688 6 ring0_trim_b[16]
port 542 nsew signal output
rlabel metal3 s 0 98744 800 98864 6 ring0_trim_b[17]
port 543 nsew signal output
rlabel metal3 s 0 100920 800 101040 6 ring0_trim_b[18]
port 544 nsew signal output
rlabel metal3 s 0 103096 800 103216 6 ring0_trim_b[19]
port 545 nsew signal output
rlabel metal3 s 0 63928 800 64048 6 ring0_trim_b[1]
port 546 nsew signal output
rlabel metal3 s 0 105272 800 105392 6 ring0_trim_b[20]
port 547 nsew signal output
rlabel metal3 s 0 107448 800 107568 6 ring0_trim_b[21]
port 548 nsew signal output
rlabel metal3 s 0 109624 800 109744 6 ring0_trim_b[22]
port 549 nsew signal output
rlabel metal3 s 0 111800 800 111920 6 ring0_trim_b[23]
port 550 nsew signal output
rlabel metal3 s 0 113976 800 114096 6 ring0_trim_b[24]
port 551 nsew signal output
rlabel metal3 s 0 116152 800 116272 6 ring0_trim_b[25]
port 552 nsew signal output
rlabel metal3 s 0 118328 800 118448 6 ring0_trim_b[26]
port 553 nsew signal output
rlabel metal3 s 0 120504 800 120624 6 ring0_trim_b[27]
port 554 nsew signal output
rlabel metal3 s 0 66104 800 66224 6 ring0_trim_b[2]
port 555 nsew signal output
rlabel metal3 s 0 68280 800 68400 6 ring0_trim_b[3]
port 556 nsew signal output
rlabel metal3 s 0 70456 800 70576 6 ring0_trim_b[4]
port 557 nsew signal output
rlabel metal3 s 0 72632 800 72752 6 ring0_trim_b[5]
port 558 nsew signal output
rlabel metal3 s 0 74808 800 74928 6 ring0_trim_b[6]
port 559 nsew signal output
rlabel metal3 s 0 76984 800 77104 6 ring0_trim_b[7]
port 560 nsew signal output
rlabel metal3 s 0 79160 800 79280 6 ring0_trim_b[8]
port 561 nsew signal output
rlabel metal3 s 0 81336 800 81456 6 ring0_trim_b[9]
port 562 nsew signal output
rlabel metal2 s 99470 0 99526 800 6 ring1_clk
port 563 nsew signal input
rlabel metal3 s 0 187960 800 188080 6 ring1_clkmux[0]
port 564 nsew signal output
rlabel metal3 s 0 190136 800 190256 6 ring1_clkmux[1]
port 565 nsew signal output
rlabel metal3 s 0 192312 800 192432 6 ring1_clkmux[2]
port 566 nsew signal output
rlabel metal3 s 0 194488 800 194608 6 ring1_start
port 567 nsew signal output
rlabel metal3 s 0 131384 800 131504 6 ring1_trim_a[0]
port 568 nsew signal output
rlabel metal3 s 0 153144 800 153264 6 ring1_trim_a[10]
port 569 nsew signal output
rlabel metal3 s 0 155320 800 155440 6 ring1_trim_a[11]
port 570 nsew signal output
rlabel metal3 s 0 157496 800 157616 6 ring1_trim_a[12]
port 571 nsew signal output
rlabel metal3 s 0 159672 800 159792 6 ring1_trim_a[13]
port 572 nsew signal output
rlabel metal3 s 0 161848 800 161968 6 ring1_trim_a[14]
port 573 nsew signal output
rlabel metal3 s 0 164024 800 164144 6 ring1_trim_a[15]
port 574 nsew signal output
rlabel metal3 s 0 166200 800 166320 6 ring1_trim_a[16]
port 575 nsew signal output
rlabel metal3 s 0 168376 800 168496 6 ring1_trim_a[17]
port 576 nsew signal output
rlabel metal3 s 0 170552 800 170672 6 ring1_trim_a[18]
port 577 nsew signal output
rlabel metal3 s 0 172728 800 172848 6 ring1_trim_a[19]
port 578 nsew signal output
rlabel metal3 s 0 133560 800 133680 6 ring1_trim_a[1]
port 579 nsew signal output
rlabel metal3 s 0 174904 800 175024 6 ring1_trim_a[20]
port 580 nsew signal output
rlabel metal3 s 0 177080 800 177200 6 ring1_trim_a[21]
port 581 nsew signal output
rlabel metal3 s 0 179256 800 179376 6 ring1_trim_a[22]
port 582 nsew signal output
rlabel metal3 s 0 181432 800 181552 6 ring1_trim_a[23]
port 583 nsew signal output
rlabel metal3 s 0 183608 800 183728 6 ring1_trim_a[24]
port 584 nsew signal output
rlabel metal3 s 0 185784 800 185904 6 ring1_trim_a[25]
port 585 nsew signal output
rlabel metal3 s 0 135736 800 135856 6 ring1_trim_a[2]
port 586 nsew signal output
rlabel metal3 s 0 137912 800 138032 6 ring1_trim_a[3]
port 587 nsew signal output
rlabel metal3 s 0 140088 800 140208 6 ring1_trim_a[4]
port 588 nsew signal output
rlabel metal3 s 0 142264 800 142384 6 ring1_trim_a[5]
port 589 nsew signal output
rlabel metal3 s 0 144440 800 144560 6 ring1_trim_a[6]
port 590 nsew signal output
rlabel metal3 s 0 146616 800 146736 6 ring1_trim_a[7]
port 591 nsew signal output
rlabel metal3 s 0 148792 800 148912 6 ring1_trim_a[8]
port 592 nsew signal output
rlabel metal3 s 0 150968 800 151088 6 ring1_trim_a[9]
port 593 nsew signal output
rlabel metal3 s 99200 191904 100000 192024 6 ring2_clk
port 594 nsew signal input
rlabel metal3 s 99200 179256 100000 179376 6 ring2_clkmux[0]
port 595 nsew signal output
rlabel metal3 s 99200 182384 100000 182504 6 ring2_clkmux[1]
port 596 nsew signal output
rlabel metal3 s 99200 185648 100000 185768 6 ring2_clkmux[2]
port 597 nsew signal output
rlabel metal3 s 99200 188776 100000 188896 6 ring2_start
port 598 nsew signal output
rlabel metal3 s 99200 1504 100000 1624 6 ring2_trim_a[0]
port 599 nsew signal output
rlabel metal3 s 99200 33192 100000 33312 6 ring2_trim_a[10]
port 600 nsew signal output
rlabel metal3 s 99200 36320 100000 36440 6 ring2_trim_a[11]
port 601 nsew signal output
rlabel metal3 s 99200 39584 100000 39704 6 ring2_trim_a[12]
port 602 nsew signal output
rlabel metal3 s 99200 42712 100000 42832 6 ring2_trim_a[13]
port 603 nsew signal output
rlabel metal3 s 99200 45840 100000 45960 6 ring2_trim_a[14]
port 604 nsew signal output
rlabel metal3 s 99200 49104 100000 49224 6 ring2_trim_a[15]
port 605 nsew signal output
rlabel metal3 s 99200 52232 100000 52352 6 ring2_trim_a[16]
port 606 nsew signal output
rlabel metal3 s 99200 55360 100000 55480 6 ring2_trim_a[17]
port 607 nsew signal output
rlabel metal3 s 99200 58624 100000 58744 6 ring2_trim_a[18]
port 608 nsew signal output
rlabel metal3 s 99200 61752 100000 61872 6 ring2_trim_a[19]
port 609 nsew signal output
rlabel metal3 s 99200 4632 100000 4752 6 ring2_trim_a[1]
port 610 nsew signal output
rlabel metal3 s 99200 64880 100000 65000 6 ring2_trim_a[20]
port 611 nsew signal output
rlabel metal3 s 99200 68144 100000 68264 6 ring2_trim_a[21]
port 612 nsew signal output
rlabel metal3 s 99200 71272 100000 71392 6 ring2_trim_a[22]
port 613 nsew signal output
rlabel metal3 s 99200 74536 100000 74656 6 ring2_trim_a[23]
port 614 nsew signal output
rlabel metal3 s 99200 77664 100000 77784 6 ring2_trim_a[24]
port 615 nsew signal output
rlabel metal3 s 99200 80792 100000 80912 6 ring2_trim_a[25]
port 616 nsew signal output
rlabel metal3 s 99200 84056 100000 84176 6 ring2_trim_a[26]
port 617 nsew signal output
rlabel metal3 s 99200 87184 100000 87304 6 ring2_trim_a[27]
port 618 nsew signal output
rlabel metal3 s 99200 7760 100000 7880 6 ring2_trim_a[2]
port 619 nsew signal output
rlabel metal3 s 99200 11024 100000 11144 6 ring2_trim_a[3]
port 620 nsew signal output
rlabel metal3 s 99200 14152 100000 14272 6 ring2_trim_a[4]
port 621 nsew signal output
rlabel metal3 s 99200 17280 100000 17400 6 ring2_trim_a[5]
port 622 nsew signal output
rlabel metal3 s 99200 20544 100000 20664 6 ring2_trim_a[6]
port 623 nsew signal output
rlabel metal3 s 99200 23672 100000 23792 6 ring2_trim_a[7]
port 624 nsew signal output
rlabel metal3 s 99200 26800 100000 26920 6 ring2_trim_a[8]
port 625 nsew signal output
rlabel metal3 s 99200 30064 100000 30184 6 ring2_trim_a[9]
port 626 nsew signal output
rlabel metal3 s 99200 90312 100000 90432 6 ring2_trim_b[0]
port 627 nsew signal output
rlabel metal3 s 99200 122136 100000 122256 6 ring2_trim_b[10]
port 628 nsew signal output
rlabel metal3 s 99200 125264 100000 125384 6 ring2_trim_b[11]
port 629 nsew signal output
rlabel metal3 s 99200 128392 100000 128512 6 ring2_trim_b[12]
port 630 nsew signal output
rlabel metal3 s 99200 131656 100000 131776 6 ring2_trim_b[13]
port 631 nsew signal output
rlabel metal3 s 99200 134784 100000 134904 6 ring2_trim_b[14]
port 632 nsew signal output
rlabel metal3 s 99200 138048 100000 138168 6 ring2_trim_b[15]
port 633 nsew signal output
rlabel metal3 s 99200 141176 100000 141296 6 ring2_trim_b[16]
port 634 nsew signal output
rlabel metal3 s 99200 144304 100000 144424 6 ring2_trim_b[17]
port 635 nsew signal output
rlabel metal3 s 99200 147568 100000 147688 6 ring2_trim_b[18]
port 636 nsew signal output
rlabel metal3 s 99200 150696 100000 150816 6 ring2_trim_b[19]
port 637 nsew signal output
rlabel metal3 s 99200 93576 100000 93696 6 ring2_trim_b[1]
port 638 nsew signal output
rlabel metal3 s 99200 153824 100000 153944 6 ring2_trim_b[20]
port 639 nsew signal output
rlabel metal3 s 99200 157088 100000 157208 6 ring2_trim_b[21]
port 640 nsew signal output
rlabel metal3 s 99200 160216 100000 160336 6 ring2_trim_b[22]
port 641 nsew signal output
rlabel metal3 s 99200 163344 100000 163464 6 ring2_trim_b[23]
port 642 nsew signal output
rlabel metal3 s 99200 166608 100000 166728 6 ring2_trim_b[24]
port 643 nsew signal output
rlabel metal3 s 99200 169736 100000 169856 6 ring2_trim_b[25]
port 644 nsew signal output
rlabel metal3 s 99200 172864 100000 172984 6 ring2_trim_b[26]
port 645 nsew signal output
rlabel metal3 s 99200 176128 100000 176248 6 ring2_trim_b[27]
port 646 nsew signal output
rlabel metal3 s 99200 96704 100000 96824 6 ring2_trim_b[2]
port 647 nsew signal output
rlabel metal3 s 99200 99832 100000 99952 6 ring2_trim_b[3]
port 648 nsew signal output
rlabel metal3 s 99200 103096 100000 103216 6 ring2_trim_b[4]
port 649 nsew signal output
rlabel metal3 s 99200 106224 100000 106344 6 ring2_trim_b[5]
port 650 nsew signal output
rlabel metal3 s 99200 109352 100000 109472 6 ring2_trim_b[6]
port 651 nsew signal output
rlabel metal3 s 99200 112616 100000 112736 6 ring2_trim_b[7]
port 652 nsew signal output
rlabel metal3 s 99200 115744 100000 115864 6 ring2_trim_b[8]
port 653 nsew signal output
rlabel metal3 s 99200 118872 100000 118992 6 ring2_trim_b[9]
port 654 nsew signal output
rlabel metal3 s 0 196664 800 196784 6 ring3_clk
port 655 nsew signal input
rlabel metal2 s 99470 199200 99526 200000 6 ring4_clk
port 656 nsew signal input
rlabel metal3 s 0 198840 800 198960 6 ring5_clk
port 657 nsew signal input
rlabel metal3 s 99200 195168 100000 195288 6 ring6_clk
port 658 nsew signal input
rlabel metal3 s 99200 198296 100000 198416 6 ring7_clk
port 659 nsew signal input
rlabel metal2 s 99654 0 99710 800 6 ring8_clk
port 660 nsew signal input
rlabel metal2 s 99838 0 99894 800 6 ring9_clk
port 661 nsew signal input
rlabel metal4 s 4208 2128 4528 197520 6 vccd1
port 662 nsew power input
rlabel metal4 s 34928 2128 35248 197520 6 vccd1
port 662 nsew power input
rlabel metal4 s 65648 2128 65968 197520 6 vccd1
port 662 nsew power input
rlabel metal4 s 96368 2128 96688 197520 6 vccd1
port 662 nsew power input
rlabel metal4 s 19568 2128 19888 197520 6 vssd1
port 663 nsew ground input
rlabel metal4 s 50288 2128 50608 197520 6 vssd1
port 663 nsew ground input
rlabel metal4 s 81008 2128 81328 197520 6 vssd1
port 663 nsew ground input
rlabel metal2 s 110 0 166 800 6 wb_clk_i
port 664 nsew signal input
rlabel metal2 s 294 0 350 800 6 wb_rst_i
port 665 nsew signal input
rlabel metal2 s 478 0 534 800 6 wbs_ack_o
port 666 nsew signal output
rlabel metal2 s 1306 0 1362 800 6 wbs_adr_i[0]
port 667 nsew signal input
rlabel metal2 s 8114 0 8170 800 6 wbs_adr_i[10]
port 668 nsew signal input
rlabel metal2 s 8758 0 8814 800 6 wbs_adr_i[11]
port 669 nsew signal input
rlabel metal2 s 9310 0 9366 800 6 wbs_adr_i[12]
port 670 nsew signal input
rlabel metal2 s 9954 0 10010 800 6 wbs_adr_i[13]
port 671 nsew signal input
rlabel metal2 s 10506 0 10562 800 6 wbs_adr_i[14]
port 672 nsew signal input
rlabel metal2 s 11150 0 11206 800 6 wbs_adr_i[15]
port 673 nsew signal input
rlabel metal2 s 11794 0 11850 800 6 wbs_adr_i[16]
port 674 nsew signal input
rlabel metal2 s 12346 0 12402 800 6 wbs_adr_i[17]
port 675 nsew signal input
rlabel metal2 s 12990 0 13046 800 6 wbs_adr_i[18]
port 676 nsew signal input
rlabel metal2 s 13542 0 13598 800 6 wbs_adr_i[19]
port 677 nsew signal input
rlabel metal2 s 2042 0 2098 800 6 wbs_adr_i[1]
port 678 nsew signal input
rlabel metal2 s 14186 0 14242 800 6 wbs_adr_i[20]
port 679 nsew signal input
rlabel metal2 s 14738 0 14794 800 6 wbs_adr_i[21]
port 680 nsew signal input
rlabel metal2 s 15382 0 15438 800 6 wbs_adr_i[22]
port 681 nsew signal input
rlabel metal2 s 16026 0 16082 800 6 wbs_adr_i[23]
port 682 nsew signal input
rlabel metal2 s 16578 0 16634 800 6 wbs_adr_i[24]
port 683 nsew signal input
rlabel metal2 s 17222 0 17278 800 6 wbs_adr_i[25]
port 684 nsew signal input
rlabel metal2 s 17774 0 17830 800 6 wbs_adr_i[26]
port 685 nsew signal input
rlabel metal2 s 18418 0 18474 800 6 wbs_adr_i[27]
port 686 nsew signal input
rlabel metal2 s 19062 0 19118 800 6 wbs_adr_i[28]
port 687 nsew signal input
rlabel metal2 s 19614 0 19670 800 6 wbs_adr_i[29]
port 688 nsew signal input
rlabel metal2 s 2870 0 2926 800 6 wbs_adr_i[2]
port 689 nsew signal input
rlabel metal2 s 20258 0 20314 800 6 wbs_adr_i[30]
port 690 nsew signal input
rlabel metal2 s 20810 0 20866 800 6 wbs_adr_i[31]
port 691 nsew signal input
rlabel metal2 s 3698 0 3754 800 6 wbs_adr_i[3]
port 692 nsew signal input
rlabel metal2 s 4526 0 4582 800 6 wbs_adr_i[4]
port 693 nsew signal input
rlabel metal2 s 5078 0 5134 800 6 wbs_adr_i[5]
port 694 nsew signal input
rlabel metal2 s 5722 0 5778 800 6 wbs_adr_i[6]
port 695 nsew signal input
rlabel metal2 s 6274 0 6330 800 6 wbs_adr_i[7]
port 696 nsew signal input
rlabel metal2 s 6918 0 6974 800 6 wbs_adr_i[8]
port 697 nsew signal input
rlabel metal2 s 7562 0 7618 800 6 wbs_adr_i[9]
port 698 nsew signal input
rlabel metal2 s 662 0 718 800 6 wbs_cyc_i
port 699 nsew signal input
rlabel metal2 s 1490 0 1546 800 6 wbs_dat_i[0]
port 700 nsew signal input
rlabel metal2 s 8298 0 8354 800 6 wbs_dat_i[10]
port 701 nsew signal input
rlabel metal2 s 8942 0 8998 800 6 wbs_dat_i[11]
port 702 nsew signal input
rlabel metal2 s 9586 0 9642 800 6 wbs_dat_i[12]
port 703 nsew signal input
rlabel metal2 s 10138 0 10194 800 6 wbs_dat_i[13]
port 704 nsew signal input
rlabel metal2 s 10782 0 10838 800 6 wbs_dat_i[14]
port 705 nsew signal input
rlabel metal2 s 11334 0 11390 800 6 wbs_dat_i[15]
port 706 nsew signal input
rlabel metal2 s 11978 0 12034 800 6 wbs_dat_i[16]
port 707 nsew signal input
rlabel metal2 s 12530 0 12586 800 6 wbs_dat_i[17]
port 708 nsew signal input
rlabel metal2 s 13174 0 13230 800 6 wbs_dat_i[18]
port 709 nsew signal input
rlabel metal2 s 13818 0 13874 800 6 wbs_dat_i[19]
port 710 nsew signal input
rlabel metal2 s 2318 0 2374 800 6 wbs_dat_i[1]
port 711 nsew signal input
rlabel metal2 s 14370 0 14426 800 6 wbs_dat_i[20]
port 712 nsew signal input
rlabel metal2 s 15014 0 15070 800 6 wbs_dat_i[21]
port 713 nsew signal input
rlabel metal2 s 15566 0 15622 800 6 wbs_dat_i[22]
port 714 nsew signal input
rlabel metal2 s 16210 0 16266 800 6 wbs_dat_i[23]
port 715 nsew signal input
rlabel metal2 s 16762 0 16818 800 6 wbs_dat_i[24]
port 716 nsew signal input
rlabel metal2 s 17406 0 17462 800 6 wbs_dat_i[25]
port 717 nsew signal input
rlabel metal2 s 18050 0 18106 800 6 wbs_dat_i[26]
port 718 nsew signal input
rlabel metal2 s 18602 0 18658 800 6 wbs_dat_i[27]
port 719 nsew signal input
rlabel metal2 s 19246 0 19302 800 6 wbs_dat_i[28]
port 720 nsew signal input
rlabel metal2 s 19798 0 19854 800 6 wbs_dat_i[29]
port 721 nsew signal input
rlabel metal2 s 3054 0 3110 800 6 wbs_dat_i[2]
port 722 nsew signal input
rlabel metal2 s 20442 0 20498 800 6 wbs_dat_i[30]
port 723 nsew signal input
rlabel metal2 s 20994 0 21050 800 6 wbs_dat_i[31]
port 724 nsew signal input
rlabel metal2 s 3882 0 3938 800 6 wbs_dat_i[3]
port 725 nsew signal input
rlabel metal2 s 4710 0 4766 800 6 wbs_dat_i[4]
port 726 nsew signal input
rlabel metal2 s 5262 0 5318 800 6 wbs_dat_i[5]
port 727 nsew signal input
rlabel metal2 s 5906 0 5962 800 6 wbs_dat_i[6]
port 728 nsew signal input
rlabel metal2 s 6550 0 6606 800 6 wbs_dat_i[7]
port 729 nsew signal input
rlabel metal2 s 7102 0 7158 800 6 wbs_dat_i[8]
port 730 nsew signal input
rlabel metal2 s 7746 0 7802 800 6 wbs_dat_i[9]
port 731 nsew signal input
rlabel metal2 s 1674 0 1730 800 6 wbs_dat_o[0]
port 732 nsew signal output
rlabel metal2 s 8574 0 8630 800 6 wbs_dat_o[10]
port 733 nsew signal output
rlabel metal2 s 9126 0 9182 800 6 wbs_dat_o[11]
port 734 nsew signal output
rlabel metal2 s 9770 0 9826 800 6 wbs_dat_o[12]
port 735 nsew signal output
rlabel metal2 s 10322 0 10378 800 6 wbs_dat_o[13]
port 736 nsew signal output
rlabel metal2 s 10966 0 11022 800 6 wbs_dat_o[14]
port 737 nsew signal output
rlabel metal2 s 11518 0 11574 800 6 wbs_dat_o[15]
port 738 nsew signal output
rlabel metal2 s 12162 0 12218 800 6 wbs_dat_o[16]
port 739 nsew signal output
rlabel metal2 s 12806 0 12862 800 6 wbs_dat_o[17]
port 740 nsew signal output
rlabel metal2 s 13358 0 13414 800 6 wbs_dat_o[18]
port 741 nsew signal output
rlabel metal2 s 14002 0 14058 800 6 wbs_dat_o[19]
port 742 nsew signal output
rlabel metal2 s 2502 0 2558 800 6 wbs_dat_o[1]
port 743 nsew signal output
rlabel metal2 s 14554 0 14610 800 6 wbs_dat_o[20]
port 744 nsew signal output
rlabel metal2 s 15198 0 15254 800 6 wbs_dat_o[21]
port 745 nsew signal output
rlabel metal2 s 15750 0 15806 800 6 wbs_dat_o[22]
port 746 nsew signal output
rlabel metal2 s 16394 0 16450 800 6 wbs_dat_o[23]
port 747 nsew signal output
rlabel metal2 s 17038 0 17094 800 6 wbs_dat_o[24]
port 748 nsew signal output
rlabel metal2 s 17590 0 17646 800 6 wbs_dat_o[25]
port 749 nsew signal output
rlabel metal2 s 18234 0 18290 800 6 wbs_dat_o[26]
port 750 nsew signal output
rlabel metal2 s 18786 0 18842 800 6 wbs_dat_o[27]
port 751 nsew signal output
rlabel metal2 s 19430 0 19486 800 6 wbs_dat_o[28]
port 752 nsew signal output
rlabel metal2 s 19982 0 20038 800 6 wbs_dat_o[29]
port 753 nsew signal output
rlabel metal2 s 3330 0 3386 800 6 wbs_dat_o[2]
port 754 nsew signal output
rlabel metal2 s 20626 0 20682 800 6 wbs_dat_o[30]
port 755 nsew signal output
rlabel metal2 s 21270 0 21326 800 6 wbs_dat_o[31]
port 756 nsew signal output
rlabel metal2 s 4066 0 4122 800 6 wbs_dat_o[3]
port 757 nsew signal output
rlabel metal2 s 4894 0 4950 800 6 wbs_dat_o[4]
port 758 nsew signal output
rlabel metal2 s 5538 0 5594 800 6 wbs_dat_o[5]
port 759 nsew signal output
rlabel metal2 s 6090 0 6146 800 6 wbs_dat_o[6]
port 760 nsew signal output
rlabel metal2 s 6734 0 6790 800 6 wbs_dat_o[7]
port 761 nsew signal output
rlabel metal2 s 7286 0 7342 800 6 wbs_dat_o[8]
port 762 nsew signal output
rlabel metal2 s 7930 0 7986 800 6 wbs_dat_o[9]
port 763 nsew signal output
rlabel metal2 s 1858 0 1914 800 6 wbs_sel_i[0]
port 764 nsew signal input
rlabel metal2 s 2686 0 2742 800 6 wbs_sel_i[1]
port 765 nsew signal input
rlabel metal2 s 3514 0 3570 800 6 wbs_sel_i[2]
port 766 nsew signal input
rlabel metal2 s 4342 0 4398 800 6 wbs_sel_i[3]
port 767 nsew signal input
rlabel metal2 s 846 0 902 800 6 wbs_stb_i
port 768 nsew signal input
rlabel metal2 s 1030 0 1086 800 6 wbs_we_i
port 769 nsew signal input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 100000 200000
string LEFview TRUE
string GDS_FILE /project/openlane/digitalcore_macro/runs/digitalcore_macro/results/magic/digitalcore_macro.gds
string GDS_END 24103584
string GDS_START 756152
<< end >>

