magic
tech sky130A
magscale 1 2
timestamp 1636592110
<< obsli1 >>
rect 1104 2159 98963 197489
<< obsm1 >>
rect 14 1300 99898 197520
<< metal2 >>
rect 386 199200 442 200000
rect 1214 199200 1270 200000
rect 2134 199200 2190 200000
rect 2962 199200 3018 200000
rect 3882 199200 3938 200000
rect 4710 199200 4766 200000
rect 5630 199200 5686 200000
rect 6458 199200 6514 200000
rect 7378 199200 7434 200000
rect 8206 199200 8262 200000
rect 9126 199200 9182 200000
rect 9954 199200 10010 200000
rect 10874 199200 10930 200000
rect 11702 199200 11758 200000
rect 12622 199200 12678 200000
rect 13542 199200 13598 200000
rect 14370 199200 14426 200000
rect 15290 199200 15346 200000
rect 16118 199200 16174 200000
rect 17038 199200 17094 200000
rect 17866 199200 17922 200000
rect 18786 199200 18842 200000
rect 19614 199200 19670 200000
rect 20534 199200 20590 200000
rect 21362 199200 21418 200000
rect 22282 199200 22338 200000
rect 23110 199200 23166 200000
rect 24030 199200 24086 200000
rect 24858 199200 24914 200000
rect 25778 199200 25834 200000
rect 26698 199200 26754 200000
rect 27526 199200 27582 200000
rect 28446 199200 28502 200000
rect 29274 199200 29330 200000
rect 30194 199200 30250 200000
rect 31022 199200 31078 200000
rect 31942 199200 31998 200000
rect 32770 199200 32826 200000
rect 33690 199200 33746 200000
rect 34518 199200 34574 200000
rect 35438 199200 35494 200000
rect 36266 199200 36322 200000
rect 37186 199200 37242 200000
rect 38106 199200 38162 200000
rect 38934 199200 38990 200000
rect 39854 199200 39910 200000
rect 40682 199200 40738 200000
rect 41602 199200 41658 200000
rect 42430 199200 42486 200000
rect 43350 199200 43406 200000
rect 44178 199200 44234 200000
rect 45098 199200 45154 200000
rect 45926 199200 45982 200000
rect 46846 199200 46902 200000
rect 47674 199200 47730 200000
rect 48594 199200 48650 200000
rect 49422 199200 49478 200000
rect 50342 199200 50398 200000
rect 51262 199200 51318 200000
rect 52090 199200 52146 200000
rect 53010 199200 53066 200000
rect 53838 199200 53894 200000
rect 54758 199200 54814 200000
rect 55586 199200 55642 200000
rect 56506 199200 56562 200000
rect 57334 199200 57390 200000
rect 58254 199200 58310 200000
rect 59082 199200 59138 200000
rect 60002 199200 60058 200000
rect 60830 199200 60886 200000
rect 61750 199200 61806 200000
rect 62578 199200 62634 200000
rect 63498 199200 63554 200000
rect 64418 199200 64474 200000
rect 65246 199200 65302 200000
rect 66166 199200 66222 200000
rect 66994 199200 67050 200000
rect 67914 199200 67970 200000
rect 68742 199200 68798 200000
rect 69662 199200 69718 200000
rect 70490 199200 70546 200000
rect 71410 199200 71466 200000
rect 72238 199200 72294 200000
rect 73158 199200 73214 200000
rect 73986 199200 74042 200000
rect 74906 199200 74962 200000
rect 75826 199200 75882 200000
rect 76654 199200 76710 200000
rect 77574 199200 77630 200000
rect 78402 199200 78458 200000
rect 79322 199200 79378 200000
rect 80150 199200 80206 200000
rect 81070 199200 81126 200000
rect 81898 199200 81954 200000
rect 82818 199200 82874 200000
rect 83646 199200 83702 200000
rect 84566 199200 84622 200000
rect 85394 199200 85450 200000
rect 86314 199200 86370 200000
rect 87142 199200 87198 200000
rect 88062 199200 88118 200000
rect 88982 199200 89038 200000
rect 89810 199200 89866 200000
rect 90730 199200 90786 200000
rect 91558 199200 91614 200000
rect 92478 199200 92534 200000
rect 93306 199200 93362 200000
rect 94226 199200 94282 200000
rect 95054 199200 95110 200000
rect 95974 199200 96030 200000
rect 96802 199200 96858 200000
rect 97722 199200 97778 200000
rect 98550 199200 98606 200000
rect 99470 199200 99526 200000
rect 110 0 166 800
rect 294 0 350 800
rect 478 0 534 800
rect 662 0 718 800
rect 846 0 902 800
rect 1122 0 1178 800
rect 1306 0 1362 800
rect 1490 0 1546 800
rect 1674 0 1730 800
rect 1858 0 1914 800
rect 2134 0 2190 800
rect 2318 0 2374 800
rect 2502 0 2558 800
rect 2686 0 2742 800
rect 2870 0 2926 800
rect 3146 0 3202 800
rect 3330 0 3386 800
rect 3514 0 3570 800
rect 3698 0 3754 800
rect 3882 0 3938 800
rect 4158 0 4214 800
rect 4342 0 4398 800
rect 4526 0 4582 800
rect 4710 0 4766 800
rect 4894 0 4950 800
rect 5170 0 5226 800
rect 5354 0 5410 800
rect 5538 0 5594 800
rect 5722 0 5778 800
rect 5906 0 5962 800
rect 6182 0 6238 800
rect 6366 0 6422 800
rect 6550 0 6606 800
rect 6734 0 6790 800
rect 6918 0 6974 800
rect 7194 0 7250 800
rect 7378 0 7434 800
rect 7562 0 7618 800
rect 7746 0 7802 800
rect 7930 0 7986 800
rect 8206 0 8262 800
rect 8390 0 8446 800
rect 8574 0 8630 800
rect 8758 0 8814 800
rect 8942 0 8998 800
rect 9218 0 9274 800
rect 9402 0 9458 800
rect 9586 0 9642 800
rect 9770 0 9826 800
rect 9954 0 10010 800
rect 10230 0 10286 800
rect 10414 0 10470 800
rect 10598 0 10654 800
rect 10782 0 10838 800
rect 10966 0 11022 800
rect 11242 0 11298 800
rect 11426 0 11482 800
rect 11610 0 11666 800
rect 11794 0 11850 800
rect 11978 0 12034 800
rect 12254 0 12310 800
rect 12438 0 12494 800
rect 12622 0 12678 800
rect 12806 0 12862 800
rect 12990 0 13046 800
rect 13266 0 13322 800
rect 13450 0 13506 800
rect 13634 0 13690 800
rect 13818 0 13874 800
rect 14002 0 14058 800
rect 14278 0 14334 800
rect 14462 0 14518 800
rect 14646 0 14702 800
rect 14830 0 14886 800
rect 15014 0 15070 800
rect 15290 0 15346 800
rect 15474 0 15530 800
rect 15658 0 15714 800
rect 15842 0 15898 800
rect 16026 0 16082 800
rect 16302 0 16358 800
rect 16486 0 16542 800
rect 16670 0 16726 800
rect 16854 0 16910 800
rect 17038 0 17094 800
rect 17314 0 17370 800
rect 17498 0 17554 800
rect 17682 0 17738 800
rect 17866 0 17922 800
rect 18050 0 18106 800
rect 18326 0 18382 800
rect 18510 0 18566 800
rect 18694 0 18750 800
rect 18878 0 18934 800
rect 19062 0 19118 800
rect 19338 0 19394 800
rect 19522 0 19578 800
rect 19706 0 19762 800
rect 19890 0 19946 800
rect 20074 0 20130 800
rect 20350 0 20406 800
rect 20534 0 20590 800
rect 20718 0 20774 800
rect 20902 0 20958 800
rect 21086 0 21142 800
rect 21362 0 21418 800
rect 21546 0 21602 800
rect 21730 0 21786 800
rect 21914 0 21970 800
rect 22098 0 22154 800
rect 22374 0 22430 800
rect 22558 0 22614 800
rect 22742 0 22798 800
rect 22926 0 22982 800
rect 23110 0 23166 800
rect 23386 0 23442 800
rect 23570 0 23626 800
rect 23754 0 23810 800
rect 23938 0 23994 800
rect 24122 0 24178 800
rect 24398 0 24454 800
rect 24582 0 24638 800
rect 24766 0 24822 800
rect 24950 0 25006 800
rect 25134 0 25190 800
rect 25410 0 25466 800
rect 25594 0 25650 800
rect 25778 0 25834 800
rect 25962 0 26018 800
rect 26146 0 26202 800
rect 26422 0 26478 800
rect 26606 0 26662 800
rect 26790 0 26846 800
rect 26974 0 27030 800
rect 27158 0 27214 800
rect 27434 0 27490 800
rect 27618 0 27674 800
rect 27802 0 27858 800
rect 27986 0 28042 800
rect 28170 0 28226 800
rect 28446 0 28502 800
rect 28630 0 28686 800
rect 28814 0 28870 800
rect 28998 0 29054 800
rect 29182 0 29238 800
rect 29458 0 29514 800
rect 29642 0 29698 800
rect 29826 0 29882 800
rect 30010 0 30066 800
rect 30194 0 30250 800
rect 30470 0 30526 800
rect 30654 0 30710 800
rect 30838 0 30894 800
rect 31022 0 31078 800
rect 31206 0 31262 800
rect 31482 0 31538 800
rect 31666 0 31722 800
rect 31850 0 31906 800
rect 32034 0 32090 800
rect 32218 0 32274 800
rect 32494 0 32550 800
rect 32678 0 32734 800
rect 32862 0 32918 800
rect 33046 0 33102 800
rect 33230 0 33286 800
rect 33506 0 33562 800
rect 33690 0 33746 800
rect 33874 0 33930 800
rect 34058 0 34114 800
rect 34242 0 34298 800
rect 34518 0 34574 800
rect 34702 0 34758 800
rect 34886 0 34942 800
rect 35070 0 35126 800
rect 35254 0 35310 800
rect 35530 0 35586 800
rect 35714 0 35770 800
rect 35898 0 35954 800
rect 36082 0 36138 800
rect 36266 0 36322 800
rect 36542 0 36598 800
rect 36726 0 36782 800
rect 36910 0 36966 800
rect 37094 0 37150 800
rect 37278 0 37334 800
rect 37554 0 37610 800
rect 37738 0 37794 800
rect 37922 0 37978 800
rect 38106 0 38162 800
rect 38290 0 38346 800
rect 38566 0 38622 800
rect 38750 0 38806 800
rect 38934 0 38990 800
rect 39118 0 39174 800
rect 39302 0 39358 800
rect 39578 0 39634 800
rect 39762 0 39818 800
rect 39946 0 40002 800
rect 40130 0 40186 800
rect 40314 0 40370 800
rect 40590 0 40646 800
rect 40774 0 40830 800
rect 40958 0 41014 800
rect 41142 0 41198 800
rect 41326 0 41382 800
rect 41602 0 41658 800
rect 41786 0 41842 800
rect 41970 0 42026 800
rect 42154 0 42210 800
rect 42338 0 42394 800
rect 42614 0 42670 800
rect 42798 0 42854 800
rect 42982 0 43038 800
rect 43166 0 43222 800
rect 43350 0 43406 800
rect 43626 0 43682 800
rect 43810 0 43866 800
rect 43994 0 44050 800
rect 44178 0 44234 800
rect 44362 0 44418 800
rect 44638 0 44694 800
rect 44822 0 44878 800
rect 45006 0 45062 800
rect 45190 0 45246 800
rect 45374 0 45430 800
rect 45650 0 45706 800
rect 45834 0 45890 800
rect 46018 0 46074 800
rect 46202 0 46258 800
rect 46386 0 46442 800
rect 46662 0 46718 800
rect 46846 0 46902 800
rect 47030 0 47086 800
rect 47214 0 47270 800
rect 47398 0 47454 800
rect 47674 0 47730 800
rect 47858 0 47914 800
rect 48042 0 48098 800
rect 48226 0 48282 800
rect 48410 0 48466 800
rect 48686 0 48742 800
rect 48870 0 48926 800
rect 49054 0 49110 800
rect 49238 0 49294 800
rect 49422 0 49478 800
rect 49698 0 49754 800
rect 49882 0 49938 800
rect 50066 0 50122 800
rect 50250 0 50306 800
rect 50434 0 50490 800
rect 50710 0 50766 800
rect 50894 0 50950 800
rect 51078 0 51134 800
rect 51262 0 51318 800
rect 51446 0 51502 800
rect 51722 0 51778 800
rect 51906 0 51962 800
rect 52090 0 52146 800
rect 52274 0 52330 800
rect 52458 0 52514 800
rect 52734 0 52790 800
rect 52918 0 52974 800
rect 53102 0 53158 800
rect 53286 0 53342 800
rect 53470 0 53526 800
rect 53746 0 53802 800
rect 53930 0 53986 800
rect 54114 0 54170 800
rect 54298 0 54354 800
rect 54482 0 54538 800
rect 54758 0 54814 800
rect 54942 0 54998 800
rect 55126 0 55182 800
rect 55310 0 55366 800
rect 55494 0 55550 800
rect 55770 0 55826 800
rect 55954 0 56010 800
rect 56138 0 56194 800
rect 56322 0 56378 800
rect 56506 0 56562 800
rect 56782 0 56838 800
rect 56966 0 57022 800
rect 57150 0 57206 800
rect 57334 0 57390 800
rect 57518 0 57574 800
rect 57794 0 57850 800
rect 57978 0 58034 800
rect 58162 0 58218 800
rect 58346 0 58402 800
rect 58530 0 58586 800
rect 58806 0 58862 800
rect 58990 0 59046 800
rect 59174 0 59230 800
rect 59358 0 59414 800
rect 59542 0 59598 800
rect 59818 0 59874 800
rect 60002 0 60058 800
rect 60186 0 60242 800
rect 60370 0 60426 800
rect 60554 0 60610 800
rect 60830 0 60886 800
rect 61014 0 61070 800
rect 61198 0 61254 800
rect 61382 0 61438 800
rect 61566 0 61622 800
rect 61842 0 61898 800
rect 62026 0 62082 800
rect 62210 0 62266 800
rect 62394 0 62450 800
rect 62578 0 62634 800
rect 62854 0 62910 800
rect 63038 0 63094 800
rect 63222 0 63278 800
rect 63406 0 63462 800
rect 63590 0 63646 800
rect 63866 0 63922 800
rect 64050 0 64106 800
rect 64234 0 64290 800
rect 64418 0 64474 800
rect 64602 0 64658 800
rect 64878 0 64934 800
rect 65062 0 65118 800
rect 65246 0 65302 800
rect 65430 0 65486 800
rect 65614 0 65670 800
rect 65890 0 65946 800
rect 66074 0 66130 800
rect 66258 0 66314 800
rect 66442 0 66498 800
rect 66626 0 66682 800
rect 66902 0 66958 800
rect 67086 0 67142 800
rect 67270 0 67326 800
rect 67454 0 67510 800
rect 67638 0 67694 800
rect 67914 0 67970 800
rect 68098 0 68154 800
rect 68282 0 68338 800
rect 68466 0 68522 800
rect 68650 0 68706 800
rect 68926 0 68982 800
rect 69110 0 69166 800
rect 69294 0 69350 800
rect 69478 0 69534 800
rect 69662 0 69718 800
rect 69938 0 69994 800
rect 70122 0 70178 800
rect 70306 0 70362 800
rect 70490 0 70546 800
rect 70674 0 70730 800
rect 70950 0 71006 800
rect 71134 0 71190 800
rect 71318 0 71374 800
rect 71502 0 71558 800
rect 71686 0 71742 800
rect 71962 0 72018 800
rect 72146 0 72202 800
rect 72330 0 72386 800
rect 72514 0 72570 800
rect 72698 0 72754 800
rect 72974 0 73030 800
rect 73158 0 73214 800
rect 73342 0 73398 800
rect 73526 0 73582 800
rect 73710 0 73766 800
rect 73986 0 74042 800
rect 74170 0 74226 800
rect 74354 0 74410 800
rect 74538 0 74594 800
rect 74722 0 74778 800
rect 74998 0 75054 800
rect 75182 0 75238 800
rect 75366 0 75422 800
rect 75550 0 75606 800
rect 75734 0 75790 800
rect 76010 0 76066 800
rect 76194 0 76250 800
rect 76378 0 76434 800
rect 76562 0 76618 800
rect 76746 0 76802 800
rect 77022 0 77078 800
rect 77206 0 77262 800
rect 77390 0 77446 800
rect 77574 0 77630 800
rect 77758 0 77814 800
rect 78034 0 78090 800
rect 78218 0 78274 800
rect 78402 0 78458 800
rect 78586 0 78642 800
rect 78770 0 78826 800
rect 79046 0 79102 800
rect 79230 0 79286 800
rect 79414 0 79470 800
rect 79598 0 79654 800
rect 79782 0 79838 800
rect 80058 0 80114 800
rect 80242 0 80298 800
rect 80426 0 80482 800
rect 80610 0 80666 800
rect 80794 0 80850 800
rect 81070 0 81126 800
rect 81254 0 81310 800
rect 81438 0 81494 800
rect 81622 0 81678 800
rect 81806 0 81862 800
rect 82082 0 82138 800
rect 82266 0 82322 800
rect 82450 0 82506 800
rect 82634 0 82690 800
rect 82818 0 82874 800
rect 83094 0 83150 800
rect 83278 0 83334 800
rect 83462 0 83518 800
rect 83646 0 83702 800
rect 83830 0 83886 800
rect 84106 0 84162 800
rect 84290 0 84346 800
rect 84474 0 84530 800
rect 84658 0 84714 800
rect 84842 0 84898 800
rect 85118 0 85174 800
rect 85302 0 85358 800
rect 85486 0 85542 800
rect 85670 0 85726 800
rect 85854 0 85910 800
rect 86130 0 86186 800
rect 86314 0 86370 800
rect 86498 0 86554 800
rect 86682 0 86738 800
rect 86866 0 86922 800
rect 87142 0 87198 800
rect 87326 0 87382 800
rect 87510 0 87566 800
rect 87694 0 87750 800
rect 87878 0 87934 800
rect 88154 0 88210 800
rect 88338 0 88394 800
rect 88522 0 88578 800
rect 88706 0 88762 800
rect 88890 0 88946 800
rect 89166 0 89222 800
rect 89350 0 89406 800
rect 89534 0 89590 800
rect 89718 0 89774 800
rect 89902 0 89958 800
rect 90178 0 90234 800
rect 90362 0 90418 800
rect 90546 0 90602 800
rect 90730 0 90786 800
rect 90914 0 90970 800
rect 91190 0 91246 800
rect 91374 0 91430 800
rect 91558 0 91614 800
rect 91742 0 91798 800
rect 91926 0 91982 800
rect 92202 0 92258 800
rect 92386 0 92442 800
rect 92570 0 92626 800
rect 92754 0 92810 800
rect 92938 0 92994 800
rect 93214 0 93270 800
rect 93398 0 93454 800
rect 93582 0 93638 800
rect 93766 0 93822 800
rect 93950 0 94006 800
rect 94226 0 94282 800
rect 94410 0 94466 800
rect 94594 0 94650 800
rect 94778 0 94834 800
rect 94962 0 95018 800
rect 95238 0 95294 800
rect 95422 0 95478 800
rect 95606 0 95662 800
rect 95790 0 95846 800
rect 95974 0 96030 800
rect 96250 0 96306 800
rect 96434 0 96490 800
rect 96618 0 96674 800
rect 96802 0 96858 800
rect 96986 0 97042 800
rect 97262 0 97318 800
rect 97446 0 97502 800
rect 97630 0 97686 800
rect 97814 0 97870 800
rect 97998 0 98054 800
rect 98274 0 98330 800
rect 98458 0 98514 800
rect 98642 0 98698 800
rect 98826 0 98882 800
rect 99010 0 99066 800
rect 99286 0 99342 800
rect 99470 0 99526 800
rect 99654 0 99710 800
rect 99838 0 99894 800
<< obsm2 >>
rect 20 199144 330 199200
rect 498 199144 1158 199200
rect 1326 199144 2078 199200
rect 2246 199144 2906 199200
rect 3074 199144 3826 199200
rect 3994 199144 4654 199200
rect 4822 199144 5574 199200
rect 5742 199144 6402 199200
rect 6570 199144 7322 199200
rect 7490 199144 8150 199200
rect 8318 199144 9070 199200
rect 9238 199144 9898 199200
rect 10066 199144 10818 199200
rect 10986 199144 11646 199200
rect 11814 199144 12566 199200
rect 12734 199144 13486 199200
rect 13654 199144 14314 199200
rect 14482 199144 15234 199200
rect 15402 199144 16062 199200
rect 16230 199144 16982 199200
rect 17150 199144 17810 199200
rect 17978 199144 18730 199200
rect 18898 199144 19558 199200
rect 19726 199144 20478 199200
rect 20646 199144 21306 199200
rect 21474 199144 22226 199200
rect 22394 199144 23054 199200
rect 23222 199144 23974 199200
rect 24142 199144 24802 199200
rect 24970 199144 25722 199200
rect 25890 199144 26642 199200
rect 26810 199144 27470 199200
rect 27638 199144 28390 199200
rect 28558 199144 29218 199200
rect 29386 199144 30138 199200
rect 30306 199144 30966 199200
rect 31134 199144 31886 199200
rect 32054 199144 32714 199200
rect 32882 199144 33634 199200
rect 33802 199144 34462 199200
rect 34630 199144 35382 199200
rect 35550 199144 36210 199200
rect 36378 199144 37130 199200
rect 37298 199144 38050 199200
rect 38218 199144 38878 199200
rect 39046 199144 39798 199200
rect 39966 199144 40626 199200
rect 40794 199144 41546 199200
rect 41714 199144 42374 199200
rect 42542 199144 43294 199200
rect 43462 199144 44122 199200
rect 44290 199144 45042 199200
rect 45210 199144 45870 199200
rect 46038 199144 46790 199200
rect 46958 199144 47618 199200
rect 47786 199144 48538 199200
rect 48706 199144 49366 199200
rect 49534 199144 50286 199200
rect 50454 199144 51206 199200
rect 51374 199144 52034 199200
rect 52202 199144 52954 199200
rect 53122 199144 53782 199200
rect 53950 199144 54702 199200
rect 54870 199144 55530 199200
rect 55698 199144 56450 199200
rect 56618 199144 57278 199200
rect 57446 199144 58198 199200
rect 58366 199144 59026 199200
rect 59194 199144 59946 199200
rect 60114 199144 60774 199200
rect 60942 199144 61694 199200
rect 61862 199144 62522 199200
rect 62690 199144 63442 199200
rect 63610 199144 64362 199200
rect 64530 199144 65190 199200
rect 65358 199144 66110 199200
rect 66278 199144 66938 199200
rect 67106 199144 67858 199200
rect 68026 199144 68686 199200
rect 68854 199144 69606 199200
rect 69774 199144 70434 199200
rect 70602 199144 71354 199200
rect 71522 199144 72182 199200
rect 72350 199144 73102 199200
rect 73270 199144 73930 199200
rect 74098 199144 74850 199200
rect 75018 199144 75770 199200
rect 75938 199144 76598 199200
rect 76766 199144 77518 199200
rect 77686 199144 78346 199200
rect 78514 199144 79266 199200
rect 79434 199144 80094 199200
rect 80262 199144 81014 199200
rect 81182 199144 81842 199200
rect 82010 199144 82762 199200
rect 82930 199144 83590 199200
rect 83758 199144 84510 199200
rect 84678 199144 85338 199200
rect 85506 199144 86258 199200
rect 86426 199144 87086 199200
rect 87254 199144 88006 199200
rect 88174 199144 88926 199200
rect 89094 199144 89754 199200
rect 89922 199144 90674 199200
rect 90842 199144 91502 199200
rect 91670 199144 92422 199200
rect 92590 199144 93250 199200
rect 93418 199144 94170 199200
rect 94338 199144 94998 199200
rect 95166 199144 95918 199200
rect 96086 199144 96746 199200
rect 96914 199144 97666 199200
rect 97834 199144 98494 199200
rect 98662 199144 99414 199200
rect 99582 199144 99892 199200
rect 20 856 99892 199144
rect 20 800 54 856
rect 222 800 238 856
rect 406 800 422 856
rect 590 800 606 856
rect 774 800 790 856
rect 958 800 1066 856
rect 1234 800 1250 856
rect 1418 800 1434 856
rect 1602 800 1618 856
rect 1786 800 1802 856
rect 1970 800 2078 856
rect 2246 800 2262 856
rect 2430 800 2446 856
rect 2614 800 2630 856
rect 2798 800 2814 856
rect 2982 800 3090 856
rect 3258 800 3274 856
rect 3442 800 3458 856
rect 3626 800 3642 856
rect 3810 800 3826 856
rect 3994 800 4102 856
rect 4270 800 4286 856
rect 4454 800 4470 856
rect 4638 800 4654 856
rect 4822 800 4838 856
rect 5006 800 5114 856
rect 5282 800 5298 856
rect 5466 800 5482 856
rect 5650 800 5666 856
rect 5834 800 5850 856
rect 6018 800 6126 856
rect 6294 800 6310 856
rect 6478 800 6494 856
rect 6662 800 6678 856
rect 6846 800 6862 856
rect 7030 800 7138 856
rect 7306 800 7322 856
rect 7490 800 7506 856
rect 7674 800 7690 856
rect 7858 800 7874 856
rect 8042 800 8150 856
rect 8318 800 8334 856
rect 8502 800 8518 856
rect 8686 800 8702 856
rect 8870 800 8886 856
rect 9054 800 9162 856
rect 9330 800 9346 856
rect 9514 800 9530 856
rect 9698 800 9714 856
rect 9882 800 9898 856
rect 10066 800 10174 856
rect 10342 800 10358 856
rect 10526 800 10542 856
rect 10710 800 10726 856
rect 10894 800 10910 856
rect 11078 800 11186 856
rect 11354 800 11370 856
rect 11538 800 11554 856
rect 11722 800 11738 856
rect 11906 800 11922 856
rect 12090 800 12198 856
rect 12366 800 12382 856
rect 12550 800 12566 856
rect 12734 800 12750 856
rect 12918 800 12934 856
rect 13102 800 13210 856
rect 13378 800 13394 856
rect 13562 800 13578 856
rect 13746 800 13762 856
rect 13930 800 13946 856
rect 14114 800 14222 856
rect 14390 800 14406 856
rect 14574 800 14590 856
rect 14758 800 14774 856
rect 14942 800 14958 856
rect 15126 800 15234 856
rect 15402 800 15418 856
rect 15586 800 15602 856
rect 15770 800 15786 856
rect 15954 800 15970 856
rect 16138 800 16246 856
rect 16414 800 16430 856
rect 16598 800 16614 856
rect 16782 800 16798 856
rect 16966 800 16982 856
rect 17150 800 17258 856
rect 17426 800 17442 856
rect 17610 800 17626 856
rect 17794 800 17810 856
rect 17978 800 17994 856
rect 18162 800 18270 856
rect 18438 800 18454 856
rect 18622 800 18638 856
rect 18806 800 18822 856
rect 18990 800 19006 856
rect 19174 800 19282 856
rect 19450 800 19466 856
rect 19634 800 19650 856
rect 19818 800 19834 856
rect 20002 800 20018 856
rect 20186 800 20294 856
rect 20462 800 20478 856
rect 20646 800 20662 856
rect 20830 800 20846 856
rect 21014 800 21030 856
rect 21198 800 21306 856
rect 21474 800 21490 856
rect 21658 800 21674 856
rect 21842 800 21858 856
rect 22026 800 22042 856
rect 22210 800 22318 856
rect 22486 800 22502 856
rect 22670 800 22686 856
rect 22854 800 22870 856
rect 23038 800 23054 856
rect 23222 800 23330 856
rect 23498 800 23514 856
rect 23682 800 23698 856
rect 23866 800 23882 856
rect 24050 800 24066 856
rect 24234 800 24342 856
rect 24510 800 24526 856
rect 24694 800 24710 856
rect 24878 800 24894 856
rect 25062 800 25078 856
rect 25246 800 25354 856
rect 25522 800 25538 856
rect 25706 800 25722 856
rect 25890 800 25906 856
rect 26074 800 26090 856
rect 26258 800 26366 856
rect 26534 800 26550 856
rect 26718 800 26734 856
rect 26902 800 26918 856
rect 27086 800 27102 856
rect 27270 800 27378 856
rect 27546 800 27562 856
rect 27730 800 27746 856
rect 27914 800 27930 856
rect 28098 800 28114 856
rect 28282 800 28390 856
rect 28558 800 28574 856
rect 28742 800 28758 856
rect 28926 800 28942 856
rect 29110 800 29126 856
rect 29294 800 29402 856
rect 29570 800 29586 856
rect 29754 800 29770 856
rect 29938 800 29954 856
rect 30122 800 30138 856
rect 30306 800 30414 856
rect 30582 800 30598 856
rect 30766 800 30782 856
rect 30950 800 30966 856
rect 31134 800 31150 856
rect 31318 800 31426 856
rect 31594 800 31610 856
rect 31778 800 31794 856
rect 31962 800 31978 856
rect 32146 800 32162 856
rect 32330 800 32438 856
rect 32606 800 32622 856
rect 32790 800 32806 856
rect 32974 800 32990 856
rect 33158 800 33174 856
rect 33342 800 33450 856
rect 33618 800 33634 856
rect 33802 800 33818 856
rect 33986 800 34002 856
rect 34170 800 34186 856
rect 34354 800 34462 856
rect 34630 800 34646 856
rect 34814 800 34830 856
rect 34998 800 35014 856
rect 35182 800 35198 856
rect 35366 800 35474 856
rect 35642 800 35658 856
rect 35826 800 35842 856
rect 36010 800 36026 856
rect 36194 800 36210 856
rect 36378 800 36486 856
rect 36654 800 36670 856
rect 36838 800 36854 856
rect 37022 800 37038 856
rect 37206 800 37222 856
rect 37390 800 37498 856
rect 37666 800 37682 856
rect 37850 800 37866 856
rect 38034 800 38050 856
rect 38218 800 38234 856
rect 38402 800 38510 856
rect 38678 800 38694 856
rect 38862 800 38878 856
rect 39046 800 39062 856
rect 39230 800 39246 856
rect 39414 800 39522 856
rect 39690 800 39706 856
rect 39874 800 39890 856
rect 40058 800 40074 856
rect 40242 800 40258 856
rect 40426 800 40534 856
rect 40702 800 40718 856
rect 40886 800 40902 856
rect 41070 800 41086 856
rect 41254 800 41270 856
rect 41438 800 41546 856
rect 41714 800 41730 856
rect 41898 800 41914 856
rect 42082 800 42098 856
rect 42266 800 42282 856
rect 42450 800 42558 856
rect 42726 800 42742 856
rect 42910 800 42926 856
rect 43094 800 43110 856
rect 43278 800 43294 856
rect 43462 800 43570 856
rect 43738 800 43754 856
rect 43922 800 43938 856
rect 44106 800 44122 856
rect 44290 800 44306 856
rect 44474 800 44582 856
rect 44750 800 44766 856
rect 44934 800 44950 856
rect 45118 800 45134 856
rect 45302 800 45318 856
rect 45486 800 45594 856
rect 45762 800 45778 856
rect 45946 800 45962 856
rect 46130 800 46146 856
rect 46314 800 46330 856
rect 46498 800 46606 856
rect 46774 800 46790 856
rect 46958 800 46974 856
rect 47142 800 47158 856
rect 47326 800 47342 856
rect 47510 800 47618 856
rect 47786 800 47802 856
rect 47970 800 47986 856
rect 48154 800 48170 856
rect 48338 800 48354 856
rect 48522 800 48630 856
rect 48798 800 48814 856
rect 48982 800 48998 856
rect 49166 800 49182 856
rect 49350 800 49366 856
rect 49534 800 49642 856
rect 49810 800 49826 856
rect 49994 800 50010 856
rect 50178 800 50194 856
rect 50362 800 50378 856
rect 50546 800 50654 856
rect 50822 800 50838 856
rect 51006 800 51022 856
rect 51190 800 51206 856
rect 51374 800 51390 856
rect 51558 800 51666 856
rect 51834 800 51850 856
rect 52018 800 52034 856
rect 52202 800 52218 856
rect 52386 800 52402 856
rect 52570 800 52678 856
rect 52846 800 52862 856
rect 53030 800 53046 856
rect 53214 800 53230 856
rect 53398 800 53414 856
rect 53582 800 53690 856
rect 53858 800 53874 856
rect 54042 800 54058 856
rect 54226 800 54242 856
rect 54410 800 54426 856
rect 54594 800 54702 856
rect 54870 800 54886 856
rect 55054 800 55070 856
rect 55238 800 55254 856
rect 55422 800 55438 856
rect 55606 800 55714 856
rect 55882 800 55898 856
rect 56066 800 56082 856
rect 56250 800 56266 856
rect 56434 800 56450 856
rect 56618 800 56726 856
rect 56894 800 56910 856
rect 57078 800 57094 856
rect 57262 800 57278 856
rect 57446 800 57462 856
rect 57630 800 57738 856
rect 57906 800 57922 856
rect 58090 800 58106 856
rect 58274 800 58290 856
rect 58458 800 58474 856
rect 58642 800 58750 856
rect 58918 800 58934 856
rect 59102 800 59118 856
rect 59286 800 59302 856
rect 59470 800 59486 856
rect 59654 800 59762 856
rect 59930 800 59946 856
rect 60114 800 60130 856
rect 60298 800 60314 856
rect 60482 800 60498 856
rect 60666 800 60774 856
rect 60942 800 60958 856
rect 61126 800 61142 856
rect 61310 800 61326 856
rect 61494 800 61510 856
rect 61678 800 61786 856
rect 61954 800 61970 856
rect 62138 800 62154 856
rect 62322 800 62338 856
rect 62506 800 62522 856
rect 62690 800 62798 856
rect 62966 800 62982 856
rect 63150 800 63166 856
rect 63334 800 63350 856
rect 63518 800 63534 856
rect 63702 800 63810 856
rect 63978 800 63994 856
rect 64162 800 64178 856
rect 64346 800 64362 856
rect 64530 800 64546 856
rect 64714 800 64822 856
rect 64990 800 65006 856
rect 65174 800 65190 856
rect 65358 800 65374 856
rect 65542 800 65558 856
rect 65726 800 65834 856
rect 66002 800 66018 856
rect 66186 800 66202 856
rect 66370 800 66386 856
rect 66554 800 66570 856
rect 66738 800 66846 856
rect 67014 800 67030 856
rect 67198 800 67214 856
rect 67382 800 67398 856
rect 67566 800 67582 856
rect 67750 800 67858 856
rect 68026 800 68042 856
rect 68210 800 68226 856
rect 68394 800 68410 856
rect 68578 800 68594 856
rect 68762 800 68870 856
rect 69038 800 69054 856
rect 69222 800 69238 856
rect 69406 800 69422 856
rect 69590 800 69606 856
rect 69774 800 69882 856
rect 70050 800 70066 856
rect 70234 800 70250 856
rect 70418 800 70434 856
rect 70602 800 70618 856
rect 70786 800 70894 856
rect 71062 800 71078 856
rect 71246 800 71262 856
rect 71430 800 71446 856
rect 71614 800 71630 856
rect 71798 800 71906 856
rect 72074 800 72090 856
rect 72258 800 72274 856
rect 72442 800 72458 856
rect 72626 800 72642 856
rect 72810 800 72918 856
rect 73086 800 73102 856
rect 73270 800 73286 856
rect 73454 800 73470 856
rect 73638 800 73654 856
rect 73822 800 73930 856
rect 74098 800 74114 856
rect 74282 800 74298 856
rect 74466 800 74482 856
rect 74650 800 74666 856
rect 74834 800 74942 856
rect 75110 800 75126 856
rect 75294 800 75310 856
rect 75478 800 75494 856
rect 75662 800 75678 856
rect 75846 800 75954 856
rect 76122 800 76138 856
rect 76306 800 76322 856
rect 76490 800 76506 856
rect 76674 800 76690 856
rect 76858 800 76966 856
rect 77134 800 77150 856
rect 77318 800 77334 856
rect 77502 800 77518 856
rect 77686 800 77702 856
rect 77870 800 77978 856
rect 78146 800 78162 856
rect 78330 800 78346 856
rect 78514 800 78530 856
rect 78698 800 78714 856
rect 78882 800 78990 856
rect 79158 800 79174 856
rect 79342 800 79358 856
rect 79526 800 79542 856
rect 79710 800 79726 856
rect 79894 800 80002 856
rect 80170 800 80186 856
rect 80354 800 80370 856
rect 80538 800 80554 856
rect 80722 800 80738 856
rect 80906 800 81014 856
rect 81182 800 81198 856
rect 81366 800 81382 856
rect 81550 800 81566 856
rect 81734 800 81750 856
rect 81918 800 82026 856
rect 82194 800 82210 856
rect 82378 800 82394 856
rect 82562 800 82578 856
rect 82746 800 82762 856
rect 82930 800 83038 856
rect 83206 800 83222 856
rect 83390 800 83406 856
rect 83574 800 83590 856
rect 83758 800 83774 856
rect 83942 800 84050 856
rect 84218 800 84234 856
rect 84402 800 84418 856
rect 84586 800 84602 856
rect 84770 800 84786 856
rect 84954 800 85062 856
rect 85230 800 85246 856
rect 85414 800 85430 856
rect 85598 800 85614 856
rect 85782 800 85798 856
rect 85966 800 86074 856
rect 86242 800 86258 856
rect 86426 800 86442 856
rect 86610 800 86626 856
rect 86794 800 86810 856
rect 86978 800 87086 856
rect 87254 800 87270 856
rect 87438 800 87454 856
rect 87622 800 87638 856
rect 87806 800 87822 856
rect 87990 800 88098 856
rect 88266 800 88282 856
rect 88450 800 88466 856
rect 88634 800 88650 856
rect 88818 800 88834 856
rect 89002 800 89110 856
rect 89278 800 89294 856
rect 89462 800 89478 856
rect 89646 800 89662 856
rect 89830 800 89846 856
rect 90014 800 90122 856
rect 90290 800 90306 856
rect 90474 800 90490 856
rect 90658 800 90674 856
rect 90842 800 90858 856
rect 91026 800 91134 856
rect 91302 800 91318 856
rect 91486 800 91502 856
rect 91670 800 91686 856
rect 91854 800 91870 856
rect 92038 800 92146 856
rect 92314 800 92330 856
rect 92498 800 92514 856
rect 92682 800 92698 856
rect 92866 800 92882 856
rect 93050 800 93158 856
rect 93326 800 93342 856
rect 93510 800 93526 856
rect 93694 800 93710 856
rect 93878 800 93894 856
rect 94062 800 94170 856
rect 94338 800 94354 856
rect 94522 800 94538 856
rect 94706 800 94722 856
rect 94890 800 94906 856
rect 95074 800 95182 856
rect 95350 800 95366 856
rect 95534 800 95550 856
rect 95718 800 95734 856
rect 95902 800 95918 856
rect 96086 800 96194 856
rect 96362 800 96378 856
rect 96546 800 96562 856
rect 96730 800 96746 856
rect 96914 800 96930 856
rect 97098 800 97206 856
rect 97374 800 97390 856
rect 97558 800 97574 856
rect 97742 800 97758 856
rect 97926 800 97942 856
rect 98110 800 98218 856
rect 98386 800 98402 856
rect 98570 800 98586 856
rect 98754 800 98770 856
rect 98938 800 98954 856
rect 99122 800 99230 856
rect 99398 800 99414 856
rect 99582 800 99598 856
rect 99766 800 99782 856
<< metal3 >>
rect 0 198840 800 198960
rect 0 196664 800 196784
rect 0 194352 800 194472
rect 0 192176 800 192296
rect 0 190000 800 190120
rect 0 187688 800 187808
rect 0 185512 800 185632
rect 0 183336 800 183456
rect 0 181024 800 181144
rect 0 178848 800 178968
rect 0 176672 800 176792
rect 0 174360 800 174480
rect 0 172184 800 172304
rect 0 170008 800 170128
rect 0 167696 800 167816
rect 0 165520 800 165640
rect 0 163344 800 163464
rect 0 161032 800 161152
rect 0 158856 800 158976
rect 0 156680 800 156800
rect 0 154368 800 154488
rect 0 152192 800 152312
rect 0 150016 800 150136
rect 0 147704 800 147824
rect 0 145528 800 145648
rect 0 143352 800 143472
rect 0 141040 800 141160
rect 0 138864 800 138984
rect 0 136688 800 136808
rect 0 134376 800 134496
rect 0 132200 800 132320
rect 0 129888 800 130008
rect 0 127712 800 127832
rect 0 125536 800 125656
rect 0 123224 800 123344
rect 0 121048 800 121168
rect 0 118872 800 118992
rect 0 116560 800 116680
rect 0 114384 800 114504
rect 0 112208 800 112328
rect 0 109896 800 110016
rect 0 107720 800 107840
rect 0 105544 800 105664
rect 0 103232 800 103352
rect 0 101056 800 101176
rect 99200 99968 100000 100088
rect 0 98880 800 99000
rect 0 96568 800 96688
rect 0 94392 800 94512
rect 0 92216 800 92336
rect 0 89904 800 90024
rect 0 87728 800 87848
rect 0 85552 800 85672
rect 0 83240 800 83360
rect 0 81064 800 81184
rect 0 78888 800 79008
rect 0 76576 800 76696
rect 0 74400 800 74520
rect 0 72224 800 72344
rect 0 69912 800 70032
rect 0 67736 800 67856
rect 0 65424 800 65544
rect 0 63248 800 63368
rect 0 61072 800 61192
rect 0 58760 800 58880
rect 0 56584 800 56704
rect 0 54408 800 54528
rect 0 52096 800 52216
rect 0 49920 800 50040
rect 0 47744 800 47864
rect 0 45432 800 45552
rect 0 43256 800 43376
rect 0 41080 800 41200
rect 0 38768 800 38888
rect 0 36592 800 36712
rect 0 34416 800 34536
rect 0 32104 800 32224
rect 0 29928 800 30048
rect 0 27752 800 27872
rect 0 25440 800 25560
rect 0 23264 800 23384
rect 0 21088 800 21208
rect 0 18776 800 18896
rect 0 16600 800 16720
rect 0 14424 800 14544
rect 0 12112 800 12232
rect 0 9936 800 10056
rect 0 7760 800 7880
rect 0 5448 800 5568
rect 0 3272 800 3392
rect 0 1096 800 1216
<< obsm3 >>
rect 880 198760 99200 198933
rect 800 196864 99200 198760
rect 880 196584 99200 196864
rect 800 194552 99200 196584
rect 880 194272 99200 194552
rect 800 192376 99200 194272
rect 880 192096 99200 192376
rect 800 190200 99200 192096
rect 880 189920 99200 190200
rect 800 187888 99200 189920
rect 880 187608 99200 187888
rect 800 185712 99200 187608
rect 880 185432 99200 185712
rect 800 183536 99200 185432
rect 880 183256 99200 183536
rect 800 181224 99200 183256
rect 880 180944 99200 181224
rect 800 179048 99200 180944
rect 880 178768 99200 179048
rect 800 176872 99200 178768
rect 880 176592 99200 176872
rect 800 174560 99200 176592
rect 880 174280 99200 174560
rect 800 172384 99200 174280
rect 880 172104 99200 172384
rect 800 170208 99200 172104
rect 880 169928 99200 170208
rect 800 167896 99200 169928
rect 880 167616 99200 167896
rect 800 165720 99200 167616
rect 880 165440 99200 165720
rect 800 163544 99200 165440
rect 880 163264 99200 163544
rect 800 161232 99200 163264
rect 880 160952 99200 161232
rect 800 159056 99200 160952
rect 880 158776 99200 159056
rect 800 156880 99200 158776
rect 880 156600 99200 156880
rect 800 154568 99200 156600
rect 880 154288 99200 154568
rect 800 152392 99200 154288
rect 880 152112 99200 152392
rect 800 150216 99200 152112
rect 880 149936 99200 150216
rect 800 147904 99200 149936
rect 880 147624 99200 147904
rect 800 145728 99200 147624
rect 880 145448 99200 145728
rect 800 143552 99200 145448
rect 880 143272 99200 143552
rect 800 141240 99200 143272
rect 880 140960 99200 141240
rect 800 139064 99200 140960
rect 880 138784 99200 139064
rect 800 136888 99200 138784
rect 880 136608 99200 136888
rect 800 134576 99200 136608
rect 880 134296 99200 134576
rect 800 132400 99200 134296
rect 880 132120 99200 132400
rect 800 130088 99200 132120
rect 880 129808 99200 130088
rect 800 127912 99200 129808
rect 880 127632 99200 127912
rect 800 125736 99200 127632
rect 880 125456 99200 125736
rect 800 123424 99200 125456
rect 880 123144 99200 123424
rect 800 121248 99200 123144
rect 880 120968 99200 121248
rect 800 119072 99200 120968
rect 880 118792 99200 119072
rect 800 116760 99200 118792
rect 880 116480 99200 116760
rect 800 114584 99200 116480
rect 880 114304 99200 114584
rect 800 112408 99200 114304
rect 880 112128 99200 112408
rect 800 110096 99200 112128
rect 880 109816 99200 110096
rect 800 107920 99200 109816
rect 880 107640 99200 107920
rect 800 105744 99200 107640
rect 880 105464 99200 105744
rect 800 103432 99200 105464
rect 880 103152 99200 103432
rect 800 101256 99200 103152
rect 880 100976 99200 101256
rect 800 100168 99200 100976
rect 800 99888 99120 100168
rect 800 99080 99200 99888
rect 880 98800 99200 99080
rect 800 96768 99200 98800
rect 880 96488 99200 96768
rect 800 94592 99200 96488
rect 880 94312 99200 94592
rect 800 92416 99200 94312
rect 880 92136 99200 92416
rect 800 90104 99200 92136
rect 880 89824 99200 90104
rect 800 87928 99200 89824
rect 880 87648 99200 87928
rect 800 85752 99200 87648
rect 880 85472 99200 85752
rect 800 83440 99200 85472
rect 880 83160 99200 83440
rect 800 81264 99200 83160
rect 880 80984 99200 81264
rect 800 79088 99200 80984
rect 880 78808 99200 79088
rect 800 76776 99200 78808
rect 880 76496 99200 76776
rect 800 74600 99200 76496
rect 880 74320 99200 74600
rect 800 72424 99200 74320
rect 880 72144 99200 72424
rect 800 70112 99200 72144
rect 880 69832 99200 70112
rect 800 67936 99200 69832
rect 880 67656 99200 67936
rect 800 65624 99200 67656
rect 880 65344 99200 65624
rect 800 63448 99200 65344
rect 880 63168 99200 63448
rect 800 61272 99200 63168
rect 880 60992 99200 61272
rect 800 58960 99200 60992
rect 880 58680 99200 58960
rect 800 56784 99200 58680
rect 880 56504 99200 56784
rect 800 54608 99200 56504
rect 880 54328 99200 54608
rect 800 52296 99200 54328
rect 880 52016 99200 52296
rect 800 50120 99200 52016
rect 880 49840 99200 50120
rect 800 47944 99200 49840
rect 880 47664 99200 47944
rect 800 45632 99200 47664
rect 880 45352 99200 45632
rect 800 43456 99200 45352
rect 880 43176 99200 43456
rect 800 41280 99200 43176
rect 880 41000 99200 41280
rect 800 38968 99200 41000
rect 880 38688 99200 38968
rect 800 36792 99200 38688
rect 880 36512 99200 36792
rect 800 34616 99200 36512
rect 880 34336 99200 34616
rect 800 32304 99200 34336
rect 880 32024 99200 32304
rect 800 30128 99200 32024
rect 880 29848 99200 30128
rect 800 27952 99200 29848
rect 880 27672 99200 27952
rect 800 25640 99200 27672
rect 880 25360 99200 25640
rect 800 23464 99200 25360
rect 880 23184 99200 23464
rect 800 21288 99200 23184
rect 880 21008 99200 21288
rect 800 18976 99200 21008
rect 880 18696 99200 18976
rect 800 16800 99200 18696
rect 880 16520 99200 16800
rect 800 14624 99200 16520
rect 880 14344 99200 14624
rect 800 12312 99200 14344
rect 880 12032 99200 12312
rect 800 10136 99200 12032
rect 880 9856 99200 10136
rect 800 7960 99200 9856
rect 880 7680 99200 7960
rect 800 5648 99200 7680
rect 880 5368 99200 5648
rect 800 3472 99200 5368
rect 880 3192 99200 3472
rect 800 1296 99200 3192
rect 880 1123 99200 1296
<< metal4 >>
rect 4208 2128 4528 197520
rect 19568 2128 19888 197520
rect 34928 2128 35248 197520
rect 50288 2128 50608 197520
rect 65648 2128 65968 197520
rect 81008 2128 81328 197520
rect 96368 2128 96688 197520
<< obsm4 >>
rect 1715 2347 4128 186421
rect 4608 2347 19488 186421
rect 19968 2347 29013 186421
<< labels >>
rlabel metal2 s 386 199200 442 200000 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 26698 199200 26754 200000 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 29274 199200 29330 200000 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 31942 199200 31998 200000 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 34518 199200 34574 200000 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 37186 199200 37242 200000 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 39854 199200 39910 200000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 42430 199200 42486 200000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 45098 199200 45154 200000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 47674 199200 47730 200000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 50342 199200 50398 200000 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 2962 199200 3018 200000 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 53010 199200 53066 200000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 55586 199200 55642 200000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 58254 199200 58310 200000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 60830 199200 60886 200000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 63498 199200 63554 200000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 66166 199200 66222 200000 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 68742 199200 68798 200000 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 71410 199200 71466 200000 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 73986 199200 74042 200000 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 76654 199200 76710 200000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 5630 199200 5686 200000 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 79322 199200 79378 200000 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 81898 199200 81954 200000 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 84566 199200 84622 200000 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 87142 199200 87198 200000 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 89810 199200 89866 200000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 92478 199200 92534 200000 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 95054 199200 95110 200000 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 97722 199200 97778 200000 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 8206 199200 8262 200000 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 10874 199200 10930 200000 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 13542 199200 13598 200000 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 16118 199200 16174 200000 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 18786 199200 18842 200000 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 21362 199200 21418 200000 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 24030 199200 24086 200000 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 1214 199200 1270 200000 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 27526 199200 27582 200000 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 30194 199200 30250 200000 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 32770 199200 32826 200000 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 35438 199200 35494 200000 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 38106 199200 38162 200000 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 40682 199200 40738 200000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 43350 199200 43406 200000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 45926 199200 45982 200000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 48594 199200 48650 200000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 51262 199200 51318 200000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 3882 199200 3938 200000 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 53838 199200 53894 200000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 56506 199200 56562 200000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 59082 199200 59138 200000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 61750 199200 61806 200000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 64418 199200 64474 200000 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 66994 199200 67050 200000 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 69662 199200 69718 200000 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 72238 199200 72294 200000 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 74906 199200 74962 200000 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 77574 199200 77630 200000 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 6458 199200 6514 200000 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 80150 199200 80206 200000 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 82818 199200 82874 200000 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 85394 199200 85450 200000 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 88062 199200 88118 200000 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 90730 199200 90786 200000 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 93306 199200 93362 200000 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 95974 199200 96030 200000 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 98550 199200 98606 200000 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 9126 199200 9182 200000 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 11702 199200 11758 200000 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 14370 199200 14426 200000 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 17038 199200 17094 200000 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 19614 199200 19670 200000 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 22282 199200 22338 200000 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 24858 199200 24914 200000 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 2134 199200 2190 200000 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 28446 199200 28502 200000 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 31022 199200 31078 200000 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 33690 199200 33746 200000 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 36266 199200 36322 200000 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 38934 199200 38990 200000 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 41602 199200 41658 200000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 44178 199200 44234 200000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 46846 199200 46902 200000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 49422 199200 49478 200000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 52090 199200 52146 200000 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 4710 199200 4766 200000 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 54758 199200 54814 200000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 57334 199200 57390 200000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 60002 199200 60058 200000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 62578 199200 62634 200000 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 65246 199200 65302 200000 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 67914 199200 67970 200000 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 70490 199200 70546 200000 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 73158 199200 73214 200000 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 75826 199200 75882 200000 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 78402 199200 78458 200000 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 7378 199200 7434 200000 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 81070 199200 81126 200000 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 83646 199200 83702 200000 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 86314 199200 86370 200000 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 88982 199200 89038 200000 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 91558 199200 91614 200000 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 94226 199200 94282 200000 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 96802 199200 96858 200000 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 99470 199200 99526 200000 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 9954 199200 10010 200000 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 12622 199200 12678 200000 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 15290 199200 15346 200000 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 17866 199200 17922 200000 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 20534 199200 20590 200000 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 23110 199200 23166 200000 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 25778 199200 25834 200000 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 99286 0 99342 800 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 99470 0 99526 800 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 99654 0 99710 800 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 21546 0 21602 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 82266 0 82322 800 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 82818 0 82874 800 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 83462 0 83518 800 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 84106 0 84162 800 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 84658 0 84714 800 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 85302 0 85358 800 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 85854 0 85910 800 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 86498 0 86554 800 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 87142 0 87198 800 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 87694 0 87750 800 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 27618 0 27674 800 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 88338 0 88394 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 88890 0 88946 800 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 89534 0 89590 800 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 90178 0 90234 800 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 90730 0 90786 800 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 91374 0 91430 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 91926 0 91982 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 92570 0 92626 800 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 93214 0 93270 800 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 93766 0 93822 800 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 28170 0 28226 800 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 94410 0 94466 800 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 94962 0 95018 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 95606 0 95662 800 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 96250 0 96306 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 96802 0 96858 800 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 97446 0 97502 800 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 97998 0 98054 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 98642 0 98698 800 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 28814 0 28870 800 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 29458 0 29514 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 30010 0 30066 800 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 30654 0 30710 800 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 31206 0 31262 800 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 31850 0 31906 800 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 32494 0 32550 800 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 33046 0 33102 800 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 22098 0 22154 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 33690 0 33746 800 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 34242 0 34298 800 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 34886 0 34942 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 35530 0 35586 800 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 36082 0 36138 800 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 36726 0 36782 800 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 37278 0 37334 800 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 37922 0 37978 800 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 38566 0 38622 800 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 39118 0 39174 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 22742 0 22798 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 39762 0 39818 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 40314 0 40370 800 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 40958 0 41014 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 41602 0 41658 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 42154 0 42210 800 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 42798 0 42854 800 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 43350 0 43406 800 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 43994 0 44050 800 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 44638 0 44694 800 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 45190 0 45246 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 23386 0 23442 800 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 45834 0 45890 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 46386 0 46442 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 47030 0 47086 800 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 47674 0 47730 800 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 48226 0 48282 800 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 48870 0 48926 800 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 49422 0 49478 800 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 50066 0 50122 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 50710 0 50766 800 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 51262 0 51318 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 23938 0 23994 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 51906 0 51962 800 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 52458 0 52514 800 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 53102 0 53158 800 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 53746 0 53802 800 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 54298 0 54354 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 54942 0 54998 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 55494 0 55550 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 56138 0 56194 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 56782 0 56838 800 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 57334 0 57390 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 24582 0 24638 800 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 57978 0 58034 800 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 58530 0 58586 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 59174 0 59230 800 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 59818 0 59874 800 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 60370 0 60426 800 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 61014 0 61070 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 61566 0 61622 800 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 62210 0 62266 800 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 62854 0 62910 800 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 63406 0 63462 800 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 25134 0 25190 800 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 64050 0 64106 800 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 64602 0 64658 800 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 65246 0 65302 800 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 65890 0 65946 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 66442 0 66498 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 67086 0 67142 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 67638 0 67694 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 68282 0 68338 800 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 68926 0 68982 800 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 69478 0 69534 800 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 25778 0 25834 800 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 70122 0 70178 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 70674 0 70730 800 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 71318 0 71374 800 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 71962 0 72018 800 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 72514 0 72570 800 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 73158 0 73214 800 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 73710 0 73766 800 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 74354 0 74410 800 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 74998 0 75054 800 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 75550 0 75606 800 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 26422 0 26478 800 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 76194 0 76250 800 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 76746 0 76802 800 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 77390 0 77446 800 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 78034 0 78090 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 78586 0 78642 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 79230 0 79286 800 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 79782 0 79838 800 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 80426 0 80482 800 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 81070 0 81126 800 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 81622 0 81678 800 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 26974 0 27030 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 21730 0 21786 800 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 82450 0 82506 800 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 83094 0 83150 800 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 83646 0 83702 800 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 84290 0 84346 800 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 84842 0 84898 800 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 85486 0 85542 800 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 86130 0 86186 800 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 86682 0 86738 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 87326 0 87382 800 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 87878 0 87934 800 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 27802 0 27858 800 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 88522 0 88578 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 89166 0 89222 800 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 89718 0 89774 800 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 90362 0 90418 800 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 90914 0 90970 800 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 91558 0 91614 800 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 92202 0 92258 800 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 92754 0 92810 800 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 93398 0 93454 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 93950 0 94006 800 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 28446 0 28502 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 94594 0 94650 800 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 95238 0 95294 800 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 95790 0 95846 800 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 96434 0 96490 800 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 96986 0 97042 800 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 97630 0 97686 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 98274 0 98330 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 98826 0 98882 800 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 28998 0 29054 800 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 29642 0 29698 800 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 30194 0 30250 800 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 30838 0 30894 800 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 31482 0 31538 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 32034 0 32090 800 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 32678 0 32734 800 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 33230 0 33286 800 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 22374 0 22430 800 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 33874 0 33930 800 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 34518 0 34574 800 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 35070 0 35126 800 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 35714 0 35770 800 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 36266 0 36322 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 36910 0 36966 800 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 37554 0 37610 800 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 38106 0 38162 800 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 38750 0 38806 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 39302 0 39358 800 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 22926 0 22982 800 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 39946 0 40002 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 40590 0 40646 800 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 41142 0 41198 800 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 41786 0 41842 800 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 42338 0 42394 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 42982 0 43038 800 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 43626 0 43682 800 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 44178 0 44234 800 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 44822 0 44878 800 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 45374 0 45430 800 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 23570 0 23626 800 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 46018 0 46074 800 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 46662 0 46718 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 47214 0 47270 800 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 47858 0 47914 800 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 48410 0 48466 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 49054 0 49110 800 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 49698 0 49754 800 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 50250 0 50306 800 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 50894 0 50950 800 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 51446 0 51502 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 24122 0 24178 800 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 52090 0 52146 800 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 52734 0 52790 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 53286 0 53342 800 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 53930 0 53986 800 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 54482 0 54538 800 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 55126 0 55182 800 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 55770 0 55826 800 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 56322 0 56378 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 56966 0 57022 800 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 57518 0 57574 800 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 24766 0 24822 800 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 58162 0 58218 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 58806 0 58862 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 59358 0 59414 800 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 60002 0 60058 800 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 60554 0 60610 800 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 61198 0 61254 800 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 61842 0 61898 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 62394 0 62450 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 63038 0 63094 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 63590 0 63646 800 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 25410 0 25466 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 64234 0 64290 800 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 64878 0 64934 800 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 65430 0 65486 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 66074 0 66130 800 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 66626 0 66682 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 67270 0 67326 800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 67914 0 67970 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 68466 0 68522 800 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 69110 0 69166 800 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 69662 0 69718 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 25962 0 26018 800 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 70306 0 70362 800 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 70950 0 71006 800 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 71502 0 71558 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 72146 0 72202 800 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 72698 0 72754 800 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 73342 0 73398 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 73986 0 74042 800 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 74538 0 74594 800 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 75182 0 75238 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 75734 0 75790 800 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 26606 0 26662 800 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 76378 0 76434 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 77022 0 77078 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 77574 0 77630 800 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 78218 0 78274 800 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 78770 0 78826 800 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 79414 0 79470 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 80058 0 80114 800 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 80610 0 80666 800 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 81254 0 81310 800 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 81806 0 81862 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 27158 0 27214 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 21914 0 21970 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 82634 0 82690 800 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 83278 0 83334 800 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 83830 0 83886 800 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 84474 0 84530 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 85118 0 85174 800 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 85670 0 85726 800 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 86314 0 86370 800 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 86866 0 86922 800 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 87510 0 87566 800 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 88154 0 88210 800 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 27986 0 28042 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 88706 0 88762 800 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 89350 0 89406 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 89902 0 89958 800 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 90546 0 90602 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 91190 0 91246 800 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 91742 0 91798 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 92386 0 92442 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 92938 0 92994 800 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 93582 0 93638 800 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 94226 0 94282 800 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 28630 0 28686 800 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 94778 0 94834 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 95422 0 95478 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 95974 0 96030 800 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 96618 0 96674 800 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 97262 0 97318 800 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 97814 0 97870 800 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 98458 0 98514 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 99010 0 99066 800 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 29182 0 29238 800 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 29826 0 29882 800 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 30470 0 30526 800 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 31022 0 31078 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 31666 0 31722 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 32218 0 32274 800 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 32862 0 32918 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 33506 0 33562 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 22558 0 22614 800 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 34058 0 34114 800 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 34702 0 34758 800 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 35254 0 35310 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 35898 0 35954 800 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 36542 0 36598 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 37094 0 37150 800 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 37738 0 37794 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 38290 0 38346 800 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 38934 0 38990 800 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 39578 0 39634 800 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 23110 0 23166 800 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 40130 0 40186 800 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 40774 0 40830 800 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 41326 0 41382 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 41970 0 42026 800 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 42614 0 42670 800 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 43166 0 43222 800 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 43810 0 43866 800 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 44362 0 44418 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 45006 0 45062 800 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 45650 0 45706 800 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 23754 0 23810 800 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 46202 0 46258 800 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 46846 0 46902 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 47398 0 47454 800 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 48042 0 48098 800 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 48686 0 48742 800 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 49238 0 49294 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 49882 0 49938 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 50434 0 50490 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 51078 0 51134 800 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 51722 0 51778 800 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 24398 0 24454 800 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 52274 0 52330 800 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 52918 0 52974 800 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 53470 0 53526 800 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 54114 0 54170 800 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 54758 0 54814 800 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 55310 0 55366 800 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 55954 0 56010 800 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 56506 0 56562 800 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 57150 0 57206 800 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 57794 0 57850 800 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 24950 0 25006 800 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 58346 0 58402 800 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 58990 0 59046 800 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 59542 0 59598 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 60186 0 60242 800 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 60830 0 60886 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 61382 0 61438 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 62026 0 62082 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 62578 0 62634 800 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 63222 0 63278 800 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 63866 0 63922 800 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 25594 0 25650 800 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 64418 0 64474 800 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 65062 0 65118 800 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 65614 0 65670 800 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 66258 0 66314 800 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 66902 0 66958 800 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 67454 0 67510 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 68098 0 68154 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 68650 0 68706 800 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 69294 0 69350 800 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 69938 0 69994 800 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 26146 0 26202 800 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 70490 0 70546 800 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 71134 0 71190 800 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 71686 0 71742 800 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 72330 0 72386 800 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 72974 0 73030 800 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 73526 0 73582 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 74170 0 74226 800 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 74722 0 74778 800 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 75366 0 75422 800 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 76010 0 76066 800 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 26790 0 26846 800 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 76562 0 76618 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 77206 0 77262 800 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 77758 0 77814 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 78402 0 78458 800 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 79046 0 79102 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 79598 0 79654 800 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 80242 0 80298 800 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 80794 0 80850 800 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 81438 0 81494 800 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 82082 0 82138 800 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 27434 0 27490 800 6 la_oenb[9]
port 501 nsew signal input
rlabel metal2 s 99838 0 99894 800 6 ring0_clk
port 502 nsew signal input
rlabel metal3 s 0 183336 800 183456 6 ring0_clkmux[0]
port 503 nsew signal output
rlabel metal3 s 0 187688 800 187808 6 ring0_clkmux[1]
port 504 nsew signal output
rlabel metal3 s 0 192176 800 192296 6 ring0_clkmux[2]
port 505 nsew signal output
rlabel metal3 s 0 196664 800 196784 6 ring0_start
port 506 nsew signal output
rlabel metal3 s 0 1096 800 1216 6 ring0_trim_a[0]
port 507 nsew signal output
rlabel metal3 s 0 45432 800 45552 6 ring0_trim_a[10]
port 508 nsew signal output
rlabel metal3 s 0 49920 800 50040 6 ring0_trim_a[11]
port 509 nsew signal output
rlabel metal3 s 0 54408 800 54528 6 ring0_trim_a[12]
port 510 nsew signal output
rlabel metal3 s 0 58760 800 58880 6 ring0_trim_a[13]
port 511 nsew signal output
rlabel metal3 s 0 63248 800 63368 6 ring0_trim_a[14]
port 512 nsew signal output
rlabel metal3 s 0 67736 800 67856 6 ring0_trim_a[15]
port 513 nsew signal output
rlabel metal3 s 0 72224 800 72344 6 ring0_trim_a[16]
port 514 nsew signal output
rlabel metal3 s 0 76576 800 76696 6 ring0_trim_a[17]
port 515 nsew signal output
rlabel metal3 s 0 81064 800 81184 6 ring0_trim_a[18]
port 516 nsew signal output
rlabel metal3 s 0 85552 800 85672 6 ring0_trim_a[19]
port 517 nsew signal output
rlabel metal3 s 0 5448 800 5568 6 ring0_trim_a[1]
port 518 nsew signal output
rlabel metal3 s 0 89904 800 90024 6 ring0_trim_a[20]
port 519 nsew signal output
rlabel metal3 s 0 94392 800 94512 6 ring0_trim_a[21]
port 520 nsew signal output
rlabel metal3 s 0 98880 800 99000 6 ring0_trim_a[22]
port 521 nsew signal output
rlabel metal3 s 0 103232 800 103352 6 ring0_trim_a[23]
port 522 nsew signal output
rlabel metal3 s 0 107720 800 107840 6 ring0_trim_a[24]
port 523 nsew signal output
rlabel metal3 s 0 112208 800 112328 6 ring0_trim_a[25]
port 524 nsew signal output
rlabel metal3 s 0 116560 800 116680 6 ring0_trim_a[26]
port 525 nsew signal output
rlabel metal3 s 0 118872 800 118992 6 ring0_trim_a[27]
port 526 nsew signal output
rlabel metal3 s 0 9936 800 10056 6 ring0_trim_a[2]
port 527 nsew signal output
rlabel metal3 s 0 14424 800 14544 6 ring0_trim_a[3]
port 528 nsew signal output
rlabel metal3 s 0 18776 800 18896 6 ring0_trim_a[4]
port 529 nsew signal output
rlabel metal3 s 0 23264 800 23384 6 ring0_trim_a[5]
port 530 nsew signal output
rlabel metal3 s 0 27752 800 27872 6 ring0_trim_a[6]
port 531 nsew signal output
rlabel metal3 s 0 32104 800 32224 6 ring0_trim_a[7]
port 532 nsew signal output
rlabel metal3 s 0 36592 800 36712 6 ring0_trim_a[8]
port 533 nsew signal output
rlabel metal3 s 0 41080 800 41200 6 ring0_trim_a[9]
port 534 nsew signal output
rlabel metal3 s 0 121048 800 121168 6 ring0_trim_b[0]
port 535 nsew signal output
rlabel metal3 s 0 143352 800 143472 6 ring0_trim_b[10]
port 536 nsew signal output
rlabel metal3 s 0 145528 800 145648 6 ring0_trim_b[11]
port 537 nsew signal output
rlabel metal3 s 0 147704 800 147824 6 ring0_trim_b[12]
port 538 nsew signal output
rlabel metal3 s 0 150016 800 150136 6 ring0_trim_b[13]
port 539 nsew signal output
rlabel metal3 s 0 152192 800 152312 6 ring0_trim_b[14]
port 540 nsew signal output
rlabel metal3 s 0 154368 800 154488 6 ring0_trim_b[15]
port 541 nsew signal output
rlabel metal3 s 0 156680 800 156800 6 ring0_trim_b[16]
port 542 nsew signal output
rlabel metal3 s 0 158856 800 158976 6 ring0_trim_b[17]
port 543 nsew signal output
rlabel metal3 s 0 161032 800 161152 6 ring0_trim_b[18]
port 544 nsew signal output
rlabel metal3 s 0 163344 800 163464 6 ring0_trim_b[19]
port 545 nsew signal output
rlabel metal3 s 0 123224 800 123344 6 ring0_trim_b[1]
port 546 nsew signal output
rlabel metal3 s 0 165520 800 165640 6 ring0_trim_b[20]
port 547 nsew signal output
rlabel metal3 s 0 167696 800 167816 6 ring0_trim_b[21]
port 548 nsew signal output
rlabel metal3 s 0 170008 800 170128 6 ring0_trim_b[22]
port 549 nsew signal output
rlabel metal3 s 0 172184 800 172304 6 ring0_trim_b[23]
port 550 nsew signal output
rlabel metal3 s 0 174360 800 174480 6 ring0_trim_b[24]
port 551 nsew signal output
rlabel metal3 s 0 176672 800 176792 6 ring0_trim_b[25]
port 552 nsew signal output
rlabel metal3 s 0 178848 800 178968 6 ring0_trim_b[26]
port 553 nsew signal output
rlabel metal3 s 0 181024 800 181144 6 ring0_trim_b[27]
port 554 nsew signal output
rlabel metal3 s 0 125536 800 125656 6 ring0_trim_b[2]
port 555 nsew signal output
rlabel metal3 s 0 127712 800 127832 6 ring0_trim_b[3]
port 556 nsew signal output
rlabel metal3 s 0 129888 800 130008 6 ring0_trim_b[4]
port 557 nsew signal output
rlabel metal3 s 0 132200 800 132320 6 ring0_trim_b[5]
port 558 nsew signal output
rlabel metal3 s 0 134376 800 134496 6 ring0_trim_b[6]
port 559 nsew signal output
rlabel metal3 s 0 136688 800 136808 6 ring0_trim_b[7]
port 560 nsew signal output
rlabel metal3 s 0 138864 800 138984 6 ring0_trim_b[8]
port 561 nsew signal output
rlabel metal3 s 0 141040 800 141160 6 ring0_trim_b[9]
port 562 nsew signal output
rlabel metal3 s 99200 99968 100000 100088 6 ring1_clk
port 563 nsew signal input
rlabel metal3 s 0 185512 800 185632 6 ring1_clkmux[0]
port 564 nsew signal output
rlabel metal3 s 0 190000 800 190120 6 ring1_clkmux[1]
port 565 nsew signal output
rlabel metal3 s 0 194352 800 194472 6 ring1_clkmux[2]
port 566 nsew signal output
rlabel metal3 s 0 198840 800 198960 6 ring1_start
port 567 nsew signal output
rlabel metal3 s 0 3272 800 3392 6 ring1_trim_a[0]
port 568 nsew signal output
rlabel metal3 s 0 47744 800 47864 6 ring1_trim_a[10]
port 569 nsew signal output
rlabel metal3 s 0 52096 800 52216 6 ring1_trim_a[11]
port 570 nsew signal output
rlabel metal3 s 0 56584 800 56704 6 ring1_trim_a[12]
port 571 nsew signal output
rlabel metal3 s 0 61072 800 61192 6 ring1_trim_a[13]
port 572 nsew signal output
rlabel metal3 s 0 65424 800 65544 6 ring1_trim_a[14]
port 573 nsew signal output
rlabel metal3 s 0 69912 800 70032 6 ring1_trim_a[15]
port 574 nsew signal output
rlabel metal3 s 0 74400 800 74520 6 ring1_trim_a[16]
port 575 nsew signal output
rlabel metal3 s 0 78888 800 79008 6 ring1_trim_a[17]
port 576 nsew signal output
rlabel metal3 s 0 83240 800 83360 6 ring1_trim_a[18]
port 577 nsew signal output
rlabel metal3 s 0 87728 800 87848 6 ring1_trim_a[19]
port 578 nsew signal output
rlabel metal3 s 0 7760 800 7880 6 ring1_trim_a[1]
port 579 nsew signal output
rlabel metal3 s 0 92216 800 92336 6 ring1_trim_a[20]
port 580 nsew signal output
rlabel metal3 s 0 96568 800 96688 6 ring1_trim_a[21]
port 581 nsew signal output
rlabel metal3 s 0 101056 800 101176 6 ring1_trim_a[22]
port 582 nsew signal output
rlabel metal3 s 0 105544 800 105664 6 ring1_trim_a[23]
port 583 nsew signal output
rlabel metal3 s 0 109896 800 110016 6 ring1_trim_a[24]
port 584 nsew signal output
rlabel metal3 s 0 114384 800 114504 6 ring1_trim_a[25]
port 585 nsew signal output
rlabel metal3 s 0 12112 800 12232 6 ring1_trim_a[2]
port 586 nsew signal output
rlabel metal3 s 0 16600 800 16720 6 ring1_trim_a[3]
port 587 nsew signal output
rlabel metal3 s 0 21088 800 21208 6 ring1_trim_a[4]
port 588 nsew signal output
rlabel metal3 s 0 25440 800 25560 6 ring1_trim_a[5]
port 589 nsew signal output
rlabel metal3 s 0 29928 800 30048 6 ring1_trim_a[6]
port 590 nsew signal output
rlabel metal3 s 0 34416 800 34536 6 ring1_trim_a[7]
port 591 nsew signal output
rlabel metal3 s 0 38768 800 38888 6 ring1_trim_a[8]
port 592 nsew signal output
rlabel metal3 s 0 43256 800 43376 6 ring1_trim_a[9]
port 593 nsew signal output
rlabel metal4 s 4208 2128 4528 197520 6 vccd1
port 594 nsew power input
rlabel metal4 s 34928 2128 35248 197520 6 vccd1
port 594 nsew power input
rlabel metal4 s 65648 2128 65968 197520 6 vccd1
port 594 nsew power input
rlabel metal4 s 96368 2128 96688 197520 6 vccd1
port 594 nsew power input
rlabel metal4 s 19568 2128 19888 197520 6 vssd1
port 595 nsew ground input
rlabel metal4 s 50288 2128 50608 197520 6 vssd1
port 595 nsew ground input
rlabel metal4 s 81008 2128 81328 197520 6 vssd1
port 595 nsew ground input
rlabel metal2 s 110 0 166 800 6 wb_clk_i
port 596 nsew signal input
rlabel metal2 s 294 0 350 800 6 wb_rst_i
port 597 nsew signal input
rlabel metal2 s 478 0 534 800 6 wbs_ack_o
port 598 nsew signal output
rlabel metal2 s 1306 0 1362 800 6 wbs_adr_i[0]
port 599 nsew signal input
rlabel metal2 s 8206 0 8262 800 6 wbs_adr_i[10]
port 600 nsew signal input
rlabel metal2 s 8758 0 8814 800 6 wbs_adr_i[11]
port 601 nsew signal input
rlabel metal2 s 9402 0 9458 800 6 wbs_adr_i[12]
port 602 nsew signal input
rlabel metal2 s 9954 0 10010 800 6 wbs_adr_i[13]
port 603 nsew signal input
rlabel metal2 s 10598 0 10654 800 6 wbs_adr_i[14]
port 604 nsew signal input
rlabel metal2 s 11242 0 11298 800 6 wbs_adr_i[15]
port 605 nsew signal input
rlabel metal2 s 11794 0 11850 800 6 wbs_adr_i[16]
port 606 nsew signal input
rlabel metal2 s 12438 0 12494 800 6 wbs_adr_i[17]
port 607 nsew signal input
rlabel metal2 s 12990 0 13046 800 6 wbs_adr_i[18]
port 608 nsew signal input
rlabel metal2 s 13634 0 13690 800 6 wbs_adr_i[19]
port 609 nsew signal input
rlabel metal2 s 2134 0 2190 800 6 wbs_adr_i[1]
port 610 nsew signal input
rlabel metal2 s 14278 0 14334 800 6 wbs_adr_i[20]
port 611 nsew signal input
rlabel metal2 s 14830 0 14886 800 6 wbs_adr_i[21]
port 612 nsew signal input
rlabel metal2 s 15474 0 15530 800 6 wbs_adr_i[22]
port 613 nsew signal input
rlabel metal2 s 16026 0 16082 800 6 wbs_adr_i[23]
port 614 nsew signal input
rlabel metal2 s 16670 0 16726 800 6 wbs_adr_i[24]
port 615 nsew signal input
rlabel metal2 s 17314 0 17370 800 6 wbs_adr_i[25]
port 616 nsew signal input
rlabel metal2 s 17866 0 17922 800 6 wbs_adr_i[26]
port 617 nsew signal input
rlabel metal2 s 18510 0 18566 800 6 wbs_adr_i[27]
port 618 nsew signal input
rlabel metal2 s 19062 0 19118 800 6 wbs_adr_i[28]
port 619 nsew signal input
rlabel metal2 s 19706 0 19762 800 6 wbs_adr_i[29]
port 620 nsew signal input
rlabel metal2 s 2870 0 2926 800 6 wbs_adr_i[2]
port 621 nsew signal input
rlabel metal2 s 20350 0 20406 800 6 wbs_adr_i[30]
port 622 nsew signal input
rlabel metal2 s 20902 0 20958 800 6 wbs_adr_i[31]
port 623 nsew signal input
rlabel metal2 s 3698 0 3754 800 6 wbs_adr_i[3]
port 624 nsew signal input
rlabel metal2 s 4526 0 4582 800 6 wbs_adr_i[4]
port 625 nsew signal input
rlabel metal2 s 5170 0 5226 800 6 wbs_adr_i[5]
port 626 nsew signal input
rlabel metal2 s 5722 0 5778 800 6 wbs_adr_i[6]
port 627 nsew signal input
rlabel metal2 s 6366 0 6422 800 6 wbs_adr_i[7]
port 628 nsew signal input
rlabel metal2 s 6918 0 6974 800 6 wbs_adr_i[8]
port 629 nsew signal input
rlabel metal2 s 7562 0 7618 800 6 wbs_adr_i[9]
port 630 nsew signal input
rlabel metal2 s 662 0 718 800 6 wbs_cyc_i
port 631 nsew signal input
rlabel metal2 s 1490 0 1546 800 6 wbs_dat_i[0]
port 632 nsew signal input
rlabel metal2 s 8390 0 8446 800 6 wbs_dat_i[10]
port 633 nsew signal input
rlabel metal2 s 8942 0 8998 800 6 wbs_dat_i[11]
port 634 nsew signal input
rlabel metal2 s 9586 0 9642 800 6 wbs_dat_i[12]
port 635 nsew signal input
rlabel metal2 s 10230 0 10286 800 6 wbs_dat_i[13]
port 636 nsew signal input
rlabel metal2 s 10782 0 10838 800 6 wbs_dat_i[14]
port 637 nsew signal input
rlabel metal2 s 11426 0 11482 800 6 wbs_dat_i[15]
port 638 nsew signal input
rlabel metal2 s 11978 0 12034 800 6 wbs_dat_i[16]
port 639 nsew signal input
rlabel metal2 s 12622 0 12678 800 6 wbs_dat_i[17]
port 640 nsew signal input
rlabel metal2 s 13266 0 13322 800 6 wbs_dat_i[18]
port 641 nsew signal input
rlabel metal2 s 13818 0 13874 800 6 wbs_dat_i[19]
port 642 nsew signal input
rlabel metal2 s 2318 0 2374 800 6 wbs_dat_i[1]
port 643 nsew signal input
rlabel metal2 s 14462 0 14518 800 6 wbs_dat_i[20]
port 644 nsew signal input
rlabel metal2 s 15014 0 15070 800 6 wbs_dat_i[21]
port 645 nsew signal input
rlabel metal2 s 15658 0 15714 800 6 wbs_dat_i[22]
port 646 nsew signal input
rlabel metal2 s 16302 0 16358 800 6 wbs_dat_i[23]
port 647 nsew signal input
rlabel metal2 s 16854 0 16910 800 6 wbs_dat_i[24]
port 648 nsew signal input
rlabel metal2 s 17498 0 17554 800 6 wbs_dat_i[25]
port 649 nsew signal input
rlabel metal2 s 18050 0 18106 800 6 wbs_dat_i[26]
port 650 nsew signal input
rlabel metal2 s 18694 0 18750 800 6 wbs_dat_i[27]
port 651 nsew signal input
rlabel metal2 s 19338 0 19394 800 6 wbs_dat_i[28]
port 652 nsew signal input
rlabel metal2 s 19890 0 19946 800 6 wbs_dat_i[29]
port 653 nsew signal input
rlabel metal2 s 3146 0 3202 800 6 wbs_dat_i[2]
port 654 nsew signal input
rlabel metal2 s 20534 0 20590 800 6 wbs_dat_i[30]
port 655 nsew signal input
rlabel metal2 s 21086 0 21142 800 6 wbs_dat_i[31]
port 656 nsew signal input
rlabel metal2 s 3882 0 3938 800 6 wbs_dat_i[3]
port 657 nsew signal input
rlabel metal2 s 4710 0 4766 800 6 wbs_dat_i[4]
port 658 nsew signal input
rlabel metal2 s 5354 0 5410 800 6 wbs_dat_i[5]
port 659 nsew signal input
rlabel metal2 s 5906 0 5962 800 6 wbs_dat_i[6]
port 660 nsew signal input
rlabel metal2 s 6550 0 6606 800 6 wbs_dat_i[7]
port 661 nsew signal input
rlabel metal2 s 7194 0 7250 800 6 wbs_dat_i[8]
port 662 nsew signal input
rlabel metal2 s 7746 0 7802 800 6 wbs_dat_i[9]
port 663 nsew signal input
rlabel metal2 s 1674 0 1730 800 6 wbs_dat_o[0]
port 664 nsew signal output
rlabel metal2 s 8574 0 8630 800 6 wbs_dat_o[10]
port 665 nsew signal output
rlabel metal2 s 9218 0 9274 800 6 wbs_dat_o[11]
port 666 nsew signal output
rlabel metal2 s 9770 0 9826 800 6 wbs_dat_o[12]
port 667 nsew signal output
rlabel metal2 s 10414 0 10470 800 6 wbs_dat_o[13]
port 668 nsew signal output
rlabel metal2 s 10966 0 11022 800 6 wbs_dat_o[14]
port 669 nsew signal output
rlabel metal2 s 11610 0 11666 800 6 wbs_dat_o[15]
port 670 nsew signal output
rlabel metal2 s 12254 0 12310 800 6 wbs_dat_o[16]
port 671 nsew signal output
rlabel metal2 s 12806 0 12862 800 6 wbs_dat_o[17]
port 672 nsew signal output
rlabel metal2 s 13450 0 13506 800 6 wbs_dat_o[18]
port 673 nsew signal output
rlabel metal2 s 14002 0 14058 800 6 wbs_dat_o[19]
port 674 nsew signal output
rlabel metal2 s 2502 0 2558 800 6 wbs_dat_o[1]
port 675 nsew signal output
rlabel metal2 s 14646 0 14702 800 6 wbs_dat_o[20]
port 676 nsew signal output
rlabel metal2 s 15290 0 15346 800 6 wbs_dat_o[21]
port 677 nsew signal output
rlabel metal2 s 15842 0 15898 800 6 wbs_dat_o[22]
port 678 nsew signal output
rlabel metal2 s 16486 0 16542 800 6 wbs_dat_o[23]
port 679 nsew signal output
rlabel metal2 s 17038 0 17094 800 6 wbs_dat_o[24]
port 680 nsew signal output
rlabel metal2 s 17682 0 17738 800 6 wbs_dat_o[25]
port 681 nsew signal output
rlabel metal2 s 18326 0 18382 800 6 wbs_dat_o[26]
port 682 nsew signal output
rlabel metal2 s 18878 0 18934 800 6 wbs_dat_o[27]
port 683 nsew signal output
rlabel metal2 s 19522 0 19578 800 6 wbs_dat_o[28]
port 684 nsew signal output
rlabel metal2 s 20074 0 20130 800 6 wbs_dat_o[29]
port 685 nsew signal output
rlabel metal2 s 3330 0 3386 800 6 wbs_dat_o[2]
port 686 nsew signal output
rlabel metal2 s 20718 0 20774 800 6 wbs_dat_o[30]
port 687 nsew signal output
rlabel metal2 s 21362 0 21418 800 6 wbs_dat_o[31]
port 688 nsew signal output
rlabel metal2 s 4158 0 4214 800 6 wbs_dat_o[3]
port 689 nsew signal output
rlabel metal2 s 4894 0 4950 800 6 wbs_dat_o[4]
port 690 nsew signal output
rlabel metal2 s 5538 0 5594 800 6 wbs_dat_o[5]
port 691 nsew signal output
rlabel metal2 s 6182 0 6238 800 6 wbs_dat_o[6]
port 692 nsew signal output
rlabel metal2 s 6734 0 6790 800 6 wbs_dat_o[7]
port 693 nsew signal output
rlabel metal2 s 7378 0 7434 800 6 wbs_dat_o[8]
port 694 nsew signal output
rlabel metal2 s 7930 0 7986 800 6 wbs_dat_o[9]
port 695 nsew signal output
rlabel metal2 s 1858 0 1914 800 6 wbs_sel_i[0]
port 696 nsew signal input
rlabel metal2 s 2686 0 2742 800 6 wbs_sel_i[1]
port 697 nsew signal input
rlabel metal2 s 3514 0 3570 800 6 wbs_sel_i[2]
port 698 nsew signal input
rlabel metal2 s 4342 0 4398 800 6 wbs_sel_i[3]
port 699 nsew signal input
rlabel metal2 s 846 0 902 800 6 wbs_stb_i
port 700 nsew signal input
rlabel metal2 s 1122 0 1178 800 6 wbs_we_i
port 701 nsew signal input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 100000 200000
string LEFview TRUE
string GDS_FILE /project/openlane/digitalcore_macro/runs/digitalcore_macro/results/magic/digitalcore_macro.gds
string GDS_END 19806606
string GDS_START 747928
<< end >>

