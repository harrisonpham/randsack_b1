magic
tech sky130A
magscale 1 2
timestamp 1641031085
<< metal1 >>
rect 218974 700952 218980 701004
rect 219032 700992 219038 701004
rect 252554 700992 252560 701004
rect 219032 700964 252560 700992
rect 219032 700952 219038 700964
rect 252554 700952 252560 700964
rect 252612 700952 252618 701004
rect 249610 700884 249616 700936
rect 249668 700924 249674 700936
rect 348786 700924 348792 700936
rect 249668 700896 348792 700924
rect 249668 700884 249674 700896
rect 348786 700884 348792 700896
rect 348844 700884 348850 700936
rect 154114 700816 154120 700868
rect 154172 700856 154178 700868
rect 255314 700856 255320 700868
rect 154172 700828 255320 700856
rect 154172 700816 154178 700828
rect 255314 700816 255320 700828
rect 255372 700816 255378 700868
rect 137830 700748 137836 700800
rect 137888 700788 137894 700800
rect 255406 700788 255412 700800
rect 137888 700760 255412 700788
rect 137888 700748 137894 700760
rect 255406 700748 255412 700760
rect 255464 700748 255470 700800
rect 246942 700680 246948 700732
rect 247000 700720 247006 700732
rect 413646 700720 413652 700732
rect 247000 700692 413652 700720
rect 247000 700680 247006 700692
rect 413646 700680 413652 700692
rect 413704 700680 413710 700732
rect 89162 700612 89168 700664
rect 89220 700652 89226 700664
rect 258074 700652 258080 700664
rect 89220 700624 258080 700652
rect 89220 700612 89226 700624
rect 258074 700612 258080 700624
rect 258132 700612 258138 700664
rect 72970 700544 72976 700596
rect 73028 700584 73034 700596
rect 258166 700584 258172 700596
rect 73028 700556 258172 700584
rect 73028 700544 73034 700556
rect 258166 700544 258172 700556
rect 258224 700544 258230 700596
rect 40494 700476 40500 700528
rect 40552 700516 40558 700528
rect 41322 700516 41328 700528
rect 40552 700488 41328 700516
rect 40552 700476 40558 700488
rect 41322 700476 41328 700488
rect 41380 700476 41386 700528
rect 244182 700476 244188 700528
rect 244240 700516 244246 700528
rect 478506 700516 478512 700528
rect 244240 700488 478512 700516
rect 244240 700476 244246 700488
rect 478506 700476 478512 700488
rect 478564 700476 478570 700528
rect 24302 700408 24308 700460
rect 24360 700448 24366 700460
rect 260834 700448 260840 700460
rect 24360 700420 260840 700448
rect 24360 700408 24366 700420
rect 260834 700408 260840 700420
rect 260892 700408 260898 700460
rect 8110 700340 8116 700392
rect 8168 700380 8174 700392
rect 259454 700380 259460 700392
rect 8168 700352 259460 700380
rect 8168 700340 8174 700352
rect 259454 700340 259460 700352
rect 259512 700340 259518 700392
rect 284938 700340 284944 700392
rect 284996 700380 285002 700392
rect 332502 700380 332508 700392
rect 284996 700352 332508 700380
rect 284996 700340 285002 700352
rect 332502 700340 332508 700352
rect 332560 700340 332566 700392
rect 241422 700272 241428 700324
rect 241480 700312 241486 700324
rect 543458 700312 543464 700324
rect 241480 700284 543464 700312
rect 241480 700272 241486 700284
rect 543458 700272 543464 700284
rect 543516 700272 543522 700324
rect 252462 700204 252468 700256
rect 252520 700244 252526 700256
rect 283834 700244 283840 700256
rect 252520 700216 283840 700244
rect 252520 700204 252526 700216
rect 283834 700204 283840 700216
rect 283892 700204 283898 700256
rect 251082 700136 251088 700188
rect 251140 700176 251146 700188
rect 267642 700176 267648 700188
rect 251140 700148 267648 700176
rect 251140 700136 251146 700148
rect 267642 700136 267648 700148
rect 267700 700136 267706 700188
rect 105446 699660 105452 699712
rect 105504 699700 105510 699712
rect 106182 699700 106188 699712
rect 105504 699672 106188 699700
rect 105504 699660 105510 699672
rect 106182 699660 106188 699672
rect 106240 699660 106246 699712
rect 170306 699660 170312 699712
rect 170364 699700 170370 699712
rect 171042 699700 171048 699712
rect 170364 699672 171048 699700
rect 170364 699660 170370 699672
rect 171042 699660 171048 699672
rect 171100 699660 171106 699712
rect 235166 699660 235172 699712
rect 235224 699700 235230 699712
rect 240778 699700 240784 699712
rect 235224 699672 240784 699700
rect 235224 699660 235230 699672
rect 240778 699660 240784 699672
rect 240836 699660 240842 699712
rect 298738 699660 298744 699712
rect 298796 699700 298802 699712
rect 300118 699700 300124 699712
rect 298796 699672 300124 699700
rect 298796 699660 298802 699672
rect 300118 699660 300124 699672
rect 300176 699660 300182 699712
rect 359458 699660 359464 699712
rect 359516 699700 359522 699712
rect 364978 699700 364984 699712
rect 359516 699672 364984 699700
rect 359516 699660 359522 699672
rect 364978 699660 364984 699672
rect 365036 699660 365042 699712
rect 396718 699660 396724 699712
rect 396776 699700 396782 699712
rect 397454 699700 397460 699712
rect 396776 699672 397460 699700
rect 396776 699660 396782 699672
rect 397454 699660 397460 699672
rect 397512 699660 397518 699712
rect 461578 699660 461584 699712
rect 461636 699700 461642 699712
rect 462314 699700 462320 699712
rect 461636 699672 462320 699700
rect 461636 699660 461642 699672
rect 462314 699660 462320 699672
rect 462372 699660 462378 699712
rect 526438 699660 526444 699712
rect 526496 699700 526502 699712
rect 527174 699700 527180 699712
rect 526496 699672 527180 699700
rect 526496 699660 526502 699672
rect 527174 699660 527180 699672
rect 527232 699660 527238 699712
rect 238662 696940 238668 696992
rect 238720 696980 238726 696992
rect 580166 696980 580172 696992
rect 238720 696952 580172 696980
rect 238720 696940 238726 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 3418 683204 3424 683256
rect 3476 683244 3482 683256
rect 262214 683244 262220 683256
rect 3476 683216 262220 683244
rect 3476 683204 3482 683216
rect 262214 683204 262220 683216
rect 262272 683204 262278 683256
rect 238570 683136 238576 683188
rect 238628 683176 238634 683188
rect 580166 683176 580172 683188
rect 238628 683148 580172 683176
rect 238628 683136 238634 683148
rect 580166 683136 580172 683148
rect 580224 683136 580230 683188
rect 3418 670760 3424 670812
rect 3476 670800 3482 670812
rect 263594 670800 263600 670812
rect 3476 670772 263600 670800
rect 3476 670760 3482 670772
rect 263594 670760 263600 670772
rect 263652 670760 263658 670812
rect 237282 670692 237288 670744
rect 237340 670732 237346 670744
rect 580166 670732 580172 670744
rect 237340 670704 580172 670732
rect 237340 670692 237346 670704
rect 580166 670692 580172 670704
rect 580224 670692 580230 670744
rect 3418 656888 3424 656940
rect 3476 656928 3482 656940
rect 262306 656928 262312 656940
rect 3476 656900 262312 656928
rect 3476 656888 3482 656900
rect 262306 656888 262312 656900
rect 262364 656888 262370 656940
rect 235902 643084 235908 643136
rect 235960 643124 235966 643136
rect 580166 643124 580172 643136
rect 235960 643096 580172 643124
rect 235960 643084 235966 643096
rect 580166 643084 580172 643096
rect 580224 643084 580230 643136
rect 3418 632068 3424 632120
rect 3476 632108 3482 632120
rect 264974 632108 264980 632120
rect 3476 632080 264980 632108
rect 3476 632068 3482 632080
rect 264974 632068 264980 632080
rect 265032 632068 265038 632120
rect 235810 630640 235816 630692
rect 235868 630680 235874 630692
rect 580166 630680 580172 630692
rect 235868 630652 580172 630680
rect 235868 630640 235874 630652
rect 580166 630640 580172 630652
rect 580224 630640 580230 630692
rect 3142 618264 3148 618316
rect 3200 618304 3206 618316
rect 266354 618304 266360 618316
rect 3200 618276 266360 618304
rect 3200 618264 3206 618276
rect 266354 618264 266360 618276
rect 266412 618264 266418 618316
rect 234522 616836 234528 616888
rect 234580 616876 234586 616888
rect 580166 616876 580172 616888
rect 234580 616848 580172 616876
rect 234580 616836 234586 616848
rect 580166 616836 580172 616848
rect 580224 616836 580230 616888
rect 3234 605820 3240 605872
rect 3292 605860 3298 605872
rect 265066 605860 265072 605872
rect 3292 605832 265072 605860
rect 3292 605820 3298 605832
rect 265066 605820 265072 605832
rect 265124 605820 265130 605872
rect 233142 590656 233148 590708
rect 233200 590696 233206 590708
rect 579798 590696 579804 590708
rect 233200 590668 579804 590696
rect 233200 590656 233206 590668
rect 579798 590656 579804 590668
rect 579856 590656 579862 590708
rect 3326 579640 3332 579692
rect 3384 579680 3390 579692
rect 266446 579680 266452 579692
rect 3384 579652 266452 579680
rect 3384 579640 3390 579652
rect 266446 579640 266452 579652
rect 266504 579640 266510 579692
rect 233050 576852 233056 576904
rect 233108 576892 233114 576904
rect 580166 576892 580172 576904
rect 233108 576864 580172 576892
rect 233108 576852 233114 576864
rect 580166 576852 580172 576864
rect 580224 576852 580230 576904
rect 3418 565836 3424 565888
rect 3476 565876 3482 565888
rect 269114 565876 269120 565888
rect 3476 565848 269120 565876
rect 3476 565836 3482 565848
rect 269114 565836 269120 565848
rect 269172 565836 269178 565888
rect 231762 563048 231768 563100
rect 231820 563088 231826 563100
rect 579798 563088 579804 563100
rect 231820 563060 579804 563088
rect 231820 563048 231826 563060
rect 579798 563048 579804 563060
rect 579856 563048 579862 563100
rect 3418 553392 3424 553444
rect 3476 553432 3482 553444
rect 267734 553432 267740 553444
rect 3476 553404 267740 553432
rect 3476 553392 3482 553404
rect 267734 553392 267740 553404
rect 267792 553392 267798 553444
rect 230382 536800 230388 536852
rect 230440 536840 230446 536852
rect 580166 536840 580172 536852
rect 230440 536812 580172 536840
rect 230440 536800 230446 536812
rect 580166 536800 580172 536812
rect 580224 536800 580230 536852
rect 3418 527144 3424 527196
rect 3476 527184 3482 527196
rect 269206 527184 269212 527196
rect 3476 527156 269212 527184
rect 3476 527144 3482 527156
rect 269206 527144 269212 527156
rect 269264 527144 269270 527196
rect 231670 524424 231676 524476
rect 231728 524464 231734 524476
rect 580166 524464 580172 524476
rect 231728 524436 580172 524464
rect 231728 524424 231734 524436
rect 580166 524424 580172 524436
rect 580224 524424 580230 524476
rect 3418 514768 3424 514820
rect 3476 514808 3482 514820
rect 271874 514808 271880 514820
rect 3476 514780 271880 514808
rect 3476 514768 3482 514780
rect 271874 514768 271880 514780
rect 271932 514768 271938 514820
rect 229002 510620 229008 510672
rect 229060 510660 229066 510672
rect 580166 510660 580172 510672
rect 229060 510632 580172 510660
rect 229060 510620 229066 510632
rect 580166 510620 580172 510632
rect 580224 510620 580230 510672
rect 3050 500964 3056 501016
rect 3108 501004 3114 501016
rect 270494 501004 270500 501016
rect 3108 500976 270500 501004
rect 3108 500964 3114 500976
rect 270494 500964 270500 500976
rect 270552 500964 270558 501016
rect 227622 484372 227628 484424
rect 227680 484412 227686 484424
rect 580166 484412 580172 484424
rect 227680 484384 580172 484412
rect 227680 484372 227686 484384
rect 580166 484372 580172 484384
rect 580224 484372 580230 484424
rect 3418 474716 3424 474768
rect 3476 474756 3482 474768
rect 271966 474756 271972 474768
rect 3476 474728 271972 474756
rect 3476 474716 3482 474728
rect 271966 474716 271972 474728
rect 272024 474716 272030 474768
rect 228910 470568 228916 470620
rect 228968 470608 228974 470620
rect 579982 470608 579988 470620
rect 228968 470580 579988 470608
rect 228968 470568 228974 470580
rect 579982 470568 579988 470580
rect 580040 470568 580046 470620
rect 3234 462340 3240 462392
rect 3292 462380 3298 462392
rect 273254 462380 273260 462392
rect 3292 462352 273260 462380
rect 3292 462340 3298 462352
rect 273254 462340 273260 462352
rect 273312 462340 273318 462392
rect 226242 456764 226248 456816
rect 226300 456804 226306 456816
rect 580166 456804 580172 456816
rect 226300 456776 580172 456804
rect 226300 456764 226306 456776
rect 580166 456764 580172 456776
rect 580224 456764 580230 456816
rect 3142 448536 3148 448588
rect 3200 448576 3206 448588
rect 273346 448576 273352 448588
rect 3200 448548 273352 448576
rect 3200 448536 3206 448548
rect 273346 448536 273352 448548
rect 273404 448536 273410 448588
rect 224862 430584 224868 430636
rect 224920 430624 224926 430636
rect 580166 430624 580172 430636
rect 224920 430596 580172 430624
rect 224920 430584 224926 430596
rect 580166 430584 580172 430596
rect 580224 430584 580230 430636
rect 3418 422288 3424 422340
rect 3476 422328 3482 422340
rect 274634 422328 274640 422340
rect 3476 422300 274640 422328
rect 3476 422288 3482 422300
rect 274634 422288 274640 422300
rect 274692 422288 274698 422340
rect 226150 418140 226156 418192
rect 226208 418180 226214 418192
rect 580166 418180 580172 418192
rect 226208 418152 580172 418180
rect 226208 418140 226214 418152
rect 580166 418140 580172 418152
rect 580224 418140 580230 418192
rect 3142 409844 3148 409896
rect 3200 409884 3206 409896
rect 276014 409884 276020 409896
rect 3200 409856 276020 409884
rect 3200 409844 3206 409856
rect 276014 409844 276020 409856
rect 276072 409844 276078 409896
rect 224770 404336 224776 404388
rect 224828 404376 224834 404388
rect 580166 404376 580172 404388
rect 224828 404348 580172 404376
rect 224828 404336 224834 404348
rect 580166 404336 580172 404348
rect 580224 404336 580230 404388
rect 3418 397468 3424 397520
rect 3476 397508 3482 397520
rect 276106 397508 276112 397520
rect 3476 397480 276112 397508
rect 3476 397468 3482 397480
rect 276106 397468 276112 397480
rect 276164 397468 276170 397520
rect 222010 378156 222016 378208
rect 222068 378196 222074 378208
rect 580166 378196 580172 378208
rect 222068 378168 580172 378196
rect 222068 378156 222074 378168
rect 580166 378156 580172 378168
rect 580224 378156 580230 378208
rect 3418 371220 3424 371272
rect 3476 371260 3482 371272
rect 277394 371260 277400 371272
rect 3476 371232 277400 371260
rect 3476 371220 3482 371232
rect 277394 371220 277400 371232
rect 277452 371220 277458 371272
rect 371602 368568 371608 368620
rect 371660 368608 371666 368620
rect 376754 368608 376760 368620
rect 371660 368580 376760 368608
rect 371660 368568 371666 368580
rect 376754 368568 376760 368580
rect 376812 368568 376818 368620
rect 371694 368500 371700 368552
rect 371752 368540 371758 368552
rect 381078 368540 381084 368552
rect 371752 368512 381084 368540
rect 371752 368500 371758 368512
rect 381078 368500 381084 368512
rect 381136 368500 381142 368552
rect 445202 368500 445208 368552
rect 445260 368540 445266 368552
rect 452838 368540 452844 368552
rect 445260 368512 452844 368540
rect 445260 368500 445266 368512
rect 452838 368500 452844 368512
rect 452896 368500 452902 368552
rect 371602 367480 371608 367532
rect 371660 367520 371666 367532
rect 373994 367520 374000 367532
rect 371660 367492 374000 367520
rect 371660 367480 371666 367492
rect 373994 367480 374000 367492
rect 374052 367480 374058 367532
rect 445662 367208 445668 367260
rect 445720 367248 445726 367260
rect 452654 367248 452660 367260
rect 445720 367220 452660 367248
rect 445720 367208 445726 367220
rect 452654 367208 452660 367220
rect 452712 367208 452718 367260
rect 371510 367072 371516 367124
rect 371568 367112 371574 367124
rect 380986 367112 380992 367124
rect 371568 367084 380992 367112
rect 371568 367072 371574 367084
rect 380986 367072 380992 367084
rect 381044 367072 381050 367124
rect 371602 365848 371608 365900
rect 371660 365888 371666 365900
rect 378226 365888 378232 365900
rect 371660 365860 378232 365888
rect 371660 365848 371666 365860
rect 378226 365848 378232 365860
rect 378284 365848 378290 365900
rect 371234 365780 371240 365832
rect 371292 365820 371298 365832
rect 375374 365820 375380 365832
rect 371292 365792 375380 365820
rect 371292 365780 371298 365792
rect 375374 365780 375380 365792
rect 375432 365780 375438 365832
rect 444926 365712 444932 365764
rect 444984 365752 444990 365764
rect 448606 365752 448612 365764
rect 444984 365724 448612 365752
rect 444984 365712 444990 365724
rect 448606 365712 448612 365724
rect 448664 365712 448670 365764
rect 371234 364692 371240 364744
rect 371292 364732 371298 364744
rect 374454 364732 374460 364744
rect 371292 364704 374460 364732
rect 371292 364692 371298 364704
rect 374454 364692 374460 364704
rect 374512 364692 374518 364744
rect 444926 364624 444932 364676
rect 444984 364664 444990 364676
rect 449986 364664 449992 364676
rect 444984 364636 449992 364664
rect 444984 364624 444990 364636
rect 449986 364624 449992 364636
rect 450044 364624 450050 364676
rect 371602 364352 371608 364404
rect 371660 364392 371666 364404
rect 378318 364392 378324 364404
rect 371660 364364 378324 364392
rect 371660 364352 371666 364364
rect 378318 364352 378324 364364
rect 378376 364352 378382 364404
rect 371602 363672 371608 363724
rect 371660 363712 371666 363724
rect 375742 363712 375748 363724
rect 371660 363684 375748 363712
rect 371660 363672 371666 363684
rect 375742 363672 375748 363684
rect 375800 363672 375806 363724
rect 444558 363128 444564 363180
rect 444616 363168 444622 363180
rect 447410 363168 447416 363180
rect 444616 363140 447416 363168
rect 444616 363128 444622 363140
rect 447410 363128 447416 363140
rect 447468 363128 447474 363180
rect 371418 362992 371424 363044
rect 371476 363032 371482 363044
rect 377030 363032 377036 363044
rect 371476 363004 377036 363032
rect 371476 362992 371482 363004
rect 377030 362992 377036 363004
rect 377088 362992 377094 363044
rect 371694 362924 371700 362976
rect 371752 362964 371758 362976
rect 378410 362964 378416 362976
rect 371752 362936 378416 362964
rect 371752 362924 371758 362936
rect 378410 362924 378416 362936
rect 378468 362924 378474 362976
rect 371418 361564 371424 361616
rect 371476 361604 371482 361616
rect 376846 361604 376852 361616
rect 371476 361576 376852 361604
rect 371476 361564 371482 361576
rect 376846 361564 376852 361576
rect 376904 361564 376910 361616
rect 444926 361564 444932 361616
rect 444984 361604 444990 361616
rect 450078 361604 450084 361616
rect 444984 361576 450084 361604
rect 444984 361564 444990 361576
rect 450078 361564 450084 361576
rect 450136 361564 450142 361616
rect 371602 360408 371608 360460
rect 371660 360448 371666 360460
rect 375558 360448 375564 360460
rect 371660 360420 375564 360448
rect 371660 360408 371666 360420
rect 375558 360408 375564 360420
rect 375616 360408 375622 360460
rect 371694 360340 371700 360392
rect 371752 360380 371758 360392
rect 374270 360380 374276 360392
rect 371752 360352 374276 360380
rect 371752 360340 371758 360352
rect 374270 360340 374276 360352
rect 374328 360340 374334 360392
rect 371510 360204 371516 360256
rect 371568 360244 371574 360256
rect 375466 360244 375472 360256
rect 371568 360216 375472 360244
rect 371568 360204 371574 360216
rect 375466 360204 375472 360216
rect 375524 360204 375530 360256
rect 445662 360204 445668 360256
rect 445720 360244 445726 360256
rect 449894 360244 449900 360256
rect 445720 360216 449900 360244
rect 445720 360204 445726 360216
rect 449894 360204 449900 360216
rect 449952 360204 449958 360256
rect 371878 359456 371884 359508
rect 371936 359496 371942 359508
rect 379514 359496 379520 359508
rect 371936 359468 379520 359496
rect 371936 359456 371942 359468
rect 379514 359456 379520 359468
rect 379572 359456 379578 359508
rect 371326 358776 371332 358828
rect 371384 358816 371390 358828
rect 383654 358816 383660 358828
rect 371384 358788 383660 358816
rect 371384 358776 371390 358788
rect 383654 358776 383660 358788
rect 383712 358776 383718 358828
rect 444466 358776 444472 358828
rect 444524 358816 444530 358828
rect 447226 358816 447232 358828
rect 444524 358788 447232 358816
rect 444524 358776 444530 358788
rect 447226 358776 447232 358788
rect 447284 358776 447290 358828
rect 371418 357688 371424 357740
rect 371476 357728 371482 357740
rect 375650 357728 375656 357740
rect 371476 357700 375656 357728
rect 371476 357688 371482 357700
rect 375650 357688 375656 357700
rect 375708 357688 375714 357740
rect 3142 357416 3148 357468
rect 3200 357456 3206 357468
rect 278774 357456 278780 357468
rect 3200 357428 278780 357456
rect 3200 357416 3206 357428
rect 278774 357416 278780 357428
rect 278832 357416 278838 357468
rect 371510 357416 371516 357468
rect 371568 357456 371574 357468
rect 382458 357456 382464 357468
rect 371568 357428 382464 357456
rect 371568 357416 371574 357428
rect 382458 357416 382464 357428
rect 382516 357416 382522 357468
rect 444926 357416 444932 357468
rect 444984 357456 444990 357468
rect 448882 357456 448888 357468
rect 444984 357428 448888 357456
rect 444984 357416 444990 357428
rect 448882 357416 448888 357428
rect 448940 357416 448946 357468
rect 444558 356736 444564 356788
rect 444616 356776 444622 356788
rect 448698 356776 448704 356788
rect 444616 356748 448704 356776
rect 444616 356736 444622 356748
rect 448698 356736 448704 356748
rect 448756 356736 448762 356788
rect 371326 356192 371332 356244
rect 371384 356232 371390 356244
rect 378134 356232 378140 356244
rect 371384 356204 378140 356232
rect 371384 356192 371390 356204
rect 378134 356192 378140 356204
rect 378192 356192 378198 356244
rect 371234 356124 371240 356176
rect 371292 356164 371298 356176
rect 381170 356164 381176 356176
rect 371292 356136 381176 356164
rect 371292 356124 371298 356136
rect 381170 356124 381176 356136
rect 381228 356124 381234 356176
rect 371418 356056 371424 356108
rect 371476 356096 371482 356108
rect 382274 356096 382280 356108
rect 371476 356068 382280 356096
rect 371476 356056 371482 356068
rect 382274 356056 382280 356068
rect 382332 356056 382338 356108
rect 444374 355104 444380 355156
rect 444432 355144 444438 355156
rect 446030 355144 446036 355156
rect 444432 355116 446036 355144
rect 444432 355104 444438 355116
rect 446030 355104 446036 355116
rect 446088 355104 446094 355156
rect 371234 354968 371240 355020
rect 371292 355008 371298 355020
rect 372890 355008 372896 355020
rect 371292 354980 372896 355008
rect 371292 354968 371298 354980
rect 372890 354968 372896 354980
rect 372948 354968 372954 355020
rect 371694 354764 371700 354816
rect 371752 354804 371758 354816
rect 376938 354804 376944 354816
rect 371752 354776 376944 354804
rect 371752 354764 371758 354776
rect 376938 354764 376944 354776
rect 376996 354764 377002 354816
rect 371510 354152 371516 354204
rect 371568 354192 371574 354204
rect 374178 354192 374184 354204
rect 371568 354164 374184 354192
rect 371568 354152 371574 354164
rect 374178 354152 374184 354164
rect 374236 354152 374242 354204
rect 444466 353336 444472 353388
rect 444524 353376 444530 353388
rect 447318 353376 447324 353388
rect 444524 353348 447324 353376
rect 444524 353336 444530 353348
rect 447318 353336 447324 353348
rect 447376 353336 447382 353388
rect 371694 353268 371700 353320
rect 371752 353308 371758 353320
rect 374086 353308 374092 353320
rect 371752 353280 374092 353308
rect 371752 353268 371758 353280
rect 374086 353268 374092 353280
rect 374144 353268 374150 353320
rect 372062 352588 372068 352640
rect 372120 352628 372126 352640
rect 377122 352628 377128 352640
rect 372120 352600 377128 352628
rect 372120 352588 372126 352600
rect 377122 352588 377128 352600
rect 377180 352588 377186 352640
rect 372246 352520 372252 352572
rect 372304 352560 372310 352572
rect 379606 352560 379612 352572
rect 372304 352532 379612 352560
rect 372304 352520 372310 352532
rect 379606 352520 379612 352532
rect 379664 352520 379670 352572
rect 444374 351976 444380 352028
rect 444432 352016 444438 352028
rect 447134 352016 447140 352028
rect 444432 351988 447140 352016
rect 444432 351976 444438 351988
rect 447134 351976 447140 351988
rect 447192 351976 447198 352028
rect 371602 348168 371608 348220
rect 371660 348208 371666 348220
rect 374362 348208 374368 348220
rect 371660 348180 374368 348208
rect 371660 348168 371666 348180
rect 374362 348168 374368 348180
rect 374420 348168 374426 348220
rect 445202 345584 445208 345636
rect 445260 345624 445266 345636
rect 450170 345624 450176 345636
rect 445260 345596 450176 345624
rect 445260 345584 445266 345596
rect 450170 345584 450176 345596
rect 450228 345584 450234 345636
rect 445662 345108 445668 345160
rect 445720 345148 445726 345160
rect 452746 345148 452752 345160
rect 445720 345120 452752 345148
rect 445720 345108 445726 345120
rect 452746 345108 452752 345120
rect 452804 345108 452810 345160
rect 3326 345040 3332 345092
rect 3384 345080 3390 345092
rect 278866 345080 278872 345092
rect 3384 345052 278872 345080
rect 3384 345040 3390 345052
rect 278866 345040 278872 345052
rect 278924 345040 278930 345092
rect 445662 343612 445668 343664
rect 445720 343652 445726 343664
rect 454034 343652 454040 343664
rect 445720 343624 454040 343652
rect 445720 343612 445726 343624
rect 454034 343612 454040 343624
rect 454092 343612 454098 343664
rect 445662 342252 445668 342304
rect 445720 342292 445726 342304
rect 451366 342292 451372 342304
rect 445720 342264 451372 342292
rect 445720 342252 445726 342264
rect 451366 342252 451372 342264
rect 451424 342252 451430 342304
rect 445110 340960 445116 341012
rect 445168 341000 445174 341012
rect 448790 341000 448796 341012
rect 445168 340972 448796 341000
rect 445168 340960 445174 340972
rect 448790 340960 448796 340972
rect 448848 340960 448854 341012
rect 444742 340212 444748 340264
rect 444800 340252 444806 340264
rect 446122 340252 446128 340264
rect 444800 340224 446128 340252
rect 444800 340212 444806 340224
rect 446122 340212 446128 340224
rect 446180 340212 446186 340264
rect 299934 337424 299940 337476
rect 299992 337464 299998 337476
rect 438946 337464 438952 337476
rect 299992 337436 438952 337464
rect 299992 337424 299998 337436
rect 438946 337424 438952 337436
rect 439004 337424 439010 337476
rect 198550 337356 198556 337408
rect 198608 337396 198614 337408
rect 366910 337396 366916 337408
rect 198608 337368 366916 337396
rect 198608 337356 198614 337368
rect 366910 337356 366916 337368
rect 366968 337356 366974 337408
rect 441246 336744 441252 336796
rect 441304 336784 441310 336796
rect 441614 336784 441620 336796
rect 441304 336756 441620 336784
rect 441304 336744 441310 336756
rect 441614 336744 441620 336756
rect 441672 336744 441678 336796
rect 368934 335316 368940 335368
rect 368992 335356 368998 335368
rect 369118 335356 369124 335368
rect 368992 335328 369124 335356
rect 368992 335316 368998 335328
rect 369118 335316 369124 335328
rect 369176 335316 369182 335368
rect 245562 327700 245568 327752
rect 245620 327740 245626 327752
rect 396718 327740 396724 327752
rect 245620 327712 396724 327740
rect 245620 327700 245626 327712
rect 396718 327700 396724 327712
rect 396776 327700 396782 327752
rect 219342 324300 219348 324352
rect 219400 324340 219406 324352
rect 580166 324340 580172 324352
rect 219400 324312 580172 324340
rect 219400 324300 219406 324312
rect 580166 324300 580172 324312
rect 580224 324300 580230 324352
rect 242710 323552 242716 323604
rect 242768 323592 242774 323604
rect 461578 323592 461584 323604
rect 242768 323564 461584 323592
rect 242768 323552 242774 323564
rect 461578 323552 461584 323564
rect 461636 323552 461642 323604
rect 3418 318792 3424 318844
rect 3476 318832 3482 318844
rect 280246 318832 280252 318844
rect 3476 318804 280252 318832
rect 3476 318792 3482 318804
rect 280246 318792 280252 318804
rect 280304 318792 280310 318844
rect 220630 311856 220636 311908
rect 220688 311896 220694 311908
rect 580166 311896 580172 311908
rect 220688 311868 580172 311896
rect 220688 311856 220694 311868
rect 580166 311856 580172 311868
rect 580224 311856 580230 311908
rect 202782 305872 202788 305924
rect 202840 305912 202846 305924
rect 252922 305912 252928 305924
rect 202840 305884 252928 305912
rect 202840 305872 202846 305884
rect 252922 305872 252928 305884
rect 252980 305872 252986 305924
rect 246850 305804 246856 305856
rect 246908 305844 246914 305856
rect 359458 305844 359464 305856
rect 246908 305816 359464 305844
rect 246908 305804 246914 305816
rect 359458 305804 359464 305816
rect 359516 305804 359522 305856
rect 244274 305736 244280 305788
rect 244332 305776 244338 305788
rect 429194 305776 429200 305788
rect 244332 305748 429200 305776
rect 244332 305736 244338 305748
rect 429194 305736 429200 305748
rect 429252 305736 429258 305788
rect 41322 305668 41328 305720
rect 41380 305708 41386 305720
rect 259822 305708 259828 305720
rect 41380 305680 259828 305708
rect 41380 305668 41386 305680
rect 259822 305668 259828 305680
rect 259880 305668 259886 305720
rect 240042 305600 240048 305652
rect 240100 305640 240106 305652
rect 526438 305640 526444 305652
rect 240100 305612 526444 305640
rect 240100 305600 240106 305612
rect 526438 305600 526444 305612
rect 526496 305600 526502 305652
rect 3234 304988 3240 305040
rect 3292 305028 3298 305040
rect 282270 305028 282276 305040
rect 3292 305000 282276 305028
rect 3292 304988 3298 305000
rect 282270 304988 282276 305000
rect 282328 304988 282334 305040
rect 240778 304784 240784 304836
rect 240836 304824 240842 304836
rect 252094 304824 252100 304836
rect 240836 304796 252100 304824
rect 240836 304784 240842 304796
rect 252094 304784 252100 304796
rect 252152 304784 252158 304836
rect 247770 304716 247776 304768
rect 247828 304756 247834 304768
rect 284938 304756 284944 304768
rect 247828 304728 284944 304756
rect 247828 304716 247834 304728
rect 284938 304716 284944 304728
rect 284996 304716 285002 304768
rect 249518 304648 249524 304700
rect 249576 304688 249582 304700
rect 298738 304688 298744 304700
rect 249576 304660 298744 304688
rect 249576 304648 249582 304660
rect 298738 304648 298744 304660
rect 298796 304648 298802 304700
rect 171042 304580 171048 304632
rect 171100 304620 171106 304632
rect 254670 304620 254676 304632
rect 171100 304592 254676 304620
rect 171100 304580 171106 304592
rect 254670 304580 254676 304592
rect 254728 304580 254734 304632
rect 106182 304512 106188 304564
rect 106240 304552 106246 304564
rect 257246 304552 257252 304564
rect 106240 304524 257252 304552
rect 106240 304512 106246 304524
rect 257246 304512 257252 304524
rect 257304 304512 257310 304564
rect 241698 304444 241704 304496
rect 241756 304484 241762 304496
rect 494054 304484 494060 304496
rect 241756 304456 494060 304484
rect 241756 304444 241762 304456
rect 494054 304444 494060 304456
rect 494112 304444 494118 304496
rect 239122 304376 239128 304428
rect 239180 304416 239186 304428
rect 558914 304416 558920 304428
rect 239180 304388 558920 304416
rect 239180 304376 239186 304388
rect 558914 304376 558920 304388
rect 558972 304376 558978 304428
rect 222746 304308 222752 304360
rect 222804 304348 222810 304360
rect 580258 304348 580264 304360
rect 222804 304320 580264 304348
rect 222804 304308 222810 304320
rect 580258 304308 580264 304320
rect 580316 304308 580322 304360
rect 220998 304240 221004 304292
rect 221056 304280 221062 304292
rect 580350 304280 580356 304292
rect 221056 304252 580356 304280
rect 221056 304240 221062 304252
rect 580350 304240 580356 304252
rect 580408 304240 580414 304292
rect 237374 303016 237380 303068
rect 237432 303056 237438 303068
rect 238662 303056 238668 303068
rect 237432 303028 238668 303056
rect 237432 303016 237438 303028
rect 238662 303016 238668 303028
rect 238720 303016 238726 303068
rect 243446 303016 243452 303068
rect 243504 303056 243510 303068
rect 244182 303056 244188 303068
rect 243504 303028 244188 303056
rect 243504 303016 243510 303028
rect 244182 303016 244188 303028
rect 244240 303016 244246 303068
rect 246022 303016 246028 303068
rect 246080 303056 246086 303068
rect 246942 303056 246948 303068
rect 246080 303028 246948 303056
rect 246080 303016 246086 303028
rect 246942 303016 246948 303028
rect 247000 303016 247006 303068
rect 248598 303016 248604 303068
rect 248656 303056 248662 303068
rect 249610 303056 249616 303068
rect 248656 303028 249616 303056
rect 248656 303016 248662 303028
rect 249610 303016 249616 303028
rect 249668 303016 249674 303068
rect 251174 303016 251180 303068
rect 251232 303056 251238 303068
rect 252462 303056 252468 303068
rect 251232 303028 252468 303056
rect 251232 303016 251238 303028
rect 252462 303016 252468 303028
rect 252520 303016 252526 303068
rect 255314 303016 255320 303068
rect 255372 303056 255378 303068
rect 256142 303056 256148 303068
rect 255372 303028 256148 303056
rect 255372 303016 255378 303028
rect 256142 303016 256148 303028
rect 256200 303016 256206 303068
rect 273254 303016 273260 303068
rect 273312 303056 273318 303068
rect 274174 303056 274180 303068
rect 273312 303028 274180 303056
rect 273312 303016 273318 303028
rect 274174 303016 274180 303028
rect 274232 303016 274238 303068
rect 215018 302948 215024 303000
rect 215076 302988 215082 303000
rect 316678 302988 316684 303000
rect 215076 302960 316684 302988
rect 215076 302948 215082 302960
rect 316678 302948 316684 302960
rect 316736 302948 316742 303000
rect 177390 302880 177396 302932
rect 177448 302920 177454 302932
rect 287422 302920 287428 302932
rect 177448 302892 287428 302920
rect 177448 302880 177454 302892
rect 287422 302880 287428 302892
rect 287480 302880 287486 302932
rect 178678 302812 178684 302864
rect 178736 302852 178742 302864
rect 298646 302852 298652 302864
rect 178736 302824 298652 302852
rect 178736 302812 178742 302824
rect 298646 302812 298652 302824
rect 298704 302812 298710 302864
rect 214098 302744 214104 302796
rect 214156 302784 214162 302796
rect 447962 302784 447968 302796
rect 214156 302756 447968 302784
rect 214156 302744 214162 302756
rect 447962 302744 447968 302756
rect 448020 302744 448026 302796
rect 211522 302676 211528 302728
rect 211580 302716 211586 302728
rect 446398 302716 446404 302728
rect 211580 302688 446404 302716
rect 211580 302676 211586 302688
rect 446398 302676 446404 302688
rect 446456 302676 446462 302728
rect 217594 302608 217600 302660
rect 217652 302648 217658 302660
rect 464338 302648 464344 302660
rect 217652 302620 464344 302648
rect 217652 302608 217658 302620
rect 464338 302608 464344 302620
rect 464396 302608 464402 302660
rect 212442 302540 212448 302592
rect 212500 302580 212506 302592
rect 461578 302580 461584 302592
rect 212500 302552 461584 302580
rect 212500 302540 212506 302552
rect 461578 302540 461584 302552
rect 461636 302540 461642 302592
rect 207198 302472 207204 302524
rect 207256 302512 207262 302524
rect 457438 302512 457444 302524
rect 207256 302484 457444 302512
rect 207256 302472 207262 302484
rect 457438 302472 457444 302484
rect 457496 302472 457502 302524
rect 204622 302404 204628 302456
rect 204680 302444 204686 302456
rect 454678 302444 454684 302456
rect 204680 302416 454684 302444
rect 204680 302404 204686 302416
rect 454678 302404 454684 302416
rect 454736 302404 454742 302456
rect 202046 302336 202052 302388
rect 202104 302376 202110 302388
rect 453298 302376 453304 302388
rect 202104 302348 453304 302376
rect 202104 302336 202110 302348
rect 453298 302336 453304 302348
rect 453356 302336 453362 302388
rect 14458 302268 14464 302320
rect 14516 302308 14522 302320
rect 292574 302308 292580 302320
rect 14516 302280 292580 302308
rect 14516 302268 14522 302280
rect 292574 302268 292580 302280
rect 292632 302268 292638 302320
rect 11698 302200 11704 302252
rect 11756 302240 11762 302252
rect 289998 302240 290004 302252
rect 11756 302212 290004 302240
rect 11756 302200 11762 302212
rect 289998 302200 290004 302212
rect 290056 302200 290062 302252
rect 230474 302132 230480 302184
rect 230532 302172 230538 302184
rect 231670 302172 231676 302184
rect 230532 302144 231676 302172
rect 230532 302132 230538 302144
rect 231670 302132 231676 302144
rect 231728 302132 231734 302184
rect 229646 302064 229652 302116
rect 229704 302104 229710 302116
rect 230382 302104 230388 302116
rect 229704 302076 230388 302104
rect 229704 302064 229710 302076
rect 230382 302064 230388 302076
rect 230440 302064 230446 302116
rect 232222 302064 232228 302116
rect 232280 302104 232286 302116
rect 233142 302104 233148 302116
rect 232280 302076 233148 302104
rect 232280 302064 232286 302076
rect 233142 302064 233148 302076
rect 233200 302064 233206 302116
rect 258074 302064 258080 302116
rect 258132 302104 258138 302116
rect 258994 302104 259000 302116
rect 258132 302076 259000 302104
rect 258132 302064 258138 302076
rect 258994 302064 259000 302076
rect 259052 302064 259058 302116
rect 278774 302064 278780 302116
rect 278832 302104 278838 302116
rect 279694 302104 279700 302116
rect 278832 302076 279700 302104
rect 278832 302064 278838 302076
rect 279694 302064 279700 302076
rect 279752 302064 279758 302116
rect 276014 301792 276020 301844
rect 276072 301832 276078 301844
rect 277026 301832 277032 301844
rect 276072 301804 277032 301832
rect 276072 301792 276078 301804
rect 277026 301792 277032 301804
rect 277084 301792 277090 301844
rect 196618 301656 196624 301708
rect 196676 301696 196682 301708
rect 281350 301696 281356 301708
rect 196676 301668 281356 301696
rect 196676 301656 196682 301668
rect 281350 301656 281356 301668
rect 281408 301656 281414 301708
rect 199378 301588 199384 301640
rect 199436 301628 199442 301640
rect 285674 301628 285680 301640
rect 199436 301600 285680 301628
rect 199436 301588 199442 301600
rect 285674 301588 285680 301600
rect 285732 301588 285738 301640
rect 215846 301520 215852 301572
rect 215904 301560 215910 301572
rect 304258 301560 304264 301572
rect 215904 301532 304264 301560
rect 215904 301520 215910 301532
rect 304258 301520 304264 301532
rect 304316 301520 304322 301572
rect 210694 301452 210700 301504
rect 210752 301492 210758 301504
rect 301498 301492 301504 301504
rect 210752 301464 301504 301492
rect 210752 301452 210758 301464
rect 301498 301452 301504 301464
rect 301556 301452 301562 301504
rect 203794 301384 203800 301436
rect 203852 301424 203858 301436
rect 309778 301424 309784 301436
rect 203852 301396 309784 301424
rect 203852 301384 203858 301396
rect 309778 301384 309784 301396
rect 309836 301384 309842 301436
rect 159358 301316 159364 301368
rect 159416 301356 159422 301368
rect 288250 301356 288256 301368
rect 159416 301328 288256 301356
rect 159416 301316 159422 301328
rect 288250 301316 288256 301328
rect 288308 301316 288314 301368
rect 151078 301248 151084 301300
rect 151136 301288 151142 301300
rect 291746 301288 291752 301300
rect 151136 301260 291752 301288
rect 151136 301248 151142 301260
rect 291746 301248 291752 301260
rect 291804 301248 291810 301300
rect 146938 301180 146944 301232
rect 146996 301220 147002 301232
rect 295150 301220 295156 301232
rect 146996 301192 295156 301220
rect 146996 301180 147002 301192
rect 295150 301180 295156 301192
rect 295208 301180 295214 301232
rect 209866 301112 209872 301164
rect 209924 301152 209930 301164
rect 465718 301152 465724 301164
rect 209924 301124 465724 301152
rect 209924 301112 209930 301124
rect 465718 301112 465724 301124
rect 465776 301112 465782 301164
rect 17218 301044 17224 301096
rect 17276 301084 17282 301096
rect 283098 301084 283104 301096
rect 17276 301056 283104 301084
rect 17276 301044 17282 301056
rect 283098 301044 283104 301056
rect 283156 301044 283162 301096
rect 7558 300976 7564 301028
rect 7616 301016 7622 301028
rect 296898 301016 296904 301028
rect 7616 300988 296904 301016
rect 7616 300976 7622 300988
rect 296898 300976 296904 300988
rect 296956 300976 296962 301028
rect 202966 300908 202972 300960
rect 203024 300948 203030 300960
rect 582466 300948 582472 300960
rect 203024 300920 582472 300948
rect 203024 300908 203030 300920
rect 582466 300908 582472 300920
rect 582524 300908 582530 300960
rect 200390 300840 200396 300892
rect 200448 300880 200454 300892
rect 582374 300880 582380 300892
rect 200448 300852 582380 300880
rect 200448 300840 200454 300852
rect 582374 300840 582380 300852
rect 582432 300840 582438 300892
rect 234798 300432 234804 300484
rect 234856 300472 234862 300484
rect 235902 300472 235908 300484
rect 234856 300444 235908 300472
rect 234856 300432 234862 300444
rect 235902 300432 235908 300444
rect 235960 300432 235966 300484
rect 223666 300296 223672 300348
rect 223724 300336 223730 300348
rect 224770 300336 224776 300348
rect 223724 300308 224776 300336
rect 223724 300296 223730 300308
rect 224770 300296 224776 300308
rect 224828 300296 224834 300348
rect 225322 300296 225328 300348
rect 225380 300336 225386 300348
rect 226150 300336 226156 300348
rect 225380 300308 226156 300336
rect 225380 300296 225386 300308
rect 226150 300296 226156 300308
rect 226208 300296 226214 300348
rect 227898 300296 227904 300348
rect 227956 300336 227962 300348
rect 228910 300336 228916 300348
rect 227956 300308 228916 300336
rect 227956 300296 227962 300308
rect 228910 300296 228916 300308
rect 228968 300296 228974 300348
rect 205542 300228 205548 300280
rect 205600 300268 205606 300280
rect 307018 300268 307024 300280
rect 205600 300240 307024 300268
rect 205600 300228 205606 300240
rect 307018 300228 307024 300240
rect 307076 300228 307082 300280
rect 201218 300160 201224 300212
rect 201276 300200 201282 300212
rect 305638 300200 305644 300212
rect 201276 300172 305644 300200
rect 201276 300160 201282 300172
rect 305638 300160 305644 300172
rect 305696 300160 305702 300212
rect 206370 300092 206376 300144
rect 206428 300132 206434 300144
rect 313918 300132 313924 300144
rect 206428 300104 313924 300132
rect 206428 300092 206434 300104
rect 313918 300092 313924 300104
rect 313976 300092 313982 300144
rect 170398 300024 170404 300076
rect 170456 300064 170462 300076
rect 290550 300064 290556 300076
rect 170456 300036 290556 300064
rect 170456 300024 170462 300036
rect 290550 300024 290556 300036
rect 290608 300024 290614 300076
rect 152458 299956 152464 300008
rect 152516 299996 152522 300008
rect 288894 299996 288900 300008
rect 152516 299968 288900 299996
rect 152516 299956 152522 299968
rect 288894 299956 288900 299968
rect 288952 299956 288958 300008
rect 155218 299888 155224 299940
rect 155276 299928 155282 299940
rect 295702 299928 295708 299940
rect 155276 299900 295708 299928
rect 155276 299888 155282 299900
rect 295702 299888 295708 299900
rect 295760 299888 295766 299940
rect 148318 299820 148324 299872
rect 148376 299860 148382 299872
rect 294046 299860 294052 299872
rect 148376 299832 294052 299860
rect 148376 299820 148382 299832
rect 294046 299820 294052 299832
rect 294104 299820 294110 299872
rect 144178 299752 144184 299804
rect 144236 299792 144242 299804
rect 297358 299792 297364 299804
rect 144236 299764 297364 299792
rect 144236 299752 144242 299764
rect 297358 299752 297364 299764
rect 297416 299752 297422 299804
rect 209314 299684 209320 299736
rect 209372 299724 209378 299736
rect 443638 299724 443644 299736
rect 209372 299696 443644 299724
rect 209372 299684 209378 299696
rect 443638 299684 443644 299696
rect 443696 299684 443702 299736
rect 213546 299616 213552 299668
rect 213604 299656 213610 299668
rect 450538 299656 450544 299668
rect 213604 299628 450544 299656
rect 213604 299616 213610 299628
rect 450538 299616 450544 299628
rect 450596 299616 450602 299668
rect 208302 299548 208308 299600
rect 208360 299588 208366 299600
rect 449158 299588 449164 299600
rect 208360 299560 449164 299588
rect 208360 299548 208366 299560
rect 449158 299548 449164 299560
rect 449216 299548 449222 299600
rect 4798 299480 4804 299532
rect 4856 299520 4862 299532
rect 293126 299520 293132 299532
rect 4856 299492 293132 299520
rect 4856 299480 4862 299492
rect 293126 299480 293132 299492
rect 293184 299480 293190 299532
rect 216674 299412 216680 299464
rect 216732 299452 216738 299464
rect 220078 299452 220084 299464
rect 216732 299424 220084 299452
rect 216732 299412 216738 299424
rect 220078 299412 220084 299424
rect 220136 299412 220142 299464
rect 237190 299412 237196 299464
rect 237248 299452 237254 299464
rect 237248 299424 244274 299452
rect 237248 299412 237254 299424
rect 212506 299356 242296 299384
rect 199838 298460 199844 298512
rect 199896 298500 199902 298512
rect 212506 298500 212534 299356
rect 216674 299316 216680 299328
rect 216646 299276 216680 299316
rect 216732 299276 216738 299328
rect 217134 299276 217140 299328
rect 217192 299276 217198 299328
rect 218054 299276 218060 299328
rect 218112 299276 218118 299328
rect 218146 299276 218152 299328
rect 218204 299276 218210 299328
rect 218698 299276 218704 299328
rect 218756 299276 218762 299328
rect 218790 299276 218796 299328
rect 218848 299276 218854 299328
rect 219894 299276 219900 299328
rect 219952 299276 219958 299328
rect 220078 299276 220084 299328
rect 220136 299316 220142 299328
rect 237190 299316 237196 299328
rect 220136 299288 232544 299316
rect 220136 299276 220142 299288
rect 216646 298704 216674 299276
rect 199896 298472 212534 298500
rect 214576 298676 216674 298704
rect 199896 298460 199902 298472
rect 3510 298392 3516 298444
rect 3568 298432 3574 298444
rect 214576 298432 214604 298676
rect 217152 298636 217180 299276
rect 216646 298608 217180 298636
rect 216646 298500 216674 298608
rect 3568 298404 214604 298432
rect 214668 298472 216674 298500
rect 3568 298392 3574 298404
rect 3602 298324 3608 298376
rect 3660 298364 3666 298376
rect 214668 298364 214696 298472
rect 3660 298336 214696 298364
rect 3660 298324 3666 298336
rect 3418 298256 3424 298308
rect 3476 298296 3482 298308
rect 3476 298268 209774 298296
rect 3476 298256 3482 298268
rect 209746 297616 209774 298268
rect 218072 298160 218100 299276
rect 218164 299112 218192 299276
rect 218164 299084 218652 299112
rect 218624 298772 218652 299084
rect 218716 298976 218744 299276
rect 218808 299044 218836 299276
rect 219912 299248 219940 299276
rect 219912 299220 231854 299248
rect 218808 299016 222194 299044
rect 218716 298948 220814 298976
rect 220786 298840 220814 298948
rect 220786 298812 222056 298840
rect 218624 298744 220814 298772
rect 220786 298568 220814 298744
rect 222028 298636 222056 298812
rect 222166 298772 222194 299016
rect 222166 298744 223436 298772
rect 222166 298676 223252 298704
rect 222166 298636 222194 298676
rect 222028 298608 222194 298636
rect 220786 298540 222194 298568
rect 222166 298296 222194 298540
rect 223224 298432 223252 298676
rect 223408 298500 223436 298744
rect 223546 298540 224954 298568
rect 223546 298500 223574 298540
rect 223408 298472 223574 298500
rect 224926 298500 224954 298540
rect 224926 298472 226334 298500
rect 223224 298404 225828 298432
rect 222166 298268 222884 298296
rect 222856 298228 222884 298268
rect 222856 298200 223344 298228
rect 217888 298132 218100 298160
rect 217888 297616 217916 298132
rect 223316 298092 223344 298200
rect 223316 298064 223574 298092
rect 223546 298024 223574 298064
rect 225800 298024 225828 298404
rect 226306 298364 226334 298472
rect 231826 298364 231854 299220
rect 232516 298432 232544 299288
rect 234586 299288 237196 299316
rect 234586 298432 234614 299288
rect 237190 299276 237196 299288
rect 237248 299276 237254 299328
rect 242158 299316 242164 299328
rect 237346 299288 242164 299316
rect 232516 298404 234614 298432
rect 237346 298364 237374 299288
rect 242158 299276 242164 299288
rect 242216 299276 242222 299328
rect 242268 299248 242296 299356
rect 242342 299276 242348 299328
rect 242400 299276 242406 299328
rect 226306 298336 227714 298364
rect 227686 298296 227714 298336
rect 229066 298336 230474 298364
rect 231826 298336 237374 298364
rect 242084 299220 242296 299248
rect 242084 298364 242112 299220
rect 242360 298704 242388 299276
rect 244246 298772 244274 299424
rect 284588 299356 289814 299384
rect 283558 299316 283564 299328
rect 263566 299288 283564 299316
rect 263566 299112 263594 299288
rect 283558 299276 283564 299288
rect 283616 299276 283622 299328
rect 284478 299276 284484 299328
rect 284536 299276 284542 299328
rect 253906 299084 260834 299112
rect 253906 298772 253934 299084
rect 260806 299044 260834 299084
rect 262186 299084 263594 299112
rect 269086 299152 270494 299180
rect 262186 299044 262214 299084
rect 244246 298744 253934 298772
rect 258046 299016 259454 299044
rect 260806 299016 262214 299044
rect 258046 298704 258074 299016
rect 259426 298772 259454 299016
rect 263566 298948 266354 298976
rect 259426 298744 260834 298772
rect 242360 298676 258074 298704
rect 260806 298636 260834 298744
rect 263566 298704 263594 298948
rect 266326 298908 266354 298948
rect 269086 298908 269114 299152
rect 270466 298976 270494 299152
rect 274606 299084 276014 299112
rect 270466 298948 271874 298976
rect 266326 298880 269114 298908
rect 271846 298908 271874 298948
rect 274606 298908 274634 299084
rect 275986 299044 276014 299084
rect 284496 299044 284524 299276
rect 275986 299016 284524 299044
rect 284588 298908 284616 299356
rect 286502 299276 286508 299328
rect 286560 299276 286566 299328
rect 271846 298880 274634 298908
rect 280126 298880 284616 298908
rect 267706 298812 269114 298840
rect 267706 298772 267734 298812
rect 262186 298676 263594 298704
rect 266326 298744 267734 298772
rect 269086 298772 269114 298812
rect 270466 298812 271874 298840
rect 270466 298772 270494 298812
rect 269086 298744 270494 298772
rect 262186 298636 262214 298676
rect 258046 298608 259454 298636
rect 260806 298608 262214 298636
rect 247006 298404 247172 298432
rect 247006 298364 247034 298404
rect 242084 298336 247034 298364
rect 247144 298364 247172 298404
rect 258046 298364 258074 298608
rect 259426 298568 259454 298608
rect 259426 298540 262214 298568
rect 262186 298500 262214 298540
rect 263566 298540 264974 298568
rect 263566 298500 263594 298540
rect 262186 298472 263594 298500
rect 264946 298500 264974 298540
rect 266326 298500 266354 298744
rect 271846 298636 271874 298812
rect 273226 298676 274634 298704
rect 273226 298636 273254 298676
rect 271846 298608 273254 298636
rect 274606 298568 274634 298676
rect 280126 298636 280154 298880
rect 275986 298608 280154 298636
rect 275986 298568 276014 298608
rect 274606 298540 276014 298568
rect 264946 298472 266354 298500
rect 247144 298336 258074 298364
rect 229066 298296 229094 298336
rect 227686 298268 229094 298296
rect 230446 298296 230474 298336
rect 286520 298296 286548 299276
rect 230446 298268 286548 298296
rect 289786 298296 289814 299356
rect 299842 299276 299848 299328
rect 299900 299316 299906 299328
rect 300118 299316 300124 299328
rect 299900 299288 300124 299316
rect 299900 299276 299906 299288
rect 300118 299276 300124 299288
rect 300176 299276 300182 299328
rect 434714 299072 434720 299124
rect 434772 299112 434778 299124
rect 441706 299112 441712 299124
rect 434772 299084 441712 299112
rect 434772 299072 434778 299084
rect 441706 299072 441712 299084
rect 441764 299072 441770 299124
rect 318058 298500 318064 298512
rect 292546 298472 318064 298500
rect 292546 298296 292574 298472
rect 318058 298460 318064 298472
rect 318116 298460 318122 298512
rect 289786 298268 292574 298296
rect 302786 298256 302792 298308
rect 302844 298296 302850 298308
rect 322198 298296 322204 298308
rect 302844 298268 322204 298296
rect 302844 298256 302850 298268
rect 322198 298256 322204 298268
rect 322256 298256 322262 298308
rect 580166 298228 580172 298240
rect 226306 298200 229094 298228
rect 226306 298024 226334 298200
rect 229066 298160 229094 298200
rect 230446 298200 231854 298228
rect 230446 298160 230474 298200
rect 229066 298132 230474 298160
rect 231826 298092 231854 298200
rect 235966 298200 580172 298228
rect 235966 298092 235994 298200
rect 580166 298188 580172 298200
rect 580224 298188 580230 298240
rect 580258 298160 580264 298172
rect 231826 298064 235994 298092
rect 237346 298132 252554 298160
rect 223546 297996 224954 298024
rect 225800 297996 226334 298024
rect 209746 297588 217916 297616
rect 224926 297616 224954 297996
rect 237346 297684 237374 298132
rect 252526 298092 252554 298132
rect 275986 298132 580264 298160
rect 275986 298092 276014 298132
rect 580258 298120 580264 298132
rect 580316 298120 580322 298172
rect 252526 298064 276014 298092
rect 371234 298052 371240 298104
rect 371292 298092 371298 298104
rect 381078 298092 381084 298104
rect 371292 298064 381084 298092
rect 371292 298052 371298 298064
rect 381078 298052 381084 298064
rect 381136 298052 381142 298104
rect 229066 297656 237374 297684
rect 229066 297616 229094 297656
rect 224926 297588 229094 297616
rect 436094 297576 436100 297628
rect 436152 297616 436158 297628
rect 441798 297616 441804 297628
rect 436152 297588 441804 297616
rect 436152 297576 436158 297588
rect 441798 297576 441804 297588
rect 441856 297576 441862 297628
rect 381078 297440 381084 297492
rect 381136 297480 381142 297492
rect 382366 297480 382372 297492
rect 381136 297452 382372 297480
rect 381136 297440 381142 297452
rect 382366 297440 382372 297452
rect 382424 297440 382430 297492
rect 371234 297372 371240 297424
rect 371292 297412 371298 297424
rect 379514 297412 379520 297424
rect 371292 297384 379520 297412
rect 371292 297372 371298 297384
rect 379514 297372 379520 297384
rect 379572 297372 379578 297424
rect 445662 296964 445668 297016
rect 445720 297004 445726 297016
rect 447778 297004 447784 297016
rect 445720 296976 447784 297004
rect 445720 296964 445726 296976
rect 447778 296964 447784 296976
rect 447836 296964 447842 297016
rect 447778 296828 447784 296880
rect 447836 296868 447842 296880
rect 452838 296868 452844 296880
rect 447836 296840 452844 296868
rect 447836 296828 447842 296840
rect 452838 296828 452844 296840
rect 452896 296828 452902 296880
rect 303062 296760 303068 296812
rect 303120 296800 303126 296812
rect 369394 296800 369400 296812
rect 303120 296772 369400 296800
rect 303120 296760 303126 296772
rect 369394 296760 369400 296772
rect 369452 296760 369458 296812
rect 302878 296692 302884 296744
rect 302936 296732 302942 296744
rect 369302 296732 369308 296744
rect 302936 296704 369308 296732
rect 302936 296692 302942 296704
rect 369302 296692 369308 296704
rect 369360 296692 369366 296744
rect 371234 296624 371240 296676
rect 371292 296664 371298 296676
rect 376754 296664 376760 296676
rect 371292 296636 376760 296664
rect 371292 296624 371298 296636
rect 376754 296624 376760 296636
rect 376812 296624 376818 296676
rect 445662 295944 445668 295996
rect 445720 295984 445726 295996
rect 452654 295984 452660 295996
rect 445720 295956 452660 295984
rect 445720 295944 445726 295956
rect 452654 295944 452660 295956
rect 452712 295944 452718 295996
rect 324958 295876 324964 295928
rect 325016 295916 325022 295928
rect 371234 295916 371240 295928
rect 325016 295888 371240 295916
rect 325016 295876 325022 295888
rect 371234 295876 371240 295888
rect 371292 295876 371298 295928
rect 352558 295808 352564 295860
rect 352616 295848 352622 295860
rect 369302 295848 369308 295860
rect 352616 295820 369308 295848
rect 352616 295808 352622 295820
rect 369302 295808 369308 295820
rect 369360 295808 369366 295860
rect 371234 295536 371240 295588
rect 371292 295576 371298 295588
rect 373350 295576 373356 295588
rect 371292 295548 373356 295576
rect 371292 295536 371298 295548
rect 373350 295536 373356 295548
rect 373408 295576 373414 295588
rect 373994 295576 374000 295588
rect 373408 295548 374000 295576
rect 373408 295536 373414 295548
rect 373994 295536 374000 295548
rect 374052 295536 374058 295588
rect 376754 295400 376760 295452
rect 376812 295440 376818 295452
rect 380894 295440 380900 295452
rect 376812 295412 380900 295440
rect 376812 295400 376818 295412
rect 380894 295400 380900 295412
rect 380952 295400 380958 295452
rect 370222 295332 370228 295384
rect 370280 295372 370286 295384
rect 377398 295372 377404 295384
rect 370280 295344 377404 295372
rect 370280 295332 370286 295344
rect 377398 295332 377404 295344
rect 377456 295372 377462 295384
rect 380986 295372 380992 295384
rect 377456 295344 380992 295372
rect 377456 295332 377462 295344
rect 380986 295332 380992 295344
rect 381044 295332 381050 295384
rect 452654 295332 452660 295384
rect 452712 295372 452718 295384
rect 454126 295372 454132 295384
rect 452712 295344 454132 295372
rect 452712 295332 452718 295344
rect 454126 295332 454132 295344
rect 454184 295332 454190 295384
rect 370130 295196 370136 295248
rect 370188 295236 370194 295248
rect 378226 295236 378232 295248
rect 370188 295208 378232 295236
rect 370188 295196 370194 295208
rect 378226 295196 378232 295208
rect 378284 295196 378290 295248
rect 445662 295196 445668 295248
rect 445720 295236 445726 295248
rect 448606 295236 448612 295248
rect 445720 295208 448612 295236
rect 445720 295196 445726 295208
rect 448606 295196 448612 295208
rect 448664 295196 448670 295248
rect 378226 294720 378232 294772
rect 378284 294760 378290 294772
rect 381078 294760 381084 294772
rect 378284 294732 381084 294760
rect 378284 294720 378290 294732
rect 381078 294720 381084 294732
rect 381136 294720 381142 294772
rect 372338 294584 372344 294636
rect 372396 294624 372402 294636
rect 372614 294624 372620 294636
rect 372396 294596 372620 294624
rect 372396 294584 372402 294596
rect 372614 294584 372620 294596
rect 372672 294624 372678 294636
rect 378226 294624 378232 294636
rect 372672 294596 378232 294624
rect 372672 294584 372678 294596
rect 378226 294584 378232 294596
rect 378284 294584 378290 294636
rect 448606 294040 448612 294092
rect 448664 294080 448670 294092
rect 452654 294080 452660 294092
rect 448664 294052 452660 294080
rect 448664 294040 448670 294052
rect 452654 294040 452660 294052
rect 452712 294040 452718 294092
rect 180058 293972 180064 294024
rect 180116 294012 180122 294024
rect 197906 294012 197912 294024
rect 180116 293984 197912 294012
rect 180116 293972 180122 293984
rect 197906 293972 197912 293984
rect 197964 293972 197970 294024
rect 302418 293972 302424 294024
rect 302476 294012 302482 294024
rect 320818 294012 320824 294024
rect 302476 293984 320824 294012
rect 302476 293972 302482 293984
rect 320818 293972 320824 293984
rect 320876 293972 320882 294024
rect 371234 293972 371240 294024
rect 371292 294012 371298 294024
rect 375374 294012 375380 294024
rect 371292 293984 375380 294012
rect 371292 293972 371298 293984
rect 375374 293972 375380 293984
rect 375432 293972 375438 294024
rect 445754 293972 445760 294024
rect 445812 294012 445818 294024
rect 450262 294012 450268 294024
rect 445812 293984 450268 294012
rect 445812 293972 445818 293984
rect 450262 293972 450268 293984
rect 450320 293972 450326 294024
rect 2866 293904 2872 293956
rect 2924 293944 2930 293956
rect 196618 293944 196624 293956
rect 2924 293916 196624 293944
rect 2924 293904 2930 293916
rect 196618 293904 196624 293916
rect 196676 293904 196682 293956
rect 371234 293224 371240 293276
rect 371292 293264 371298 293276
rect 378318 293264 378324 293276
rect 371292 293236 378324 293264
rect 371292 293224 371298 293236
rect 378318 293224 378324 293236
rect 378376 293224 378382 293276
rect 371234 292884 371240 292936
rect 371292 292924 371298 292936
rect 374454 292924 374460 292936
rect 371292 292896 374460 292924
rect 371292 292884 371298 292896
rect 374454 292884 374460 292896
rect 374512 292924 374518 292936
rect 374914 292924 374920 292936
rect 374512 292896 374920 292924
rect 374512 292884 374518 292896
rect 374914 292884 374920 292896
rect 374972 292884 374978 292936
rect 445662 292884 445668 292936
rect 445720 292924 445726 292936
rect 446490 292924 446496 292936
rect 445720 292896 446496 292924
rect 445720 292884 445726 292896
rect 446490 292884 446496 292896
rect 446548 292924 446554 292936
rect 449986 292924 449992 292936
rect 446548 292896 449992 292924
rect 446548 292884 446554 292896
rect 449986 292884 449992 292896
rect 450044 292884 450050 292936
rect 378318 292544 378324 292596
rect 378376 292584 378382 292596
rect 378502 292584 378508 292596
rect 378376 292556 378508 292584
rect 378376 292544 378382 292556
rect 378502 292544 378508 292556
rect 378560 292544 378566 292596
rect 371234 291864 371240 291916
rect 371292 291904 371298 291916
rect 375742 291904 375748 291916
rect 371292 291876 375748 291904
rect 371292 291864 371298 291876
rect 375742 291864 375748 291876
rect 375800 291904 375806 291916
rect 378318 291904 378324 291916
rect 375800 291876 378324 291904
rect 375800 291864 375806 291876
rect 378318 291864 378324 291876
rect 378376 291864 378382 291916
rect 195238 291796 195244 291848
rect 195296 291836 195302 291848
rect 198090 291836 198096 291848
rect 195296 291808 198096 291836
rect 195296 291796 195302 291808
rect 198090 291796 198096 291808
rect 198148 291796 198154 291848
rect 372338 291796 372344 291848
rect 372396 291836 372402 291848
rect 373258 291836 373264 291848
rect 372396 291808 373264 291836
rect 372396 291796 372402 291808
rect 373258 291796 373264 291808
rect 373316 291836 373322 291848
rect 378410 291836 378416 291848
rect 373316 291808 378416 291836
rect 373316 291796 373322 291808
rect 378410 291796 378416 291808
rect 378468 291796 378474 291848
rect 302326 291184 302332 291236
rect 302384 291224 302390 291236
rect 359458 291224 359464 291236
rect 302384 291196 359464 291224
rect 302384 291184 302390 291196
rect 359458 291184 359464 291196
rect 359516 291184 359522 291236
rect 371234 291184 371240 291236
rect 371292 291224 371298 291236
rect 376018 291224 376024 291236
rect 371292 291196 376024 291224
rect 371292 291184 371298 291196
rect 376018 291184 376024 291196
rect 376076 291224 376082 291236
rect 377030 291224 377036 291236
rect 376076 291196 377036 291224
rect 376076 291184 376082 291196
rect 377030 291184 377036 291196
rect 377088 291184 377094 291236
rect 445662 291184 445668 291236
rect 445720 291224 445726 291236
rect 447410 291224 447416 291236
rect 445720 291196 447416 291224
rect 445720 291184 445726 291196
rect 447410 291184 447416 291196
rect 447468 291224 447474 291236
rect 451274 291224 451280 291236
rect 447468 291196 451280 291224
rect 447468 291184 447474 291196
rect 451274 291184 451280 291196
rect 451332 291184 451338 291236
rect 448606 291116 448612 291168
rect 448664 291156 448670 291168
rect 450078 291156 450084 291168
rect 448664 291128 450084 291156
rect 448664 291116 448670 291128
rect 450078 291116 450084 291128
rect 450136 291116 450142 291168
rect 445662 290572 445668 290624
rect 445720 290612 445726 290624
rect 448606 290612 448612 290624
rect 445720 290584 448612 290612
rect 445720 290572 445726 290584
rect 448606 290572 448612 290584
rect 448664 290572 448670 290624
rect 372338 290504 372344 290556
rect 372396 290544 372402 290556
rect 372798 290544 372804 290556
rect 372396 290516 372804 290544
rect 372396 290504 372402 290516
rect 372798 290504 372804 290516
rect 372856 290544 372862 290556
rect 376754 290544 376760 290556
rect 372856 290516 376760 290544
rect 372856 290504 372862 290516
rect 376754 290504 376760 290516
rect 376812 290504 376818 290556
rect 371234 290436 371240 290488
rect 371292 290476 371298 290488
rect 376846 290476 376852 290488
rect 371292 290448 376852 290476
rect 371292 290436 371298 290448
rect 376846 290436 376852 290448
rect 376904 290436 376910 290488
rect 184198 289824 184204 289876
rect 184256 289864 184262 289876
rect 197354 289864 197360 289876
rect 184256 289836 197360 289864
rect 184256 289824 184262 289836
rect 197354 289824 197360 289836
rect 197412 289824 197418 289876
rect 445662 289416 445668 289468
rect 445720 289456 445726 289468
rect 445846 289456 445852 289468
rect 445720 289428 445852 289456
rect 445720 289416 445726 289428
rect 445846 289416 445852 289428
rect 445904 289456 445910 289468
rect 450078 289456 450084 289468
rect 445904 289428 450084 289456
rect 445904 289416 445910 289428
rect 450078 289416 450084 289428
rect 450136 289416 450142 289468
rect 371234 289008 371240 289060
rect 371292 289048 371298 289060
rect 374270 289048 374276 289060
rect 371292 289020 374276 289048
rect 371292 289008 371298 289020
rect 374270 289008 374276 289020
rect 374328 289048 374334 289060
rect 375742 289048 375748 289060
rect 374328 289020 375748 289048
rect 374328 289008 374334 289020
rect 375742 289008 375748 289020
rect 375800 289008 375806 289060
rect 372338 288940 372344 288992
rect 372396 288980 372402 288992
rect 374730 288980 374736 288992
rect 372396 288952 374736 288980
rect 372396 288940 372402 288952
rect 374730 288940 374736 288952
rect 374788 288980 374794 288992
rect 375466 288980 375472 288992
rect 374788 288952 375472 288980
rect 374788 288940 374794 288952
rect 375466 288940 375472 288952
rect 375524 288940 375530 288992
rect 372798 288532 372804 288584
rect 372856 288572 372862 288584
rect 375558 288572 375564 288584
rect 372856 288544 375564 288572
rect 372856 288532 372862 288544
rect 375558 288532 375564 288544
rect 375616 288532 375622 288584
rect 371234 288328 371240 288380
rect 371292 288368 371298 288380
rect 377122 288368 377128 288380
rect 371292 288340 377128 288368
rect 371292 288328 371298 288340
rect 377122 288328 377128 288340
rect 377180 288368 377186 288380
rect 383654 288368 383660 288380
rect 377180 288340 383660 288368
rect 377180 288328 377186 288340
rect 383654 288328 383660 288340
rect 383712 288328 383718 288380
rect 445662 288328 445668 288380
rect 445720 288368 445726 288380
rect 447870 288368 447876 288380
rect 445720 288340 447876 288368
rect 445720 288328 445726 288340
rect 447870 288328 447876 288340
rect 447928 288368 447934 288380
rect 449894 288368 449900 288380
rect 447928 288340 449900 288368
rect 447928 288328 447934 288340
rect 449894 288328 449900 288340
rect 449952 288328 449958 288380
rect 445110 288056 445116 288108
rect 445168 288096 445174 288108
rect 447226 288096 447232 288108
rect 445168 288068 447232 288096
rect 445168 288056 445174 288068
rect 447226 288056 447232 288068
rect 447284 288096 447290 288108
rect 448514 288096 448520 288108
rect 447284 288068 448520 288096
rect 447284 288056 447290 288068
rect 448514 288056 448520 288068
rect 448572 288056 448578 288108
rect 160094 287036 160100 287088
rect 160152 287076 160158 287088
rect 197630 287076 197636 287088
rect 160152 287048 197636 287076
rect 160152 287036 160158 287048
rect 197630 287036 197636 287048
rect 197688 287036 197694 287088
rect 372338 287036 372344 287088
rect 372396 287076 372402 287088
rect 382642 287076 382648 287088
rect 372396 287048 382648 287076
rect 372396 287036 372402 287048
rect 382642 287036 382648 287048
rect 382700 287076 382706 287088
rect 383562 287076 383568 287088
rect 382700 287048 383568 287076
rect 382700 287036 382706 287048
rect 383562 287036 383568 287048
rect 383620 287036 383626 287088
rect 371878 286560 371884 286612
rect 371936 286600 371942 286612
rect 372338 286600 372344 286612
rect 371936 286572 372344 286600
rect 371936 286560 371942 286572
rect 372338 286560 372344 286572
rect 372396 286560 372402 286612
rect 371326 286424 371332 286476
rect 371384 286464 371390 286476
rect 375650 286464 375656 286476
rect 371384 286436 375656 286464
rect 371384 286424 371390 286436
rect 375650 286424 375656 286436
rect 375708 286424 375714 286476
rect 371878 286356 371884 286408
rect 371936 286396 371942 286408
rect 376110 286396 376116 286408
rect 371936 286368 376116 286396
rect 371936 286356 371942 286368
rect 376110 286356 376116 286368
rect 376168 286396 376174 286408
rect 382458 286396 382464 286408
rect 376168 286368 382464 286396
rect 376168 286356 376174 286368
rect 382458 286356 382464 286368
rect 382516 286356 382522 286408
rect 372522 286288 372528 286340
rect 372580 286328 372586 286340
rect 379606 286328 379612 286340
rect 372580 286300 379612 286328
rect 372580 286288 372586 286300
rect 379606 286288 379612 286300
rect 379664 286288 379670 286340
rect 188338 285676 188344 285728
rect 188396 285716 188402 285728
rect 197354 285716 197360 285728
rect 188396 285688 197360 285716
rect 188396 285676 188402 285688
rect 197354 285676 197360 285688
rect 197412 285676 197418 285728
rect 302786 285676 302792 285728
rect 302844 285716 302850 285728
rect 353938 285716 353944 285728
rect 302844 285688 353944 285716
rect 302844 285676 302850 285688
rect 353938 285676 353944 285688
rect 353996 285676 354002 285728
rect 375650 285676 375656 285728
rect 375708 285716 375714 285728
rect 380894 285716 380900 285728
rect 375708 285688 380900 285716
rect 375708 285676 375714 285688
rect 380894 285676 380900 285688
rect 380952 285676 380958 285728
rect 445662 285676 445668 285728
rect 445720 285716 445726 285728
rect 448882 285716 448888 285728
rect 445720 285688 448888 285716
rect 445720 285676 445726 285688
rect 448882 285676 448888 285688
rect 448940 285716 448946 285728
rect 449894 285716 449900 285728
rect 448940 285688 449900 285716
rect 448940 285676 448946 285688
rect 449894 285676 449900 285688
rect 449952 285676 449958 285728
rect 371878 285608 371884 285660
rect 371936 285648 371942 285660
rect 381170 285648 381176 285660
rect 371936 285620 381176 285648
rect 371936 285608 371942 285620
rect 381170 285608 381176 285620
rect 381228 285608 381234 285660
rect 371878 285064 371884 285116
rect 371936 285104 371942 285116
rect 374638 285104 374644 285116
rect 371936 285076 374644 285104
rect 371936 285064 371942 285076
rect 374638 285064 374644 285076
rect 374696 285104 374702 285116
rect 378134 285104 378140 285116
rect 374696 285076 378140 285104
rect 374696 285064 374702 285076
rect 378134 285064 378140 285076
rect 378192 285064 378198 285116
rect 445662 284860 445668 284912
rect 445720 284900 445726 284912
rect 446674 284900 446680 284912
rect 445720 284872 446680 284900
rect 445720 284860 445726 284872
rect 446674 284860 446680 284872
rect 446732 284900 446738 284912
rect 448698 284900 448704 284912
rect 446732 284872 448704 284900
rect 446732 284860 446738 284872
rect 448698 284860 448704 284872
rect 448756 284860 448762 284912
rect 381170 284384 381176 284436
rect 381228 284424 381234 284436
rect 382550 284424 382556 284436
rect 381228 284396 382556 284424
rect 381228 284384 381234 284396
rect 382550 284384 382556 284396
rect 382608 284384 382614 284436
rect 371878 284316 371884 284368
rect 371936 284356 371942 284368
rect 378134 284356 378140 284368
rect 371936 284328 378140 284356
rect 371936 284316 371942 284328
rect 378134 284316 378140 284328
rect 378192 284356 378198 284368
rect 382274 284356 382280 284368
rect 378192 284328 382280 284356
rect 378192 284316 378198 284328
rect 382274 284316 382280 284328
rect 382332 284316 382338 284368
rect 445478 283636 445484 283688
rect 445536 283676 445542 283688
rect 446030 283676 446036 283688
rect 445536 283648 446036 283676
rect 445536 283636 445542 283648
rect 446030 283636 446036 283648
rect 446088 283636 446094 283688
rect 371878 283568 371884 283620
rect 371936 283608 371942 283620
rect 376938 283608 376944 283620
rect 371936 283580 376944 283608
rect 371936 283568 371942 283580
rect 376938 283568 376944 283580
rect 376996 283608 377002 283620
rect 377214 283608 377220 283620
rect 376996 283580 377220 283608
rect 376996 283568 377002 283580
rect 377214 283568 377220 283580
rect 377272 283568 377278 283620
rect 371878 283160 371884 283212
rect 371936 283200 371942 283212
rect 372890 283200 372896 283212
rect 371936 283172 372896 283200
rect 371936 283160 371942 283172
rect 372890 283160 372896 283172
rect 372948 283200 372954 283212
rect 375466 283200 375472 283212
rect 372948 283172 375472 283200
rect 372948 283160 372954 283172
rect 375466 283160 375472 283172
rect 375524 283160 375530 283212
rect 184290 282888 184296 282940
rect 184348 282928 184354 282940
rect 197354 282928 197360 282940
rect 184348 282900 197360 282928
rect 184348 282888 184354 282900
rect 197354 282888 197360 282900
rect 197412 282888 197418 282940
rect 446030 282888 446036 282940
rect 446088 282928 446094 282940
rect 448698 282928 448704 282940
rect 446088 282900 448704 282928
rect 446088 282888 446094 282900
rect 448698 282888 448704 282900
rect 448756 282888 448762 282940
rect 371878 282684 371884 282736
rect 371936 282724 371942 282736
rect 374178 282724 374184 282736
rect 371936 282696 374184 282724
rect 371936 282684 371942 282696
rect 374178 282684 374184 282696
rect 374236 282724 374242 282736
rect 374546 282724 374552 282736
rect 374236 282696 374552 282724
rect 374236 282684 374242 282696
rect 374546 282684 374552 282696
rect 374604 282684 374610 282736
rect 445386 282480 445392 282532
rect 445444 282520 445450 282532
rect 447226 282520 447232 282532
rect 445444 282492 447232 282520
rect 445444 282480 445450 282492
rect 447226 282480 447232 282492
rect 447284 282480 447290 282532
rect 371878 282140 371884 282192
rect 371936 282180 371942 282192
rect 374086 282180 374092 282192
rect 371936 282152 374092 282180
rect 371936 282140 371942 282152
rect 374086 282140 374092 282152
rect 374144 282180 374150 282192
rect 374270 282180 374276 282192
rect 374144 282152 374276 282180
rect 374144 282140 374150 282152
rect 374270 282140 374276 282152
rect 374328 282140 374334 282192
rect 302418 281528 302424 281580
rect 302476 281568 302482 281580
rect 356698 281568 356704 281580
rect 302476 281540 356704 281568
rect 302476 281528 302482 281540
rect 356698 281528 356704 281540
rect 356756 281528 356762 281580
rect 445110 281460 445116 281512
rect 445168 281500 445174 281512
rect 446582 281500 446588 281512
rect 445168 281472 446588 281500
rect 445168 281460 445174 281472
rect 446582 281460 446588 281472
rect 446640 281500 446646 281512
rect 447134 281500 447140 281512
rect 446640 281472 447140 281500
rect 446640 281460 446646 281472
rect 447134 281460 447140 281472
rect 447192 281460 447198 281512
rect 444742 280576 444748 280628
rect 444800 280616 444806 280628
rect 445938 280616 445944 280628
rect 444800 280588 445944 280616
rect 444800 280576 444806 280588
rect 445938 280576 445944 280588
rect 445996 280616 446002 280628
rect 447134 280616 447140 280628
rect 445996 280588 447140 280616
rect 445996 280576 446002 280588
rect 447134 280576 447140 280588
rect 447192 280576 447198 280628
rect 186958 280168 186964 280220
rect 187016 280208 187022 280220
rect 197354 280208 197360 280220
rect 187016 280180 197360 280208
rect 187016 280168 187022 280180
rect 197354 280168 197360 280180
rect 197412 280168 197418 280220
rect 358078 280100 358084 280152
rect 358136 280140 358142 280152
rect 360194 280140 360200 280152
rect 358136 280112 360200 280140
rect 358136 280100 358142 280112
rect 360194 280100 360200 280112
rect 360252 280100 360258 280152
rect 444558 280032 444564 280084
rect 444616 280072 444622 280084
rect 444834 280072 444840 280084
rect 444616 280044 444840 280072
rect 444616 280032 444622 280044
rect 444834 280032 444840 280044
rect 444892 280032 444898 280084
rect 193950 278944 193956 278996
rect 194008 278984 194014 278996
rect 197354 278984 197360 278996
rect 194008 278956 197360 278984
rect 194008 278944 194014 278956
rect 197354 278944 197360 278956
rect 197412 278944 197418 278996
rect 302602 278740 302608 278792
rect 302660 278780 302666 278792
rect 358078 278780 358084 278792
rect 302660 278752 358084 278780
rect 302660 278740 302666 278752
rect 358078 278740 358084 278752
rect 358136 278740 358142 278792
rect 372154 278672 372160 278724
rect 372212 278712 372218 278724
rect 372982 278712 372988 278724
rect 372212 278684 372988 278712
rect 372212 278672 372218 278684
rect 372982 278672 372988 278684
rect 373040 278672 373046 278724
rect 444374 278672 444380 278724
rect 444432 278712 444438 278724
rect 445110 278712 445116 278724
rect 444432 278684 445116 278712
rect 444432 278672 444438 278684
rect 445110 278672 445116 278684
rect 445168 278672 445174 278724
rect 372338 277448 372344 277500
rect 372396 277488 372402 277500
rect 374178 277488 374184 277500
rect 372396 277460 374184 277488
rect 372396 277448 372402 277460
rect 374178 277448 374184 277460
rect 374236 277448 374242 277500
rect 369118 277176 369124 277228
rect 369176 277216 369182 277228
rect 369302 277216 369308 277228
rect 369176 277188 369308 277216
rect 369176 277176 369182 277188
rect 369302 277176 369308 277188
rect 369360 277176 369366 277228
rect 371602 276360 371608 276412
rect 371660 276400 371666 276412
rect 372154 276400 372160 276412
rect 371660 276372 372160 276400
rect 371660 276360 371666 276372
rect 372154 276360 372160 276372
rect 372212 276360 372218 276412
rect 182818 276020 182824 276072
rect 182876 276060 182882 276072
rect 197538 276060 197544 276072
rect 182876 276032 197544 276060
rect 182876 276020 182882 276032
rect 197538 276020 197544 276032
rect 197596 276020 197602 276072
rect 371602 276020 371608 276072
rect 371660 276060 371666 276072
rect 373994 276060 374000 276072
rect 371660 276032 374000 276060
rect 371660 276020 371666 276032
rect 373994 276020 374000 276032
rect 374052 276060 374058 276072
rect 374362 276060 374368 276072
rect 374052 276032 374368 276060
rect 374052 276020 374058 276032
rect 374362 276020 374368 276032
rect 374420 276020 374426 276072
rect 196618 274864 196624 274916
rect 196676 274904 196682 274916
rect 198366 274904 198372 274916
rect 196676 274876 198372 274904
rect 196676 274864 196682 274876
rect 198366 274864 198372 274876
rect 198424 274864 198430 274916
rect 445570 274592 445576 274644
rect 445628 274632 445634 274644
rect 449250 274632 449256 274644
rect 445628 274604 449256 274632
rect 445628 274592 445634 274604
rect 449250 274592 449256 274604
rect 449308 274632 449314 274644
rect 452746 274632 452752 274644
rect 449308 274604 452752 274632
rect 449308 274592 449314 274604
rect 452746 274592 452752 274604
rect 452804 274592 452810 274644
rect 445662 273232 445668 273284
rect 445720 273272 445726 273284
rect 450170 273272 450176 273284
rect 445720 273244 450176 273272
rect 445720 273232 445726 273244
rect 450170 273232 450176 273244
rect 450228 273272 450234 273284
rect 452930 273272 452936 273284
rect 450228 273244 452936 273272
rect 450228 273232 450234 273244
rect 452930 273232 452936 273244
rect 452988 273232 452994 273284
rect 371050 273164 371056 273216
rect 371108 273204 371114 273216
rect 374362 273204 374368 273216
rect 371108 273176 374368 273204
rect 371108 273164 371114 273176
rect 374362 273164 374368 273176
rect 374420 273164 374426 273216
rect 445662 272484 445668 272536
rect 445720 272524 445726 272536
rect 454034 272524 454040 272536
rect 445720 272496 454040 272524
rect 445720 272484 445726 272496
rect 454034 272484 454040 272496
rect 454092 272484 454098 272536
rect 181438 271872 181444 271924
rect 181496 271912 181502 271924
rect 197354 271912 197360 271924
rect 181496 271884 197360 271912
rect 181496 271872 181502 271884
rect 197354 271872 197360 271884
rect 197412 271872 197418 271924
rect 371510 271464 371516 271516
rect 371568 271464 371574 271516
rect 371528 271176 371556 271464
rect 371510 271124 371516 271176
rect 371568 271124 371574 271176
rect 371786 271124 371792 271176
rect 371844 271164 371850 271176
rect 371970 271164 371976 271176
rect 371844 271136 371976 271164
rect 371844 271124 371850 271136
rect 371970 271124 371976 271136
rect 372028 271124 372034 271176
rect 358078 271056 358084 271108
rect 358136 271096 358142 271108
rect 360654 271096 360660 271108
rect 358136 271068 360660 271096
rect 358136 271056 358142 271068
rect 360654 271056 360660 271068
rect 360712 271056 360718 271108
rect 445662 270580 445668 270632
rect 445720 270620 445726 270632
rect 451366 270620 451372 270632
rect 445720 270592 451372 270620
rect 445720 270580 445726 270592
rect 451366 270580 451372 270592
rect 451424 270580 451430 270632
rect 178770 270512 178776 270564
rect 178828 270552 178834 270564
rect 197354 270552 197360 270564
rect 178828 270524 197360 270552
rect 178828 270512 178834 270524
rect 197354 270512 197360 270524
rect 197412 270512 197418 270564
rect 302326 270444 302332 270496
rect 302384 270484 302390 270496
rect 352558 270484 352564 270496
rect 302384 270456 352564 270484
rect 302384 270444 302390 270456
rect 352558 270444 352564 270456
rect 352616 270444 352622 270496
rect 445662 269084 445668 269136
rect 445720 269124 445726 269136
rect 448790 269124 448796 269136
rect 445720 269096 448796 269124
rect 445720 269084 445726 269096
rect 448790 269084 448796 269096
rect 448848 269124 448854 269136
rect 452838 269124 452844 269136
rect 448848 269096 452844 269124
rect 448848 269084 448854 269096
rect 452838 269084 452844 269096
rect 452896 269084 452902 269136
rect 372154 268336 372160 268388
rect 372212 268376 372218 268388
rect 372890 268376 372896 268388
rect 372212 268348 372896 268376
rect 372212 268336 372218 268348
rect 372890 268336 372896 268348
rect 372948 268336 372954 268388
rect 175918 267724 175924 267776
rect 175976 267764 175982 267776
rect 197722 267764 197728 267776
rect 175976 267736 197728 267764
rect 175976 267724 175982 267736
rect 197722 267724 197728 267736
rect 197780 267724 197786 267776
rect 3234 267656 3240 267708
rect 3292 267696 3298 267708
rect 17218 267696 17224 267708
rect 3292 267668 17224 267696
rect 3292 267656 3298 267668
rect 17218 267656 17224 267668
rect 17276 267656 17282 267708
rect 302418 267656 302424 267708
rect 302476 267696 302482 267708
rect 324958 267696 324964 267708
rect 302476 267668 324964 267696
rect 302476 267656 302482 267668
rect 324958 267656 324964 267668
rect 325016 267656 325022 267708
rect 302510 266976 302516 267028
rect 302568 267016 302574 267028
rect 370222 267016 370228 267028
rect 302568 266988 370228 267016
rect 302568 266976 302574 266988
rect 370222 266976 370228 266988
rect 370280 266976 370286 267028
rect 362862 266296 362868 266348
rect 362920 266336 362926 266348
rect 435174 266336 435180 266348
rect 362920 266308 435180 266336
rect 362920 266296 362926 266308
rect 435174 266296 435180 266308
rect 435232 266336 435238 266348
rect 436002 266336 436008 266348
rect 435232 266308 436008 266336
rect 435232 266296 435238 266308
rect 436002 266296 436008 266308
rect 436060 266336 436066 266348
rect 441706 266336 441712 266348
rect 436060 266308 441712 266336
rect 436060 266296 436066 266308
rect 441706 266296 441712 266308
rect 441764 266296 441770 266348
rect 364886 266228 364892 266280
rect 364944 266268 364950 266280
rect 437382 266268 437388 266280
rect 364944 266240 437388 266268
rect 364944 266228 364950 266240
rect 437382 266228 437388 266240
rect 437440 266268 437446 266280
rect 441798 266268 441804 266280
rect 437440 266240 441804 266268
rect 437440 266228 437446 266240
rect 441798 266228 441804 266240
rect 441856 266228 441862 266280
rect 302970 266160 302976 266212
rect 303028 266200 303034 266212
rect 368934 266200 368940 266212
rect 303028 266172 368940 266200
rect 303028 266160 303034 266172
rect 368934 266160 368940 266172
rect 368992 266200 368998 266212
rect 369118 266200 369124 266212
rect 368992 266172 369124 266200
rect 368992 266160 368998 266172
rect 369118 266160 369124 266172
rect 369176 266200 369182 266212
rect 441338 266200 441344 266212
rect 369176 266172 441344 266200
rect 369176 266160 369182 266172
rect 441338 266160 441344 266172
rect 441396 266200 441402 266212
rect 441522 266200 441528 266212
rect 441396 266172 441528 266200
rect 441396 266160 441402 266172
rect 441522 266160 441528 266172
rect 441580 266160 441586 266212
rect 300118 266092 300124 266144
rect 300176 266132 300182 266144
rect 366910 266132 366916 266144
rect 300176 266104 366916 266132
rect 300176 266092 300182 266104
rect 366910 266092 366916 266104
rect 366968 266092 366974 266144
rect 360930 265684 360936 265736
rect 360988 265724 360994 265736
rect 431954 265724 431960 265736
rect 360988 265696 431960 265724
rect 360988 265684 360994 265696
rect 431954 265684 431960 265696
rect 432012 265724 432018 265736
rect 432598 265724 432604 265736
rect 432012 265696 432604 265724
rect 432012 265684 432018 265696
rect 432598 265684 432604 265696
rect 432656 265684 432662 265736
rect 300026 265616 300032 265668
rect 300084 265656 300090 265668
rect 438854 265656 438860 265668
rect 300084 265628 438860 265656
rect 300084 265616 300090 265628
rect 438854 265616 438860 265628
rect 438912 265616 438918 265668
rect 174538 264936 174544 264988
rect 174596 264976 174602 264988
rect 197354 264976 197360 264988
rect 174596 264948 197360 264976
rect 174596 264936 174602 264948
rect 197354 264936 197360 264948
rect 197412 264936 197418 264988
rect 360194 264936 360200 264988
rect 360252 264976 360258 264988
rect 360930 264976 360936 264988
rect 360252 264948 360936 264976
rect 360252 264936 360258 264948
rect 360930 264936 360936 264948
rect 360988 264936 360994 264988
rect 180150 263576 180156 263628
rect 180208 263616 180214 263628
rect 197906 263616 197912 263628
rect 180208 263588 197912 263616
rect 180208 263576 180214 263588
rect 197906 263576 197912 263588
rect 197964 263576 197970 263628
rect 196710 261808 196716 261860
rect 196768 261848 196774 261860
rect 198642 261848 198648 261860
rect 196768 261820 198648 261848
rect 196768 261808 196774 261820
rect 198642 261808 198648 261820
rect 198700 261808 198706 261860
rect 302786 260788 302792 260840
rect 302844 260828 302850 260840
rect 370130 260828 370136 260840
rect 302844 260800 370136 260828
rect 302844 260788 302850 260800
rect 370130 260788 370136 260800
rect 370188 260788 370194 260840
rect 195330 259496 195336 259548
rect 195388 259536 195394 259548
rect 197722 259536 197728 259548
rect 195388 259508 197728 259536
rect 195388 259496 195394 259508
rect 197722 259496 197728 259508
rect 197780 259496 197786 259548
rect 464338 259360 464344 259412
rect 464396 259400 464402 259412
rect 580166 259400 580172 259412
rect 464396 259372 580172 259400
rect 464396 259360 464402 259372
rect 580166 259360 580172 259372
rect 580224 259360 580230 259412
rect 191098 256708 191104 256760
rect 191156 256748 191162 256760
rect 198090 256748 198096 256760
rect 191156 256720 198096 256748
rect 191156 256708 191162 256720
rect 198090 256708 198096 256720
rect 198148 256708 198154 256760
rect 302786 256708 302792 256760
rect 302844 256748 302850 256760
rect 370866 256748 370872 256760
rect 302844 256720 370872 256748
rect 302844 256708 302850 256720
rect 370866 256708 370872 256720
rect 370924 256708 370930 256760
rect 188430 255280 188436 255332
rect 188488 255320 188494 255332
rect 197354 255320 197360 255332
rect 188488 255292 197360 255320
rect 188488 255280 188494 255292
rect 197354 255280 197360 255292
rect 197412 255280 197418 255332
rect 187050 252560 187056 252612
rect 187108 252600 187114 252612
rect 197354 252600 197360 252612
rect 187108 252572 197360 252600
rect 187108 252560 187114 252572
rect 197354 252560 197360 252572
rect 197412 252560 197418 252612
rect 171778 248412 171784 248464
rect 171836 248452 171842 248464
rect 198182 248452 198188 248464
rect 171836 248424 198188 248452
rect 171836 248412 171842 248424
rect 198182 248412 198188 248424
rect 198240 248412 198246 248464
rect 302878 247664 302884 247716
rect 302936 247704 302942 247716
rect 370498 247704 370504 247716
rect 302936 247676 370504 247704
rect 302936 247664 302942 247676
rect 370498 247664 370504 247676
rect 370556 247664 370562 247716
rect 304258 245556 304264 245608
rect 304316 245596 304322 245608
rect 580166 245596 580172 245608
rect 304316 245568 580172 245596
rect 304316 245556 304322 245568
rect 580166 245556 580172 245568
rect 580224 245556 580230 245608
rect 171870 244264 171876 244316
rect 171928 244304 171934 244316
rect 197354 244304 197360 244316
rect 171928 244276 197360 244304
rect 171928 244264 171934 244276
rect 197354 244264 197360 244276
rect 197412 244264 197418 244316
rect 192478 241544 192484 241596
rect 192536 241584 192542 241596
rect 197722 241584 197728 241596
rect 192536 241556 197728 241584
rect 192536 241544 192542 241556
rect 197722 241544 197728 241556
rect 197780 241544 197786 241596
rect 370498 241476 370504 241528
rect 370556 241516 370562 241528
rect 375374 241516 375380 241528
rect 370556 241488 375380 241516
rect 370556 241476 370562 241488
rect 375374 241476 375380 241488
rect 375432 241476 375438 241528
rect 303154 240728 303160 240780
rect 303212 240768 303218 240780
rect 370314 240768 370320 240780
rect 303212 240740 370320 240768
rect 303212 240728 303218 240740
rect 370314 240728 370320 240740
rect 370372 240728 370378 240780
rect 171962 238756 171968 238808
rect 172020 238796 172026 238808
rect 197354 238796 197360 238808
rect 172020 238768 197360 238796
rect 172020 238756 172026 238768
rect 197354 238756 197360 238768
rect 197412 238756 197418 238808
rect 184382 237396 184388 237448
rect 184440 237436 184446 237448
rect 197354 237436 197360 237448
rect 184440 237408 197360 237436
rect 184440 237396 184446 237408
rect 197354 237396 197360 237408
rect 197412 237396 197418 237448
rect 303062 235220 303068 235272
rect 303120 235260 303126 235272
rect 369210 235260 369216 235272
rect 303120 235232 369216 235260
rect 303120 235220 303126 235232
rect 369210 235220 369216 235232
rect 369268 235220 369274 235272
rect 172054 234608 172060 234660
rect 172112 234648 172118 234660
rect 197538 234648 197544 234660
rect 172112 234620 197544 234648
rect 172112 234608 172118 234620
rect 197538 234608 197544 234620
rect 197596 234608 197602 234660
rect 191190 233384 191196 233436
rect 191248 233424 191254 233436
rect 198182 233424 198188 233436
rect 191248 233396 198188 233424
rect 191248 233384 191254 233396
rect 198182 233384 198188 233396
rect 198240 233384 198246 233436
rect 447962 233180 447968 233232
rect 448020 233220 448026 233232
rect 579982 233220 579988 233232
rect 448020 233192 579988 233220
rect 448020 233180 448026 233192
rect 579982 233180 579988 233192
rect 580040 233180 580046 233232
rect 369210 231684 369216 231736
rect 369268 231724 369274 231736
rect 374914 231724 374920 231736
rect 369268 231696 374920 231724
rect 369268 231684 369274 231696
rect 374914 231684 374920 231696
rect 374972 231684 374978 231736
rect 177482 230460 177488 230512
rect 177540 230500 177546 230512
rect 197630 230500 197636 230512
rect 177540 230472 197636 230500
rect 177540 230460 177546 230472
rect 197630 230460 197636 230472
rect 197688 230460 197694 230512
rect 302970 229712 302976 229764
rect 303028 229752 303034 229764
rect 369394 229752 369400 229764
rect 303028 229724 369400 229752
rect 303028 229712 303034 229724
rect 369394 229712 369400 229724
rect 369452 229712 369458 229764
rect 177298 229100 177304 229152
rect 177356 229140 177362 229152
rect 197354 229140 197360 229152
rect 177356 229112 197360 229140
rect 177356 229100 177362 229112
rect 197354 229100 197360 229112
rect 197412 229100 197418 229152
rect 369394 229100 369400 229152
rect 369452 229140 369458 229152
rect 373258 229140 373264 229152
rect 369452 229112 373264 229140
rect 369452 229100 369458 229112
rect 373258 229100 373264 229112
rect 373316 229100 373322 229152
rect 303154 228352 303160 228404
rect 303212 228392 303218 228404
rect 370222 228392 370228 228404
rect 303212 228364 370228 228392
rect 303212 228352 303218 228364
rect 370222 228352 370228 228364
rect 370280 228352 370286 228404
rect 436002 227740 436008 227792
rect 436060 227780 436066 227792
rect 441890 227780 441896 227792
rect 436060 227752 441896 227780
rect 436060 227740 436066 227752
rect 441890 227740 441896 227752
rect 441948 227740 441954 227792
rect 316678 226992 316684 227044
rect 316736 227032 316742 227044
rect 580258 227032 580264 227044
rect 316736 227004 580264 227032
rect 316736 226992 316742 227004
rect 580258 226992 580264 227004
rect 580316 226992 580322 227044
rect 437382 226244 437388 226296
rect 437440 226284 437446 226296
rect 441706 226284 441712 226296
rect 437440 226256 441712 226284
rect 437440 226244 437446 226256
rect 441706 226244 441712 226256
rect 441764 226244 441770 226296
rect 303246 225632 303252 225684
rect 303304 225672 303310 225684
rect 369946 225672 369952 225684
rect 303304 225644 369952 225672
rect 303304 225632 303310 225644
rect 369946 225632 369952 225644
rect 370004 225632 370010 225684
rect 302786 225564 302792 225616
rect 302844 225604 302850 225616
rect 370130 225604 370136 225616
rect 302844 225576 370136 225604
rect 302844 225564 302850 225576
rect 370130 225564 370136 225576
rect 370188 225564 370194 225616
rect 371602 225564 371608 225616
rect 371660 225604 371666 225616
rect 382366 225604 382372 225616
rect 371660 225576 382372 225604
rect 371660 225564 371666 225576
rect 382366 225564 382372 225576
rect 382424 225564 382430 225616
rect 445570 225564 445576 225616
rect 445628 225604 445634 225616
rect 447778 225604 447784 225616
rect 445628 225576 447784 225604
rect 445628 225564 445634 225576
rect 447778 225564 447784 225576
rect 447836 225604 447842 225616
rect 454218 225604 454224 225616
rect 447836 225576 454224 225604
rect 447836 225564 447842 225576
rect 454218 225564 454224 225576
rect 454276 225564 454282 225616
rect 372706 225020 372712 225072
rect 372764 225060 372770 225072
rect 372764 225032 383654 225060
rect 372764 225020 372770 225032
rect 371602 224952 371608 225004
rect 371660 224992 371666 225004
rect 374454 224992 374460 225004
rect 371660 224964 374460 224992
rect 371660 224952 371666 224964
rect 374454 224952 374460 224964
rect 374512 224992 374518 225004
rect 379514 224992 379520 225004
rect 374512 224964 379520 224992
rect 374512 224952 374518 224964
rect 379514 224952 379520 224964
rect 379572 224952 379578 225004
rect 383626 224992 383654 225032
rect 441798 224992 441804 225004
rect 383626 224964 441804 224992
rect 441798 224952 441804 224964
rect 441856 224952 441862 225004
rect 302694 224340 302700 224392
rect 302752 224380 302758 224392
rect 369854 224380 369860 224392
rect 302752 224352 369860 224380
rect 302752 224340 302758 224352
rect 369854 224340 369860 224352
rect 369912 224340 369918 224392
rect 302878 224272 302884 224324
rect 302936 224312 302942 224324
rect 370038 224312 370044 224324
rect 302936 224284 370044 224312
rect 302936 224272 302942 224284
rect 370038 224272 370044 224284
rect 370096 224272 370102 224324
rect 302786 224204 302792 224256
rect 302844 224244 302850 224256
rect 370314 224244 370320 224256
rect 302844 224216 370320 224244
rect 302844 224204 302850 224216
rect 370314 224204 370320 224216
rect 370372 224204 370378 224256
rect 372246 224204 372252 224256
rect 372304 224244 372310 224256
rect 373350 224244 373356 224256
rect 372304 224216 373356 224244
rect 372304 224204 372310 224216
rect 373350 224204 373356 224216
rect 373408 224244 373414 224256
rect 377122 224244 377128 224256
rect 373408 224216 377128 224244
rect 373408 224204 373414 224216
rect 377122 224204 377128 224216
rect 377180 224204 377186 224256
rect 379606 224244 379612 224256
rect 377232 224216 379612 224244
rect 376938 224176 376944 224188
rect 373966 224148 376944 224176
rect 359550 224068 359556 224120
rect 359608 224108 359614 224120
rect 373966 224108 373994 224148
rect 376938 224136 376944 224148
rect 376996 224176 377002 224188
rect 377232 224176 377260 224216
rect 379606 224204 379612 224216
rect 379664 224204 379670 224256
rect 382458 224176 382464 224188
rect 376996 224148 377260 224176
rect 379348 224148 382464 224176
rect 376996 224136 377002 224148
rect 359608 224080 373994 224108
rect 359608 224068 359614 224080
rect 359734 224000 359740 224052
rect 359792 224040 359798 224052
rect 379348 224040 379376 224148
rect 382458 224136 382464 224148
rect 382516 224176 382522 224188
rect 382642 224176 382648 224188
rect 382516 224148 382648 224176
rect 382516 224136 382522 224148
rect 382642 224136 382648 224148
rect 382700 224136 382706 224188
rect 359792 224012 379376 224040
rect 359792 224000 359798 224012
rect 379514 224000 379520 224052
rect 379572 224040 379578 224052
rect 380986 224040 380992 224052
rect 379572 224012 380992 224040
rect 379572 224000 379578 224012
rect 380986 224000 380992 224012
rect 381044 224000 381050 224052
rect 359642 223932 359648 223984
rect 359700 223972 359706 223984
rect 383654 223972 383660 223984
rect 359700 223944 383660 223972
rect 359700 223932 359706 223944
rect 383654 223932 383660 223944
rect 383712 223932 383718 223984
rect 358906 223864 358912 223916
rect 358964 223904 358970 223916
rect 358964 223876 369992 223904
rect 358964 223864 358970 223876
rect 369964 223836 369992 223876
rect 372706 223864 372712 223916
rect 372764 223904 372770 223916
rect 441798 223904 441804 223916
rect 372764 223876 441804 223904
rect 372764 223864 372770 223876
rect 441798 223864 441804 223876
rect 441856 223904 441862 223916
rect 452746 223904 452752 223916
rect 441856 223876 452752 223904
rect 441856 223864 441862 223876
rect 452746 223864 452752 223876
rect 452804 223904 452810 223916
rect 454126 223904 454132 223916
rect 452804 223876 454132 223904
rect 452804 223864 452810 223876
rect 454126 223864 454132 223876
rect 454184 223864 454190 223916
rect 372798 223836 372804 223848
rect 369964 223808 372804 223836
rect 372798 223796 372804 223808
rect 372856 223796 372862 223848
rect 371602 223728 371608 223780
rect 371660 223768 371666 223780
rect 379514 223768 379520 223780
rect 371660 223740 379520 223768
rect 371660 223728 371666 223740
rect 379514 223728 379520 223740
rect 379572 223728 379578 223780
rect 193858 223592 193864 223644
rect 193916 223632 193922 223644
rect 198274 223632 198280 223644
rect 193916 223604 198280 223632
rect 193916 223592 193922 223604
rect 198274 223592 198280 223604
rect 198332 223592 198338 223644
rect 441706 223592 441712 223644
rect 441764 223632 441770 223644
rect 441890 223632 441896 223644
rect 441764 223604 441896 223632
rect 441764 223592 441770 223604
rect 441890 223592 441896 223604
rect 441948 223592 441954 223644
rect 370866 223524 370872 223576
rect 370924 223564 370930 223576
rect 371418 223564 371424 223576
rect 370924 223536 371424 223564
rect 370924 223524 370930 223536
rect 371418 223524 371424 223536
rect 371476 223564 371482 223576
rect 378226 223564 378232 223576
rect 371476 223536 378232 223564
rect 371476 223524 371482 223536
rect 378226 223524 378232 223536
rect 378284 223564 378290 223576
rect 380986 223564 380992 223576
rect 378284 223536 380992 223564
rect 378284 223524 378290 223536
rect 380986 223524 380992 223536
rect 381044 223524 381050 223576
rect 447502 223524 447508 223576
rect 447560 223564 447566 223576
rect 450262 223564 450268 223576
rect 447560 223536 450268 223564
rect 447560 223524 447566 223536
rect 450262 223524 450268 223536
rect 450320 223524 450326 223576
rect 371602 223456 371608 223508
rect 371660 223496 371666 223508
rect 377398 223496 377404 223508
rect 371660 223468 377404 223496
rect 371660 223456 371666 223468
rect 377398 223456 377404 223468
rect 377456 223496 377462 223508
rect 381170 223496 381176 223508
rect 377456 223468 381176 223496
rect 377456 223456 377462 223468
rect 381170 223456 381176 223468
rect 381228 223456 381234 223508
rect 445662 223116 445668 223168
rect 445720 223156 445726 223168
rect 447502 223156 447508 223168
rect 445720 223128 447508 223156
rect 445720 223116 445726 223128
rect 447502 223116 447508 223128
rect 447560 223116 447566 223168
rect 371602 222640 371608 222692
rect 371660 222680 371666 222692
rect 375558 222680 375564 222692
rect 371660 222652 375564 222680
rect 371660 222640 371666 222652
rect 375558 222640 375564 222652
rect 375616 222680 375622 222692
rect 381078 222680 381084 222692
rect 375616 222652 381084 222680
rect 375616 222640 375622 222652
rect 381078 222640 381084 222652
rect 381136 222640 381142 222692
rect 170490 222164 170496 222216
rect 170548 222204 170554 222216
rect 197354 222204 197360 222216
rect 170548 222176 197360 222204
rect 170548 222164 170554 222176
rect 197354 222164 197360 222176
rect 197412 222164 197418 222216
rect 302786 222096 302792 222148
rect 302844 222136 302850 222148
rect 358906 222136 358912 222148
rect 302844 222108 358912 222136
rect 302844 222096 302850 222108
rect 358906 222096 358912 222108
rect 358964 222096 358970 222148
rect 375374 222096 375380 222148
rect 375432 222136 375438 222148
rect 378410 222136 378416 222148
rect 375432 222108 378416 222136
rect 375432 222096 375438 222108
rect 378410 222096 378416 222108
rect 378468 222096 378474 222148
rect 377030 222028 377036 222080
rect 377088 222068 377094 222080
rect 378502 222068 378508 222080
rect 377088 222040 378508 222068
rect 377088 222028 377094 222040
rect 378502 222028 378508 222040
rect 378560 222028 378566 222080
rect 445662 221212 445668 221264
rect 445720 221252 445726 221264
rect 451458 221252 451464 221264
rect 445720 221224 451464 221252
rect 445720 221212 445726 221224
rect 451458 221212 451464 221224
rect 451516 221252 451522 221264
rect 452654 221252 452660 221264
rect 451516 221224 452660 221252
rect 451516 221212 451522 221224
rect 452654 221212 452660 221224
rect 452712 221212 452718 221264
rect 370406 220872 370412 220924
rect 370464 220912 370470 220924
rect 377030 220912 377036 220924
rect 370464 220884 377036 220912
rect 370464 220872 370470 220884
rect 377030 220872 377036 220884
rect 377088 220872 377094 220924
rect 374914 220736 374920 220788
rect 374972 220776 374978 220788
rect 378318 220776 378324 220788
rect 374972 220748 378324 220776
rect 374972 220736 374978 220748
rect 378318 220736 378324 220748
rect 378376 220736 378382 220788
rect 445662 220736 445668 220788
rect 445720 220776 445726 220788
rect 446490 220776 446496 220788
rect 445720 220748 446496 220776
rect 445720 220736 445726 220748
rect 446490 220736 446496 220748
rect 446548 220776 446554 220788
rect 448882 220776 448888 220788
rect 446548 220748 448888 220776
rect 446548 220736 446554 220748
rect 448882 220736 448888 220748
rect 448940 220736 448946 220788
rect 375650 220668 375656 220720
rect 375708 220708 375714 220720
rect 378226 220708 378232 220720
rect 375708 220680 378232 220708
rect 375708 220668 375714 220680
rect 378226 220668 378232 220680
rect 378284 220668 378290 220720
rect 450170 219988 450176 220040
rect 450228 220028 450234 220040
rect 451274 220028 451280 220040
rect 450228 220000 451280 220028
rect 450228 219988 450234 220000
rect 451274 219988 451280 220000
rect 451332 219988 451338 220040
rect 369854 219648 369860 219700
rect 369912 219688 369918 219700
rect 375650 219688 375656 219700
rect 369912 219660 375656 219688
rect 369912 219648 369918 219660
rect 375650 219648 375656 219660
rect 375708 219648 375714 219700
rect 445662 219580 445668 219632
rect 445720 219620 445726 219632
rect 450170 219620 450176 219632
rect 445720 219592 450176 219620
rect 445720 219580 445726 219592
rect 450170 219580 450176 219592
rect 450228 219580 450234 219632
rect 369854 219512 369860 219564
rect 369912 219552 369918 219564
rect 370222 219552 370228 219564
rect 369912 219524 370228 219552
rect 369912 219512 369918 219524
rect 370222 219512 370228 219524
rect 370280 219512 370286 219564
rect 180242 219444 180248 219496
rect 180300 219484 180306 219496
rect 197538 219484 197544 219496
rect 180300 219456 197544 219484
rect 180300 219444 180306 219456
rect 197538 219444 197544 219456
rect 197596 219444 197602 219496
rect 373258 219444 373264 219496
rect 373316 219484 373322 219496
rect 374822 219484 374828 219496
rect 373316 219456 374828 219484
rect 373316 219444 373322 219456
rect 374822 219444 374828 219456
rect 374880 219444 374886 219496
rect 302786 219376 302792 219428
rect 302844 219416 302850 219428
rect 359734 219416 359740 219428
rect 302844 219388 359740 219416
rect 302844 219376 302850 219388
rect 359734 219376 359740 219388
rect 359792 219376 359798 219428
rect 369854 219376 369860 219428
rect 369912 219416 369918 219428
rect 376018 219416 376024 219428
rect 369912 219388 376024 219416
rect 369912 219376 369918 219388
rect 376018 219376 376024 219388
rect 376076 219376 376082 219428
rect 446122 218900 446128 218952
rect 446180 218940 446186 218952
rect 448606 218940 448612 218952
rect 446180 218912 448612 218940
rect 446180 218900 446186 218912
rect 448606 218900 448612 218912
rect 448664 218900 448670 218952
rect 369946 218832 369952 218884
rect 370004 218872 370010 218884
rect 373350 218872 373356 218884
rect 370004 218844 373356 218872
rect 370004 218832 370010 218844
rect 373350 218832 373356 218844
rect 373408 218872 373414 218884
rect 376754 218872 376760 218884
rect 373408 218844 376760 218872
rect 373408 218832 373414 218844
rect 376754 218832 376760 218844
rect 376812 218832 376818 218884
rect 370038 218696 370044 218748
rect 370096 218736 370102 218748
rect 376846 218736 376852 218748
rect 370096 218708 376852 218736
rect 370096 218696 370102 218708
rect 376846 218696 376852 218708
rect 376904 218696 376910 218748
rect 445478 218424 445484 218476
rect 445536 218464 445542 218476
rect 446122 218464 446128 218476
rect 445536 218436 446128 218464
rect 445536 218424 445542 218436
rect 446122 218424 446128 218436
rect 446180 218424 446186 218476
rect 196802 218152 196808 218204
rect 196860 218192 196866 218204
rect 198458 218192 198464 218204
rect 196860 218164 198464 218192
rect 196860 218152 196866 218164
rect 198458 218152 198464 218164
rect 198516 218152 198522 218204
rect 376018 218016 376024 218068
rect 376076 218056 376082 218068
rect 378226 218056 378232 218068
rect 376076 218028 378232 218056
rect 376076 218016 376082 218028
rect 378226 218016 378232 218028
rect 378284 218016 378290 218068
rect 370130 217948 370136 218000
rect 370188 217988 370194 218000
rect 370406 217988 370412 218000
rect 370188 217960 370412 217988
rect 370188 217948 370194 217960
rect 370406 217948 370412 217960
rect 370464 217988 370470 218000
rect 374730 217988 374736 218000
rect 370464 217960 374736 217988
rect 370464 217948 370470 217960
rect 374730 217948 374736 217960
rect 374788 217988 374794 218000
rect 376846 217988 376852 218000
rect 374788 217960 376852 217988
rect 374788 217948 374794 217960
rect 376846 217948 376852 217960
rect 376904 217948 376910 218000
rect 445662 217336 445668 217388
rect 445720 217376 445726 217388
rect 449986 217376 449992 217388
rect 445720 217348 449992 217376
rect 445720 217336 445726 217348
rect 449986 217336 449992 217348
rect 450044 217336 450050 217388
rect 370314 216928 370320 216980
rect 370372 216968 370378 216980
rect 374914 216968 374920 216980
rect 370372 216940 374920 216968
rect 370372 216928 370378 216940
rect 374914 216928 374920 216940
rect 374972 216968 374978 216980
rect 375742 216968 375748 216980
rect 374972 216940 375748 216968
rect 374972 216928 374978 216940
rect 375742 216928 375748 216940
rect 375800 216928 375806 216980
rect 302786 216588 302792 216640
rect 302844 216628 302850 216640
rect 359642 216628 359648 216640
rect 302844 216600 359648 216628
rect 302844 216588 302850 216600
rect 359642 216588 359648 216600
rect 359700 216588 359706 216640
rect 382642 216588 382648 216640
rect 382700 216628 382706 216640
rect 383654 216628 383660 216640
rect 382700 216600 383660 216628
rect 382700 216588 382706 216600
rect 383654 216588 383660 216600
rect 383712 216588 383718 216640
rect 371602 216520 371608 216572
rect 371660 216560 371666 216572
rect 382458 216560 382464 216572
rect 371660 216532 382464 216560
rect 371660 216520 371666 216532
rect 382458 216520 382464 216532
rect 382516 216560 382522 216572
rect 383746 216560 383752 216572
rect 382516 216532 383752 216560
rect 382516 216520 382522 216532
rect 383746 216520 383752 216532
rect 383804 216520 383810 216572
rect 372062 216384 372068 216436
rect 372120 216424 372126 216436
rect 372798 216424 372804 216436
rect 372120 216396 372804 216424
rect 372120 216384 372126 216396
rect 372798 216384 372804 216396
rect 372856 216424 372862 216436
rect 375834 216424 375840 216436
rect 372856 216396 375840 216424
rect 372856 216384 372862 216396
rect 375834 216384 375840 216396
rect 375892 216384 375898 216436
rect 445662 216112 445668 216164
rect 445720 216152 445726 216164
rect 447870 216152 447876 216164
rect 445720 216124 447876 216152
rect 445720 216112 445726 216124
rect 447870 216112 447876 216124
rect 447928 216112 447934 216164
rect 195422 215296 195428 215348
rect 195480 215336 195486 215348
rect 197906 215336 197912 215348
rect 195480 215308 197912 215336
rect 195480 215296 195486 215308
rect 197906 215296 197912 215308
rect 197964 215296 197970 215348
rect 371602 215296 371608 215348
rect 371660 215336 371666 215348
rect 382274 215336 382280 215348
rect 371660 215308 382280 215336
rect 371660 215296 371666 215308
rect 382274 215296 382280 215308
rect 382332 215336 382338 215348
rect 382642 215336 382648 215348
rect 382332 215308 382648 215336
rect 382332 215296 382338 215308
rect 382642 215296 382648 215308
rect 382700 215296 382706 215348
rect 447870 215296 447876 215348
rect 447928 215336 447934 215348
rect 448790 215336 448796 215348
rect 447928 215308 448796 215336
rect 447928 215296 447934 215308
rect 448790 215296 448796 215308
rect 448848 215296 448854 215348
rect 3326 215228 3332 215280
rect 3384 215268 3390 215280
rect 199378 215268 199384 215280
rect 3384 215240 199384 215268
rect 3384 215228 3390 215240
rect 199378 215228 199384 215240
rect 199436 215228 199442 215280
rect 445478 214752 445484 214804
rect 445536 214792 445542 214804
rect 448514 214792 448520 214804
rect 445536 214764 448520 214792
rect 445536 214752 445542 214764
rect 448514 214752 448520 214764
rect 448572 214792 448578 214804
rect 450078 214792 450084 214804
rect 448572 214764 450084 214792
rect 448572 214752 448578 214764
rect 450078 214752 450084 214764
rect 450136 214752 450142 214804
rect 371602 214616 371608 214668
rect 371660 214656 371666 214668
rect 376110 214656 376116 214668
rect 371660 214628 376116 214656
rect 371660 214616 371666 214628
rect 376110 214616 376116 214628
rect 376168 214656 376174 214668
rect 379606 214656 379612 214668
rect 376168 214628 379612 214656
rect 376168 214616 376174 214628
rect 379606 214616 379612 214628
rect 379664 214616 379670 214668
rect 371694 214548 371700 214600
rect 371752 214588 371758 214600
rect 376938 214588 376944 214600
rect 371752 214560 376944 214588
rect 371752 214548 371758 214560
rect 376938 214548 376944 214560
rect 376996 214548 377002 214600
rect 191282 213936 191288 213988
rect 191340 213976 191346 213988
rect 197354 213976 197360 213988
rect 191340 213948 197360 213976
rect 191340 213936 191346 213948
rect 197354 213936 197360 213948
rect 197412 213936 197418 213988
rect 302786 213868 302792 213920
rect 302844 213908 302850 213920
rect 359550 213908 359556 213920
rect 302844 213880 359556 213908
rect 302844 213868 302850 213880
rect 359550 213868 359556 213880
rect 359608 213868 359614 213920
rect 445662 213868 445668 213920
rect 445720 213908 445726 213920
rect 447318 213908 447324 213920
rect 445720 213880 447324 213908
rect 445720 213868 445726 213880
rect 447318 213868 447324 213880
rect 447376 213908 447382 213920
rect 449894 213908 449900 213920
rect 447376 213880 449900 213908
rect 447376 213868 447382 213880
rect 449894 213868 449900 213880
rect 449952 213868 449958 213920
rect 371694 213256 371700 213308
rect 371752 213296 371758 213308
rect 374638 213296 374644 213308
rect 371752 213268 374644 213296
rect 371752 213256 371758 213268
rect 374638 213256 374644 213268
rect 374696 213296 374702 213308
rect 380894 213296 380900 213308
rect 374696 213268 380900 213296
rect 374696 213256 374702 213268
rect 380894 213256 380900 213268
rect 380952 213256 380958 213308
rect 371602 213188 371608 213240
rect 371660 213228 371666 213240
rect 382550 213228 382556 213240
rect 371660 213200 382556 213228
rect 371660 213188 371666 213200
rect 382550 213188 382556 213200
rect 382608 213188 382614 213240
rect 371418 213052 371424 213104
rect 371476 213092 371482 213104
rect 375742 213092 375748 213104
rect 371476 213064 375748 213092
rect 371476 213052 371482 213064
rect 375742 213052 375748 213064
rect 375800 213092 375806 213104
rect 380802 213092 380808 213104
rect 375800 213064 380808 213092
rect 375800 213052 375806 213064
rect 380802 213052 380808 213064
rect 380860 213052 380866 213104
rect 445662 212712 445668 212764
rect 445720 212752 445726 212764
rect 446674 212752 446680 212764
rect 445720 212724 446680 212752
rect 445720 212712 445726 212724
rect 446674 212712 446680 212724
rect 446732 212752 446738 212764
rect 448606 212752 448612 212764
rect 446732 212724 448612 212752
rect 446732 212712 446738 212724
rect 448606 212712 448612 212724
rect 448664 212712 448670 212764
rect 446030 212440 446036 212492
rect 446088 212480 446094 212492
rect 448698 212480 448704 212492
rect 446088 212452 448704 212480
rect 446088 212440 446094 212452
rect 448698 212440 448704 212452
rect 448756 212440 448762 212492
rect 373166 211964 373172 212016
rect 373224 212004 373230 212016
rect 375466 212004 375472 212016
rect 373224 211976 375472 212004
rect 373224 211964 373230 211976
rect 375466 211964 375472 211976
rect 375524 211964 375530 212016
rect 371418 211828 371424 211880
rect 371476 211868 371482 211880
rect 377214 211868 377220 211880
rect 371476 211840 377220 211868
rect 371476 211828 371482 211840
rect 377214 211828 377220 211840
rect 377272 211828 377278 211880
rect 370222 211760 370228 211812
rect 370280 211800 370286 211812
rect 378134 211800 378140 211812
rect 370280 211772 378140 211800
rect 370280 211760 370286 211772
rect 378134 211760 378140 211772
rect 378192 211760 378198 211812
rect 445478 211556 445484 211608
rect 445536 211596 445542 211608
rect 446030 211596 446036 211608
rect 445536 211568 446036 211596
rect 445536 211556 445542 211568
rect 446030 211556 446036 211568
rect 446088 211556 446094 211608
rect 188522 211148 188528 211200
rect 188580 211188 188586 211200
rect 197722 211188 197728 211200
rect 188580 211160 197728 211188
rect 188580 211148 188586 211160
rect 197722 211148 197728 211160
rect 197780 211148 197786 211200
rect 373074 210604 373080 210656
rect 373132 210644 373138 210656
rect 374546 210644 374552 210656
rect 373132 210616 374552 210644
rect 373132 210604 373138 210616
rect 374546 210604 374552 210616
rect 374604 210604 374610 210656
rect 445386 210468 445392 210520
rect 445444 210508 445450 210520
rect 447226 210508 447232 210520
rect 445444 210480 447232 210508
rect 445444 210468 445450 210480
rect 447226 210468 447232 210480
rect 447284 210468 447290 210520
rect 445202 209176 445208 209228
rect 445260 209216 445266 209228
rect 446582 209216 446588 209228
rect 445260 209188 446588 209216
rect 445260 209176 445266 209188
rect 446582 209176 446588 209188
rect 446640 209176 446646 209228
rect 187142 208360 187148 208412
rect 187200 208400 187206 208412
rect 197354 208400 197360 208412
rect 187200 208372 197360 208400
rect 187200 208360 187206 208372
rect 197354 208360 197360 208372
rect 197412 208360 197418 208412
rect 446582 208360 446588 208412
rect 446640 208400 446646 208412
rect 447410 208400 447416 208412
rect 446640 208372 447416 208400
rect 446640 208360 446646 208372
rect 447410 208360 447416 208372
rect 447468 208360 447474 208412
rect 444742 207884 444748 207936
rect 444800 207924 444806 207936
rect 445938 207924 445944 207936
rect 444800 207896 445944 207924
rect 444800 207884 444806 207896
rect 445938 207884 445944 207896
rect 445996 207924 446002 207936
rect 447134 207924 447140 207936
rect 445996 207896 447140 207924
rect 445996 207884 446002 207896
rect 447134 207884 447140 207896
rect 447192 207884 447198 207936
rect 173158 207000 173164 207052
rect 173216 207040 173222 207052
rect 197354 207040 197360 207052
rect 173216 207012 197360 207040
rect 173216 207000 173222 207012
rect 197354 207000 197360 207012
rect 197412 207000 197418 207052
rect 450538 206932 450544 206984
rect 450596 206972 450602 206984
rect 579798 206972 579804 206984
rect 450596 206944 579804 206972
rect 450596 206932 450602 206944
rect 579798 206932 579804 206944
rect 579856 206932 579862 206984
rect 371602 206252 371608 206304
rect 371660 206292 371666 206304
rect 374178 206292 374184 206304
rect 371660 206264 374184 206292
rect 371660 206252 371666 206264
rect 374178 206252 374184 206264
rect 374236 206252 374242 206304
rect 371694 205776 371700 205828
rect 371752 205816 371758 205828
rect 372982 205816 372988 205828
rect 371752 205788 372988 205816
rect 371752 205776 371758 205788
rect 372982 205776 372988 205788
rect 373040 205776 373046 205828
rect 302326 205640 302332 205692
rect 302384 205680 302390 205692
rect 359550 205680 359556 205692
rect 302384 205652 359556 205680
rect 302384 205640 302390 205652
rect 359550 205640 359556 205652
rect 359608 205640 359614 205692
rect 373810 205572 373816 205624
rect 373868 205612 373874 205624
rect 374178 205612 374184 205624
rect 373868 205584 374184 205612
rect 373868 205572 373874 205584
rect 374178 205572 374184 205584
rect 374236 205572 374242 205624
rect 369118 205164 369124 205216
rect 369176 205204 369182 205216
rect 369302 205204 369308 205216
rect 369176 205176 369308 205204
rect 369176 205164 369182 205176
rect 369302 205164 369308 205176
rect 369360 205164 369366 205216
rect 173250 204280 173256 204332
rect 173308 204320 173314 204332
rect 197538 204320 197544 204332
rect 173308 204292 197544 204320
rect 173308 204280 173314 204292
rect 197538 204280 197544 204292
rect 197596 204280 197602 204332
rect 372062 204212 372068 204264
rect 372120 204252 372126 204264
rect 373994 204252 374000 204264
rect 372120 204224 374000 204252
rect 372120 204212 372126 204224
rect 373994 204212 374000 204224
rect 374052 204212 374058 204264
rect 173342 202852 173348 202904
rect 173400 202892 173406 202904
rect 197354 202892 197360 202904
rect 173400 202864 197360 202892
rect 173400 202852 173406 202864
rect 197354 202852 197360 202864
rect 197412 202852 197418 202904
rect 302786 202852 302792 202904
rect 302844 202892 302850 202904
rect 359642 202892 359648 202904
rect 302844 202864 359648 202892
rect 302844 202852 302850 202864
rect 359642 202852 359648 202864
rect 359700 202852 359706 202904
rect 3050 202784 3056 202836
rect 3108 202824 3114 202836
rect 177390 202824 177396 202836
rect 3108 202796 177396 202824
rect 3108 202784 3114 202796
rect 177390 202784 177396 202796
rect 177448 202784 177454 202836
rect 370130 202716 370136 202768
rect 370188 202756 370194 202768
rect 374270 202756 374276 202768
rect 370188 202728 374276 202756
rect 370188 202716 370194 202728
rect 374270 202716 374276 202728
rect 374328 202716 374334 202768
rect 373166 202648 373172 202700
rect 373224 202688 373230 202700
rect 375374 202688 375380 202700
rect 373224 202660 375380 202688
rect 373224 202648 373230 202660
rect 375374 202648 375380 202660
rect 375432 202648 375438 202700
rect 372614 202512 372620 202564
rect 372672 202552 372678 202564
rect 373258 202552 373264 202564
rect 372672 202524 373264 202552
rect 372672 202512 372678 202524
rect 373258 202512 373264 202524
rect 373316 202512 373322 202564
rect 371602 201560 371608 201612
rect 371660 201600 371666 201612
rect 373994 201600 374000 201612
rect 371660 201572 374000 201600
rect 371660 201560 371666 201572
rect 373994 201560 374000 201572
rect 374052 201600 374058 201612
rect 374362 201600 374368 201612
rect 374052 201572 374368 201600
rect 374052 201560 374058 201572
rect 374362 201560 374368 201572
rect 374420 201560 374426 201612
rect 445662 201492 445668 201544
rect 445720 201532 445726 201544
rect 448514 201532 448520 201544
rect 445720 201504 448520 201532
rect 445720 201492 445726 201504
rect 448514 201492 448520 201504
rect 448572 201532 448578 201544
rect 452930 201532 452936 201544
rect 448572 201504 452936 201532
rect 448572 201492 448578 201504
rect 452930 201492 452936 201504
rect 452988 201492 452994 201544
rect 173434 200132 173440 200184
rect 173492 200172 173498 200184
rect 197354 200172 197360 200184
rect 173492 200144 197360 200172
rect 173492 200132 173498 200144
rect 197354 200132 197360 200144
rect 197412 200132 197418 200184
rect 445662 200132 445668 200184
rect 445720 200172 445726 200184
rect 449250 200172 449256 200184
rect 445720 200144 449256 200172
rect 445720 200132 445726 200144
rect 449250 200132 449256 200144
rect 449308 200172 449314 200184
rect 452654 200172 452660 200184
rect 449308 200144 452660 200172
rect 449308 200132 449314 200144
rect 452654 200132 452660 200144
rect 452712 200132 452718 200184
rect 445662 199452 445668 199504
rect 445720 199492 445726 199504
rect 449894 199492 449900 199504
rect 445720 199464 449900 199492
rect 445720 199452 445726 199464
rect 449894 199452 449900 199464
rect 449952 199492 449958 199504
rect 454034 199492 454040 199504
rect 449952 199464 454040 199492
rect 449952 199452 449958 199464
rect 454034 199452 454040 199464
rect 454092 199452 454098 199504
rect 445662 198772 445668 198824
rect 445720 198812 445726 198824
rect 451366 198812 451372 198824
rect 445720 198784 451372 198812
rect 445720 198772 445726 198784
rect 451366 198772 451372 198784
rect 451424 198772 451430 198824
rect 173526 198704 173532 198756
rect 173584 198744 173590 198756
rect 197354 198744 197360 198756
rect 173584 198716 197360 198744
rect 173584 198704 173590 198716
rect 197354 198704 197360 198716
rect 197412 198704 197418 198756
rect 302510 198704 302516 198756
rect 302568 198744 302574 198756
rect 359366 198744 359372 198756
rect 302568 198716 359372 198744
rect 302568 198704 302574 198716
rect 359366 198704 359372 198716
rect 359424 198704 359430 198756
rect 445662 197752 445668 197804
rect 445720 197792 445726 197804
rect 447134 197792 447140 197804
rect 445720 197764 447140 197792
rect 445720 197752 445726 197764
rect 447134 197752 447140 197764
rect 447192 197792 447198 197804
rect 452838 197792 452844 197804
rect 447192 197764 452844 197792
rect 447192 197752 447198 197764
rect 452838 197752 452844 197764
rect 452896 197752 452902 197804
rect 302878 197208 302884 197260
rect 302936 197248 302942 197260
rect 379606 197248 379612 197260
rect 302936 197220 379612 197248
rect 302936 197208 302942 197220
rect 379606 197208 379612 197220
rect 379664 197208 379670 197260
rect 302694 197140 302700 197192
rect 302752 197180 302758 197192
rect 370314 197180 370320 197192
rect 302752 197152 370320 197180
rect 302752 197140 302758 197152
rect 370314 197140 370320 197152
rect 370372 197140 370378 197192
rect 359642 197072 359648 197124
rect 359700 197112 359706 197124
rect 382458 197112 382464 197124
rect 359700 197084 382464 197112
rect 359700 197072 359706 197084
rect 382458 197072 382464 197084
rect 382516 197072 382522 197124
rect 359366 197004 359372 197056
rect 359424 197044 359430 197056
rect 380894 197044 380900 197056
rect 359424 197016 380900 197044
rect 359424 197004 359430 197016
rect 380894 197004 380900 197016
rect 380952 197004 380958 197056
rect 359550 196936 359556 196988
rect 359608 196976 359614 196988
rect 375742 196976 375748 196988
rect 359608 196948 375748 196976
rect 359608 196936 359614 196948
rect 375742 196936 375748 196948
rect 375800 196936 375806 196988
rect 302970 196664 302976 196716
rect 303028 196704 303034 196716
rect 369854 196704 369860 196716
rect 303028 196676 369860 196704
rect 303028 196664 303034 196676
rect 369854 196664 369860 196676
rect 369912 196664 369918 196716
rect 303062 196596 303068 196648
rect 303120 196636 303126 196648
rect 375374 196636 375380 196648
rect 303120 196608 375380 196636
rect 303120 196596 303126 196608
rect 375374 196596 375380 196608
rect 375432 196596 375438 196648
rect 369854 196052 369860 196104
rect 369912 196092 369918 196104
rect 371142 196092 371148 196104
rect 369912 196064 371148 196092
rect 369912 196052 369918 196064
rect 371142 196052 371148 196064
rect 371200 196052 371206 196104
rect 173618 195984 173624 196036
rect 173676 196024 173682 196036
rect 197354 196024 197360 196036
rect 173676 195996 197360 196024
rect 173676 195984 173682 195996
rect 197354 195984 197360 195996
rect 197412 195984 197418 196036
rect 322198 195916 322204 195968
rect 322256 195956 322262 195968
rect 438762 195956 438768 195968
rect 322256 195928 438768 195956
rect 322256 195916 322262 195928
rect 438762 195916 438768 195928
rect 438820 195916 438826 195968
rect 302878 195236 302884 195288
rect 302936 195276 302942 195288
rect 370498 195276 370504 195288
rect 302936 195248 370504 195276
rect 302936 195236 302942 195248
rect 370498 195236 370504 195248
rect 370556 195236 370562 195288
rect 302418 194488 302424 194540
rect 302476 194528 302482 194540
rect 370958 194528 370964 194540
rect 302476 194500 370964 194528
rect 302476 194488 302482 194500
rect 370958 194488 370964 194500
rect 371016 194528 371022 194540
rect 372706 194528 372712 194540
rect 371016 194500 372712 194528
rect 371016 194488 371022 194500
rect 372706 194488 372712 194500
rect 372764 194488 372770 194540
rect 437382 194488 437388 194540
rect 437440 194528 437446 194540
rect 441798 194528 441804 194540
rect 437440 194500 441804 194528
rect 437440 194488 437446 194500
rect 441798 194488 441804 194500
rect 441856 194488 441862 194540
rect 318058 194420 318064 194472
rect 318116 194460 318122 194472
rect 366910 194460 366916 194472
rect 318116 194432 366916 194460
rect 318116 194420 318122 194432
rect 366910 194420 366916 194432
rect 366968 194420 366974 194472
rect 436002 194420 436008 194472
rect 436060 194460 436066 194472
rect 441706 194460 441712 194472
rect 436060 194432 441712 194460
rect 436060 194420 436066 194432
rect 441706 194420 441712 194432
rect 441764 194420 441770 194472
rect 196894 194352 196900 194404
rect 196952 194392 196958 194404
rect 198642 194392 198648 194404
rect 196952 194364 198648 194392
rect 196952 194352 196958 194364
rect 198642 194352 198648 194364
rect 198700 194352 198706 194404
rect 435174 193604 435180 193656
rect 435232 193644 435238 193656
rect 436002 193644 436008 193656
rect 435232 193616 436008 193644
rect 435232 193604 435238 193616
rect 436002 193604 436008 193616
rect 436060 193604 436066 193656
rect 373074 193196 373080 193248
rect 373132 193236 373138 193248
rect 374086 193236 374092 193248
rect 373132 193208 374092 193236
rect 373132 193196 373138 193208
rect 374086 193196 374092 193208
rect 374144 193196 374150 193248
rect 446398 193128 446404 193180
rect 446456 193168 446462 193180
rect 580166 193168 580172 193180
rect 446456 193140 580172 193168
rect 446456 193128 446462 193140
rect 580166 193128 580172 193140
rect 580224 193128 580230 193180
rect 176010 191836 176016 191888
rect 176068 191876 176074 191888
rect 197354 191876 197360 191888
rect 176068 191848 197360 191876
rect 176068 191836 176074 191848
rect 197354 191836 197360 191848
rect 197412 191836 197418 191888
rect 172422 190408 172428 190460
rect 172480 190448 172486 190460
rect 188338 190448 188344 190460
rect 172480 190420 188344 190448
rect 172480 190408 172486 190420
rect 188338 190408 188344 190420
rect 188396 190408 188402 190460
rect 172422 188980 172428 189032
rect 172480 189020 172486 189032
rect 184290 189020 184296 189032
rect 172480 188992 184296 189020
rect 172480 188980 172486 188992
rect 184290 188980 184296 188992
rect 184348 188980 184354 189032
rect 181530 187688 181536 187740
rect 181588 187728 181594 187740
rect 197354 187728 197360 187740
rect 181588 187700 197360 187728
rect 181588 187688 181594 187700
rect 197354 187688 197360 187700
rect 197412 187688 197418 187740
rect 172422 187620 172428 187672
rect 172480 187660 172486 187672
rect 186958 187660 186964 187672
rect 172480 187632 186964 187660
rect 172480 187620 172486 187632
rect 186958 187620 186964 187632
rect 187016 187620 187022 187672
rect 302694 187620 302700 187672
rect 302752 187660 302758 187672
rect 374086 187660 374092 187672
rect 302752 187632 374092 187660
rect 302752 187620 302758 187632
rect 374086 187620 374092 187632
rect 374144 187620 374150 187672
rect 172422 186260 172428 186312
rect 172480 186300 172486 186312
rect 193950 186300 193956 186312
rect 172480 186272 193956 186300
rect 172480 186260 172486 186272
rect 193950 186260 193956 186272
rect 194008 186260 194014 186312
rect 182910 184900 182916 184952
rect 182968 184940 182974 184952
rect 197354 184940 197360 184952
rect 182968 184912 197360 184940
rect 182968 184900 182974 184912
rect 197354 184900 197360 184912
rect 197412 184900 197418 184952
rect 172330 184832 172336 184884
rect 172388 184872 172394 184884
rect 196618 184872 196624 184884
rect 172388 184844 196624 184872
rect 172388 184832 172394 184844
rect 196618 184832 196624 184844
rect 196676 184832 196682 184884
rect 302786 184832 302792 184884
rect 302844 184872 302850 184884
rect 370130 184872 370136 184884
rect 302844 184844 370136 184872
rect 302844 184832 302850 184844
rect 370130 184832 370136 184844
rect 370188 184872 370194 184884
rect 374270 184872 374276 184884
rect 370188 184844 374276 184872
rect 370188 184832 370194 184844
rect 374270 184832 374276 184844
rect 374328 184832 374334 184884
rect 172422 184764 172428 184816
rect 172480 184804 172486 184816
rect 182818 184804 182824 184816
rect 172480 184776 182824 184804
rect 172480 184764 172486 184776
rect 182818 184764 182824 184776
rect 182876 184764 182882 184816
rect 172422 183472 172428 183524
rect 172480 183512 172486 183524
rect 181438 183512 181444 183524
rect 172480 183484 181444 183512
rect 172480 183472 172486 183484
rect 181438 183472 181444 183484
rect 181496 183472 181502 183524
rect 178862 182792 178868 182844
rect 178920 182832 178926 182844
rect 197538 182832 197544 182844
rect 178920 182804 197544 182832
rect 178920 182792 178926 182804
rect 197538 182792 197544 182804
rect 197596 182792 197602 182844
rect 172422 182044 172428 182096
rect 172480 182084 172486 182096
rect 178770 182084 178776 182096
rect 172480 182056 178776 182084
rect 172480 182044 172486 182056
rect 178770 182044 178776 182056
rect 178828 182044 178834 182096
rect 172146 180820 172152 180872
rect 172204 180860 172210 180872
rect 197354 180860 197360 180872
rect 172204 180832 197360 180860
rect 172204 180820 172210 180832
rect 197354 180820 197360 180832
rect 197412 180820 197418 180872
rect 172422 180548 172428 180600
rect 172480 180588 172486 180600
rect 175918 180588 175924 180600
rect 172480 180560 175924 180588
rect 172480 180548 172486 180560
rect 175918 180548 175924 180560
rect 175976 180548 175982 180600
rect 461578 179324 461584 179376
rect 461636 179364 461642 179376
rect 580166 179364 580172 179376
rect 461636 179336 580172 179364
rect 461636 179324 461642 179336
rect 580166 179324 580172 179336
rect 580224 179324 580230 179376
rect 172422 179188 172428 179240
rect 172480 179228 172486 179240
rect 174538 179228 174544 179240
rect 172480 179200 174544 179228
rect 172480 179188 172486 179200
rect 174538 179188 174544 179200
rect 174596 179188 174602 179240
rect 191374 178032 191380 178084
rect 191432 178072 191438 178084
rect 197538 178072 197544 178084
rect 191432 178044 197544 178072
rect 191432 178032 191438 178044
rect 197538 178032 197544 178044
rect 197596 178032 197602 178084
rect 172422 177964 172428 178016
rect 172480 178004 172486 178016
rect 196710 178004 196716 178016
rect 172480 177976 196716 178004
rect 172480 177964 172486 177976
rect 196710 177964 196716 177976
rect 196768 177964 196774 178016
rect 172330 177896 172336 177948
rect 172388 177936 172394 177948
rect 180150 177936 180156 177948
rect 172388 177908 180156 177936
rect 172388 177896 172394 177908
rect 180150 177896 180156 177908
rect 180208 177896 180214 177948
rect 180334 176672 180340 176724
rect 180392 176712 180398 176724
rect 197354 176712 197360 176724
rect 180392 176684 197360 176712
rect 180392 176672 180398 176684
rect 197354 176672 197360 176684
rect 197412 176672 197418 176724
rect 172422 176604 172428 176656
rect 172480 176644 172486 176656
rect 195330 176644 195336 176656
rect 172480 176616 195336 176644
rect 172480 176604 172486 176616
rect 195330 176604 195336 176616
rect 195388 176604 195394 176656
rect 171686 175176 171692 175228
rect 171744 175216 171750 175228
rect 191098 175216 191104 175228
rect 171744 175188 191104 175216
rect 171744 175176 171750 175188
rect 191098 175176 191104 175188
rect 191156 175176 191162 175228
rect 302234 175176 302240 175228
rect 302292 175216 302298 175228
rect 370866 175216 370872 175228
rect 302292 175188 370872 175216
rect 302292 175176 302298 175188
rect 370866 175176 370872 175188
rect 370924 175176 370930 175228
rect 446122 175216 446128 175228
rect 373966 175188 446128 175216
rect 369762 175108 369768 175160
rect 369820 175148 369826 175160
rect 373810 175148 373816 175160
rect 369820 175120 373816 175148
rect 369820 175108 369826 175120
rect 373810 175108 373816 175120
rect 373868 175148 373874 175160
rect 373966 175148 373994 175188
rect 446122 175176 446128 175188
rect 446180 175176 446186 175228
rect 373868 175120 373994 175148
rect 373868 175108 373874 175120
rect 188338 173884 188344 173936
rect 188396 173924 188402 173936
rect 197630 173924 197636 173936
rect 188396 173896 197636 173924
rect 188396 173884 188402 173896
rect 197630 173884 197636 173896
rect 197688 173884 197694 173936
rect 171502 173816 171508 173868
rect 171560 173856 171566 173868
rect 188430 173856 188436 173868
rect 171560 173828 188436 173856
rect 171560 173816 171566 173828
rect 188430 173816 188436 173828
rect 188488 173816 188494 173868
rect 174538 172524 174544 172576
rect 174596 172564 174602 172576
rect 197354 172564 197360 172576
rect 174596 172536 197360 172564
rect 174596 172524 174602 172536
rect 197354 172524 197360 172536
rect 197412 172524 197418 172576
rect 172422 172456 172428 172508
rect 172480 172496 172486 172508
rect 187050 172496 187056 172508
rect 172480 172468 187056 172496
rect 172480 172456 172486 172468
rect 187050 172456 187056 172468
rect 187108 172456 187114 172508
rect 370130 172456 370136 172508
rect 370188 172496 370194 172508
rect 371694 172496 371700 172508
rect 370188 172468 371700 172496
rect 370188 172456 370194 172468
rect 371694 172456 371700 172468
rect 371752 172456 371758 172508
rect 302786 171096 302792 171148
rect 302844 171136 302850 171148
rect 370130 171136 370136 171148
rect 302844 171108 370136 171136
rect 302844 171096 302850 171108
rect 370130 171096 370136 171108
rect 370188 171096 370194 171148
rect 172422 171028 172428 171080
rect 172480 171068 172486 171080
rect 197998 171068 198004 171080
rect 172480 171040 198004 171068
rect 172480 171028 172486 171040
rect 197998 171028 198004 171040
rect 198056 171028 198062 171080
rect 186958 169736 186964 169788
rect 187016 169776 187022 169788
rect 197354 169776 197360 169788
rect 187016 169748 197360 169776
rect 187016 169736 187022 169748
rect 197354 169736 197360 169748
rect 197412 169736 197418 169788
rect 172422 169668 172428 169720
rect 172480 169708 172486 169720
rect 198090 169708 198096 169720
rect 172480 169680 198096 169708
rect 172480 169668 172486 169680
rect 198090 169668 198096 169680
rect 198148 169668 198154 169720
rect 369670 169668 369676 169720
rect 369728 169708 369734 169720
rect 374730 169708 374736 169720
rect 369728 169680 374736 169708
rect 369728 169668 369734 169680
rect 374730 169668 374736 169680
rect 374788 169708 374794 169720
rect 448698 169708 448704 169720
rect 374788 169680 448704 169708
rect 374788 169668 374794 169680
rect 448698 169668 448704 169680
rect 448756 169668 448762 169720
rect 369578 168308 369584 168360
rect 369636 168348 369642 168360
rect 374638 168348 374644 168360
rect 369636 168320 374644 168348
rect 369636 168308 369642 168320
rect 374638 168308 374644 168320
rect 374696 168348 374702 168360
rect 450078 168348 450084 168360
rect 374696 168320 450084 168348
rect 374696 168308 374702 168320
rect 450078 168308 450084 168320
rect 450136 168308 450142 168360
rect 195330 167016 195336 167068
rect 195388 167056 195394 167068
rect 197906 167056 197912 167068
rect 195388 167028 197912 167056
rect 195388 167016 195394 167028
rect 197906 167016 197912 167028
rect 197964 167016 197970 167068
rect 172422 166948 172428 167000
rect 172480 166988 172486 167000
rect 192478 166988 192484 167000
rect 172480 166960 192484 166988
rect 172480 166948 172486 166960
rect 192478 166948 192484 166960
rect 192536 166948 192542 167000
rect 301498 166948 301504 167000
rect 301556 166988 301562 167000
rect 580166 166988 580172 167000
rect 301556 166960 580172 166988
rect 301556 166948 301562 166960
rect 580166 166948 580172 166960
rect 580224 166948 580230 167000
rect 191098 166064 191104 166116
rect 191156 166104 191162 166116
rect 198458 166104 198464 166116
rect 191156 166076 198464 166104
rect 191156 166064 191162 166076
rect 198458 166064 198464 166076
rect 198516 166064 198522 166116
rect 171778 164840 171784 164892
rect 171836 164880 171842 164892
rect 191190 164880 191196 164892
rect 171836 164852 191196 164880
rect 171836 164840 171842 164852
rect 191190 164840 191196 164852
rect 191248 164840 191254 164892
rect 447410 164268 447416 164280
rect 370516 164240 447416 164268
rect 370516 164212 370544 164240
rect 447410 164228 447416 164240
rect 447468 164228 447474 164280
rect 3234 164160 3240 164212
rect 3292 164200 3298 164212
rect 159358 164200 159364 164212
rect 3292 164172 159364 164200
rect 3292 164160 3298 164172
rect 159358 164160 159364 164172
rect 159416 164160 159422 164212
rect 172422 164160 172428 164212
rect 172480 164200 172486 164212
rect 184382 164200 184388 164212
rect 172480 164172 184388 164200
rect 172480 164160 172486 164172
rect 184382 164160 184388 164172
rect 184440 164160 184446 164212
rect 370038 164160 370044 164212
rect 370096 164200 370102 164212
rect 370498 164200 370504 164212
rect 370096 164172 370504 164200
rect 370096 164160 370102 164172
rect 370498 164160 370504 164172
rect 370556 164160 370562 164212
rect 370590 164160 370596 164212
rect 370648 164200 370654 164212
rect 372982 164200 372988 164212
rect 370648 164172 372988 164200
rect 370648 164160 370654 164172
rect 372982 164160 372988 164172
rect 373040 164200 373046 164212
rect 449986 164200 449992 164212
rect 373040 164172 449992 164200
rect 373040 164160 373046 164172
rect 449986 164160 449992 164172
rect 450044 164160 450050 164212
rect 370222 162664 370228 162716
rect 370280 162704 370286 162716
rect 371142 162704 371148 162716
rect 370280 162676 371148 162704
rect 370280 162664 370286 162676
rect 371142 162664 371148 162676
rect 371200 162664 371206 162716
rect 372062 162188 372068 162240
rect 372120 162228 372126 162240
rect 444650 162228 444656 162240
rect 372120 162200 444656 162228
rect 372120 162188 372126 162200
rect 444650 162188 444656 162200
rect 444708 162188 444714 162240
rect 171778 162120 171784 162172
rect 171836 162160 171842 162172
rect 191374 162160 191380 162172
rect 171836 162132 191380 162160
rect 171836 162120 171842 162132
rect 191374 162120 191380 162132
rect 191432 162120 191438 162172
rect 302694 162120 302700 162172
rect 302752 162160 302758 162172
rect 370222 162160 370228 162172
rect 302752 162132 370228 162160
rect 302752 162120 302758 162132
rect 370222 162120 370228 162132
rect 370280 162120 370286 162172
rect 373258 162120 373264 162172
rect 373316 162160 373322 162172
rect 447226 162160 447232 162172
rect 373316 162132 447232 162160
rect 373316 162120 373322 162132
rect 447226 162120 447232 162132
rect 447284 162120 447290 162172
rect 184290 161440 184296 161492
rect 184348 161480 184354 161492
rect 197354 161480 197360 161492
rect 184348 161452 197360 161480
rect 184348 161440 184354 161452
rect 197354 161440 197360 161452
rect 197412 161440 197418 161492
rect 172238 161100 172244 161152
rect 172296 161140 172302 161152
rect 177482 161140 177488 161152
rect 172296 161112 177488 161140
rect 172296 161100 172302 161112
rect 177482 161100 177488 161112
rect 177540 161100 177546 161152
rect 169202 160760 169208 160812
rect 169260 160800 169266 160812
rect 180058 160800 180064 160812
rect 169260 160772 180064 160800
rect 169260 160760 169266 160772
rect 180058 160760 180064 160772
rect 180116 160760 180122 160812
rect 195238 160732 195244 160744
rect 171106 160704 195244 160732
rect 165154 160488 165160 160540
rect 165212 160528 165218 160540
rect 171106 160528 171134 160704
rect 195238 160692 195244 160704
rect 195296 160692 195302 160744
rect 165212 160500 171134 160528
rect 165212 160488 165218 160500
rect 446030 160120 446036 160132
rect 371252 160092 446036 160120
rect 369854 160012 369860 160064
rect 369912 160052 369918 160064
rect 371252 160052 371280 160092
rect 446030 160080 446036 160092
rect 446088 160080 446094 160132
rect 447318 160052 447324 160064
rect 369912 160024 371280 160052
rect 373966 160024 447324 160052
rect 369912 160012 369918 160024
rect 373966 159996 373994 160024
rect 447318 160012 447324 160024
rect 447376 160012 447382 160064
rect 369394 159944 369400 159996
rect 369452 159984 369458 159996
rect 373902 159984 373908 159996
rect 369452 159956 373908 159984
rect 369452 159944 369458 159956
rect 373902 159944 373908 159956
rect 373960 159956 373994 159996
rect 373960 159944 373966 159956
rect 180058 158720 180064 158772
rect 180116 158760 180122 158772
rect 197354 158760 197360 158772
rect 180116 158732 197360 158760
rect 180116 158720 180122 158732
rect 197354 158720 197360 158732
rect 197412 158720 197418 158772
rect 162854 158652 162860 158704
rect 162912 158692 162918 158704
rect 184198 158692 184204 158704
rect 162912 158664 184204 158692
rect 162912 158652 162918 158664
rect 184198 158652 184204 158664
rect 184256 158652 184262 158704
rect 166902 157972 166908 158024
rect 166960 158012 166966 158024
rect 196618 158012 196624 158024
rect 166960 157984 196624 158012
rect 166960 157972 166966 157984
rect 196618 157972 196624 157984
rect 196676 157972 196682 158024
rect 371878 157972 371884 158024
rect 371936 158012 371942 158024
rect 444466 158012 444472 158024
rect 371936 157984 444472 158012
rect 371936 157972 371942 157984
rect 444466 157972 444472 157984
rect 444524 157972 444530 158024
rect 177390 157360 177396 157412
rect 177448 157400 177454 157412
rect 197354 157400 197360 157412
rect 177448 157372 197360 157400
rect 177448 157360 177454 157372
rect 197354 157360 197360 157372
rect 197412 157360 197418 157412
rect 369486 156612 369492 156664
rect 369544 156652 369550 156664
rect 374546 156652 374552 156664
rect 369544 156624 374552 156652
rect 369544 156612 369550 156624
rect 374546 156612 374552 156624
rect 374604 156652 374610 156664
rect 444742 156652 444748 156664
rect 374604 156624 444748 156652
rect 374604 156612 374610 156624
rect 444742 156612 444748 156624
rect 444800 156652 444806 156664
rect 448606 156652 448612 156664
rect 444800 156624 448612 156652
rect 444800 156612 444806 156624
rect 448606 156612 448612 156624
rect 448664 156612 448670 156664
rect 436002 155864 436008 155916
rect 436060 155904 436066 155916
rect 441706 155904 441712 155916
rect 436060 155876 441712 155904
rect 436060 155864 436066 155876
rect 441706 155864 441712 155876
rect 441764 155864 441770 155916
rect 188430 155184 188436 155236
rect 188488 155224 188494 155236
rect 198182 155224 198188 155236
rect 188488 155196 198188 155224
rect 188488 155184 188494 155196
rect 198182 155184 198188 155196
rect 198240 155184 198246 155236
rect 372154 155184 372160 155236
rect 372212 155224 372218 155236
rect 444558 155224 444564 155236
rect 372212 155196 444564 155224
rect 372212 155184 372218 155196
rect 444558 155184 444564 155196
rect 444616 155184 444622 155236
rect 171226 154504 171232 154556
rect 171284 154544 171290 154556
rect 196802 154544 196808 154556
rect 171284 154516 196808 154544
rect 171284 154504 171290 154516
rect 196802 154504 196808 154516
rect 196860 154504 196866 154556
rect 302786 154504 302792 154556
rect 302844 154544 302850 154556
rect 370038 154544 370044 154556
rect 302844 154516 370044 154544
rect 302844 154504 302850 154516
rect 370038 154504 370044 154516
rect 370096 154544 370102 154556
rect 370590 154544 370596 154556
rect 370096 154516 370596 154544
rect 370096 154504 370102 154516
rect 370590 154504 370596 154516
rect 370648 154504 370654 154556
rect 371694 154504 371700 154556
rect 371752 154544 371758 154556
rect 382366 154544 382372 154556
rect 371752 154516 382372 154544
rect 371752 154504 371758 154516
rect 382366 154504 382372 154516
rect 382424 154504 382430 154556
rect 445662 154504 445668 154556
rect 445720 154544 445726 154556
rect 454218 154544 454224 154556
rect 445720 154516 454224 154544
rect 445720 154504 445726 154516
rect 454218 154504 454224 154516
rect 454276 154504 454282 154556
rect 171594 153960 171600 154012
rect 171652 154000 171658 154012
rect 180242 154000 180248 154012
rect 171652 153972 180248 154000
rect 171652 153960 171658 153972
rect 180242 153960 180248 153972
rect 180300 153960 180306 154012
rect 370130 153824 370136 153876
rect 370188 153864 370194 153876
rect 444926 153864 444932 153876
rect 370188 153836 444932 153864
rect 370188 153824 370194 153836
rect 444926 153824 444932 153836
rect 444984 153864 444990 153876
rect 451458 153864 451464 153876
rect 444984 153836 451464 153864
rect 444984 153824 444990 153836
rect 451458 153824 451464 153836
rect 451516 153824 451522 153876
rect 437382 153552 437388 153604
rect 437440 153592 437446 153604
rect 441890 153592 441896 153604
rect 437440 153564 441896 153592
rect 437440 153552 437446 153564
rect 441890 153552 441896 153564
rect 441948 153552 441954 153604
rect 371694 153348 371700 153400
rect 371752 153388 371758 153400
rect 374454 153388 374460 153400
rect 371752 153360 374460 153388
rect 371752 153348 371758 153360
rect 374454 153348 374460 153360
rect 374512 153348 374518 153400
rect 172422 153144 172428 153196
rect 172480 153184 172486 153196
rect 195422 153184 195428 153196
rect 172480 153156 195428 153184
rect 172480 153144 172486 153156
rect 195422 153144 195428 153156
rect 195480 153144 195486 153196
rect 302970 153144 302976 153196
rect 303028 153184 303034 153196
rect 369762 153184 369768 153196
rect 303028 153156 369768 153184
rect 303028 153144 303034 153156
rect 369762 153144 369768 153156
rect 369820 153144 369826 153196
rect 371510 153144 371516 153196
rect 371568 153184 371574 153196
rect 379514 153184 379520 153196
rect 371568 153156 379520 153184
rect 371568 153144 371574 153156
rect 379514 153144 379520 153156
rect 379572 153144 379578 153196
rect 443638 153144 443644 153196
rect 443696 153184 443702 153196
rect 580166 153184 580172 153196
rect 443696 153156 580172 153184
rect 443696 153144 443702 153156
rect 580166 153144 580172 153156
rect 580224 153144 580230 153196
rect 172330 153076 172336 153128
rect 172388 153116 172394 153128
rect 191282 153116 191288 153128
rect 172388 153088 191288 153116
rect 172388 153076 172394 153088
rect 191282 153076 191288 153088
rect 191340 153076 191346 153128
rect 302878 153076 302884 153128
rect 302936 153116 302942 153128
rect 369670 153116 369676 153128
rect 302936 153088 369676 153116
rect 302936 153076 302942 153088
rect 369670 153076 369676 153088
rect 369728 153076 369734 153128
rect 371694 153076 371700 153128
rect 371752 153116 371758 153128
rect 377122 153116 377128 153128
rect 371752 153088 377128 153116
rect 371752 153076 371758 153088
rect 377122 153076 377128 153088
rect 377180 153076 377186 153128
rect 302786 153008 302792 153060
rect 302844 153048 302850 153060
rect 369578 153048 369584 153060
rect 302844 153020 369584 153048
rect 302844 153008 302850 153020
rect 369578 153008 369584 153020
rect 369636 153008 369642 153060
rect 369670 152736 369676 152788
rect 369728 152776 369734 152788
rect 369946 152776 369952 152788
rect 369728 152748 369952 152776
rect 369728 152736 369734 152748
rect 369946 152736 369952 152748
rect 370004 152736 370010 152788
rect 302694 152464 302700 152516
rect 302752 152504 302758 152516
rect 369210 152504 369216 152516
rect 302752 152476 369216 152504
rect 302752 152464 302758 152476
rect 369210 152464 369216 152476
rect 369268 152464 369274 152516
rect 369578 152464 369584 152516
rect 369636 152504 369642 152516
rect 370314 152504 370320 152516
rect 369636 152476 370320 152504
rect 369636 152464 369642 152476
rect 370314 152464 370320 152476
rect 370372 152464 370378 152516
rect 359366 151988 359372 152040
rect 359424 152028 359430 152040
rect 369302 152028 369308 152040
rect 359424 152000 369308 152028
rect 359424 151988 359430 152000
rect 369302 151988 369308 152000
rect 369360 151988 369366 152040
rect 359550 151920 359556 151972
rect 359608 151960 359614 151972
rect 369118 151960 369124 151972
rect 359608 151932 369124 151960
rect 359608 151920 359614 151932
rect 369118 151920 369124 151932
rect 369176 151960 369182 151972
rect 369854 151960 369860 151972
rect 369176 151932 369860 151960
rect 369176 151920 369182 151932
rect 369854 151920 369860 151932
rect 369912 151920 369918 151972
rect 358998 151852 359004 151904
rect 359056 151892 359062 151904
rect 369486 151892 369492 151904
rect 359056 151864 369492 151892
rect 359056 151852 359062 151864
rect 369486 151852 369492 151864
rect 369544 151852 369550 151904
rect 444834 151852 444840 151904
rect 444892 151892 444898 151904
rect 452746 151892 452752 151904
rect 444892 151864 452752 151892
rect 444892 151852 444898 151864
rect 452746 151852 452752 151864
rect 452804 151852 452810 151904
rect 371694 151716 371700 151768
rect 371752 151756 371758 151768
rect 381170 151756 381176 151768
rect 371752 151728 381176 151756
rect 371752 151716 371758 151728
rect 381170 151716 381176 151728
rect 381228 151716 381234 151768
rect 172330 151648 172336 151700
rect 172388 151688 172394 151700
rect 187142 151688 187148 151700
rect 172388 151660 187148 151688
rect 172388 151648 172394 151660
rect 187142 151648 187148 151660
rect 187200 151648 187206 151700
rect 371510 151648 371516 151700
rect 371568 151688 371574 151700
rect 380986 151688 380992 151700
rect 371568 151660 380992 151688
rect 371568 151648 371574 151660
rect 380986 151648 380992 151660
rect 381044 151648 381050 151700
rect 172422 151580 172428 151632
rect 172480 151620 172486 151632
rect 188522 151620 188528 151632
rect 172480 151592 188528 151620
rect 172480 151580 172486 151592
rect 188522 151580 188528 151592
rect 188580 151580 188586 151632
rect 444834 151308 444840 151360
rect 444892 151348 444898 151360
rect 447502 151348 447508 151360
rect 444892 151320 447508 151348
rect 444892 151308 444898 151320
rect 447502 151308 447508 151320
rect 447560 151308 447566 151360
rect 187050 151036 187056 151088
rect 187108 151076 187114 151088
rect 198274 151076 198280 151088
rect 187108 151048 198280 151076
rect 187108 151036 187114 151048
rect 198274 151036 198280 151048
rect 198332 151036 198338 151088
rect 371694 151036 371700 151088
rect 371752 151076 371758 151088
rect 375558 151076 375564 151088
rect 371752 151048 375564 151076
rect 371752 151036 371758 151048
rect 375558 151036 375564 151048
rect 375616 151036 375622 151088
rect 196710 150560 196716 150612
rect 196768 150600 196774 150612
rect 198366 150600 198372 150612
rect 196768 150572 198372 150600
rect 196768 150560 196774 150572
rect 198366 150560 198372 150572
rect 198424 150560 198430 150612
rect 171870 150492 171876 150544
rect 171928 150532 171934 150544
rect 173158 150532 173164 150544
rect 171928 150504 173164 150532
rect 171928 150492 171934 150504
rect 173158 150492 173164 150504
rect 173216 150492 173222 150544
rect 3418 150356 3424 150408
rect 3476 150396 3482 150408
rect 11698 150396 11704 150408
rect 3476 150368 11704 150396
rect 3476 150356 3482 150368
rect 11698 150356 11704 150368
rect 11756 150356 11762 150408
rect 302786 150356 302792 150408
rect 302844 150396 302850 150408
rect 359366 150396 359372 150408
rect 302844 150368 359372 150396
rect 302844 150356 302850 150368
rect 359366 150356 359372 150368
rect 359424 150356 359430 150408
rect 371694 150356 371700 150408
rect 371752 150396 371758 150408
rect 378410 150396 378416 150408
rect 371752 150368 378416 150396
rect 371752 150356 371758 150368
rect 378410 150356 378416 150368
rect 378468 150356 378474 150408
rect 371510 150288 371516 150340
rect 371568 150328 371574 150340
rect 377030 150328 377036 150340
rect 371568 150300 377036 150328
rect 371568 150288 371574 150300
rect 377030 150288 377036 150300
rect 377088 150288 377094 150340
rect 171502 150016 171508 150068
rect 171560 150056 171566 150068
rect 173250 150056 173256 150068
rect 171560 150028 173256 150056
rect 171560 150016 171566 150028
rect 173250 150016 173256 150028
rect 173308 150016 173314 150068
rect 171686 149404 171692 149456
rect 171744 149444 171750 149456
rect 173342 149444 173348 149456
rect 171744 149416 173348 149444
rect 171744 149404 171750 149416
rect 173342 149404 173348 149416
rect 173400 149404 173406 149456
rect 171686 148996 171692 149048
rect 171744 149036 171750 149048
rect 173526 149036 173532 149048
rect 171744 149008 173532 149036
rect 171744 148996 171750 149008
rect 173526 148996 173532 149008
rect 173584 148996 173590 149048
rect 371694 148996 371700 149048
rect 371752 149036 371758 149048
rect 378318 149036 378324 149048
rect 371752 149008 378324 149036
rect 371752 148996 371758 149008
rect 378318 148996 378324 149008
rect 378376 148996 378382 149048
rect 171870 148860 171876 148912
rect 171928 148900 171934 148912
rect 173434 148900 173440 148912
rect 171928 148872 173440 148900
rect 171928 148860 171934 148872
rect 173434 148860 173440 148872
rect 173492 148860 173498 148912
rect 445294 148860 445300 148912
rect 445352 148900 445358 148912
rect 448882 148900 448888 148912
rect 445352 148872 448888 148900
rect 445352 148860 445358 148872
rect 448882 148860 448888 148872
rect 448940 148860 448946 148912
rect 371694 148384 371700 148436
rect 371752 148424 371758 148436
rect 374822 148424 374828 148436
rect 371752 148396 374828 148424
rect 371752 148384 371758 148396
rect 374822 148384 374828 148396
rect 374880 148384 374886 148436
rect 173158 148316 173164 148368
rect 173216 148356 173222 148368
rect 197998 148356 198004 148368
rect 173216 148328 198004 148356
rect 173216 148316 173222 148328
rect 197998 148316 198004 148328
rect 198056 148316 198062 148368
rect 171686 148180 171692 148232
rect 171744 148220 171750 148232
rect 173618 148220 173624 148232
rect 171744 148192 173624 148220
rect 171744 148180 171750 148192
rect 173618 148180 173624 148192
rect 173676 148180 173682 148232
rect 371694 148180 371700 148232
rect 371752 148220 371758 148232
rect 375650 148220 375656 148232
rect 371752 148192 375656 148220
rect 371752 148180 371758 148192
rect 375650 148180 375656 148192
rect 375708 148180 375714 148232
rect 445570 148112 445576 148164
rect 445628 148152 445634 148164
rect 450170 148152 450176 148164
rect 445628 148124 450176 148152
rect 445628 148112 445634 148124
rect 450170 148112 450176 148124
rect 450228 148112 450234 148164
rect 195238 147636 195244 147688
rect 195296 147676 195302 147688
rect 198274 147676 198280 147688
rect 195296 147648 198280 147676
rect 195296 147636 195302 147648
rect 198274 147636 198280 147648
rect 198332 147636 198338 147688
rect 172422 147568 172428 147620
rect 172480 147608 172486 147620
rect 196894 147608 196900 147620
rect 172480 147580 196900 147608
rect 172480 147568 172486 147580
rect 196894 147568 196900 147580
rect 196952 147568 196958 147620
rect 171870 147500 171876 147552
rect 171928 147540 171934 147552
rect 176010 147540 176016 147552
rect 171928 147512 176016 147540
rect 171928 147500 171934 147512
rect 176010 147500 176016 147512
rect 176068 147500 176074 147552
rect 371234 147500 371240 147552
rect 371292 147540 371298 147552
rect 378226 147540 378232 147552
rect 371292 147512 378232 147540
rect 371292 147500 371298 147512
rect 378226 147500 378232 147512
rect 378284 147500 378290 147552
rect 371234 146684 371240 146736
rect 371292 146724 371298 146736
rect 373350 146724 373356 146736
rect 371292 146696 373356 146724
rect 371292 146684 371298 146696
rect 373350 146684 373356 146696
rect 373408 146684 373414 146736
rect 444834 146548 444840 146600
rect 444892 146588 444898 146600
rect 446122 146588 446128 146600
rect 444892 146560 446128 146588
rect 444892 146548 444898 146560
rect 446122 146548 446128 146560
rect 446180 146548 446186 146600
rect 191190 146480 191196 146532
rect 191248 146520 191254 146532
rect 197722 146520 197728 146532
rect 191248 146492 197728 146520
rect 191248 146480 191254 146492
rect 197722 146480 197728 146492
rect 197780 146480 197786 146532
rect 172330 146208 172336 146260
rect 172388 146248 172394 146260
rect 182910 146248 182916 146260
rect 172388 146220 182916 146248
rect 172388 146208 172394 146220
rect 182910 146208 182916 146220
rect 182968 146208 182974 146260
rect 302786 146208 302792 146260
rect 302844 146248 302850 146260
rect 358998 146248 359004 146260
rect 302844 146220 359004 146248
rect 302844 146208 302850 146220
rect 358998 146208 359004 146220
rect 359056 146208 359062 146260
rect 172422 146140 172428 146192
rect 172480 146180 172486 146192
rect 181530 146180 181536 146192
rect 172480 146152 181536 146180
rect 172480 146140 172486 146152
rect 181530 146140 181536 146152
rect 181588 146140 181594 146192
rect 371510 146140 371516 146192
rect 371568 146180 371574 146192
rect 376846 146180 376852 146192
rect 371568 146152 376852 146180
rect 371568 146140 371574 146152
rect 376846 146140 376852 146152
rect 376904 146140 376910 146192
rect 172238 146072 172244 146124
rect 172296 146112 172302 146124
rect 178862 146112 178868 146124
rect 172296 146084 178868 146112
rect 172296 146072 172302 146084
rect 178862 146072 178868 146084
rect 178920 146072 178926 146124
rect 371694 146072 371700 146124
rect 371752 146112 371758 146124
rect 376754 146112 376760 146124
rect 371752 146084 376760 146112
rect 371752 146072 371758 146084
rect 376754 146072 376760 146084
rect 376812 146072 376818 146124
rect 445478 146004 445484 146056
rect 445536 146044 445542 146056
rect 449986 146044 449992 146056
rect 445536 146016 449992 146044
rect 445536 146004 445542 146016
rect 449986 146004 449992 146016
rect 450044 146004 450050 146056
rect 371694 145052 371700 145104
rect 371752 145092 371758 145104
rect 374914 145092 374920 145104
rect 371752 145064 374920 145092
rect 371752 145052 371758 145064
rect 374914 145052 374920 145064
rect 374972 145052 374978 145104
rect 172422 144848 172428 144900
rect 172480 144888 172486 144900
rect 188430 144888 188436 144900
rect 172480 144860 188436 144888
rect 172480 144848 172486 144860
rect 188430 144848 188436 144860
rect 188488 144848 188494 144900
rect 371510 144848 371516 144900
rect 371568 144888 371574 144900
rect 383746 144888 383752 144900
rect 371568 144860 383752 144888
rect 371568 144848 371574 144860
rect 383746 144848 383752 144860
rect 383804 144848 383810 144900
rect 372062 144780 372068 144832
rect 372120 144820 372126 144832
rect 382274 144820 382280 144832
rect 372120 144792 382280 144820
rect 372120 144780 372126 144792
rect 382274 144780 382280 144792
rect 382332 144780 382338 144832
rect 445110 144712 445116 144764
rect 445168 144752 445174 144764
rect 448698 144752 448704 144764
rect 445168 144724 448704 144752
rect 445168 144712 445174 144724
rect 448698 144712 448704 144724
rect 448756 144712 448762 144764
rect 371694 144508 371700 144560
rect 371752 144548 371758 144560
rect 375834 144548 375840 144560
rect 371752 144520 375840 144548
rect 371752 144508 371758 144520
rect 375834 144508 375840 144520
rect 375892 144508 375898 144560
rect 171686 144168 171692 144220
rect 171744 144208 171750 144220
rect 188338 144208 188344 144220
rect 171744 144180 188344 144208
rect 171744 144168 171750 144180
rect 188338 144168 188344 144180
rect 188396 144168 188402 144220
rect 188522 143556 188528 143608
rect 188580 143596 188586 143608
rect 197354 143596 197360 143608
rect 188580 143568 197360 143596
rect 188580 143556 188586 143568
rect 197354 143556 197360 143568
rect 197412 143556 197418 143608
rect 171870 143488 171876 143540
rect 171928 143528 171934 143540
rect 180334 143528 180340 143540
rect 171928 143500 180340 143528
rect 171928 143488 171934 143500
rect 180334 143488 180340 143500
rect 180392 143488 180398 143540
rect 302786 143488 302792 143540
rect 302844 143528 302850 143540
rect 359550 143528 359556 143540
rect 302844 143500 359556 143528
rect 302844 143488 302850 143500
rect 359550 143488 359556 143500
rect 359608 143488 359614 143540
rect 371234 143488 371240 143540
rect 371292 143528 371298 143540
rect 379606 143528 379612 143540
rect 371292 143500 379612 143528
rect 371292 143488 371298 143500
rect 379606 143488 379612 143500
rect 379664 143488 379670 143540
rect 371694 143420 371700 143472
rect 371752 143460 371758 143472
rect 376938 143460 376944 143472
rect 371752 143432 376944 143460
rect 371752 143420 371758 143432
rect 376938 143420 376944 143432
rect 376996 143420 377002 143472
rect 445110 143148 445116 143200
rect 445168 143188 445174 143200
rect 450078 143188 450084 143200
rect 445168 143160 450084 143188
rect 445168 143148 445174 143160
rect 450078 143148 450084 143160
rect 450136 143148 450142 143200
rect 171778 142808 171784 142860
rect 171836 142848 171842 142860
rect 186958 142848 186964 142860
rect 171836 142820 186964 142848
rect 171836 142808 171842 142820
rect 186958 142808 186964 142820
rect 187016 142808 187022 142860
rect 171502 142264 171508 142316
rect 171560 142304 171566 142316
rect 174538 142304 174544 142316
rect 171560 142276 174544 142304
rect 171560 142264 171566 142276
rect 174538 142264 174544 142276
rect 174596 142264 174602 142316
rect 187142 142128 187148 142180
rect 187200 142168 187206 142180
rect 197354 142168 197360 142180
rect 187200 142140 197360 142168
rect 187200 142128 187206 142140
rect 197354 142128 197360 142140
rect 197412 142128 197418 142180
rect 172422 142060 172428 142112
rect 172480 142100 172486 142112
rect 195330 142100 195336 142112
rect 172480 142072 195336 142100
rect 172480 142060 172486 142072
rect 195330 142060 195336 142072
rect 195388 142060 195394 142112
rect 371510 142060 371516 142112
rect 371568 142100 371574 142112
rect 382458 142100 382464 142112
rect 371568 142072 382464 142100
rect 371568 142060 371574 142072
rect 382458 142060 382464 142072
rect 382516 142060 382522 142112
rect 444374 142060 444380 142112
rect 444432 142100 444438 142112
rect 444834 142100 444840 142112
rect 444432 142072 444840 142100
rect 444432 142060 444438 142072
rect 444834 142060 444840 142072
rect 444892 142060 444898 142112
rect 371234 141992 371240 142044
rect 371292 142032 371298 142044
rect 380894 142032 380900 142044
rect 371292 142004 380900 142032
rect 371292 141992 371298 142004
rect 380894 141992 380900 142004
rect 380952 141992 380958 142044
rect 371694 141924 371700 141976
rect 371752 141964 371758 141976
rect 375742 141964 375748 141976
rect 371752 141936 375748 141964
rect 371752 141924 371758 141936
rect 375742 141924 375748 141936
rect 375800 141924 375806 141976
rect 444374 141924 444380 141976
rect 444432 141964 444438 141976
rect 447318 141964 447324 141976
rect 444432 141936 447324 141964
rect 444432 141924 444438 141936
rect 447318 141924 447324 141936
rect 447376 141924 447382 141976
rect 171686 141380 171692 141432
rect 171744 141420 171750 141432
rect 191098 141420 191104 141432
rect 171744 141392 191104 141420
rect 171744 141380 171750 141392
rect 191098 141380 191104 141392
rect 191156 141380 191162 141432
rect 371694 140632 371700 140684
rect 371752 140672 371758 140684
rect 378134 140672 378140 140684
rect 371752 140644 378140 140672
rect 371752 140632 371758 140644
rect 378134 140632 378140 140644
rect 378192 140632 378198 140684
rect 444374 140428 444380 140480
rect 444432 140468 444438 140480
rect 446030 140468 446036 140480
rect 444432 140440 446036 140468
rect 444432 140428 444438 140440
rect 446030 140428 446036 140440
rect 446088 140428 446094 140480
rect 172330 140020 172336 140072
rect 172388 140060 172394 140072
rect 198090 140060 198096 140072
rect 172388 140032 198096 140060
rect 172388 140020 172394 140032
rect 198090 140020 198096 140032
rect 198148 140020 198154 140072
rect 171686 139748 171692 139800
rect 171744 139788 171750 139800
rect 173158 139788 173164 139800
rect 171744 139760 173164 139788
rect 171744 139748 171750 139760
rect 173158 139748 173164 139760
rect 173216 139748 173222 139800
rect 172422 139340 172428 139392
rect 172480 139380 172486 139392
rect 184290 139380 184296 139392
rect 172480 139352 184296 139380
rect 172480 139340 172486 139352
rect 184290 139340 184296 139352
rect 184348 139340 184354 139392
rect 371510 139340 371516 139392
rect 371568 139380 371574 139392
rect 374270 139380 374276 139392
rect 371568 139352 374276 139380
rect 371568 139340 371574 139352
rect 374270 139340 374276 139352
rect 374328 139340 374334 139392
rect 465718 139340 465724 139392
rect 465776 139380 465782 139392
rect 580166 139380 580172 139392
rect 465776 139352 580172 139380
rect 465776 139340 465782 139352
rect 580166 139340 580172 139352
rect 580224 139340 580230 139392
rect 371694 139204 371700 139256
rect 371752 139244 371758 139256
rect 375374 139244 375380 139256
rect 371752 139216 375380 139244
rect 371752 139204 371758 139216
rect 375374 139204 375380 139216
rect 375432 139204 375438 139256
rect 171594 139068 171600 139120
rect 171652 139108 171658 139120
rect 180058 139108 180064 139120
rect 171652 139080 180064 139108
rect 171652 139068 171658 139080
rect 180058 139068 180064 139080
rect 180116 139068 180122 139120
rect 371694 138864 371700 138916
rect 371752 138904 371758 138916
rect 374086 138904 374092 138916
rect 371752 138876 374092 138904
rect 371752 138864 371758 138876
rect 374086 138864 374092 138876
rect 374144 138864 374150 138916
rect 444374 138592 444380 138644
rect 444432 138632 444438 138644
rect 447226 138632 447232 138644
rect 444432 138604 447232 138632
rect 444432 138592 444438 138604
rect 447226 138592 447232 138604
rect 447284 138592 447290 138644
rect 171502 138184 171508 138236
rect 171560 138224 171566 138236
rect 177390 138224 177396 138236
rect 171560 138196 177396 138224
rect 171560 138184 171566 138196
rect 177390 138184 177396 138196
rect 177448 138184 177454 138236
rect 3234 137912 3240 137964
rect 3292 137952 3298 137964
rect 152458 137952 152464 137964
rect 3292 137924 152464 137952
rect 3292 137912 3298 137924
rect 152458 137912 152464 137924
rect 152516 137912 152522 137964
rect 172054 137912 172060 137964
rect 172112 137952 172118 137964
rect 187050 137952 187056 137964
rect 172112 137924 187056 137952
rect 172112 137912 172118 137924
rect 187050 137912 187056 137924
rect 187108 137912 187114 137964
rect 444374 137300 444380 137352
rect 444432 137340 444438 137352
rect 447410 137340 447416 137352
rect 444432 137312 447416 137340
rect 444432 137300 444438 137312
rect 447410 137300 447416 137312
rect 447468 137300 447474 137352
rect 172422 137232 172428 137284
rect 172480 137272 172486 137284
rect 196710 137272 196716 137284
rect 172480 137244 196716 137272
rect 172480 137232 172486 137244
rect 196710 137232 196716 137244
rect 196768 137232 196774 137284
rect 172514 136620 172520 136672
rect 172572 136660 172578 136672
rect 197538 136660 197544 136672
rect 172572 136632 197544 136660
rect 172572 136620 172578 136632
rect 197538 136620 197544 136632
rect 197596 136620 197602 136672
rect 172238 136552 172244 136604
rect 172296 136592 172302 136604
rect 195238 136592 195244 136604
rect 172296 136564 195244 136592
rect 172296 136552 172302 136564
rect 195238 136552 195244 136564
rect 195296 136552 195302 136604
rect 171686 136484 171692 136536
rect 171744 136524 171750 136536
rect 191190 136524 191196 136536
rect 171744 136496 191196 136524
rect 171744 136484 171750 136496
rect 191190 136484 191196 136496
rect 191248 136484 191254 136536
rect 172330 135260 172336 135312
rect 172388 135300 172394 135312
rect 198090 135300 198096 135312
rect 172388 135272 198096 135300
rect 172388 135260 172394 135272
rect 198090 135260 198096 135272
rect 198148 135260 198154 135312
rect 171226 135192 171232 135244
rect 171284 135232 171290 135244
rect 198274 135232 198280 135244
rect 171284 135204 198280 135232
rect 171284 135192 171290 135204
rect 198274 135192 198280 135204
rect 198332 135192 198338 135244
rect 369210 135192 369216 135244
rect 369268 135232 369274 135244
rect 369394 135232 369400 135244
rect 369268 135204 369400 135232
rect 369268 135192 369274 135204
rect 369394 135192 369400 135204
rect 369452 135192 369458 135244
rect 172422 135124 172428 135176
rect 172480 135164 172486 135176
rect 188522 135164 188528 135176
rect 172480 135136 188528 135164
rect 172480 135124 172486 135136
rect 188522 135124 188528 135136
rect 188580 135124 188586 135176
rect 172238 135056 172244 135108
rect 172296 135096 172302 135108
rect 187142 135096 187148 135108
rect 172296 135068 187148 135096
rect 172296 135056 172302 135068
rect 187142 135056 187148 135068
rect 187200 135056 187206 135108
rect 171134 132472 171140 132524
rect 171192 132512 171198 132524
rect 197538 132512 197544 132524
rect 171192 132484 197544 132512
rect 171192 132472 171198 132484
rect 197538 132472 197544 132484
rect 197596 132472 197602 132524
rect 172422 131724 172428 131776
rect 172480 131764 172486 131776
rect 197906 131764 197912 131776
rect 172480 131736 197912 131764
rect 172480 131724 172486 131736
rect 197906 131724 197912 131736
rect 197964 131724 197970 131776
rect 370222 130636 370228 130688
rect 370280 130676 370286 130688
rect 373258 130676 373264 130688
rect 370280 130648 373264 130676
rect 370280 130636 370286 130648
rect 373258 130636 373264 130648
rect 373316 130636 373322 130688
rect 443914 130364 443920 130416
rect 443972 130404 443978 130416
rect 448514 130404 448520 130416
rect 443972 130376 448520 130404
rect 443972 130364 443978 130376
rect 448514 130364 448520 130376
rect 448572 130364 448578 130416
rect 171870 130024 171876 130076
rect 171928 130064 171934 130076
rect 179414 130064 179420 130076
rect 171928 130036 179420 130064
rect 171928 130024 171934 130036
rect 179414 130024 179420 130036
rect 179472 130024 179478 130076
rect 171502 129684 171508 129736
rect 171560 129724 171566 129736
rect 197354 129724 197360 129736
rect 171560 129696 197360 129724
rect 171560 129684 171566 129696
rect 197354 129684 197360 129696
rect 197412 129684 197418 129736
rect 369854 129072 369860 129124
rect 369912 129112 369918 129124
rect 373994 129112 374000 129124
rect 369912 129084 374000 129112
rect 369912 129072 369918 129084
rect 373994 129072 374000 129084
rect 374052 129112 374058 129124
rect 427814 129112 427820 129124
rect 374052 129084 427820 129112
rect 374052 129072 374058 129084
rect 427814 129072 427820 129084
rect 427872 129072 427878 129124
rect 370314 129004 370320 129056
rect 370372 129044 370378 129056
rect 371418 129044 371424 129056
rect 370372 129016 371424 129044
rect 370372 129004 370378 129016
rect 371418 129004 371424 129016
rect 371476 129044 371482 129056
rect 430574 129044 430580 129056
rect 371476 129016 430580 129044
rect 371476 129004 371482 129016
rect 430574 129004 430580 129016
rect 430632 129004 430638 129056
rect 443638 128324 443644 128376
rect 443696 128364 443702 128376
rect 452654 128364 452660 128376
rect 443696 128336 452660 128364
rect 443696 128324 443702 128336
rect 452654 128324 452660 128336
rect 452712 128324 452718 128376
rect 444374 128052 444380 128104
rect 444432 128092 444438 128104
rect 449894 128092 449900 128104
rect 444432 128064 449900 128092
rect 444432 128052 444438 128064
rect 449894 128052 449900 128064
rect 449952 128052 449958 128104
rect 172514 127576 172520 127628
rect 172572 127616 172578 127628
rect 197998 127616 198004 127628
rect 172572 127588 198004 127616
rect 172572 127576 172578 127588
rect 197998 127576 198004 127588
rect 198056 127576 198062 127628
rect 172330 126896 172336 126948
rect 172388 126936 172394 126948
rect 197354 126936 197360 126948
rect 172388 126908 197360 126936
rect 172388 126896 172394 126908
rect 197354 126896 197360 126908
rect 197412 126896 197418 126948
rect 449158 126896 449164 126948
rect 449216 126936 449222 126948
rect 580166 126936 580172 126948
rect 449216 126908 580172 126936
rect 449216 126896 449222 126908
rect 580166 126896 580172 126908
rect 580224 126896 580230 126948
rect 444374 126624 444380 126676
rect 444432 126664 444438 126676
rect 447134 126664 447140 126676
rect 444432 126636 447140 126664
rect 444432 126624 444438 126636
rect 447134 126624 447140 126636
rect 447192 126624 447198 126676
rect 372430 126012 372436 126064
rect 372488 126052 372494 126064
rect 443086 126052 443092 126064
rect 372488 126024 443092 126052
rect 372488 126012 372494 126024
rect 443086 126012 443092 126024
rect 443144 126012 443150 126064
rect 371786 125944 371792 125996
rect 371844 125984 371850 125996
rect 442994 125984 443000 125996
rect 371844 125956 443000 125984
rect 371844 125944 371850 125956
rect 442994 125944 443000 125956
rect 443052 125944 443058 125996
rect 370406 125876 370412 125928
rect 370464 125916 370470 125928
rect 371602 125916 371608 125928
rect 370464 125888 371608 125916
rect 370464 125876 370470 125888
rect 371602 125876 371608 125888
rect 371660 125916 371666 125928
rect 443638 125916 443644 125928
rect 371660 125888 443644 125916
rect 371660 125876 371666 125888
rect 443638 125876 443644 125888
rect 443696 125876 443702 125928
rect 172422 125740 172428 125792
rect 172480 125780 172486 125792
rect 186958 125780 186964 125792
rect 172480 125752 186964 125780
rect 172480 125740 172486 125752
rect 186958 125740 186964 125752
rect 187016 125740 187022 125792
rect 172330 125672 172336 125724
rect 172388 125712 172394 125724
rect 188338 125712 188344 125724
rect 172388 125684 188344 125712
rect 172388 125672 172394 125684
rect 188338 125672 188344 125684
rect 188396 125672 188402 125724
rect 172238 125604 172244 125656
rect 172296 125644 172302 125656
rect 191098 125644 191104 125656
rect 172296 125616 191104 125644
rect 172296 125604 172302 125616
rect 191098 125604 191104 125616
rect 191156 125604 191162 125656
rect 179414 125536 179420 125588
rect 179472 125576 179478 125588
rect 198550 125576 198556 125588
rect 179472 125548 198556 125576
rect 179472 125536 179478 125548
rect 198550 125536 198556 125548
rect 198608 125536 198614 125588
rect 370498 125468 370504 125520
rect 370556 125508 370562 125520
rect 372614 125508 372620 125520
rect 370556 125480 372620 125508
rect 370556 125468 370562 125480
rect 372614 125468 372620 125480
rect 372672 125508 372678 125520
rect 441614 125508 441620 125520
rect 372672 125480 441620 125508
rect 372672 125468 372678 125480
rect 441614 125468 441620 125480
rect 441672 125468 441678 125520
rect 427814 125400 427820 125452
rect 427872 125440 427878 125452
rect 444742 125440 444748 125452
rect 427872 125412 444748 125440
rect 427872 125400 427878 125412
rect 444742 125400 444748 125412
rect 444800 125400 444806 125452
rect 430574 125332 430580 125384
rect 430632 125372 430638 125384
rect 444834 125372 444840 125384
rect 430632 125344 444840 125372
rect 430632 125332 430638 125344
rect 444834 125332 444840 125344
rect 444892 125332 444898 125384
rect 371326 125264 371332 125316
rect 371384 125304 371390 125316
rect 441890 125304 441896 125316
rect 371384 125276 441896 125304
rect 371384 125264 371390 125276
rect 441890 125264 441896 125276
rect 441948 125264 441954 125316
rect 302786 125196 302792 125248
rect 302844 125236 302850 125248
rect 370314 125236 370320 125248
rect 302844 125208 370320 125236
rect 302844 125196 302850 125208
rect 370314 125196 370320 125208
rect 370372 125196 370378 125248
rect 303062 125128 303068 125180
rect 303120 125168 303126 125180
rect 369854 125168 369860 125180
rect 303120 125140 369860 125168
rect 303120 125128 303126 125140
rect 369854 125128 369860 125140
rect 369912 125128 369918 125180
rect 302878 125060 302884 125112
rect 302936 125100 302942 125112
rect 370222 125100 370228 125112
rect 302936 125072 370228 125100
rect 302936 125060 302942 125072
rect 370222 125060 370228 125072
rect 370280 125060 370286 125112
rect 302970 124992 302976 125044
rect 303028 125032 303034 125044
rect 369946 125032 369952 125044
rect 303028 125004 369952 125032
rect 303028 124992 303034 125004
rect 369946 124992 369952 125004
rect 370004 124992 370010 125044
rect 302602 124924 302608 124976
rect 302660 124964 302666 124976
rect 370038 124964 370044 124976
rect 302660 124936 370044 124964
rect 302660 124924 302666 124936
rect 370038 124924 370044 124936
rect 370096 124924 370102 124976
rect 370774 124856 370780 124908
rect 370832 124896 370838 124908
rect 441890 124896 441896 124908
rect 370832 124868 441896 124896
rect 370832 124856 370838 124868
rect 441890 124856 441896 124868
rect 441948 124896 441954 124908
rect 445846 124896 445852 124908
rect 441948 124868 445852 124896
rect 441948 124856 441954 124868
rect 445846 124856 445852 124868
rect 445904 124856 445910 124908
rect 172422 124312 172428 124364
rect 172480 124352 172486 124364
rect 184198 124352 184204 124364
rect 172480 124324 184204 124352
rect 172480 124312 172486 124324
rect 184198 124312 184204 124324
rect 184256 124312 184262 124364
rect 171686 124244 171692 124296
rect 171744 124284 171750 124296
rect 180058 124284 180064 124296
rect 171744 124256 180064 124284
rect 171744 124244 171750 124256
rect 180058 124244 180064 124256
rect 180116 124244 180122 124296
rect 172146 124176 172152 124228
rect 172204 124216 172210 124228
rect 173158 124216 173164 124228
rect 172204 124188 173164 124216
rect 172204 124176 172210 124188
rect 173158 124176 173164 124188
rect 173216 124176 173222 124228
rect 302694 124108 302700 124160
rect 302752 124148 302758 124160
rect 371234 124148 371240 124160
rect 302752 124120 371240 124148
rect 302752 124108 302758 124120
rect 371234 124108 371240 124120
rect 371292 124108 371298 124160
rect 302970 123564 302976 123616
rect 303028 123604 303034 123616
rect 370406 123604 370412 123616
rect 303028 123576 370412 123604
rect 303028 123564 303034 123576
rect 370406 123564 370412 123576
rect 370464 123564 370470 123616
rect 302878 123428 302884 123480
rect 302936 123468 302942 123480
rect 369946 123468 369952 123480
rect 302936 123440 369952 123468
rect 302936 123428 302942 123440
rect 369946 123428 369952 123440
rect 370004 123428 370010 123480
rect 160922 122952 160928 123004
rect 160980 122992 160986 123004
rect 170490 122992 170496 123004
rect 160980 122964 170496 122992
rect 160980 122952 160986 122964
rect 170490 122952 170496 122964
rect 170548 122952 170554 123004
rect 162854 122884 162860 122936
rect 162912 122924 162918 122936
rect 193858 122924 193864 122936
rect 162912 122896 193864 122924
rect 162912 122884 162918 122896
rect 193858 122884 193864 122896
rect 193916 122884 193922 122936
rect 164878 122816 164884 122868
rect 164936 122856 164942 122868
rect 198734 122856 198740 122868
rect 164936 122828 198740 122856
rect 164936 122816 164942 122828
rect 198734 122816 198740 122828
rect 198792 122816 198798 122868
rect 166902 122748 166908 122800
rect 166960 122788 166966 122800
rect 178678 122788 178684 122800
rect 166960 122760 178684 122788
rect 166960 122748 166966 122760
rect 178678 122748 178684 122760
rect 178736 122748 178742 122800
rect 320818 122748 320824 122800
rect 320876 122788 320882 122800
rect 438854 122788 438860 122800
rect 320876 122760 438860 122788
rect 320876 122748 320882 122760
rect 438854 122748 438860 122760
rect 438912 122748 438918 122800
rect 168926 122680 168932 122732
rect 168984 122720 168990 122732
rect 177298 122720 177304 122732
rect 168984 122692 177304 122720
rect 168984 122680 168990 122692
rect 177298 122680 177304 122692
rect 177356 122680 177362 122732
rect 359458 122680 359464 122732
rect 359516 122720 359522 122732
rect 366910 122720 366916 122732
rect 359516 122692 366916 122720
rect 359516 122680 359522 122692
rect 366910 122680 366916 122692
rect 366968 122680 366974 122732
rect 437198 122680 437204 122732
rect 437256 122720 437262 122732
rect 441798 122720 441804 122732
rect 437256 122692 441804 122720
rect 437256 122680 437262 122692
rect 441798 122680 441804 122692
rect 441856 122680 441862 122732
rect 435174 122612 435180 122664
rect 435232 122652 435238 122664
rect 441706 122652 441712 122664
rect 435232 122624 441712 122652
rect 435232 122612 435238 122624
rect 441706 122612 441712 122624
rect 441764 122612 441770 122664
rect 172054 121388 172060 121440
rect 172112 121428 172118 121440
rect 197538 121428 197544 121440
rect 172112 121400 197544 121428
rect 172112 121388 172118 121400
rect 197538 121388 197544 121400
rect 197596 121388 197602 121440
rect 302786 121388 302792 121440
rect 302844 121428 302850 121440
rect 370130 121428 370136 121440
rect 302844 121400 370136 121428
rect 302844 121388 302850 121400
rect 370130 121388 370136 121400
rect 370188 121388 370194 121440
rect 188338 119348 188344 119400
rect 188396 119388 188402 119400
rect 197998 119388 198004 119400
rect 188396 119360 198004 119388
rect 188396 119348 188402 119360
rect 197998 119348 198004 119360
rect 198056 119348 198062 119400
rect 171870 118600 171876 118652
rect 171928 118640 171934 118652
rect 198090 118640 198096 118652
rect 171928 118612 198096 118640
rect 171928 118600 171934 118612
rect 198090 118600 198096 118612
rect 198148 118600 198154 118652
rect 302786 118600 302792 118652
rect 302844 118640 302850 118652
rect 371786 118640 371792 118652
rect 302844 118612 371792 118640
rect 302844 118600 302850 118612
rect 371786 118600 371792 118612
rect 371844 118600 371850 118652
rect 171962 117240 171968 117292
rect 172020 117280 172026 117292
rect 197538 117280 197544 117292
rect 172020 117252 197544 117280
rect 172020 117240 172026 117252
rect 197538 117240 197544 117252
rect 197596 117240 197602 117292
rect 171778 114452 171784 114504
rect 171836 114492 171842 114504
rect 197354 114492 197360 114504
rect 171836 114464 197360 114492
rect 171836 114452 171842 114464
rect 197354 114452 197360 114464
rect 197412 114452 197418 114504
rect 313918 113092 313924 113144
rect 313976 113132 313982 113144
rect 579798 113132 579804 113144
rect 313976 113104 579804 113132
rect 313976 113092 313982 113104
rect 579798 113092 579804 113104
rect 579856 113092 579862 113144
rect 3418 111732 3424 111784
rect 3476 111772 3482 111784
rect 170398 111772 170404 111784
rect 3476 111744 170404 111772
rect 3476 111732 3482 111744
rect 170398 111732 170404 111744
rect 170456 111732 170462 111784
rect 191098 111732 191104 111784
rect 191156 111772 191162 111784
rect 197354 111772 197360 111784
rect 191156 111744 197360 111772
rect 191156 111732 191162 111744
rect 197354 111732 197360 111744
rect 197412 111732 197418 111784
rect 302326 111732 302332 111784
rect 302384 111772 302390 111784
rect 370590 111772 370596 111784
rect 302384 111744 370596 111772
rect 302384 111732 302390 111744
rect 370590 111732 370596 111744
rect 370648 111732 370654 111784
rect 302786 108944 302792 108996
rect 302844 108984 302850 108996
rect 371326 108984 371332 108996
rect 302844 108956 371332 108984
rect 302844 108944 302850 108956
rect 371326 108944 371332 108956
rect 371384 108944 371390 108996
rect 186958 107584 186964 107636
rect 187016 107624 187022 107636
rect 198550 107624 198556 107636
rect 187016 107596 198556 107624
rect 187016 107584 187022 107596
rect 198550 107584 198556 107596
rect 198608 107584 198614 107636
rect 184198 106224 184204 106276
rect 184256 106264 184262 106276
rect 197538 106264 197544 106276
rect 184256 106236 197544 106264
rect 184256 106224 184262 106236
rect 197538 106224 197544 106236
rect 197596 106224 197602 106276
rect 180058 103436 180064 103488
rect 180116 103476 180122 103488
rect 197906 103476 197912 103488
rect 180116 103448 197912 103476
rect 180116 103436 180122 103448
rect 197906 103436 197912 103448
rect 197964 103436 197970 103488
rect 173158 102076 173164 102128
rect 173216 102116 173222 102128
rect 197538 102116 197544 102128
rect 173216 102088 197544 102116
rect 173216 102076 173222 102088
rect 197538 102076 197544 102088
rect 197596 102076 197602 102128
rect 302786 102076 302792 102128
rect 302844 102116 302850 102128
rect 369854 102116 369860 102128
rect 302844 102088 369860 102116
rect 302844 102076 302850 102088
rect 369854 102076 369860 102088
rect 369912 102076 369918 102128
rect 457438 100648 457444 100700
rect 457496 100688 457502 100700
rect 580166 100688 580172 100700
rect 457496 100660 580172 100688
rect 457496 100648 457502 100660
rect 580166 100648 580172 100660
rect 580224 100648 580230 100700
rect 196618 99356 196624 99408
rect 196676 99396 196682 99408
rect 299474 99396 299480 99408
rect 196676 99368 299480 99396
rect 196676 99356 196682 99368
rect 299474 99356 299480 99368
rect 299532 99356 299538 99408
rect 112438 99288 112444 99340
rect 112496 99328 112502 99340
rect 217594 99328 217600 99340
rect 112496 99300 217600 99328
rect 112496 99288 112502 99300
rect 217594 99288 217600 99300
rect 217652 99288 217658 99340
rect 278866 99288 278872 99340
rect 278924 99328 278930 99340
rect 414658 99328 414664 99340
rect 278924 99300 414664 99328
rect 278924 99288 278930 99300
rect 414658 99288 414664 99300
rect 414716 99288 414722 99340
rect 98638 99220 98644 99272
rect 98696 99260 98702 99272
rect 213362 99260 213368 99272
rect 98696 99232 213368 99260
rect 98696 99220 98702 99232
rect 213362 99220 213368 99232
rect 213420 99220 213426 99272
rect 240502 99220 240508 99272
rect 240560 99260 240566 99272
rect 241054 99260 241060 99272
rect 240560 99232 241060 99260
rect 240560 99220 240566 99232
rect 241054 99220 241060 99232
rect 241112 99220 241118 99272
rect 271046 99220 271052 99272
rect 271104 99260 271110 99272
rect 413278 99260 413284 99272
rect 271104 99232 413284 99260
rect 271104 99220 271110 99232
rect 413278 99220 413284 99232
rect 413336 99220 413342 99272
rect 97258 99152 97264 99204
rect 97316 99192 97322 99204
rect 211522 99192 211528 99204
rect 97316 99164 211528 99192
rect 97316 99152 97322 99164
rect 211522 99152 211528 99164
rect 211580 99152 211586 99204
rect 271598 99152 271604 99204
rect 271656 99192 271662 99204
rect 417418 99192 417424 99204
rect 271656 99164 417424 99192
rect 271656 99152 271662 99164
rect 417418 99152 417424 99164
rect 417476 99152 417482 99204
rect 88978 99084 88984 99136
rect 89036 99124 89042 99136
rect 209774 99124 209780 99136
rect 89036 99096 209780 99124
rect 89036 99084 89042 99096
rect 209774 99084 209780 99096
rect 209832 99084 209838 99136
rect 272242 99084 272248 99136
rect 272300 99124 272306 99136
rect 421558 99124 421564 99136
rect 272300 99096 421564 99124
rect 272300 99084 272306 99096
rect 421558 99084 421564 99096
rect 421616 99084 421622 99136
rect 93118 99016 93124 99068
rect 93176 99056 93182 99068
rect 215386 99056 215392 99068
rect 93176 99028 215392 99056
rect 93176 99016 93182 99028
rect 215386 99016 215392 99028
rect 215444 99016 215450 99068
rect 273438 99016 273444 99068
rect 273496 99056 273502 99068
rect 430574 99056 430580 99068
rect 273496 99028 430580 99056
rect 273496 99016 273502 99028
rect 430574 99016 430580 99028
rect 430632 99016 430638 99068
rect 87598 98948 87604 99000
rect 87656 98988 87662 99000
rect 214374 98988 214380 99000
rect 87656 98960 214380 98988
rect 87656 98948 87662 98960
rect 214374 98948 214380 98960
rect 214432 98948 214438 99000
rect 274634 98948 274640 99000
rect 274692 98988 274698 99000
rect 435358 98988 435364 99000
rect 274692 98960 435364 98988
rect 274692 98948 274698 98960
rect 435358 98948 435364 98960
rect 435416 98948 435422 99000
rect 71038 98880 71044 98932
rect 71096 98920 71102 98932
rect 210326 98920 210332 98932
rect 71096 98892 210332 98920
rect 71096 98880 71102 98892
rect 210326 98880 210332 98892
rect 210384 98880 210390 98932
rect 275278 98880 275284 98932
rect 275336 98920 275342 98932
rect 439498 98920 439504 98932
rect 275336 98892 439504 98920
rect 275336 98880 275342 98892
rect 439498 98880 439504 98892
rect 439556 98880 439562 98932
rect 43438 98812 43444 98864
rect 43496 98852 43502 98864
rect 205910 98852 205916 98864
rect 43496 98824 205916 98852
rect 43496 98812 43502 98824
rect 205910 98812 205916 98824
rect 205968 98812 205974 98864
rect 276474 98812 276480 98864
rect 276532 98852 276538 98864
rect 448514 98852 448520 98864
rect 276532 98824 448520 98852
rect 276532 98812 276538 98824
rect 448514 98812 448520 98824
rect 448572 98812 448578 98864
rect 22738 98744 22744 98796
rect 22796 98784 22802 98796
rect 203058 98784 203064 98796
rect 22796 98756 203064 98784
rect 22796 98744 22802 98756
rect 203058 98744 203064 98756
rect 203116 98744 203122 98796
rect 283374 98744 283380 98796
rect 283432 98784 283438 98796
rect 486418 98784 486424 98796
rect 283432 98756 486424 98784
rect 283432 98744 283438 98756
rect 486418 98744 486424 98756
rect 486476 98744 486482 98796
rect 33778 98676 33784 98728
rect 33836 98716 33842 98728
rect 204530 98716 204536 98728
rect 33836 98688 204536 98716
rect 33836 98676 33842 98688
rect 204530 98676 204536 98688
rect 204588 98676 204594 98728
rect 289998 98676 290004 98728
rect 290056 98716 290062 98728
rect 525058 98716 525064 98728
rect 290056 98688 525064 98716
rect 290056 98676 290062 98688
rect 525058 98676 525064 98688
rect 525116 98676 525122 98728
rect 21358 98608 21364 98660
rect 21416 98648 21422 98660
rect 202874 98648 202880 98660
rect 21416 98620 202880 98648
rect 21416 98608 21422 98620
rect 202874 98608 202880 98620
rect 202932 98608 202938 98660
rect 297082 98608 297088 98660
rect 297140 98648 297146 98660
rect 568574 98648 568580 98660
rect 297140 98620 568580 98648
rect 297140 98608 297146 98620
rect 568574 98608 568580 98620
rect 568632 98608 568638 98660
rect 259914 98540 259920 98592
rect 259972 98580 259978 98592
rect 348418 98580 348424 98592
rect 259972 98552 348424 98580
rect 259972 98540 259978 98552
rect 348418 98540 348424 98552
rect 348476 98540 348482 98592
rect 259362 98472 259368 98524
rect 259420 98512 259426 98524
rect 345658 98512 345664 98524
rect 259420 98484 345664 98512
rect 259420 98472 259426 98484
rect 345658 98472 345664 98484
rect 345716 98472 345722 98524
rect 258718 98404 258724 98456
rect 258776 98444 258782 98456
rect 342898 98444 342904 98456
rect 258776 98416 342904 98444
rect 258776 98404 258782 98416
rect 342898 98404 342904 98416
rect 342956 98404 342962 98456
rect 211154 98268 211160 98320
rect 211212 98308 211218 98320
rect 211430 98308 211436 98320
rect 211212 98280 211436 98308
rect 211212 98268 211218 98280
rect 211430 98268 211436 98280
rect 211488 98268 211494 98320
rect 211614 98268 211620 98320
rect 211672 98308 211678 98320
rect 211982 98308 211988 98320
rect 211672 98280 211988 98308
rect 211672 98268 211678 98280
rect 211982 98268 211988 98280
rect 212040 98268 212046 98320
rect 216030 98268 216036 98320
rect 216088 98308 216094 98320
rect 216398 98308 216404 98320
rect 216088 98280 216404 98308
rect 216088 98268 216094 98280
rect 216398 98268 216404 98280
rect 216456 98268 216462 98320
rect 238202 98268 238208 98320
rect 238260 98308 238266 98320
rect 238478 98308 238484 98320
rect 238260 98280 238484 98308
rect 238260 98268 238266 98280
rect 238478 98268 238484 98280
rect 238536 98268 238542 98320
rect 274450 98064 274456 98116
rect 274508 98104 274514 98116
rect 278222 98104 278228 98116
rect 274508 98076 278228 98104
rect 274508 98064 274514 98076
rect 278222 98064 278228 98076
rect 278280 98064 278286 98116
rect 278130 97996 278136 98048
rect 278188 98036 278194 98048
rect 278188 98008 282500 98036
rect 278188 97996 278194 98008
rect 3418 97928 3424 97980
rect 3476 97968 3482 97980
rect 14458 97968 14464 97980
rect 3476 97940 14464 97968
rect 3476 97928 3482 97940
rect 14458 97928 14464 97940
rect 14516 97928 14522 97980
rect 150342 97928 150348 97980
rect 150400 97968 150406 97980
rect 225506 97968 225512 97980
rect 150400 97940 225512 97968
rect 150400 97928 150406 97940
rect 225506 97928 225512 97940
rect 225564 97928 225570 97980
rect 269022 97928 269028 97980
rect 269080 97968 269086 97980
rect 282362 97968 282368 97980
rect 269080 97940 282368 97968
rect 269080 97928 269086 97940
rect 282362 97928 282368 97940
rect 282420 97928 282426 97980
rect 282472 97968 282500 98008
rect 286778 97996 286784 98048
rect 286836 98036 286842 98048
rect 286962 98036 286968 98048
rect 286836 98008 286968 98036
rect 286836 97996 286842 98008
rect 286962 97996 286968 98008
rect 287020 97996 287026 98048
rect 295978 97996 295984 98048
rect 296036 98036 296042 98048
rect 296346 98036 296352 98048
rect 296036 98008 296352 98036
rect 296036 97996 296042 98008
rect 296346 97996 296352 98008
rect 296404 97996 296410 98048
rect 323670 97968 323676 97980
rect 282472 97940 323676 97968
rect 323670 97928 323676 97940
rect 323728 97928 323734 97980
rect 126882 97860 126888 97912
rect 126940 97900 126946 97912
rect 210878 97900 210884 97912
rect 126940 97872 210884 97900
rect 126940 97860 126946 97872
rect 210878 97860 210884 97872
rect 210936 97860 210942 97912
rect 231302 97860 231308 97912
rect 231360 97900 231366 97912
rect 238018 97900 238024 97912
rect 231360 97872 238024 97900
rect 231360 97860 231366 97872
rect 238018 97860 238024 97872
rect 238076 97860 238082 97912
rect 246850 97860 246856 97912
rect 246908 97900 246914 97912
rect 253198 97900 253204 97912
rect 246908 97872 253204 97900
rect 246908 97860 246914 97872
rect 253198 97860 253204 97872
rect 253256 97860 253262 97912
rect 272334 97860 272340 97912
rect 272392 97900 272398 97912
rect 309870 97900 309876 97912
rect 272392 97872 309876 97900
rect 272392 97860 272398 97872
rect 309870 97860 309876 97872
rect 309928 97860 309934 97912
rect 124858 97792 124864 97844
rect 124916 97832 124922 97844
rect 202506 97832 202512 97844
rect 124916 97804 202512 97832
rect 124916 97792 124922 97804
rect 202506 97792 202512 97804
rect 202564 97792 202570 97844
rect 202782 97792 202788 97844
rect 202840 97832 202846 97844
rect 234522 97832 234528 97844
rect 202840 97804 210372 97832
rect 202840 97792 202846 97804
rect 126238 97724 126244 97776
rect 126296 97764 126302 97776
rect 210234 97764 210240 97776
rect 126296 97736 210240 97764
rect 126296 97724 126302 97736
rect 210234 97724 210240 97736
rect 210292 97724 210298 97776
rect 210344 97764 210372 97804
rect 210804 97804 234528 97832
rect 210804 97764 210832 97804
rect 234522 97792 234528 97804
rect 234580 97792 234586 97844
rect 247678 97792 247684 97844
rect 247736 97832 247742 97844
rect 251818 97832 251824 97844
rect 247736 97804 251824 97832
rect 247736 97792 247742 97804
rect 251818 97792 251824 97804
rect 251876 97792 251882 97844
rect 272242 97792 272248 97844
rect 272300 97832 272306 97844
rect 341518 97832 341524 97844
rect 272300 97804 341524 97832
rect 272300 97792 272306 97804
rect 341518 97792 341524 97804
rect 341576 97792 341582 97844
rect 210344 97736 210832 97764
rect 210878 97724 210884 97776
rect 210936 97764 210942 97776
rect 221458 97764 221464 97776
rect 210936 97736 221464 97764
rect 210936 97724 210942 97736
rect 221458 97724 221464 97736
rect 221516 97724 221522 97776
rect 245470 97724 245476 97776
rect 245528 97764 245534 97776
rect 253014 97764 253020 97776
rect 245528 97736 253020 97764
rect 245528 97724 245534 97736
rect 253014 97724 253020 97736
rect 253072 97724 253078 97776
rect 259730 97724 259736 97776
rect 259788 97764 259794 97776
rect 259788 97736 263732 97764
rect 259788 97724 259794 97736
rect 115198 97656 115204 97708
rect 115256 97696 115262 97708
rect 219434 97696 219440 97708
rect 115256 97668 219440 97696
rect 115256 97656 115262 97668
rect 219434 97656 219440 97668
rect 219492 97656 219498 97708
rect 254118 97656 254124 97708
rect 254176 97696 254182 97708
rect 254176 97668 256924 97696
rect 254176 97656 254182 97668
rect 111058 97588 111064 97640
rect 111116 97628 111122 97640
rect 215754 97628 215760 97640
rect 111116 97600 215760 97628
rect 111116 97588 111122 97600
rect 215754 97588 215760 97600
rect 215812 97588 215818 97640
rect 241974 97588 241980 97640
rect 242032 97628 242038 97640
rect 242710 97628 242716 97640
rect 242032 97600 242716 97628
rect 242032 97588 242038 97600
rect 242710 97588 242716 97600
rect 242768 97588 242774 97640
rect 247494 97588 247500 97640
rect 247552 97628 247558 97640
rect 256786 97628 256792 97640
rect 247552 97600 256792 97628
rect 247552 97588 247558 97600
rect 256786 97588 256792 97600
rect 256844 97588 256850 97640
rect 256896 97628 256924 97668
rect 256970 97656 256976 97708
rect 257028 97696 257034 97708
rect 263134 97696 263140 97708
rect 257028 97668 263140 97696
rect 257028 97656 257034 97668
rect 263134 97656 263140 97668
rect 263192 97656 263198 97708
rect 263704 97696 263732 97736
rect 267182 97724 267188 97776
rect 267240 97764 267246 97776
rect 352558 97764 352564 97776
rect 267240 97736 352564 97764
rect 267240 97724 267246 97736
rect 352558 97724 352564 97736
rect 352616 97724 352622 97776
rect 347038 97696 347044 97708
rect 263704 97668 347044 97696
rect 347038 97656 347044 97668
rect 347096 97656 347102 97708
rect 263870 97628 263876 97640
rect 256896 97600 263876 97628
rect 263870 97588 263876 97600
rect 263928 97588 263934 97640
rect 264974 97588 264980 97640
rect 265032 97628 265038 97640
rect 268194 97628 268200 97640
rect 265032 97600 268200 97628
rect 265032 97588 265038 97600
rect 268194 97588 268200 97600
rect 268252 97588 268258 97640
rect 270218 97588 270224 97640
rect 270276 97628 270282 97640
rect 270276 97600 275324 97628
rect 270276 97588 270282 97600
rect 94498 97520 94504 97572
rect 94556 97560 94562 97572
rect 204070 97560 204076 97572
rect 94556 97532 204076 97560
rect 94556 97520 94562 97532
rect 204070 97520 204076 97532
rect 204128 97520 204134 97572
rect 217042 97560 217048 97572
rect 205606 97532 217048 97560
rect 104158 97452 104164 97504
rect 104216 97492 104222 97504
rect 205606 97492 205634 97532
rect 217042 97520 217048 97532
rect 217100 97520 217106 97572
rect 225046 97560 225052 97572
rect 220096 97532 225052 97560
rect 104216 97464 205634 97492
rect 104216 97452 104222 97464
rect 212534 97452 212540 97504
rect 212592 97492 212598 97504
rect 220096 97492 220124 97532
rect 225046 97520 225052 97532
rect 225104 97520 225110 97572
rect 248690 97520 248696 97572
rect 248748 97560 248754 97572
rect 263042 97560 263048 97572
rect 248748 97532 263048 97560
rect 248748 97520 248754 97532
rect 263042 97520 263048 97532
rect 263100 97520 263106 97572
rect 263686 97520 263692 97572
rect 263744 97560 263750 97572
rect 272334 97560 272340 97572
rect 263744 97532 272340 97560
rect 263744 97520 263750 97532
rect 272334 97520 272340 97532
rect 272392 97520 272398 97572
rect 212592 97464 220124 97492
rect 212592 97452 212598 97464
rect 220170 97452 220176 97504
rect 220228 97492 220234 97504
rect 229922 97492 229928 97504
rect 220228 97464 229928 97492
rect 220228 97452 220234 97464
rect 229922 97452 229928 97464
rect 229980 97452 229986 97504
rect 251082 97452 251088 97504
rect 251140 97492 251146 97504
rect 263594 97492 263600 97504
rect 251140 97464 263600 97492
rect 251140 97452 251146 97464
rect 263594 97452 263600 97464
rect 263652 97452 263658 97504
rect 264790 97452 264796 97504
rect 264848 97492 264854 97504
rect 272242 97492 272248 97504
rect 264848 97464 272248 97492
rect 264848 97452 264854 97464
rect 272242 97452 272248 97464
rect 272300 97452 272306 97504
rect 275296 97492 275324 97600
rect 277946 97588 277952 97640
rect 278004 97628 278010 97640
rect 369118 97628 369124 97640
rect 278004 97600 369124 97628
rect 278004 97588 278010 97600
rect 369118 97588 369124 97600
rect 369176 97588 369182 97640
rect 377398 97560 377404 97572
rect 277964 97532 377404 97560
rect 277964 97492 277992 97532
rect 377398 97520 377404 97532
rect 377456 97520 377462 97572
rect 275296 97464 277992 97492
rect 278130 97452 278136 97504
rect 278188 97492 278194 97504
rect 388438 97492 388444 97504
rect 278188 97464 388444 97492
rect 278188 97452 278194 97464
rect 388438 97452 388444 97464
rect 388496 97452 388502 97504
rect 213914 97384 213920 97436
rect 213972 97424 213978 97436
rect 232958 97424 232964 97436
rect 213972 97396 232964 97424
rect 213972 97384 213978 97396
rect 232958 97384 232964 97396
rect 233016 97384 233022 97436
rect 243814 97384 243820 97436
rect 243872 97424 243878 97436
rect 258258 97424 258264 97436
rect 243872 97396 258264 97424
rect 243872 97384 243878 97396
rect 258258 97384 258264 97396
rect 258316 97384 258322 97436
rect 262398 97384 262404 97436
rect 262456 97424 262462 97436
rect 265066 97424 265072 97436
rect 262456 97396 265072 97424
rect 262456 97384 262462 97396
rect 265066 97384 265072 97396
rect 265124 97384 265130 97436
rect 265434 97384 265440 97436
rect 265492 97424 265498 97436
rect 271046 97424 271052 97436
rect 265492 97396 271052 97424
rect 265492 97384 265498 97396
rect 271046 97384 271052 97396
rect 271104 97384 271110 97436
rect 275296 97396 277348 97424
rect 58618 97316 58624 97368
rect 58676 97356 58682 97368
rect 206738 97356 206744 97368
rect 58676 97328 206744 97356
rect 58676 97316 58682 97328
rect 206738 97316 206744 97328
rect 206796 97316 206802 97368
rect 208302 97316 208308 97368
rect 208360 97356 208366 97368
rect 227530 97356 227536 97368
rect 208360 97328 227536 97356
rect 208360 97316 208366 97328
rect 227530 97316 227536 97328
rect 227588 97316 227594 97368
rect 227622 97316 227628 97368
rect 227680 97356 227686 97368
rect 238754 97356 238760 97368
rect 227680 97328 238760 97356
rect 227680 97316 227686 97328
rect 238754 97316 238760 97328
rect 238812 97316 238818 97368
rect 263410 97316 263416 97368
rect 263468 97356 263474 97368
rect 275296 97356 275324 97396
rect 263468 97328 275324 97356
rect 263468 97316 263474 97328
rect 275646 97316 275652 97368
rect 275704 97356 275710 97368
rect 275704 97328 276704 97356
rect 275704 97316 275710 97328
rect 25498 97248 25504 97300
rect 25556 97288 25562 97300
rect 203334 97288 203340 97300
rect 25556 97260 203340 97288
rect 25556 97248 25562 97260
rect 203334 97248 203340 97260
rect 203392 97248 203398 97300
rect 204162 97248 204168 97300
rect 204220 97288 204226 97300
rect 234706 97288 234712 97300
rect 204220 97260 234712 97288
rect 204220 97248 204226 97260
rect 234706 97248 234712 97260
rect 234764 97248 234770 97300
rect 253198 97248 253204 97300
rect 253256 97288 253262 97300
rect 271138 97288 271144 97300
rect 253256 97260 271144 97288
rect 253256 97248 253262 97260
rect 271138 97248 271144 97260
rect 271196 97248 271202 97300
rect 276566 97288 276572 97300
rect 271340 97260 276572 97288
rect 191190 97180 191196 97232
rect 191248 97220 191254 97232
rect 218238 97220 218244 97232
rect 191248 97192 218244 97220
rect 191248 97180 191254 97192
rect 218238 97180 218244 97192
rect 218296 97180 218302 97232
rect 243170 97180 243176 97232
rect 243228 97220 243234 97232
rect 259454 97220 259460 97232
rect 243228 97192 259460 97220
rect 243228 97180 243234 97192
rect 259454 97180 259460 97192
rect 259512 97180 259518 97232
rect 265066 97180 265072 97232
rect 265124 97220 265130 97232
rect 265124 97192 267734 97220
rect 265124 97180 265130 97192
rect 188430 97112 188436 97164
rect 188488 97152 188494 97164
rect 207290 97152 207296 97164
rect 188488 97124 207296 97152
rect 188488 97112 188494 97124
rect 207290 97112 207296 97124
rect 207348 97112 207354 97164
rect 210970 97152 210976 97164
rect 208320 97124 210976 97152
rect 196618 97044 196624 97096
rect 196676 97084 196682 97096
rect 208320 97084 208348 97124
rect 210970 97112 210976 97124
rect 211028 97112 211034 97164
rect 211154 97112 211160 97164
rect 211212 97152 211218 97164
rect 222654 97152 222660 97164
rect 211212 97124 222660 97152
rect 211212 97112 211218 97124
rect 222654 97112 222660 97124
rect 222712 97112 222718 97164
rect 242986 97112 242992 97164
rect 243044 97152 243050 97164
rect 250254 97152 250260 97164
rect 243044 97124 250260 97152
rect 243044 97112 243050 97124
rect 250254 97112 250260 97124
rect 250312 97112 250318 97164
rect 255958 97112 255964 97164
rect 256016 97152 256022 97164
rect 256602 97152 256608 97164
rect 256016 97124 256608 97152
rect 256016 97112 256022 97124
rect 256602 97112 256608 97124
rect 256660 97112 256666 97164
rect 256786 97112 256792 97164
rect 256844 97152 256850 97164
rect 260098 97152 260104 97164
rect 256844 97124 260104 97152
rect 256844 97112 256850 97124
rect 260098 97112 260104 97124
rect 260156 97112 260162 97164
rect 261202 97112 261208 97164
rect 261260 97152 261266 97164
rect 267706 97152 267734 97192
rect 268378 97180 268384 97232
rect 268436 97220 268442 97232
rect 271340 97220 271368 97260
rect 276566 97248 276572 97260
rect 276624 97248 276630 97300
rect 276676 97288 276704 97328
rect 276842 97316 276848 97368
rect 276900 97356 276906 97368
rect 277210 97356 277216 97368
rect 276900 97328 277216 97356
rect 276900 97316 276906 97328
rect 277210 97316 277216 97328
rect 277268 97316 277274 97368
rect 277320 97356 277348 97396
rect 278314 97384 278320 97436
rect 278372 97424 278378 97436
rect 393958 97424 393964 97436
rect 278372 97396 393964 97424
rect 278372 97384 278378 97396
rect 393958 97384 393964 97396
rect 394016 97384 394022 97436
rect 277946 97356 277952 97368
rect 277320 97328 277952 97356
rect 277946 97316 277952 97328
rect 278004 97316 278010 97368
rect 282638 97356 282644 97368
rect 278516 97328 282644 97356
rect 278516 97288 278544 97328
rect 282638 97316 282644 97328
rect 282696 97316 282702 97368
rect 283650 97316 283656 97368
rect 283708 97356 283714 97368
rect 411898 97356 411904 97368
rect 283708 97328 411904 97356
rect 283708 97316 283714 97328
rect 411898 97316 411904 97328
rect 411956 97316 411962 97368
rect 276676 97260 278544 97288
rect 283006 97248 283012 97300
rect 283064 97288 283070 97300
rect 418798 97288 418804 97300
rect 283064 97260 418804 97288
rect 283064 97248 283070 97260
rect 418798 97248 418804 97260
rect 418856 97248 418862 97300
rect 268436 97192 271368 97220
rect 268436 97180 268442 97192
rect 271414 97180 271420 97232
rect 271472 97220 271478 97232
rect 278130 97220 278136 97232
rect 271472 97192 278136 97220
rect 271472 97180 271478 97192
rect 278130 97180 278136 97192
rect 278188 97180 278194 97232
rect 278222 97180 278228 97232
rect 278280 97220 278286 97232
rect 282178 97220 282184 97232
rect 278280 97192 282184 97220
rect 278280 97180 278286 97192
rect 282178 97180 282184 97192
rect 282236 97180 282242 97232
rect 304258 97220 304264 97232
rect 283116 97192 304264 97220
rect 271230 97152 271236 97164
rect 261260 97124 264376 97152
rect 267706 97124 271236 97152
rect 261260 97112 261266 97124
rect 196676 97056 208348 97084
rect 196676 97044 196682 97056
rect 210234 97044 210240 97096
rect 210292 97084 210298 97096
rect 221274 97084 221280 97096
rect 210292 97056 221280 97084
rect 210292 97044 210298 97056
rect 221274 97044 221280 97056
rect 221332 97044 221338 97096
rect 241422 97044 241428 97096
rect 241480 97084 241486 97096
rect 242158 97084 242164 97096
rect 241480 97056 242164 97084
rect 241480 97044 241486 97056
rect 242158 97044 242164 97056
rect 242216 97044 242222 97096
rect 242434 97044 242440 97096
rect 242492 97084 242498 97096
rect 246298 97084 246304 97096
rect 242492 97056 246304 97084
rect 242492 97044 242498 97056
rect 246298 97044 246304 97056
rect 246356 97044 246362 97096
rect 249702 97084 249708 97096
rect 249352 97056 249708 97084
rect 199378 96976 199384 97028
rect 199436 97016 199442 97028
rect 209130 97016 209136 97028
rect 199436 96988 209136 97016
rect 199436 96976 199442 96988
rect 209130 96976 209136 96988
rect 209188 96976 209194 97028
rect 204254 96908 204260 96960
rect 204312 96948 204318 96960
rect 207750 96948 207756 96960
rect 204312 96920 207756 96948
rect 204312 96908 204318 96920
rect 207750 96908 207756 96920
rect 207808 96908 207814 96960
rect 223574 96908 223580 96960
rect 223632 96948 223638 96960
rect 225230 96948 225236 96960
rect 223632 96920 225236 96948
rect 223632 96908 223638 96920
rect 225230 96908 225236 96920
rect 225288 96908 225294 96960
rect 244458 96908 244464 96960
rect 244516 96948 244522 96960
rect 245286 96948 245292 96960
rect 244516 96920 245292 96948
rect 244516 96908 244522 96920
rect 245286 96908 245292 96920
rect 245344 96908 245350 96960
rect 245838 96908 245844 96960
rect 245896 96948 245902 96960
rect 246482 96948 246488 96960
rect 245896 96920 246488 96948
rect 245896 96908 245902 96920
rect 246482 96908 246488 96920
rect 246540 96908 246546 96960
rect 247218 96908 247224 96960
rect 247276 96948 247282 96960
rect 248230 96948 248236 96960
rect 247276 96920 248236 96948
rect 247276 96908 247282 96920
rect 248230 96908 248236 96920
rect 248288 96908 248294 96960
rect 203886 96840 203892 96892
rect 203944 96880 203950 96892
rect 207934 96880 207940 96892
rect 203944 96852 207940 96880
rect 203944 96840 203950 96852
rect 207934 96840 207940 96852
rect 207992 96840 207998 96892
rect 237374 96840 237380 96892
rect 237432 96880 237438 96892
rect 239214 96880 239220 96892
rect 237432 96852 239220 96880
rect 237432 96840 237438 96852
rect 239214 96840 239220 96852
rect 239272 96840 239278 96892
rect 241790 96840 241796 96892
rect 241848 96880 241854 96892
rect 244366 96880 244372 96892
rect 241848 96852 244372 96880
rect 241848 96840 241854 96852
rect 244366 96840 244372 96852
rect 244424 96840 244430 96892
rect 245654 96840 245660 96892
rect 245712 96880 245718 96892
rect 246666 96880 246672 96892
rect 245712 96852 246672 96880
rect 245712 96840 245718 96852
rect 246666 96840 246672 96852
rect 246724 96840 246730 96892
rect 249352 96824 249380 97056
rect 249702 97044 249708 97056
rect 249760 97044 249766 97096
rect 256142 97044 256148 97096
rect 256200 97084 256206 97096
rect 256418 97084 256424 97096
rect 256200 97056 256424 97084
rect 256200 97044 256206 97056
rect 256418 97044 256424 97056
rect 256476 97044 256482 97096
rect 260558 97044 260564 97096
rect 260616 97084 260622 97096
rect 262858 97084 262864 97096
rect 260616 97056 262864 97084
rect 260616 97044 260622 97056
rect 262858 97044 262864 97056
rect 262916 97044 262922 97096
rect 264348 97084 264376 97124
rect 271230 97112 271236 97124
rect 271288 97112 271294 97164
rect 278682 97112 278688 97164
rect 278740 97152 278746 97164
rect 283116 97152 283144 97192
rect 304258 97180 304264 97192
rect 304316 97180 304322 97232
rect 278740 97124 283144 97152
rect 278740 97112 278746 97124
rect 287974 97112 287980 97164
rect 288032 97152 288038 97164
rect 288250 97152 288256 97164
rect 288032 97124 288256 97152
rect 288032 97112 288038 97124
rect 288250 97112 288256 97124
rect 288308 97112 288314 97164
rect 288802 97112 288808 97164
rect 288860 97152 288866 97164
rect 289722 97152 289728 97164
rect 288860 97124 289728 97152
rect 288860 97112 288866 97124
rect 289722 97112 289728 97124
rect 289780 97112 289786 97164
rect 292206 97112 292212 97164
rect 292264 97152 292270 97164
rect 292482 97152 292488 97164
rect 292264 97124 292488 97152
rect 292264 97112 292270 97124
rect 292482 97112 292488 97124
rect 292540 97112 292546 97164
rect 296070 97112 296076 97164
rect 296128 97152 296134 97164
rect 296346 97152 296352 97164
rect 296128 97124 296352 97152
rect 296128 97112 296134 97124
rect 296346 97112 296352 97124
rect 296404 97112 296410 97164
rect 296622 97112 296628 97164
rect 296680 97152 296686 97164
rect 322198 97152 322204 97164
rect 296680 97124 322204 97152
rect 296680 97112 296686 97124
rect 322198 97112 322204 97124
rect 322256 97112 322262 97164
rect 274174 97084 274180 97096
rect 264348 97056 274180 97084
rect 274174 97044 274180 97056
rect 274232 97044 274238 97096
rect 278332 97056 281672 97084
rect 250438 96976 250444 97028
rect 250496 97016 250502 97028
rect 251082 97016 251088 97028
rect 250496 96988 251088 97016
rect 250496 96976 250502 96988
rect 251082 96976 251088 96988
rect 251140 96976 251146 97028
rect 251450 96976 251456 97028
rect 251508 97016 251514 97028
rect 252278 97016 252284 97028
rect 251508 96988 252284 97016
rect 251508 96976 251514 96988
rect 252278 96976 252284 96988
rect 252336 96976 252342 97028
rect 258166 96976 258172 97028
rect 258224 97016 258230 97028
rect 258994 97016 259000 97028
rect 258224 96988 259000 97016
rect 258224 96976 258230 96988
rect 258994 96976 259000 96988
rect 259052 96976 259058 97028
rect 262766 96976 262772 97028
rect 262824 97016 262830 97028
rect 263502 97016 263508 97028
rect 262824 96988 263508 97016
rect 262824 96976 262830 96988
rect 263502 96976 263508 96988
rect 263560 96976 263566 97028
rect 265618 96976 265624 97028
rect 265676 97016 265682 97028
rect 266262 97016 266268 97028
rect 265676 96988 266268 97016
rect 265676 96976 265682 96988
rect 266262 96976 266268 96988
rect 266320 96976 266326 97028
rect 266446 96976 266452 97028
rect 266504 97016 266510 97028
rect 267458 97016 267464 97028
rect 266504 96988 267464 97016
rect 266504 96976 266510 96988
rect 267458 96976 267464 96988
rect 267516 96976 267522 97028
rect 268654 96976 268660 97028
rect 268712 97016 268718 97028
rect 269022 97016 269028 97028
rect 268712 96988 269028 97016
rect 268712 96976 268718 96988
rect 269022 96976 269028 96988
rect 269080 96976 269086 97028
rect 269206 96976 269212 97028
rect 269264 97016 269270 97028
rect 270310 97016 270316 97028
rect 269264 96988 270316 97016
rect 269264 96976 269270 96988
rect 270310 96976 270316 96988
rect 270368 96976 270374 97028
rect 272058 96976 272064 97028
rect 272116 97016 272122 97028
rect 278222 97016 278228 97028
rect 272116 96988 278228 97016
rect 272116 96976 272122 96988
rect 278222 96976 278228 96988
rect 278280 96976 278286 97028
rect 250070 96908 250076 96960
rect 250128 96948 250134 96960
rect 250990 96948 250996 96960
rect 250128 96920 250996 96948
rect 250128 96908 250134 96920
rect 250990 96908 250996 96920
rect 251048 96908 251054 96960
rect 251910 96908 251916 96960
rect 251968 96948 251974 96960
rect 252186 96948 252192 96960
rect 251968 96920 252192 96948
rect 251968 96908 251974 96920
rect 252186 96908 252192 96920
rect 252244 96908 252250 96960
rect 253106 96908 253112 96960
rect 253164 96948 253170 96960
rect 253566 96948 253572 96960
rect 253164 96920 253572 96948
rect 253164 96908 253170 96920
rect 253566 96908 253572 96920
rect 253624 96908 253630 96960
rect 254854 96908 254860 96960
rect 254912 96948 254918 96960
rect 255130 96948 255136 96960
rect 254912 96920 255136 96948
rect 254912 96908 254918 96920
rect 255130 96908 255136 96920
rect 255188 96908 255194 96960
rect 255498 96908 255504 96960
rect 255556 96948 255562 96960
rect 256326 96948 256332 96960
rect 255556 96920 256332 96948
rect 255556 96908 255562 96920
rect 256326 96908 256332 96920
rect 256384 96908 256390 96960
rect 257614 96908 257620 96960
rect 257672 96948 257678 96960
rect 257890 96948 257896 96960
rect 257672 96920 257896 96948
rect 257672 96908 257678 96920
rect 257890 96908 257896 96920
rect 257948 96908 257954 96960
rect 258534 96908 258540 96960
rect 258592 96948 258598 96960
rect 259086 96948 259092 96960
rect 258592 96920 259092 96948
rect 258592 96908 258598 96920
rect 259086 96908 259092 96920
rect 259144 96908 259150 96960
rect 260190 96908 260196 96960
rect 260248 96948 260254 96960
rect 260650 96948 260656 96960
rect 260248 96920 260656 96948
rect 260248 96908 260254 96920
rect 260650 96908 260656 96920
rect 260708 96908 260714 96960
rect 262950 96908 262956 96960
rect 263008 96948 263014 96960
rect 263410 96948 263416 96960
rect 263008 96920 263416 96948
rect 263008 96908 263014 96920
rect 263410 96908 263416 96920
rect 263468 96908 263474 96960
rect 264422 96908 264428 96960
rect 264480 96948 264486 96960
rect 264882 96948 264888 96960
rect 264480 96920 264888 96948
rect 264480 96908 264486 96920
rect 264882 96908 264888 96920
rect 264940 96908 264946 96960
rect 265802 96908 265808 96960
rect 265860 96948 265866 96960
rect 266078 96948 266084 96960
rect 265860 96920 266084 96948
rect 265860 96908 265866 96920
rect 266078 96908 266084 96920
rect 266136 96908 266142 96960
rect 266998 96908 267004 96960
rect 267056 96948 267062 96960
rect 267366 96948 267372 96960
rect 267056 96920 267372 96948
rect 267056 96908 267062 96920
rect 267366 96908 267372 96920
rect 267424 96908 267430 96960
rect 268010 96908 268016 96960
rect 268068 96948 268074 96960
rect 268930 96948 268936 96960
rect 268068 96920 268936 96948
rect 268068 96908 268074 96920
rect 268930 96908 268936 96920
rect 268988 96908 268994 96960
rect 269666 96908 269672 96960
rect 269724 96948 269730 96960
rect 270126 96948 270132 96960
rect 269724 96920 270132 96948
rect 269724 96908 269730 96920
rect 270126 96908 270132 96920
rect 270184 96908 270190 96960
rect 270862 96908 270868 96960
rect 270920 96948 270926 96960
rect 271782 96948 271788 96960
rect 270920 96920 271788 96948
rect 270920 96908 270926 96920
rect 271782 96908 271788 96920
rect 271840 96908 271846 96960
rect 272426 96908 272432 96960
rect 272484 96948 272490 96960
rect 272978 96948 272984 96960
rect 272484 96920 272984 96948
rect 272484 96908 272490 96920
rect 272978 96908 272984 96920
rect 273036 96908 273042 96960
rect 273254 96908 273260 96960
rect 273312 96948 273318 96960
rect 273898 96948 273904 96960
rect 273312 96920 273904 96948
rect 273312 96908 273318 96920
rect 273898 96908 273904 96920
rect 273956 96908 273962 96960
rect 275646 96908 275652 96960
rect 275704 96948 275710 96960
rect 275922 96948 275928 96960
rect 275704 96920 275928 96948
rect 275704 96908 275710 96920
rect 275922 96908 275928 96920
rect 275980 96908 275986 96960
rect 276290 96908 276296 96960
rect 276348 96948 276354 96960
rect 278332 96948 278360 97056
rect 279142 96976 279148 97028
rect 279200 97016 279206 97028
rect 281166 97016 281172 97028
rect 279200 96988 281172 97016
rect 279200 96976 279206 96988
rect 281166 96976 281172 96988
rect 281224 96976 281230 97028
rect 276348 96920 278360 96948
rect 276348 96908 276354 96920
rect 280154 96908 280160 96960
rect 280212 96948 280218 96960
rect 281350 96948 281356 96960
rect 280212 96920 281356 96948
rect 280212 96908 280218 96920
rect 281350 96908 281356 96920
rect 281408 96908 281414 96960
rect 281644 96948 281672 97056
rect 281718 97044 281724 97096
rect 281776 97084 281782 97096
rect 284294 97084 284300 97096
rect 281776 97056 284300 97084
rect 281776 97044 281782 97056
rect 284294 97044 284300 97056
rect 284352 97044 284358 97096
rect 286318 97044 286324 97096
rect 286376 97084 286382 97096
rect 286686 97084 286692 97096
rect 286376 97056 286692 97084
rect 286376 97044 286382 97056
rect 286686 97044 286692 97056
rect 286744 97044 286750 97096
rect 286778 97044 286784 97096
rect 286836 97084 286842 97096
rect 312538 97084 312544 97096
rect 286836 97056 312544 97084
rect 286836 97044 286842 97056
rect 312538 97044 312544 97056
rect 312596 97044 312602 97096
rect 282362 96976 282368 97028
rect 282420 97016 282426 97028
rect 282420 96988 297588 97016
rect 282420 96976 282426 96988
rect 297560 96948 297588 96988
rect 297634 96976 297640 97028
rect 297692 97016 297698 97028
rect 298002 97016 298008 97028
rect 297692 96988 298008 97016
rect 297692 96976 297698 96988
rect 298002 96976 298008 96988
rect 298060 96976 298066 97028
rect 298094 96976 298100 97028
rect 298152 97016 298158 97028
rect 299106 97016 299112 97028
rect 298152 96988 299112 97016
rect 298152 96976 298158 96988
rect 299106 96976 299112 96988
rect 299164 96976 299170 97028
rect 281644 96920 296760 96948
rect 297560 96920 297772 96948
rect 250714 96840 250720 96892
rect 250772 96880 250778 96892
rect 250898 96880 250904 96892
rect 250772 96852 250904 96880
rect 250772 96840 250778 96852
rect 250898 96840 250904 96852
rect 250956 96840 250962 96892
rect 252002 96840 252008 96892
rect 252060 96880 252066 96892
rect 252462 96880 252468 96892
rect 252060 96852 252468 96880
rect 252060 96840 252066 96852
rect 252462 96840 252468 96852
rect 252520 96840 252526 96892
rect 252646 96840 252652 96892
rect 252704 96880 252710 96892
rect 253750 96880 253756 96892
rect 252704 96852 253756 96880
rect 252704 96840 252710 96852
rect 253750 96840 253756 96852
rect 253808 96840 253814 96892
rect 253934 96840 253940 96892
rect 253992 96880 253998 96892
rect 255038 96880 255044 96892
rect 253992 96852 255044 96880
rect 253992 96840 253998 96852
rect 255038 96840 255044 96852
rect 255096 96840 255102 96892
rect 256694 96840 256700 96892
rect 256752 96880 256758 96892
rect 257798 96880 257804 96892
rect 256752 96852 257804 96880
rect 256752 96840 256758 96852
rect 257798 96840 257804 96852
rect 257856 96840 257862 96892
rect 258902 96840 258908 96892
rect 258960 96880 258966 96892
rect 259270 96880 259276 96892
rect 258960 96852 259276 96880
rect 258960 96840 258966 96852
rect 259270 96840 259276 96852
rect 259328 96840 259334 96892
rect 261570 96840 261576 96892
rect 261628 96880 261634 96892
rect 261938 96880 261944 96892
rect 261628 96852 261944 96880
rect 261628 96840 261634 96852
rect 261938 96840 261944 96852
rect 261996 96840 262002 96892
rect 262582 96840 262588 96892
rect 262640 96880 262646 96892
rect 263318 96880 263324 96892
rect 262640 96852 263324 96880
rect 262640 96840 262646 96852
rect 263318 96840 263324 96852
rect 263376 96840 263382 96892
rect 263778 96840 263784 96892
rect 263836 96880 263842 96892
rect 264606 96880 264612 96892
rect 263836 96852 264612 96880
rect 263836 96840 263842 96852
rect 264606 96840 264612 96852
rect 264664 96840 264670 96892
rect 265894 96840 265900 96892
rect 265952 96880 265958 96892
rect 266170 96880 266176 96892
rect 265952 96852 266176 96880
rect 265952 96840 265958 96852
rect 266170 96840 266176 96852
rect 266228 96840 266234 96892
rect 266814 96840 266820 96892
rect 266872 96880 266878 96892
rect 267550 96880 267556 96892
rect 266872 96852 267556 96880
rect 266872 96840 266878 96852
rect 267550 96840 267556 96852
rect 267608 96840 267614 96892
rect 267826 96840 267832 96892
rect 267884 96880 267890 96892
rect 268838 96880 268844 96892
rect 267884 96852 268844 96880
rect 267884 96840 267890 96852
rect 268838 96840 268844 96852
rect 268896 96840 268902 96892
rect 269942 96840 269948 96892
rect 270000 96880 270006 96892
rect 270402 96880 270408 96892
rect 270000 96852 270408 96880
rect 270000 96840 270006 96852
rect 270402 96840 270408 96852
rect 270460 96840 270466 96892
rect 272886 96840 272892 96892
rect 272944 96880 272950 96892
rect 273162 96880 273168 96892
rect 272944 96852 273168 96880
rect 272944 96840 272950 96852
rect 273162 96840 273168 96852
rect 273220 96840 273226 96892
rect 276658 96840 276664 96892
rect 276716 96880 276722 96892
rect 277210 96880 277216 96892
rect 276716 96852 277216 96880
rect 276716 96840 276722 96852
rect 277210 96840 277216 96852
rect 277268 96840 277274 96892
rect 280890 96840 280896 96892
rect 280948 96880 280954 96892
rect 281442 96880 281448 96892
rect 280948 96852 281448 96880
rect 280948 96840 280954 96852
rect 281442 96840 281448 96852
rect 281500 96840 281506 96892
rect 282178 96840 282184 96892
rect 282236 96880 282242 96892
rect 283650 96880 283656 96892
rect 282236 96852 283656 96880
rect 282236 96840 282242 96852
rect 283650 96840 283656 96852
rect 283708 96840 283714 96892
rect 283834 96840 283840 96892
rect 283892 96880 283898 96892
rect 284110 96880 284116 96892
rect 283892 96852 284116 96880
rect 283892 96840 283898 96852
rect 284110 96840 284116 96852
rect 284168 96840 284174 96892
rect 285122 96840 285128 96892
rect 285180 96880 285186 96892
rect 285398 96880 285404 96892
rect 285180 96852 285404 96880
rect 285180 96840 285186 96852
rect 285398 96840 285404 96852
rect 285456 96840 285462 96892
rect 285766 96840 285772 96892
rect 285824 96880 285830 96892
rect 286410 96880 286416 96892
rect 285824 96852 286416 96880
rect 285824 96840 285830 96852
rect 286410 96840 286416 96852
rect 286468 96840 286474 96892
rect 287146 96840 287152 96892
rect 287204 96880 287210 96892
rect 288158 96880 288164 96892
rect 287204 96852 288164 96880
rect 287204 96840 287210 96852
rect 288158 96840 288164 96852
rect 288216 96840 288222 96892
rect 288618 96840 288624 96892
rect 288676 96880 288682 96892
rect 289262 96880 289268 96892
rect 288676 96852 289268 96880
rect 288676 96840 288682 96852
rect 289262 96840 289268 96852
rect 289320 96840 289326 96892
rect 290550 96840 290556 96892
rect 290608 96880 290614 96892
rect 290918 96880 290924 96892
rect 290608 96852 290924 96880
rect 290608 96840 290614 96852
rect 290918 96840 290924 96852
rect 290976 96840 290982 96892
rect 291378 96840 291384 96892
rect 291436 96880 291442 96892
rect 291930 96880 291936 96892
rect 291436 96852 291936 96880
rect 291436 96840 291442 96852
rect 291930 96840 291936 96852
rect 291988 96840 291994 96892
rect 293034 96840 293040 96892
rect 293092 96880 293098 96892
rect 293402 96880 293408 96892
rect 293092 96852 293408 96880
rect 293092 96840 293098 96852
rect 293402 96840 293408 96852
rect 293460 96840 293466 96892
rect 293494 96840 293500 96892
rect 293552 96880 293558 96892
rect 293862 96880 293868 96892
rect 293552 96852 293868 96880
rect 293552 96840 293558 96852
rect 293862 96840 293868 96852
rect 293920 96840 293926 96892
rect 294598 96840 294604 96892
rect 294656 96880 294662 96892
rect 295242 96880 295248 96892
rect 294656 96852 295248 96880
rect 294656 96840 294662 96852
rect 295242 96840 295248 96852
rect 295300 96840 295306 96892
rect 295426 96840 295432 96892
rect 295484 96880 295490 96892
rect 296070 96880 296076 96892
rect 295484 96852 296076 96880
rect 295484 96840 295490 96852
rect 296070 96840 296076 96852
rect 296128 96840 296134 96892
rect 86862 96772 86868 96824
rect 86920 96812 86926 96824
rect 86920 96784 195974 96812
rect 86920 96772 86926 96784
rect 195946 96744 195974 96784
rect 235994 96772 236000 96824
rect 236052 96812 236058 96824
rect 239030 96812 239036 96824
rect 236052 96784 239036 96812
rect 236052 96772 236058 96784
rect 239030 96772 239036 96784
rect 239088 96772 239094 96824
rect 244642 96772 244648 96824
rect 244700 96812 244706 96824
rect 245378 96812 245384 96824
rect 244700 96784 245384 96812
rect 244700 96772 244706 96784
rect 245378 96772 245384 96784
rect 245436 96772 245442 96824
rect 246206 96772 246212 96824
rect 246264 96812 246270 96824
rect 246758 96812 246764 96824
rect 246264 96784 246764 96812
rect 246264 96772 246270 96784
rect 246758 96772 246764 96784
rect 246816 96772 246822 96824
rect 248414 96772 248420 96824
rect 248472 96812 248478 96824
rect 249242 96812 249248 96824
rect 248472 96784 249248 96812
rect 248472 96772 248478 96784
rect 249242 96772 249248 96784
rect 249300 96772 249306 96824
rect 249334 96772 249340 96824
rect 249392 96772 249398 96824
rect 254486 96772 254492 96824
rect 254544 96812 254550 96824
rect 255130 96812 255136 96824
rect 254544 96784 255136 96812
rect 254544 96772 254550 96784
rect 255130 96772 255136 96784
rect 255188 96772 255194 96824
rect 256050 96772 256056 96824
rect 256108 96812 256114 96824
rect 256510 96812 256516 96824
rect 256108 96784 256516 96812
rect 256108 96772 256114 96784
rect 256510 96772 256516 96784
rect 256568 96772 256574 96824
rect 257338 96772 257344 96824
rect 257396 96812 257402 96824
rect 257890 96812 257896 96824
rect 257396 96784 257896 96812
rect 257396 96772 257402 96784
rect 257890 96772 257896 96784
rect 257948 96772 257954 96824
rect 258350 96772 258356 96824
rect 258408 96812 258414 96824
rect 259362 96812 259368 96824
rect 258408 96784 259368 96812
rect 258408 96772 258414 96784
rect 259362 96772 259368 96784
rect 259420 96772 259426 96824
rect 260466 96772 260472 96824
rect 260524 96812 260530 96824
rect 260742 96812 260748 96824
rect 260524 96784 260748 96812
rect 260524 96772 260530 96784
rect 260742 96772 260748 96784
rect 260800 96772 260806 96824
rect 263962 96772 263968 96824
rect 264020 96812 264026 96824
rect 264698 96812 264704 96824
rect 264020 96784 264704 96812
rect 264020 96772 264026 96784
rect 264698 96772 264704 96784
rect 264756 96772 264762 96824
rect 266630 96772 266636 96824
rect 266688 96812 266694 96824
rect 267274 96812 267280 96824
rect 266688 96784 267280 96812
rect 266688 96772 266694 96784
rect 267274 96772 267280 96784
rect 267332 96772 267338 96824
rect 270678 96772 270684 96824
rect 270736 96812 270742 96824
rect 271598 96812 271604 96824
rect 270736 96784 271604 96812
rect 270736 96772 270742 96784
rect 271598 96772 271604 96784
rect 271656 96772 271662 96824
rect 272610 96772 272616 96824
rect 272668 96812 272674 96824
rect 272668 96784 273254 96812
rect 272668 96772 272674 96784
rect 214466 96744 214472 96756
rect 195946 96716 214472 96744
rect 214466 96704 214472 96716
rect 214524 96704 214530 96756
rect 215938 96704 215944 96756
rect 215996 96744 216002 96756
rect 218790 96744 218796 96756
rect 215996 96716 218796 96744
rect 215996 96704 216002 96716
rect 218790 96704 218796 96716
rect 218848 96704 218854 96756
rect 219434 96704 219440 96756
rect 219492 96744 219498 96756
rect 223022 96744 223028 96756
rect 219492 96716 223028 96744
rect 219492 96704 219498 96716
rect 223022 96704 223028 96716
rect 223080 96704 223086 96756
rect 233878 96704 233884 96756
rect 233936 96744 233942 96756
rect 238570 96744 238576 96756
rect 233936 96716 238576 96744
rect 233936 96704 233942 96716
rect 238570 96704 238576 96716
rect 238628 96704 238634 96756
rect 246022 96704 246028 96756
rect 246080 96744 246086 96756
rect 246850 96744 246856 96756
rect 246080 96716 246856 96744
rect 246080 96704 246086 96716
rect 246850 96704 246856 96716
rect 246908 96704 246914 96756
rect 260926 96704 260932 96756
rect 260984 96744 260990 96756
rect 261846 96744 261852 96756
rect 260984 96716 261852 96744
rect 260984 96704 260990 96716
rect 261846 96704 261852 96716
rect 261904 96704 261910 96756
rect 265158 96704 265164 96756
rect 265216 96744 265222 96756
rect 266170 96744 266176 96756
rect 265216 96716 266176 96744
rect 265216 96704 265222 96716
rect 266170 96704 266176 96716
rect 266228 96704 266234 96756
rect 269850 96704 269856 96756
rect 269908 96744 269914 96756
rect 270218 96744 270224 96756
rect 269908 96716 270224 96744
rect 269908 96704 269914 96716
rect 270218 96704 270224 96716
rect 270276 96704 270282 96756
rect 271874 96704 271880 96756
rect 271932 96744 271938 96756
rect 272886 96744 272892 96756
rect 271932 96716 272892 96744
rect 271932 96704 271938 96716
rect 272886 96704 272892 96716
rect 272944 96704 272950 96756
rect 273226 96744 273254 96784
rect 274910 96772 274916 96824
rect 274968 96812 274974 96824
rect 275922 96812 275928 96824
rect 274968 96784 275928 96812
rect 274968 96772 274974 96784
rect 275922 96772 275928 96784
rect 275980 96772 275986 96824
rect 276106 96772 276112 96824
rect 276164 96812 276170 96824
rect 277118 96812 277124 96824
rect 276164 96784 277124 96812
rect 276164 96772 276170 96784
rect 277118 96772 277124 96784
rect 277176 96772 277182 96824
rect 280338 96772 280344 96824
rect 280396 96812 280402 96824
rect 281074 96812 281080 96824
rect 280396 96784 281080 96812
rect 280396 96772 280402 96784
rect 281074 96772 281080 96784
rect 281132 96772 281138 96824
rect 281166 96772 281172 96824
rect 281224 96812 281230 96824
rect 282270 96812 282276 96824
rect 281224 96784 282276 96812
rect 281224 96772 281230 96784
rect 282270 96772 282276 96784
rect 282328 96772 282334 96824
rect 283558 96772 283564 96824
rect 283616 96812 283622 96824
rect 284018 96812 284024 96824
rect 283616 96784 284024 96812
rect 283616 96772 283622 96784
rect 284018 96772 284024 96784
rect 284076 96772 284082 96824
rect 284570 96772 284576 96824
rect 284628 96812 284634 96824
rect 285306 96812 285312 96824
rect 284628 96784 285312 96812
rect 284628 96772 284634 96784
rect 285306 96772 285312 96784
rect 285364 96772 285370 96824
rect 285950 96772 285956 96824
rect 286008 96812 286014 96824
rect 286594 96812 286600 96824
rect 286008 96784 286600 96812
rect 286008 96772 286014 96784
rect 286594 96772 286600 96784
rect 286652 96772 286658 96824
rect 287882 96772 287888 96824
rect 287940 96812 287946 96824
rect 288342 96812 288348 96824
rect 287940 96784 288348 96812
rect 287940 96772 287946 96784
rect 288342 96772 288348 96784
rect 288400 96772 288406 96824
rect 288986 96772 288992 96824
rect 289044 96812 289050 96824
rect 289538 96812 289544 96824
rect 289044 96784 289544 96812
rect 289044 96772 289050 96784
rect 289538 96772 289544 96784
rect 289596 96772 289602 96824
rect 291838 96772 291844 96824
rect 291896 96812 291902 96824
rect 292298 96812 292304 96824
rect 291896 96784 292304 96812
rect 291896 96772 291902 96784
rect 292298 96772 292304 96784
rect 292356 96772 292362 96824
rect 292574 96772 292580 96824
rect 292632 96812 292638 96824
rect 293678 96812 293684 96824
rect 292632 96784 293684 96812
rect 292632 96772 292638 96784
rect 293678 96772 293684 96784
rect 293736 96772 293742 96824
rect 295610 96772 295616 96824
rect 295668 96812 295674 96824
rect 296254 96812 296260 96824
rect 295668 96784 296260 96812
rect 295668 96772 295674 96784
rect 296254 96772 296260 96784
rect 296312 96772 296318 96824
rect 286778 96744 286784 96756
rect 273226 96716 286784 96744
rect 286778 96704 286784 96716
rect 286836 96704 286842 96756
rect 289170 96704 289176 96756
rect 289228 96744 289234 96756
rect 289630 96744 289636 96756
rect 289228 96716 289636 96744
rect 289228 96704 289234 96716
rect 289630 96704 289636 96716
rect 289688 96704 289694 96756
rect 290182 96704 290188 96756
rect 290240 96744 290246 96756
rect 290826 96744 290832 96756
rect 290240 96716 290832 96744
rect 290240 96704 290246 96716
rect 290826 96704 290832 96716
rect 290884 96704 290890 96756
rect 291194 96704 291200 96756
rect 291252 96744 291258 96756
rect 292114 96744 292120 96756
rect 291252 96716 292120 96744
rect 291252 96704 291258 96716
rect 292114 96704 292120 96716
rect 292172 96704 292178 96756
rect 294874 96704 294880 96756
rect 294932 96744 294938 96756
rect 295058 96744 295064 96756
rect 294932 96716 295064 96744
rect 294932 96704 294938 96716
rect 295058 96704 295064 96716
rect 295116 96704 295122 96756
rect 295794 96704 295800 96756
rect 295852 96744 295858 96756
rect 296530 96744 296536 96756
rect 295852 96716 296536 96744
rect 295852 96704 295858 96716
rect 296530 96704 296536 96716
rect 296588 96704 296594 96756
rect 197998 96636 198004 96688
rect 198056 96676 198062 96688
rect 200850 96676 200856 96688
rect 198056 96648 200856 96676
rect 198056 96636 198062 96648
rect 200850 96636 200856 96648
rect 200908 96636 200914 96688
rect 202138 96636 202144 96688
rect 202196 96676 202202 96688
rect 205542 96676 205548 96688
rect 202196 96648 205548 96676
rect 202196 96636 202202 96648
rect 205542 96636 205548 96648
rect 205600 96636 205606 96688
rect 209038 96636 209044 96688
rect 209096 96676 209102 96688
rect 212166 96676 212172 96688
rect 209096 96648 212172 96676
rect 209096 96636 209102 96648
rect 212166 96636 212172 96648
rect 212224 96636 212230 96688
rect 217410 96636 217416 96688
rect 217468 96676 217474 96688
rect 219986 96676 219992 96688
rect 217468 96648 219992 96676
rect 217468 96636 217474 96648
rect 219986 96636 219992 96648
rect 220044 96636 220050 96688
rect 222194 96636 222200 96688
rect 222252 96676 222258 96688
rect 224034 96676 224040 96688
rect 222252 96648 224040 96676
rect 222252 96636 222258 96648
rect 224034 96636 224040 96648
rect 224092 96636 224098 96688
rect 233970 96636 233976 96688
rect 234028 96676 234034 96688
rect 237558 96676 237564 96688
rect 234028 96648 237564 96676
rect 234028 96636 234034 96648
rect 237558 96636 237564 96648
rect 237616 96636 237622 96688
rect 238018 96636 238024 96688
rect 238076 96676 238082 96688
rect 238938 96676 238944 96688
rect 238076 96648 238944 96676
rect 238076 96636 238082 96648
rect 238938 96636 238944 96648
rect 238996 96636 239002 96688
rect 240134 96636 240140 96688
rect 240192 96676 240198 96688
rect 240962 96676 240968 96688
rect 240192 96648 240968 96676
rect 240192 96636 240198 96648
rect 240962 96636 240968 96648
rect 241020 96636 241026 96688
rect 242250 96636 242256 96688
rect 242308 96676 242314 96688
rect 242802 96676 242808 96688
rect 242308 96648 242808 96676
rect 242308 96636 242314 96648
rect 242802 96636 242808 96648
rect 242860 96636 242866 96688
rect 248874 96636 248880 96688
rect 248932 96676 248938 96688
rect 249518 96676 249524 96688
rect 248932 96648 249524 96676
rect 248932 96636 248938 96648
rect 249518 96636 249524 96648
rect 249576 96636 249582 96688
rect 259546 96636 259552 96688
rect 259604 96676 259610 96688
rect 260742 96676 260748 96688
rect 259604 96648 260748 96676
rect 259604 96636 259610 96648
rect 260742 96636 260748 96648
rect 260800 96636 260806 96688
rect 261662 96636 261668 96688
rect 261720 96676 261726 96688
rect 262122 96676 262128 96688
rect 261720 96648 262128 96676
rect 261720 96636 261726 96648
rect 262122 96636 262128 96648
rect 262180 96636 262186 96688
rect 264146 96636 264152 96688
rect 264204 96676 264210 96688
rect 266998 96676 267004 96688
rect 264204 96648 267004 96676
rect 264204 96636 264210 96648
rect 266998 96636 267004 96648
rect 267056 96636 267062 96688
rect 269390 96636 269396 96688
rect 269448 96676 269454 96688
rect 270402 96676 270408 96688
rect 269448 96648 270408 96676
rect 269448 96636 269454 96648
rect 270402 96636 270408 96648
rect 270460 96636 270466 96688
rect 274082 96636 274088 96688
rect 274140 96676 274146 96688
rect 274542 96676 274548 96688
rect 274140 96648 274548 96676
rect 274140 96636 274146 96648
rect 274542 96636 274548 96648
rect 274600 96636 274606 96688
rect 275094 96636 275100 96688
rect 275152 96676 275158 96688
rect 275738 96676 275744 96688
rect 275152 96648 275744 96676
rect 275152 96636 275158 96648
rect 275738 96636 275744 96648
rect 275796 96636 275802 96688
rect 276934 96636 276940 96688
rect 276992 96676 276998 96688
rect 277302 96676 277308 96688
rect 276992 96648 277308 96676
rect 276992 96636 276998 96648
rect 277302 96636 277308 96648
rect 277360 96636 277366 96688
rect 277486 96636 277492 96688
rect 277544 96676 277550 96688
rect 278314 96676 278320 96688
rect 277544 96648 278320 96676
rect 277544 96636 277550 96648
rect 278314 96636 278320 96648
rect 278372 96636 278378 96688
rect 278406 96636 278412 96688
rect 278464 96676 278470 96688
rect 278682 96676 278688 96688
rect 278464 96648 278688 96676
rect 278464 96636 278470 96648
rect 278682 96636 278688 96648
rect 278740 96636 278746 96688
rect 280706 96636 280712 96688
rect 280764 96676 280770 96688
rect 281166 96676 281172 96688
rect 280764 96648 281172 96676
rect 280764 96636 280770 96648
rect 281166 96636 281172 96648
rect 281224 96636 281230 96688
rect 281534 96636 281540 96688
rect 281592 96676 281598 96688
rect 282822 96676 282828 96688
rect 281592 96648 282828 96676
rect 281592 96636 281598 96648
rect 282822 96636 282828 96648
rect 282880 96636 282886 96688
rect 282914 96636 282920 96688
rect 282972 96676 282978 96688
rect 284110 96676 284116 96688
rect 282972 96648 284116 96676
rect 282972 96636 282978 96648
rect 284110 96636 284116 96648
rect 284168 96636 284174 96688
rect 284294 96636 284300 96688
rect 284352 96676 284358 96688
rect 296622 96676 296628 96688
rect 284352 96648 296628 96676
rect 284352 96636 284358 96648
rect 296622 96636 296628 96648
rect 296680 96636 296686 96688
rect 296732 96676 296760 96920
rect 296806 96772 296812 96824
rect 296864 96812 296870 96824
rect 297634 96812 297640 96824
rect 296864 96784 297640 96812
rect 296864 96772 296870 96784
rect 297634 96772 297640 96784
rect 297692 96772 297698 96824
rect 297744 96744 297772 96920
rect 298646 96908 298652 96960
rect 298704 96948 298710 96960
rect 299014 96948 299020 96960
rect 298704 96920 299020 96948
rect 298704 96908 298710 96920
rect 299014 96908 299020 96920
rect 299072 96908 299078 96960
rect 298462 96840 298468 96892
rect 298520 96880 298526 96892
rect 299198 96880 299204 96892
rect 298520 96852 299204 96880
rect 298520 96840 298526 96852
rect 299198 96840 299204 96852
rect 299256 96840 299262 96892
rect 298278 96772 298284 96824
rect 298336 96812 298342 96824
rect 299382 96812 299388 96824
rect 298336 96784 299388 96812
rect 298336 96772 298342 96784
rect 299382 96772 299388 96784
rect 299440 96772 299446 96824
rect 301498 96744 301504 96756
rect 297744 96716 301504 96744
rect 301498 96704 301504 96716
rect 301556 96704 301562 96756
rect 302878 96676 302884 96688
rect 296732 96648 302884 96676
rect 302878 96636 302884 96648
rect 302936 96636 302942 96688
rect 176562 96568 176568 96620
rect 176620 96608 176626 96620
rect 220170 96608 220176 96620
rect 176620 96580 220176 96608
rect 176620 96568 176626 96580
rect 220170 96568 220176 96580
rect 220228 96568 220234 96620
rect 254670 96568 254676 96620
rect 254728 96608 254734 96620
rect 320174 96608 320180 96620
rect 254728 96580 320180 96608
rect 254728 96568 254734 96580
rect 320174 96568 320180 96580
rect 320232 96568 320238 96620
rect 161382 96500 161388 96552
rect 161440 96540 161446 96552
rect 208302 96540 208308 96552
rect 161440 96512 208308 96540
rect 161440 96500 161446 96512
rect 208302 96500 208308 96512
rect 208360 96500 208366 96552
rect 257522 96500 257528 96552
rect 257580 96540 257586 96552
rect 335998 96540 336004 96552
rect 257580 96512 336004 96540
rect 257580 96500 257586 96512
rect 335998 96500 336004 96512
rect 336056 96500 336062 96552
rect 183462 96432 183468 96484
rect 183520 96472 183526 96484
rect 231118 96472 231124 96484
rect 183520 96444 231124 96472
rect 183520 96432 183526 96444
rect 231118 96432 231124 96444
rect 231176 96432 231182 96484
rect 271046 96432 271052 96484
rect 271104 96472 271110 96484
rect 271230 96472 271236 96484
rect 271104 96444 271236 96472
rect 271104 96432 271110 96444
rect 271230 96432 271236 96444
rect 271288 96432 271294 96484
rect 284938 96432 284944 96484
rect 284996 96472 285002 96484
rect 461578 96472 461584 96484
rect 284996 96444 461584 96472
rect 284996 96432 285002 96444
rect 461578 96432 461584 96444
rect 461636 96432 461642 96484
rect 179322 96364 179328 96416
rect 179380 96404 179386 96416
rect 230474 96404 230480 96416
rect 179380 96376 230480 96404
rect 179380 96364 179386 96376
rect 230474 96364 230480 96376
rect 230532 96364 230538 96416
rect 284386 96364 284392 96416
rect 284444 96404 284450 96416
rect 468478 96404 468484 96416
rect 284444 96376 468484 96404
rect 284444 96364 284450 96376
rect 468478 96364 468484 96376
rect 468536 96364 468542 96416
rect 173158 96296 173164 96348
rect 173216 96336 173222 96348
rect 229278 96336 229284 96348
rect 173216 96308 229284 96336
rect 173216 96296 173222 96308
rect 229278 96296 229284 96308
rect 229336 96296 229342 96348
rect 231118 96296 231124 96348
rect 231176 96336 231182 96348
rect 235350 96336 235356 96348
rect 231176 96308 235356 96336
rect 231176 96296 231182 96308
rect 235350 96296 235356 96308
rect 235408 96296 235414 96348
rect 283742 96296 283748 96348
rect 283800 96336 283806 96348
rect 472618 96336 472624 96348
rect 283800 96308 472624 96336
rect 283800 96296 283806 96308
rect 472618 96296 472624 96308
rect 472676 96296 472682 96348
rect 169662 96228 169668 96280
rect 169720 96268 169726 96280
rect 228726 96268 228732 96280
rect 169720 96240 228732 96268
rect 169720 96228 169726 96240
rect 228726 96228 228732 96240
rect 228784 96228 228790 96280
rect 281902 96228 281908 96280
rect 281960 96268 281966 96280
rect 479518 96268 479524 96280
rect 281960 96240 479524 96268
rect 281960 96228 281966 96240
rect 479518 96228 479524 96240
rect 479576 96228 479582 96280
rect 165522 96160 165528 96212
rect 165580 96200 165586 96212
rect 228082 96200 228088 96212
rect 165580 96172 228088 96200
rect 165580 96160 165586 96172
rect 228082 96160 228088 96172
rect 228140 96160 228146 96212
rect 283098 96160 283104 96212
rect 283156 96200 283162 96212
rect 475378 96200 475384 96212
rect 283156 96172 475384 96200
rect 283156 96160 283162 96172
rect 475378 96160 475384 96172
rect 475436 96160 475442 96212
rect 133782 96092 133788 96144
rect 133840 96132 133846 96144
rect 211154 96132 211160 96144
rect 133840 96104 211160 96132
rect 133840 96092 133846 96104
rect 211154 96092 211160 96104
rect 211212 96092 211218 96144
rect 282546 96092 282552 96144
rect 282604 96132 282610 96144
rect 483014 96132 483020 96144
rect 282604 96104 483020 96132
rect 282604 96092 282610 96104
rect 483014 96092 483020 96104
rect 483072 96092 483078 96144
rect 131022 96024 131028 96076
rect 131080 96064 131086 96076
rect 222286 96064 222292 96076
rect 131080 96036 222292 96064
rect 131080 96024 131086 96036
rect 222286 96024 222292 96036
rect 222344 96024 222350 96076
rect 285582 96024 285588 96076
rect 285640 96064 285646 96076
rect 500954 96064 500960 96076
rect 285640 96036 500960 96064
rect 285640 96024 285646 96036
rect 500954 96024 500960 96036
rect 501012 96024 501018 96076
rect 54478 95956 54484 96008
rect 54536 95996 54542 96008
rect 208670 95996 208676 96008
rect 54536 95968 208676 95996
rect 54536 95956 54542 95968
rect 208670 95956 208676 95968
rect 208728 95956 208734 96008
rect 245010 95956 245016 96008
rect 245068 95996 245074 96008
rect 267826 95996 267832 96008
rect 245068 95968 267832 95996
rect 245068 95956 245074 95968
rect 267826 95956 267832 95968
rect 267884 95956 267890 96008
rect 286134 95956 286140 96008
rect 286192 95996 286198 96008
rect 502978 95996 502984 96008
rect 286192 95968 502984 95996
rect 286192 95956 286198 95968
rect 502978 95956 502984 95968
rect 503036 95956 503042 96008
rect 17218 95888 17224 95940
rect 17276 95928 17282 95940
rect 202046 95928 202052 95940
rect 17276 95900 202052 95928
rect 17276 95888 17282 95900
rect 202046 95888 202052 95900
rect 202104 95888 202110 95940
rect 228358 95888 228364 95940
rect 228416 95928 228422 95940
rect 237466 95928 237472 95940
rect 228416 95900 237472 95928
rect 228416 95888 228422 95900
rect 237466 95888 237472 95900
rect 237524 95888 237530 95940
rect 248046 95888 248052 95940
rect 248104 95928 248110 95940
rect 284386 95928 284392 95940
rect 248104 95900 284392 95928
rect 248104 95888 248110 95900
rect 284386 95888 284392 95900
rect 284444 95888 284450 95940
rect 294322 95888 294328 95940
rect 294380 95928 294386 95940
rect 295058 95928 295064 95940
rect 294380 95900 295064 95928
rect 294380 95888 294386 95900
rect 295058 95888 295064 95900
rect 295116 95888 295122 95940
rect 295334 95888 295340 95940
rect 295392 95928 295398 95940
rect 511994 95928 512000 95940
rect 295392 95900 512000 95928
rect 295392 95888 295398 95900
rect 511994 95888 512000 95900
rect 512052 95888 512058 95940
rect 186958 95820 186964 95872
rect 187016 95860 187022 95872
rect 231762 95860 231768 95872
rect 187016 95832 231768 95860
rect 187016 95820 187022 95832
rect 231762 95820 231768 95832
rect 231820 95820 231826 95872
rect 253474 95820 253480 95872
rect 253532 95860 253538 95872
rect 313274 95860 313280 95872
rect 253532 95832 313280 95860
rect 253532 95820 253538 95832
rect 313274 95820 313280 95832
rect 313332 95820 313338 95872
rect 191098 95752 191104 95804
rect 191156 95792 191162 95804
rect 232314 95792 232320 95804
rect 191156 95764 232320 95792
rect 191156 95752 191162 95764
rect 232314 95752 232320 95764
rect 232372 95752 232378 95804
rect 251266 95752 251272 95804
rect 251324 95792 251330 95804
rect 302326 95792 302332 95804
rect 251324 95764 302332 95792
rect 251324 95752 251330 95764
rect 302326 95752 302332 95764
rect 302384 95752 302390 95804
rect 197262 95684 197268 95736
rect 197320 95724 197326 95736
rect 233510 95724 233516 95736
rect 197320 95696 233516 95724
rect 197320 95684 197326 95696
rect 233510 95684 233516 95696
rect 233568 95684 233574 95736
rect 251082 95684 251088 95736
rect 251140 95724 251146 95736
rect 299658 95724 299664 95736
rect 251140 95696 299664 95724
rect 251140 95684 251146 95696
rect 299658 95684 299664 95696
rect 299716 95684 299722 95736
rect 200022 95616 200028 95668
rect 200080 95656 200086 95668
rect 234154 95656 234160 95668
rect 200080 95628 234160 95656
rect 200080 95616 200086 95628
rect 234154 95616 234160 95628
rect 234212 95616 234218 95668
rect 263594 95616 263600 95668
rect 263652 95656 263658 95668
rect 299474 95656 299480 95668
rect 263652 95628 299480 95656
rect 263652 95616 263658 95628
rect 299474 95616 299480 95628
rect 299532 95616 299538 95668
rect 194502 95548 194508 95600
rect 194560 95588 194566 95600
rect 213914 95588 213920 95600
rect 194560 95560 213920 95588
rect 194560 95548 194566 95560
rect 213914 95548 213920 95560
rect 213972 95548 213978 95600
rect 249886 95548 249892 95600
rect 249944 95588 249950 95600
rect 299566 95588 299572 95600
rect 249944 95560 299572 95588
rect 249944 95548 249950 95560
rect 299566 95548 299572 95560
rect 299624 95548 299630 95600
rect 287330 95480 287336 95532
rect 287388 95520 287394 95532
rect 295334 95520 295340 95532
rect 287388 95492 295340 95520
rect 287388 95480 287394 95492
rect 295334 95480 295340 95492
rect 295392 95480 295398 95532
rect 235902 95276 235908 95328
rect 235960 95316 235966 95328
rect 240226 95316 240232 95328
rect 235960 95288 240232 95316
rect 235960 95276 235966 95288
rect 240226 95276 240232 95288
rect 240284 95276 240290 95328
rect 210510 95208 210516 95260
rect 210568 95248 210574 95260
rect 210694 95248 210700 95260
rect 210568 95220 210700 95248
rect 210568 95208 210574 95220
rect 210694 95208 210700 95220
rect 210752 95208 210758 95260
rect 238110 95208 238116 95260
rect 238168 95248 238174 95260
rect 239398 95248 239404 95260
rect 238168 95220 239404 95248
rect 238168 95208 238174 95220
rect 239398 95208 239404 95220
rect 239456 95208 239462 95260
rect 171042 95140 171048 95192
rect 171100 95180 171106 95192
rect 229094 95180 229100 95192
rect 171100 95152 229100 95180
rect 171100 95140 171106 95152
rect 229094 95140 229100 95152
rect 229152 95140 229158 95192
rect 261386 95140 261392 95192
rect 261444 95180 261450 95192
rect 358814 95180 358820 95192
rect 261444 95152 358820 95180
rect 261444 95140 261450 95152
rect 358814 95140 358820 95152
rect 358872 95140 358878 95192
rect 162762 95072 162768 95124
rect 162820 95112 162826 95124
rect 227714 95112 227720 95124
rect 162820 95084 227720 95112
rect 162820 95072 162826 95084
rect 227714 95072 227720 95084
rect 227772 95072 227778 95124
rect 295978 95072 295984 95124
rect 296036 95112 296042 95124
rect 465718 95112 465724 95124
rect 296036 95084 465724 95112
rect 296036 95072 296042 95084
rect 465718 95072 465724 95084
rect 465776 95072 465782 95124
rect 147582 95004 147588 95056
rect 147640 95044 147646 95056
rect 212534 95044 212540 95056
rect 147640 95016 212540 95044
rect 147640 95004 147646 95016
rect 212534 95004 212540 95016
rect 212592 95004 212598 95056
rect 293310 95004 293316 95056
rect 293368 95044 293374 95056
rect 485038 95044 485044 95056
rect 293368 95016 485044 95044
rect 293368 95004 293374 95016
rect 485038 95004 485044 95016
rect 485096 95004 485102 95056
rect 159358 94936 159364 94988
rect 159416 94976 159422 94988
rect 226886 94976 226892 94988
rect 159416 94948 226892 94976
rect 159416 94936 159422 94948
rect 226886 94936 226892 94948
rect 226944 94936 226950 94988
rect 288250 94936 288256 94988
rect 288308 94976 288314 94988
rect 489178 94976 489184 94988
rect 288308 94948 489184 94976
rect 288308 94936 288314 94948
rect 489178 94936 489184 94948
rect 489236 94936 489242 94988
rect 155310 94868 155316 94920
rect 155368 94908 155374 94920
rect 226242 94908 226248 94920
rect 155368 94880 226248 94908
rect 155368 94868 155374 94880
rect 226242 94868 226248 94880
rect 226300 94868 226306 94920
rect 286962 94868 286968 94920
rect 287020 94908 287026 94920
rect 507854 94908 507860 94920
rect 287020 94880 507860 94908
rect 287020 94868 287026 94880
rect 507854 94868 507860 94880
rect 507912 94868 507918 94920
rect 144822 94800 144828 94852
rect 144880 94840 144886 94852
rect 224494 94840 224500 94852
rect 144880 94812 224500 94840
rect 144880 94800 144886 94812
rect 224494 94800 224500 94812
rect 224552 94800 224558 94852
rect 230382 94800 230388 94852
rect 230440 94840 230446 94852
rect 237374 94840 237380 94852
rect 230440 94812 237380 94840
rect 230440 94800 230446 94812
rect 237374 94800 237380 94812
rect 237432 94800 237438 94852
rect 292482 94800 292488 94852
rect 292540 94840 292546 94852
rect 519538 94840 519544 94852
rect 292540 94812 519544 94840
rect 292540 94800 292546 94812
rect 519538 94800 519544 94812
rect 519596 94800 519602 94852
rect 137278 94732 137284 94784
rect 137336 94772 137342 94784
rect 223298 94772 223304 94784
rect 137336 94744 223304 94772
rect 137336 94732 137342 94744
rect 223298 94732 223304 94744
rect 223356 94732 223362 94784
rect 290366 94732 290372 94784
rect 290424 94772 290430 94784
rect 529934 94772 529940 94784
rect 290424 94744 529940 94772
rect 290424 94732 290430 94744
rect 529934 94732 529940 94744
rect 529992 94732 529998 94784
rect 128262 94664 128268 94716
rect 128320 94704 128326 94716
rect 221642 94704 221648 94716
rect 128320 94676 221648 94704
rect 128320 94664 128326 94676
rect 221642 94664 221648 94676
rect 221700 94664 221706 94716
rect 234982 94664 234988 94716
rect 235040 94704 235046 94716
rect 235166 94704 235172 94716
rect 235040 94676 235172 94704
rect 235040 94664 235046 94676
rect 235166 94664 235172 94676
rect 235224 94664 235230 94716
rect 291010 94664 291016 94716
rect 291068 94704 291074 94716
rect 532694 94704 532700 94716
rect 291068 94676 532700 94704
rect 291068 94664 291074 94676
rect 532694 94664 532700 94676
rect 532752 94664 532758 94716
rect 121362 94596 121368 94648
rect 121420 94636 121426 94648
rect 220630 94636 220636 94648
rect 121420 94608 220636 94636
rect 121420 94596 121426 94608
rect 220630 94596 220636 94608
rect 220688 94596 220694 94648
rect 232130 94596 232136 94648
rect 232188 94636 232194 94648
rect 232406 94636 232412 94648
rect 232188 94608 232412 94636
rect 232188 94596 232194 94608
rect 232406 94596 232412 94608
rect 232464 94596 232470 94648
rect 236362 94636 236368 94648
rect 234586 94608 236368 94636
rect 101398 94528 101404 94580
rect 101456 94568 101462 94580
rect 212810 94568 212816 94580
rect 101456 94540 212816 94568
rect 101456 94528 101462 94540
rect 212810 94528 212816 94540
rect 212868 94528 212874 94580
rect 212902 94528 212908 94580
rect 212960 94568 212966 94580
rect 213086 94568 213092 94580
rect 212960 94540 213092 94568
rect 212960 94528 212966 94540
rect 213086 94528 213092 94540
rect 213144 94528 213150 94580
rect 216122 94528 216128 94580
rect 216180 94568 216186 94580
rect 216490 94568 216496 94580
rect 216180 94540 216496 94568
rect 216180 94528 216186 94540
rect 216490 94528 216496 94540
rect 216548 94528 216554 94580
rect 216950 94528 216956 94580
rect 217008 94568 217014 94580
rect 217318 94568 217324 94580
rect 217008 94540 217324 94568
rect 217008 94528 217014 94540
rect 217318 94528 217324 94540
rect 217376 94528 217382 94580
rect 218514 94528 218520 94580
rect 218572 94568 218578 94580
rect 218882 94568 218888 94580
rect 218572 94540 218888 94568
rect 218572 94528 218578 94540
rect 218882 94528 218888 94540
rect 218940 94528 218946 94580
rect 219710 94528 219716 94580
rect 219768 94568 219774 94580
rect 220354 94568 220360 94580
rect 219768 94540 220360 94568
rect 219768 94528 219774 94540
rect 220354 94528 220360 94540
rect 220412 94528 220418 94580
rect 220906 94528 220912 94580
rect 220964 94568 220970 94580
rect 221550 94568 221556 94580
rect 220964 94540 221556 94568
rect 220964 94528 220970 94540
rect 221550 94528 221556 94540
rect 221608 94528 221614 94580
rect 228450 94528 228456 94580
rect 228508 94568 228514 94580
rect 234586 94568 234614 94608
rect 236362 94596 236368 94608
rect 236420 94596 236426 94648
rect 291562 94596 291568 94648
rect 291620 94636 291626 94648
rect 536834 94636 536840 94648
rect 291620 94608 536840 94636
rect 291620 94596 291626 94608
rect 536834 94596 536840 94608
rect 536892 94596 536898 94648
rect 228508 94540 234614 94568
rect 228508 94528 228514 94540
rect 234798 94528 234804 94580
rect 234856 94568 234862 94580
rect 235442 94568 235448 94580
rect 234856 94540 235448 94568
rect 234856 94528 234862 94540
rect 235442 94528 235448 94540
rect 235500 94528 235506 94580
rect 236638 94528 236644 94580
rect 236696 94568 236702 94580
rect 237098 94568 237104 94580
rect 236696 94540 237104 94568
rect 236696 94528 236702 94540
rect 237098 94528 237104 94540
rect 237156 94528 237162 94580
rect 239122 94528 239128 94580
rect 239180 94568 239186 94580
rect 239674 94568 239680 94580
rect 239180 94540 239680 94568
rect 239180 94528 239186 94540
rect 239674 94528 239680 94540
rect 239732 94528 239738 94580
rect 240318 94528 240324 94580
rect 240376 94568 240382 94580
rect 240686 94568 240692 94580
rect 240376 94540 240692 94568
rect 240376 94528 240382 94540
rect 240686 94528 240692 94540
rect 240744 94528 240750 94580
rect 278038 94528 278044 94580
rect 278096 94568 278102 94580
rect 278406 94568 278412 94580
rect 278096 94540 278412 94568
rect 278096 94528 278102 94540
rect 278406 94528 278412 94540
rect 278464 94528 278470 94580
rect 292850 94528 292856 94580
rect 292908 94568 292914 94580
rect 543734 94568 543740 94580
rect 292908 94540 543740 94568
rect 292908 94528 292914 94540
rect 543734 94528 543740 94540
rect 543792 94528 543798 94580
rect 29638 94460 29644 94512
rect 29696 94500 29702 94512
rect 199838 94500 199844 94512
rect 29696 94472 199844 94500
rect 29696 94460 29702 94472
rect 199838 94460 199844 94472
rect 199896 94460 199902 94512
rect 200206 94460 200212 94512
rect 200264 94500 200270 94512
rect 200574 94500 200580 94512
rect 200264 94472 200580 94500
rect 200264 94460 200270 94472
rect 200574 94460 200580 94472
rect 200632 94460 200638 94512
rect 201770 94460 201776 94512
rect 201828 94500 201834 94512
rect 202598 94500 202604 94512
rect 201828 94472 202604 94500
rect 201828 94460 201834 94472
rect 202598 94460 202604 94472
rect 202656 94460 202662 94512
rect 204438 94460 204444 94512
rect 204496 94500 204502 94512
rect 205174 94500 205180 94512
rect 204496 94472 205180 94500
rect 204496 94460 204502 94472
rect 205174 94460 205180 94472
rect 205232 94460 205238 94512
rect 212718 94460 212724 94512
rect 212776 94500 212782 94512
rect 213270 94500 213276 94512
rect 212776 94472 213276 94500
rect 212776 94460 212782 94472
rect 213270 94460 213276 94472
rect 213328 94460 213334 94512
rect 217134 94460 217140 94512
rect 217192 94500 217198 94512
rect 217686 94500 217692 94512
rect 217192 94472 217692 94500
rect 217192 94460 217198 94472
rect 217686 94460 217692 94472
rect 217744 94460 217750 94512
rect 221090 94460 221096 94512
rect 221148 94500 221154 94512
rect 221918 94500 221924 94512
rect 221148 94472 221924 94500
rect 221148 94460 221154 94472
rect 221918 94460 221924 94472
rect 221976 94460 221982 94512
rect 232038 94460 232044 94512
rect 232096 94500 232102 94512
rect 232406 94500 232412 94512
rect 232096 94472 232412 94500
rect 232096 94460 232102 94472
rect 232406 94460 232412 94472
rect 232464 94460 232470 94512
rect 241606 94460 241612 94512
rect 241664 94500 241670 94512
rect 242526 94500 242532 94512
rect 241664 94472 242532 94500
rect 241664 94460 241670 94472
rect 242526 94460 242532 94472
rect 242584 94460 242590 94512
rect 243630 94460 243636 94512
rect 243688 94500 243694 94512
rect 244090 94500 244096 94512
rect 243688 94472 244096 94500
rect 243688 94460 243694 94472
rect 244090 94460 244096 94472
rect 244148 94460 244154 94512
rect 247034 94460 247040 94512
rect 247092 94500 247098 94512
rect 264238 94500 264244 94512
rect 247092 94472 264244 94500
rect 247092 94460 247098 94472
rect 264238 94460 264244 94472
rect 264296 94460 264302 94512
rect 278222 94460 278228 94512
rect 278280 94500 278286 94512
rect 278590 94500 278596 94512
rect 278280 94472 278596 94500
rect 278280 94460 278286 94472
rect 278590 94460 278596 94472
rect 278648 94460 278654 94512
rect 297266 94460 297272 94512
rect 297324 94500 297330 94512
rect 565078 94500 565084 94512
rect 297324 94472 565084 94500
rect 297324 94460 297330 94472
rect 565078 94460 565084 94472
rect 565136 94460 565142 94512
rect 173802 94392 173808 94444
rect 173860 94432 173866 94444
rect 229462 94432 229468 94444
rect 173860 94404 229468 94432
rect 173860 94392 173866 94404
rect 229462 94392 229468 94404
rect 229520 94392 229526 94444
rect 255314 94392 255320 94444
rect 255372 94432 255378 94444
rect 324406 94432 324412 94444
rect 255372 94404 324412 94432
rect 255372 94392 255378 94404
rect 324406 94392 324412 94404
rect 324464 94392 324470 94444
rect 188338 94324 188344 94376
rect 188396 94364 188402 94376
rect 231486 94364 231492 94376
rect 188396 94336 231492 94364
rect 188396 94324 188402 94336
rect 231486 94324 231492 94336
rect 231544 94324 231550 94376
rect 252922 94324 252928 94376
rect 252980 94364 252986 94376
rect 309134 94364 309140 94376
rect 252980 94336 309140 94364
rect 252980 94324 252986 94336
rect 309134 94324 309140 94336
rect 309192 94324 309198 94376
rect 200206 94256 200212 94308
rect 200264 94296 200270 94308
rect 201126 94296 201132 94308
rect 200264 94268 201132 94296
rect 200264 94256 200270 94268
rect 201126 94256 201132 94268
rect 201184 94256 201190 94308
rect 233694 94296 233700 94308
rect 205606 94268 233700 94296
rect 198642 94188 198648 94240
rect 198700 94228 198706 94240
rect 205606 94228 205634 94268
rect 233694 94256 233700 94268
rect 233752 94256 233758 94308
rect 252370 94256 252376 94308
rect 252428 94296 252434 94308
rect 306374 94296 306380 94308
rect 252428 94268 306380 94296
rect 252428 94256 252434 94268
rect 306374 94256 306380 94268
rect 306432 94256 306438 94308
rect 198700 94200 205634 94228
rect 198700 94188 198706 94200
rect 212626 94188 212632 94240
rect 212684 94228 212690 94240
rect 213454 94228 213460 94240
rect 212684 94200 213460 94228
rect 212684 94188 212690 94200
rect 213454 94188 213460 94200
rect 213512 94188 213518 94240
rect 218054 94188 218060 94240
rect 218112 94228 218118 94240
rect 218330 94228 218336 94240
rect 218112 94200 218336 94228
rect 218112 94188 218118 94200
rect 218330 94188 218336 94200
rect 218388 94188 218394 94240
rect 263870 94188 263876 94240
rect 263928 94228 263934 94240
rect 316034 94228 316040 94240
rect 263928 94200 316040 94228
rect 263928 94188 263934 94200
rect 316034 94188 316040 94200
rect 316092 94188 316098 94240
rect 199838 94120 199844 94172
rect 199896 94160 199902 94172
rect 203702 94160 203708 94172
rect 199896 94132 203708 94160
rect 199896 94120 199902 94132
rect 203702 94120 203708 94132
rect 203760 94120 203766 94172
rect 212718 94120 212724 94172
rect 212776 94160 212782 94172
rect 213638 94160 213644 94172
rect 212776 94132 213644 94160
rect 212776 94120 212782 94132
rect 213638 94120 213644 94132
rect 213696 94120 213702 94172
rect 251726 94120 251732 94172
rect 251784 94160 251790 94172
rect 302234 94160 302240 94172
rect 251784 94132 302240 94160
rect 251784 94120 251790 94132
rect 302234 94120 302240 94132
rect 302292 94120 302298 94172
rect 170398 93780 170404 93832
rect 170456 93820 170462 93832
rect 170456 93792 228404 93820
rect 170456 93780 170462 93792
rect 166902 93712 166908 93764
rect 166960 93752 166966 93764
rect 228266 93752 228272 93764
rect 166960 93724 228272 93752
rect 166960 93712 166966 93724
rect 228266 93712 228272 93724
rect 228324 93712 228330 93764
rect 228376 93752 228404 93792
rect 228542 93780 228548 93832
rect 228600 93820 228606 93832
rect 234246 93820 234252 93832
rect 228600 93792 234252 93820
rect 228600 93780 228606 93792
rect 234246 93780 234252 93792
rect 234304 93780 234310 93832
rect 257706 93780 257712 93832
rect 257764 93820 257770 93832
rect 338114 93820 338120 93832
rect 257764 93792 338120 93820
rect 257764 93780 257770 93792
rect 338114 93780 338120 93792
rect 338172 93780 338178 93832
rect 228818 93752 228824 93764
rect 228376 93724 228824 93752
rect 228818 93712 228824 93724
rect 228876 93712 228882 93764
rect 262030 93712 262036 93764
rect 262088 93752 262094 93764
rect 362954 93752 362960 93764
rect 262088 93724 362960 93752
rect 262088 93712 262094 93724
rect 362954 93712 362960 93724
rect 363012 93712 363018 93764
rect 160002 93644 160008 93696
rect 160060 93684 160066 93696
rect 226978 93684 226984 93696
rect 160060 93656 226984 93684
rect 160060 93644 160066 93656
rect 226978 93644 226984 93656
rect 227036 93644 227042 93696
rect 266262 93644 266268 93696
rect 266320 93684 266326 93696
rect 382918 93684 382924 93696
rect 266320 93656 382924 93684
rect 266320 93644 266326 93656
rect 382918 93644 382924 93656
rect 382976 93644 382982 93696
rect 153102 93576 153108 93628
rect 153160 93616 153166 93628
rect 225782 93616 225788 93628
rect 153160 93588 225788 93616
rect 153160 93576 153166 93588
rect 225782 93576 225788 93588
rect 225840 93576 225846 93628
rect 270402 93576 270408 93628
rect 270460 93616 270466 93628
rect 407206 93616 407212 93628
rect 270460 93588 407212 93616
rect 270460 93576 270466 93588
rect 407206 93576 407212 93588
rect 407264 93576 407270 93628
rect 145558 93508 145564 93560
rect 145616 93548 145622 93560
rect 224586 93548 224592 93560
rect 145616 93520 224592 93548
rect 145616 93508 145622 93520
rect 224586 93508 224592 93520
rect 224644 93508 224650 93560
rect 277762 93508 277768 93560
rect 277820 93548 277826 93560
rect 454770 93548 454776 93560
rect 277820 93520 454776 93548
rect 277820 93508 277826 93520
rect 454770 93508 454776 93520
rect 454828 93508 454834 93560
rect 142062 93440 142068 93492
rect 142120 93480 142126 93492
rect 222194 93480 222200 93492
rect 142120 93452 222200 93480
rect 142120 93440 142126 93452
rect 222194 93440 222200 93452
rect 222252 93440 222258 93492
rect 293402 93440 293408 93492
rect 293460 93480 293466 93492
rect 542998 93480 543004 93492
rect 293460 93452 543004 93480
rect 293460 93440 293466 93452
rect 542998 93440 543004 93452
rect 543056 93440 543062 93492
rect 136542 93372 136548 93424
rect 136600 93412 136606 93424
rect 219434 93412 219440 93424
rect 136600 93384 219440 93412
rect 136600 93372 136606 93384
rect 219434 93372 219440 93384
rect 219492 93372 219498 93424
rect 295242 93372 295248 93424
rect 295300 93412 295306 93424
rect 554774 93412 554780 93424
rect 295300 93384 554780 93412
rect 295300 93372 295306 93384
rect 554774 93372 554780 93384
rect 554832 93372 554838 93424
rect 135162 93304 135168 93356
rect 135220 93344 135226 93356
rect 222746 93344 222752 93356
rect 135220 93316 222752 93344
rect 135220 93304 135226 93316
rect 222746 93304 222752 93316
rect 222804 93304 222810 93356
rect 295150 93304 295156 93356
rect 295208 93344 295214 93356
rect 557534 93344 557540 93356
rect 295208 93316 557540 93344
rect 295208 93304 295214 93316
rect 557534 93304 557540 93316
rect 557592 93304 557598 93356
rect 61378 93236 61384 93288
rect 61436 93276 61442 93288
rect 209222 93276 209228 93288
rect 61436 93248 209228 93276
rect 61436 93236 61442 93248
rect 209222 93236 209228 93248
rect 209280 93236 209286 93288
rect 296530 93236 296536 93288
rect 296588 93276 296594 93288
rect 561674 93276 561680 93288
rect 296588 93248 561680 93276
rect 296588 93236 296594 93248
rect 561674 93236 561680 93248
rect 561732 93236 561738 93288
rect 36538 93168 36544 93220
rect 36596 93208 36602 93220
rect 204990 93208 204996 93220
rect 36596 93180 204996 93208
rect 36596 93168 36602 93180
rect 204990 93168 204996 93180
rect 205048 93168 205054 93220
rect 246850 93168 246856 93220
rect 246908 93208 246914 93220
rect 257338 93208 257344 93220
rect 246908 93180 257344 93208
rect 246908 93168 246914 93180
rect 257338 93168 257344 93180
rect 257396 93168 257402 93220
rect 298002 93168 298008 93220
rect 298060 93208 298066 93220
rect 572806 93208 572812 93220
rect 298060 93180 572812 93208
rect 298060 93168 298066 93180
rect 572806 93168 572812 93180
rect 572864 93168 572870 93220
rect 15838 93100 15844 93152
rect 15896 93140 15902 93152
rect 201586 93140 201592 93152
rect 15896 93112 201592 93140
rect 15896 93100 15902 93112
rect 201586 93100 201592 93112
rect 201644 93100 201650 93152
rect 243906 93100 243912 93152
rect 243964 93140 243970 93152
rect 255958 93140 255964 93152
rect 243964 93112 255964 93140
rect 243964 93100 243970 93112
rect 255958 93100 255964 93112
rect 256016 93100 256022 93152
rect 299382 93100 299388 93152
rect 299440 93140 299446 93152
rect 575474 93140 575480 93152
rect 299440 93112 575480 93140
rect 299440 93100 299446 93112
rect 575474 93100 575480 93112
rect 575532 93100 575538 93152
rect 177942 93032 177948 93084
rect 178000 93072 178006 93084
rect 230014 93072 230020 93084
rect 178000 93044 230020 93072
rect 178000 93032 178006 93044
rect 230014 93032 230020 93044
rect 230072 93032 230078 93084
rect 257246 93032 257252 93084
rect 257304 93072 257310 93084
rect 333974 93072 333980 93084
rect 257304 93044 333980 93072
rect 257304 93032 257310 93044
rect 333974 93032 333980 93044
rect 334032 93032 334038 93084
rect 180702 92964 180708 93016
rect 180760 93004 180766 93016
rect 230750 93004 230756 93016
rect 180760 92976 230756 93004
rect 180760 92964 180766 92976
rect 230750 92964 230756 92976
rect 230808 92964 230814 93016
rect 256050 92964 256056 93016
rect 256108 93004 256114 93016
rect 331214 93004 331220 93016
rect 256108 92976 331220 93004
rect 256108 92964 256114 92976
rect 331214 92964 331220 92976
rect 331272 92964 331278 93016
rect 184842 92896 184848 92948
rect 184900 92936 184906 92948
rect 231394 92936 231400 92948
rect 184900 92908 231400 92936
rect 184900 92896 184906 92908
rect 231394 92896 231400 92908
rect 231452 92896 231458 92948
rect 256602 92896 256608 92948
rect 256660 92936 256666 92948
rect 327074 92936 327080 92948
rect 256660 92908 327080 92936
rect 256660 92896 256666 92908
rect 327074 92896 327080 92908
rect 327132 92896 327138 92948
rect 195882 92828 195888 92880
rect 195940 92868 195946 92880
rect 233142 92868 233148 92880
rect 195940 92840 233148 92868
rect 195940 92828 195946 92840
rect 233142 92828 233148 92840
rect 233200 92828 233206 92880
rect 229738 92556 229744 92608
rect 229796 92596 229802 92608
rect 236822 92596 236828 92608
rect 229796 92568 236828 92596
rect 229796 92556 229802 92568
rect 236822 92556 236828 92568
rect 236880 92556 236886 92608
rect 231210 92488 231216 92540
rect 231268 92528 231274 92540
rect 235626 92528 235632 92540
rect 231268 92500 235632 92528
rect 231268 92488 231274 92500
rect 235626 92488 235632 92500
rect 235684 92488 235690 92540
rect 175182 92420 175188 92472
rect 175240 92460 175246 92472
rect 229646 92460 229652 92472
rect 175240 92432 229652 92460
rect 175240 92420 175246 92432
rect 229646 92420 229652 92432
rect 229704 92420 229710 92472
rect 238202 92420 238208 92472
rect 238260 92460 238266 92472
rect 239858 92460 239864 92472
rect 238260 92432 239864 92460
rect 238260 92420 238266 92432
rect 239858 92420 239864 92432
rect 239916 92420 239922 92472
rect 263318 92420 263324 92472
rect 263376 92460 263382 92472
rect 364978 92460 364984 92472
rect 263376 92432 364984 92460
rect 263376 92420 263382 92432
rect 364978 92420 364984 92432
rect 365036 92420 365042 92472
rect 169018 92352 169024 92404
rect 169076 92392 169082 92404
rect 228634 92392 228640 92404
rect 169076 92364 228640 92392
rect 169076 92352 169082 92364
rect 228634 92352 228640 92364
rect 228692 92352 228698 92404
rect 263226 92352 263232 92404
rect 263284 92392 263290 92404
rect 369854 92392 369860 92404
rect 263284 92364 369860 92392
rect 263284 92352 263290 92364
rect 369854 92352 369860 92364
rect 369912 92352 369918 92404
rect 164142 92284 164148 92336
rect 164200 92324 164206 92336
rect 227990 92324 227996 92336
rect 164200 92296 227996 92324
rect 164200 92284 164206 92296
rect 227990 92284 227996 92296
rect 228048 92284 228054 92336
rect 264606 92284 264612 92336
rect 264664 92324 264670 92336
rect 373994 92324 374000 92336
rect 264664 92296 374000 92324
rect 264664 92284 264670 92296
rect 373994 92284 374000 92296
rect 374052 92284 374058 92336
rect 156598 92216 156604 92268
rect 156656 92256 156662 92268
rect 226518 92256 226524 92268
rect 156656 92228 226524 92256
rect 156656 92216 156662 92228
rect 226518 92216 226524 92228
rect 226576 92216 226582 92268
rect 268194 92216 268200 92268
rect 268252 92256 268258 92268
rect 380894 92256 380900 92268
rect 268252 92228 380900 92256
rect 268252 92216 268258 92228
rect 380894 92216 380900 92228
rect 380952 92216 380958 92268
rect 148962 92148 148968 92200
rect 149020 92188 149026 92200
rect 223574 92188 223580 92200
rect 149020 92160 223580 92188
rect 149020 92148 149026 92160
rect 223574 92148 223580 92160
rect 223632 92148 223638 92200
rect 265986 92148 265992 92200
rect 266044 92188 266050 92200
rect 385678 92188 385684 92200
rect 266044 92160 385684 92188
rect 266044 92148 266050 92160
rect 385678 92148 385684 92160
rect 385736 92148 385742 92200
rect 137922 92080 137928 92132
rect 137980 92120 137986 92132
rect 223390 92120 223396 92132
rect 137980 92092 223396 92120
rect 137980 92080 137986 92092
rect 223390 92080 223396 92092
rect 223448 92080 223454 92132
rect 267642 92080 267648 92132
rect 267700 92120 267706 92132
rect 396074 92120 396080 92132
rect 267700 92092 396080 92120
rect 267700 92080 267706 92092
rect 396074 92080 396080 92092
rect 396132 92080 396138 92132
rect 128170 92012 128176 92064
rect 128228 92052 128234 92064
rect 221734 92052 221740 92064
rect 128228 92024 221740 92052
rect 128228 92012 128234 92024
rect 221734 92012 221740 92024
rect 221792 92012 221798 92064
rect 275646 92012 275652 92064
rect 275704 92052 275710 92064
rect 428458 92052 428464 92064
rect 275704 92024 428464 92052
rect 275704 92012 275710 92024
rect 428458 92012 428464 92024
rect 428516 92012 428522 92064
rect 84102 91944 84108 91996
rect 84160 91984 84166 91996
rect 214190 91984 214196 91996
rect 84160 91956 214196 91984
rect 84160 91944 84166 91956
rect 214190 91944 214196 91956
rect 214248 91944 214254 91996
rect 250254 91944 250260 91996
rect 250312 91984 250318 91996
rect 251266 91984 251272 91996
rect 250312 91956 251272 91984
rect 250312 91944 250318 91956
rect 251266 91944 251272 91956
rect 251324 91944 251330 91996
rect 274542 91944 274548 91996
rect 274600 91984 274606 91996
rect 432598 91984 432604 91996
rect 274600 91956 432604 91984
rect 274600 91944 274606 91956
rect 432598 91944 432604 91956
rect 432656 91944 432662 91996
rect 70302 91876 70308 91928
rect 70360 91916 70366 91928
rect 211706 91916 211712 91928
rect 70360 91888 211712 91916
rect 70360 91876 70366 91888
rect 211706 91876 211712 91888
rect 211764 91876 211770 91928
rect 276842 91876 276848 91928
rect 276900 91916 276906 91928
rect 446398 91916 446404 91928
rect 276900 91888 446404 91916
rect 276900 91876 276906 91888
rect 446398 91876 446404 91888
rect 446456 91876 446462 91928
rect 66162 91808 66168 91860
rect 66220 91848 66226 91860
rect 211430 91848 211436 91860
rect 66220 91820 211436 91848
rect 66220 91808 66226 91820
rect 211430 91808 211436 91820
rect 211488 91808 211494 91860
rect 279602 91808 279608 91860
rect 279660 91848 279666 91860
rect 464338 91848 464344 91860
rect 279660 91820 464344 91848
rect 279660 91808 279666 91820
rect 464338 91808 464344 91820
rect 464396 91808 464402 91860
rect 45462 91740 45468 91792
rect 45520 91780 45526 91792
rect 204254 91780 204260 91792
rect 45520 91752 204260 91780
rect 45520 91740 45526 91752
rect 204254 91740 204260 91752
rect 204312 91740 204318 91792
rect 224862 91740 224868 91792
rect 224920 91780 224926 91792
rect 238478 91780 238484 91792
rect 224920 91752 238484 91780
rect 224920 91740 224926 91752
rect 238478 91740 238484 91752
rect 238536 91740 238542 91792
rect 246942 91740 246948 91792
rect 247000 91780 247006 91792
rect 264330 91780 264336 91792
rect 247000 91752 264336 91780
rect 247000 91740 247006 91752
rect 264330 91740 264336 91752
rect 264388 91740 264394 91792
rect 289722 91740 289728 91792
rect 289780 91780 289786 91792
rect 520274 91780 520280 91792
rect 289780 91752 520280 91780
rect 289780 91740 289786 91752
rect 520274 91740 520280 91752
rect 520332 91740 520338 91792
rect 182082 91672 182088 91724
rect 182140 91712 182146 91724
rect 230842 91712 230848 91724
rect 182140 91684 230848 91712
rect 182140 91672 182146 91684
rect 230842 91672 230848 91684
rect 230900 91672 230906 91724
rect 260466 91672 260472 91724
rect 260524 91712 260530 91724
rect 356054 91712 356060 91724
rect 260524 91684 356060 91712
rect 260524 91672 260530 91684
rect 356054 91672 356060 91684
rect 356112 91672 356118 91724
rect 254394 91604 254400 91656
rect 254452 91644 254458 91656
rect 317414 91644 317420 91656
rect 254452 91616 317420 91644
rect 254452 91604 254458 91616
rect 317414 91604 317420 91616
rect 317472 91604 317478 91656
rect 177850 90992 177856 91044
rect 177908 91032 177914 91044
rect 230198 91032 230204 91044
rect 177908 91004 230204 91032
rect 177908 90992 177914 91004
rect 230198 90992 230204 91004
rect 230256 90992 230262 91044
rect 260558 90992 260564 91044
rect 260616 91032 260622 91044
rect 353294 91032 353300 91044
rect 260616 91004 353300 91032
rect 260616 90992 260622 91004
rect 353294 90992 353300 91004
rect 353352 90992 353358 91044
rect 161290 90924 161296 90976
rect 161348 90964 161354 90976
rect 227162 90964 227168 90976
rect 161348 90936 227168 90964
rect 161348 90924 161354 90936
rect 227162 90924 227168 90936
rect 227220 90924 227226 90976
rect 271598 90924 271604 90976
rect 271656 90964 271662 90976
rect 406378 90964 406384 90976
rect 271656 90936 406384 90964
rect 271656 90924 271662 90936
rect 406378 90924 406384 90936
rect 406436 90924 406442 90976
rect 153010 90856 153016 90908
rect 153068 90896 153074 90908
rect 225966 90896 225972 90908
rect 153068 90868 225972 90896
rect 153068 90856 153074 90868
rect 225966 90856 225972 90868
rect 226024 90856 226030 90908
rect 278682 90856 278688 90908
rect 278740 90896 278746 90908
rect 457438 90896 457444 90908
rect 278740 90868 457444 90896
rect 278740 90856 278746 90868
rect 457438 90856 457444 90868
rect 457496 90856 457502 90908
rect 143442 90788 143448 90840
rect 143500 90828 143506 90840
rect 224126 90828 224132 90840
rect 143500 90800 224132 90828
rect 143500 90788 143506 90800
rect 224126 90788 224132 90800
rect 224184 90788 224190 90840
rect 282730 90788 282736 90840
rect 282788 90828 282794 90840
rect 471238 90828 471244 90840
rect 282788 90800 471244 90828
rect 282788 90788 282794 90800
rect 471238 90788 471244 90800
rect 471296 90788 471302 90840
rect 139302 90720 139308 90772
rect 139360 90760 139366 90772
rect 223758 90760 223764 90772
rect 139360 90732 223764 90760
rect 139360 90720 139366 90732
rect 223758 90720 223764 90732
rect 223816 90720 223822 90772
rect 282086 90720 282092 90772
rect 282144 90760 282150 90772
rect 481634 90760 481640 90772
rect 282144 90732 481640 90760
rect 282144 90720 282150 90732
rect 481634 90720 481640 90732
rect 481692 90720 481698 90772
rect 116578 90652 116584 90704
rect 116636 90692 116642 90704
rect 219618 90692 219624 90704
rect 116636 90664 219624 90692
rect 116636 90652 116642 90664
rect 219618 90652 219624 90664
rect 219676 90652 219682 90704
rect 283926 90652 283932 90704
rect 283984 90692 283990 90704
rect 490558 90692 490564 90704
rect 283984 90664 490564 90692
rect 283984 90652 283990 90664
rect 490558 90652 490564 90664
rect 490616 90652 490622 90704
rect 105538 90584 105544 90636
rect 105596 90624 105602 90636
rect 216030 90624 216036 90636
rect 105596 90596 216036 90624
rect 105596 90584 105602 90596
rect 216030 90584 216036 90596
rect 216088 90584 216094 90636
rect 285306 90584 285312 90636
rect 285364 90624 285370 90636
rect 493318 90624 493324 90636
rect 285364 90596 493324 90624
rect 285364 90584 285370 90596
rect 493318 90584 493324 90596
rect 493376 90584 493382 90636
rect 86770 90516 86776 90568
rect 86828 90556 86834 90568
rect 214650 90556 214656 90568
rect 86828 90528 214656 90556
rect 86828 90516 86834 90528
rect 214650 90516 214656 90528
rect 214708 90516 214714 90568
rect 286410 90516 286416 90568
rect 286468 90556 286474 90568
rect 500218 90556 500224 90568
rect 286468 90528 500224 90556
rect 286468 90516 286474 90528
rect 500218 90516 500224 90528
rect 500276 90516 500282 90568
rect 73062 90448 73068 90500
rect 73120 90488 73126 90500
rect 212258 90488 212264 90500
rect 73120 90460 212264 90488
rect 73120 90448 73126 90460
rect 212258 90448 212264 90460
rect 212316 90448 212322 90500
rect 287698 90448 287704 90500
rect 287756 90488 287762 90500
rect 511258 90488 511264 90500
rect 287756 90460 511264 90488
rect 287756 90448 287762 90460
rect 511258 90448 511264 90460
rect 511316 90448 511322 90500
rect 68278 90380 68284 90432
rect 68336 90420 68342 90432
rect 208210 90420 208216 90432
rect 68336 90392 208216 90420
rect 68336 90380 68342 90392
rect 208210 90380 208216 90392
rect 208268 90380 208274 90432
rect 290918 90380 290924 90432
rect 290976 90420 290982 90432
rect 529198 90420 529204 90432
rect 290976 90392 529204 90420
rect 290976 90380 290982 90392
rect 529198 90380 529204 90392
rect 529256 90380 529262 90432
rect 18598 90312 18604 90364
rect 18656 90352 18662 90364
rect 202230 90352 202236 90364
rect 18656 90324 202236 90352
rect 18656 90312 18662 90324
rect 202230 90312 202236 90324
rect 202288 90312 202294 90364
rect 248138 90312 248144 90364
rect 248196 90352 248202 90364
rect 282178 90352 282184 90364
rect 248196 90324 282184 90352
rect 248196 90312 248202 90324
rect 282178 90312 282184 90324
rect 282236 90312 282242 90364
rect 296070 90312 296076 90364
rect 296128 90352 296134 90364
rect 556798 90352 556804 90364
rect 296128 90324 556804 90352
rect 296128 90312 296134 90324
rect 556798 90312 556804 90324
rect 556856 90312 556862 90364
rect 254946 90244 254952 90296
rect 255004 90284 255010 90296
rect 321554 90284 321560 90296
rect 255004 90256 321560 90284
rect 255004 90244 255010 90256
rect 321554 90244 321560 90256
rect 321612 90244 321618 90296
rect 253566 90176 253572 90228
rect 253624 90216 253630 90228
rect 310514 90216 310520 90228
rect 253624 90188 310520 90216
rect 253624 90176 253630 90188
rect 310514 90176 310520 90188
rect 310572 90176 310578 90228
rect 252186 90108 252192 90160
rect 252244 90148 252250 90160
rect 303614 90148 303620 90160
rect 252244 90120 303620 90148
rect 252244 90108 252250 90120
rect 303614 90108 303620 90120
rect 303672 90108 303678 90160
rect 267274 89632 267280 89684
rect 267332 89672 267338 89684
rect 389818 89672 389824 89684
rect 267332 89644 389824 89672
rect 267332 89632 267338 89644
rect 389818 89632 389824 89644
rect 389876 89632 389882 89684
rect 268654 89564 268660 89616
rect 268712 89604 268718 89616
rect 398834 89604 398840 89616
rect 268712 89576 398840 89604
rect 268712 89564 268718 89576
rect 398834 89564 398840 89576
rect 398892 89564 398898 89616
rect 297818 89496 297824 89548
rect 297876 89536 297882 89548
rect 467098 89536 467104 89548
rect 297876 89508 467104 89536
rect 297876 89496 297882 89508
rect 467098 89496 467104 89508
rect 467156 89496 467162 89548
rect 157978 89428 157984 89480
rect 158036 89468 158042 89480
rect 226610 89468 226616 89480
rect 158036 89440 226616 89468
rect 158036 89428 158042 89440
rect 226610 89428 226616 89440
rect 226668 89428 226674 89480
rect 281442 89428 281448 89480
rect 281500 89468 281506 89480
rect 472710 89468 472716 89480
rect 281500 89440 472716 89468
rect 281500 89428 281506 89440
rect 472710 89428 472716 89440
rect 472768 89428 472774 89480
rect 122742 89360 122748 89412
rect 122800 89400 122806 89412
rect 221550 89400 221556 89412
rect 122800 89372 221556 89400
rect 122800 89360 122806 89372
rect 221550 89360 221556 89372
rect 221608 89360 221614 89412
rect 285398 89360 285404 89412
rect 285456 89400 285462 89412
rect 497458 89400 497464 89412
rect 285456 89372 497464 89400
rect 285456 89360 285462 89372
rect 497458 89360 497464 89372
rect 497516 89360 497522 89412
rect 119982 89292 119988 89344
rect 120040 89332 120046 89344
rect 220262 89332 220268 89344
rect 120040 89304 220268 89332
rect 120040 89292 120046 89304
rect 220262 89292 220268 89304
rect 220320 89292 220326 89344
rect 286870 89292 286876 89344
rect 286928 89332 286934 89344
rect 504358 89332 504364 89344
rect 286928 89304 504364 89332
rect 286928 89292 286934 89304
rect 504358 89292 504364 89304
rect 504416 89292 504422 89344
rect 108298 89224 108304 89276
rect 108356 89264 108362 89276
rect 214098 89264 214104 89276
rect 108356 89236 214104 89264
rect 108356 89224 108362 89236
rect 214098 89224 214104 89236
rect 214156 89224 214162 89276
rect 286686 89224 286692 89276
rect 286744 89264 286750 89276
rect 506474 89264 506480 89276
rect 286744 89236 506480 89264
rect 286744 89224 286750 89236
rect 506474 89224 506480 89236
rect 506532 89224 506538 89276
rect 53742 89156 53748 89208
rect 53800 89196 53806 89208
rect 199378 89196 199384 89208
rect 53800 89168 199384 89196
rect 53800 89156 53806 89168
rect 199378 89156 199384 89168
rect 199436 89156 199442 89208
rect 292114 89156 292120 89208
rect 292172 89196 292178 89208
rect 518158 89196 518164 89208
rect 292172 89168 518164 89196
rect 292172 89156 292178 89168
rect 518158 89156 518164 89168
rect 518216 89156 518222 89208
rect 47578 89088 47584 89140
rect 47636 89128 47642 89140
rect 205818 89128 205824 89140
rect 47636 89100 205824 89128
rect 47636 89088 47642 89100
rect 205818 89088 205824 89100
rect 205876 89088 205882 89140
rect 288066 89088 288072 89140
rect 288124 89128 288130 89140
rect 515398 89128 515404 89140
rect 288124 89100 515404 89128
rect 288124 89088 288130 89100
rect 515398 89088 515404 89100
rect 515456 89088 515462 89140
rect 43530 89020 43536 89072
rect 43588 89060 43594 89072
rect 207198 89060 207204 89072
rect 43588 89032 207204 89060
rect 43588 89020 43594 89032
rect 207198 89020 207204 89032
rect 207256 89020 207262 89072
rect 289354 89020 289360 89072
rect 289412 89060 289418 89072
rect 522298 89060 522304 89072
rect 289412 89032 522304 89060
rect 289412 89020 289418 89032
rect 522298 89020 522304 89032
rect 522356 89020 522362 89072
rect 40678 88952 40684 89004
rect 40736 88992 40742 89004
rect 205726 88992 205732 89004
rect 40736 88964 205732 88992
rect 40736 88952 40742 88964
rect 205726 88952 205732 88964
rect 205784 88952 205790 89004
rect 293586 88952 293592 89004
rect 293644 88992 293650 89004
rect 547966 88992 547972 89004
rect 293644 88964 547972 88992
rect 293644 88952 293650 88964
rect 547966 88952 547972 88964
rect 548024 88952 548030 89004
rect 257798 88884 257804 88936
rect 257856 88924 257862 88936
rect 331858 88924 331864 88936
rect 257856 88896 331864 88924
rect 257856 88884 257862 88896
rect 331858 88884 331864 88896
rect 331916 88884 331922 88936
rect 256326 88816 256332 88868
rect 256384 88856 256390 88868
rect 323578 88856 323584 88868
rect 256384 88828 323584 88856
rect 256384 88816 256390 88828
rect 323578 88816 323584 88828
rect 323636 88816 323642 88868
rect 256418 88272 256424 88324
rect 256476 88312 256482 88324
rect 328454 88312 328460 88324
rect 256476 88284 328460 88312
rect 256476 88272 256482 88284
rect 328454 88272 328460 88284
rect 328512 88272 328518 88324
rect 257890 88204 257896 88256
rect 257948 88244 257954 88256
rect 335354 88244 335360 88256
rect 257948 88216 335360 88244
rect 257948 88204 257954 88216
rect 335354 88204 335360 88216
rect 335412 88204 335418 88256
rect 261846 88136 261852 88188
rect 261904 88176 261910 88188
rect 357434 88176 357440 88188
rect 261904 88148 357440 88176
rect 261904 88136 261910 88148
rect 357434 88136 357440 88148
rect 357492 88136 357498 88188
rect 263410 88068 263416 88120
rect 263468 88108 263474 88120
rect 367738 88108 367744 88120
rect 263468 88080 367744 88108
rect 263468 88068 263474 88080
rect 367738 88068 367744 88080
rect 367796 88068 367802 88120
rect 124122 88000 124128 88052
rect 124180 88040 124186 88052
rect 221182 88040 221188 88052
rect 124180 88012 221188 88040
rect 124180 88000 124186 88012
rect 221182 88000 221188 88012
rect 221240 88000 221246 88052
rect 270034 88000 270040 88052
rect 270092 88040 270098 88052
rect 409874 88040 409880 88052
rect 270092 88012 409880 88040
rect 270092 88000 270098 88012
rect 409874 88000 409880 88012
rect 409932 88000 409938 88052
rect 117222 87932 117228 87984
rect 117280 87972 117286 87984
rect 219802 87972 219808 87984
rect 117280 87944 219808 87972
rect 117280 87932 117286 87944
rect 219802 87932 219808 87944
rect 219860 87932 219866 87984
rect 272886 87932 272892 87984
rect 272944 87972 272950 87984
rect 420914 87972 420920 87984
rect 272944 87944 420920 87972
rect 272944 87932 272950 87944
rect 420914 87932 420920 87944
rect 420972 87932 420978 87984
rect 75178 87864 75184 87916
rect 75236 87904 75242 87916
rect 211246 87904 211252 87916
rect 75236 87876 211252 87904
rect 75236 87864 75242 87876
rect 211246 87864 211252 87876
rect 211304 87864 211310 87916
rect 294966 87864 294972 87916
rect 295024 87904 295030 87916
rect 536098 87904 536104 87916
rect 295024 87876 536104 87904
rect 295024 87864 295030 87876
rect 536098 87864 536104 87876
rect 536156 87864 536162 87916
rect 57238 87796 57244 87848
rect 57296 87836 57302 87848
rect 209406 87836 209412 87848
rect 57296 87808 209412 87836
rect 57296 87796 57302 87808
rect 209406 87796 209412 87808
rect 209464 87796 209470 87848
rect 292298 87796 292304 87848
rect 292356 87836 292362 87848
rect 538214 87836 538220 87848
rect 292356 87808 538220 87836
rect 292356 87796 292362 87808
rect 538214 87796 538220 87808
rect 538272 87796 538278 87848
rect 53098 87728 53104 87780
rect 53156 87768 53162 87780
rect 206830 87768 206836 87780
rect 53156 87740 206836 87768
rect 53156 87728 53162 87740
rect 206830 87728 206836 87740
rect 206888 87728 206894 87780
rect 292206 87728 292212 87780
rect 292264 87768 292270 87780
rect 540238 87768 540244 87780
rect 292264 87740 540244 87768
rect 292264 87728 292270 87740
rect 540238 87728 540244 87740
rect 540296 87728 540302 87780
rect 46842 87660 46848 87712
rect 46900 87700 46906 87712
rect 203518 87700 203524 87712
rect 46900 87672 203524 87700
rect 46900 87660 46906 87672
rect 203518 87660 203524 87672
rect 203576 87660 203582 87712
rect 295058 87660 295064 87712
rect 295116 87700 295122 87712
rect 547138 87700 547144 87712
rect 295116 87672 547144 87700
rect 295116 87660 295122 87672
rect 547138 87660 547144 87672
rect 547196 87660 547202 87712
rect 14458 87592 14464 87644
rect 14516 87632 14522 87644
rect 201678 87632 201684 87644
rect 14516 87604 201684 87632
rect 14516 87592 14522 87604
rect 201678 87592 201684 87604
rect 201736 87592 201742 87644
rect 296346 87592 296352 87644
rect 296404 87632 296410 87644
rect 560938 87632 560944 87644
rect 296404 87604 560944 87632
rect 296404 87592 296410 87604
rect 560938 87592 560944 87604
rect 560996 87592 561002 87644
rect 253658 87524 253664 87576
rect 253716 87564 253722 87576
rect 313918 87564 313924 87576
rect 253716 87536 313924 87564
rect 253716 87524 253722 87536
rect 313918 87524 313924 87536
rect 313976 87524 313982 87576
rect 307018 86912 307024 86964
rect 307076 86952 307082 86964
rect 580166 86952 580172 86964
rect 307076 86924 580172 86952
rect 307076 86912 307082 86924
rect 580166 86912 580172 86924
rect 580224 86912 580230 86964
rect 257614 86844 257620 86896
rect 257672 86884 257678 86896
rect 339494 86884 339500 86896
rect 257672 86856 339500 86884
rect 257672 86844 257678 86856
rect 339494 86844 339500 86856
rect 339552 86844 339558 86896
rect 261938 86776 261944 86828
rect 261996 86816 262002 86828
rect 360194 86816 360200 86828
rect 261996 86788 360200 86816
rect 261996 86776 262002 86788
rect 360194 86776 360200 86788
rect 360252 86776 360258 86828
rect 261662 86708 261668 86760
rect 261720 86748 261726 86760
rect 363598 86748 363604 86760
rect 261720 86720 363604 86748
rect 261720 86708 261726 86720
rect 363598 86708 363604 86720
rect 363656 86708 363662 86760
rect 264698 86640 264704 86692
rect 264756 86680 264762 86692
rect 374086 86680 374092 86692
rect 264756 86652 374092 86680
rect 264756 86640 264762 86652
rect 374086 86640 374092 86652
rect 374144 86640 374150 86692
rect 268746 86572 268752 86624
rect 268804 86612 268810 86624
rect 402974 86612 402980 86624
rect 268804 86584 402980 86612
rect 268804 86572 268810 86584
rect 402974 86572 402980 86584
rect 403032 86572 403038 86624
rect 107562 86504 107568 86556
rect 107620 86544 107626 86556
rect 191190 86544 191196 86556
rect 107620 86516 191196 86544
rect 107620 86504 107626 86516
rect 191190 86504 191196 86516
rect 191248 86504 191254 86556
rect 271690 86504 271696 86556
rect 271748 86544 271754 86556
rect 416774 86544 416780 86556
rect 271748 86516 416780 86544
rect 271748 86504 271754 86516
rect 416774 86504 416780 86516
rect 416832 86504 416838 86556
rect 90358 86436 90364 86488
rect 90416 86476 90422 86488
rect 215110 86476 215116 86488
rect 90416 86448 215116 86476
rect 90416 86436 90422 86448
rect 215110 86436 215116 86448
rect 215168 86436 215174 86488
rect 277026 86436 277032 86488
rect 277084 86476 277090 86488
rect 425698 86476 425704 86488
rect 277084 86448 425704 86476
rect 277084 86436 277090 86448
rect 425698 86436 425704 86448
rect 425756 86436 425762 86488
rect 79318 86368 79324 86420
rect 79376 86408 79382 86420
rect 208854 86408 208860 86420
rect 79376 86380 208860 86408
rect 79376 86368 79382 86380
rect 208854 86368 208860 86380
rect 208912 86368 208918 86420
rect 278406 86368 278412 86420
rect 278464 86408 278470 86420
rect 453390 86408 453396 86420
rect 278464 86380 453396 86408
rect 278464 86368 278470 86380
rect 453390 86368 453396 86380
rect 453448 86368 453454 86420
rect 76558 86300 76564 86352
rect 76616 86340 76622 86352
rect 211614 86340 211620 86352
rect 76616 86312 211620 86340
rect 76616 86300 76622 86312
rect 211614 86300 211620 86312
rect 211672 86300 211678 86352
rect 297634 86300 297640 86352
rect 297692 86340 297698 86352
rect 566458 86340 566464 86352
rect 297692 86312 566464 86340
rect 297692 86300 297698 86312
rect 566458 86300 566464 86312
rect 566516 86300 566522 86352
rect 35158 86232 35164 86284
rect 35216 86272 35222 86284
rect 201862 86272 201868 86284
rect 35216 86244 201868 86272
rect 35216 86232 35222 86244
rect 201862 86232 201868 86244
rect 201920 86232 201926 86284
rect 248230 86232 248236 86284
rect 248288 86272 248294 86284
rect 261478 86272 261484 86284
rect 248288 86244 261484 86272
rect 248288 86232 248294 86244
rect 261478 86232 261484 86244
rect 261536 86232 261542 86284
rect 296438 86232 296444 86284
rect 296496 86272 296502 86284
rect 565814 86272 565820 86284
rect 296496 86244 565820 86272
rect 296496 86232 296502 86244
rect 565814 86232 565820 86244
rect 565872 86232 565878 86284
rect 255038 86164 255044 86216
rect 255096 86204 255102 86216
rect 316126 86204 316132 86216
rect 255096 86176 316132 86204
rect 255096 86164 255102 86176
rect 316126 86164 316132 86176
rect 316184 86164 316190 86216
rect 3142 85484 3148 85536
rect 3200 85524 3206 85536
rect 151078 85524 151084 85536
rect 3200 85496 151084 85524
rect 3200 85484 3206 85496
rect 151078 85484 151084 85496
rect 151136 85484 151142 85536
rect 253750 85416 253756 85468
rect 253808 85456 253814 85468
rect 307018 85456 307024 85468
rect 253808 85428 307024 85456
rect 253808 85416 253814 85428
rect 307018 85416 307024 85428
rect 307076 85416 307082 85468
rect 263134 85348 263140 85400
rect 263192 85388 263198 85400
rect 332686 85388 332692 85400
rect 263192 85360 332692 85388
rect 263192 85348 263198 85360
rect 332686 85348 332692 85360
rect 332744 85348 332750 85400
rect 266998 85280 267004 85332
rect 267056 85320 267062 85332
rect 375374 85320 375380 85332
rect 267056 85292 375380 85320
rect 267056 85280 267062 85292
rect 375374 85280 375380 85292
rect 375432 85280 375438 85332
rect 264790 85212 264796 85264
rect 264848 85252 264854 85264
rect 378134 85252 378140 85264
rect 264848 85224 378140 85252
rect 264848 85212 264854 85224
rect 378134 85212 378140 85224
rect 378192 85212 378198 85264
rect 272978 85144 272984 85196
rect 273036 85184 273042 85196
rect 423766 85184 423772 85196
rect 273036 85156 423772 85184
rect 273036 85144 273042 85156
rect 423766 85144 423772 85156
rect 423824 85144 423830 85196
rect 278498 85076 278504 85128
rect 278556 85116 278562 85128
rect 459554 85116 459560 85128
rect 278556 85088 459560 85116
rect 278556 85076 278562 85088
rect 459554 85076 459560 85088
rect 459612 85076 459618 85128
rect 282270 85008 282276 85060
rect 282328 85048 282334 85060
rect 463694 85048 463700 85060
rect 282328 85020 463700 85048
rect 282328 85008 282334 85020
rect 463694 85008 463700 85020
rect 463752 85008 463758 85060
rect 284110 84940 284116 84992
rect 284168 84980 284174 84992
rect 485774 84980 485780 84992
rect 284168 84952 485780 84980
rect 284168 84940 284174 84952
rect 485774 84940 485780 84952
rect 485832 84940 485838 84992
rect 284018 84872 284024 84924
rect 284076 84912 284082 84924
rect 490006 84912 490012 84924
rect 284076 84884 490012 84912
rect 284076 84872 284082 84884
rect 490006 84872 490012 84884
rect 490064 84872 490070 84924
rect 5442 84804 5448 84856
rect 5500 84844 5506 84856
rect 197998 84844 198004 84856
rect 5500 84816 198004 84844
rect 5500 84804 5506 84816
rect 197998 84804 198004 84816
rect 198056 84804 198062 84856
rect 290734 84804 290740 84856
rect 290792 84844 290798 84856
rect 530578 84844 530584 84856
rect 290792 84816 530584 84844
rect 290792 84804 290798 84816
rect 530578 84804 530584 84816
rect 530636 84804 530642 84856
rect 255130 83988 255136 84040
rect 255188 84028 255194 84040
rect 318058 84028 318064 84040
rect 255188 84000 318064 84028
rect 255188 83988 255194 84000
rect 318058 83988 318064 84000
rect 318116 83988 318122 84040
rect 256142 83920 256148 83972
rect 256200 83960 256206 83972
rect 324958 83960 324964 83972
rect 256200 83932 324964 83960
rect 256200 83920 256206 83932
rect 324958 83920 324964 83932
rect 325016 83920 325022 83972
rect 261754 83852 261760 83904
rect 261812 83892 261818 83904
rect 360838 83892 360844 83904
rect 261812 83864 360844 83892
rect 261812 83852 261818 83864
rect 360838 83852 360844 83864
rect 360896 83852 360902 83904
rect 268838 83784 268844 83836
rect 268896 83824 268902 83836
rect 395338 83824 395344 83836
rect 268896 83796 395344 83824
rect 268896 83784 268902 83796
rect 395338 83784 395344 83796
rect 395396 83784 395402 83836
rect 282730 83716 282736 83768
rect 282788 83756 282794 83768
rect 477494 83756 477500 83768
rect 282788 83728 477500 83756
rect 282788 83716 282794 83728
rect 477494 83716 477500 83728
rect 477552 83716 477558 83768
rect 283834 83648 283840 83700
rect 283892 83688 283898 83700
rect 492674 83688 492680 83700
rect 283892 83660 492680 83688
rect 283892 83648 283898 83660
rect 492674 83648 492680 83660
rect 492732 83648 492738 83700
rect 285122 83580 285128 83632
rect 285180 83620 285186 83632
rect 496814 83620 496820 83632
rect 285180 83592 496820 83620
rect 285180 83580 285186 83592
rect 496814 83580 496820 83592
rect 496872 83580 496878 83632
rect 290826 83512 290832 83564
rect 290884 83552 290890 83564
rect 528554 83552 528560 83564
rect 290884 83524 528560 83552
rect 290884 83512 290890 83524
rect 528554 83512 528560 83524
rect 528612 83512 528618 83564
rect 293678 83444 293684 83496
rect 293736 83484 293742 83496
rect 542354 83484 542360 83496
rect 293736 83456 542360 83484
rect 293736 83444 293742 83456
rect 542354 83444 542360 83456
rect 542412 83444 542418 83496
rect 271322 82492 271328 82544
rect 271380 82532 271386 82544
rect 365806 82532 365812 82544
rect 271380 82504 365812 82532
rect 271380 82492 271386 82504
rect 365806 82492 365812 82504
rect 365864 82492 365870 82544
rect 271230 82424 271236 82476
rect 271288 82464 271294 82476
rect 382274 82464 382280 82476
rect 271288 82436 382280 82464
rect 271288 82424 271294 82436
rect 382274 82424 382280 82436
rect 382332 82424 382338 82476
rect 270126 82356 270132 82408
rect 270184 82396 270190 82408
rect 392578 82396 392584 82408
rect 270184 82368 392584 82396
rect 270184 82356 270190 82368
rect 392578 82356 392584 82368
rect 392636 82356 392642 82408
rect 276658 82288 276664 82340
rect 276716 82328 276722 82340
rect 400214 82328 400220 82340
rect 276716 82300 400220 82328
rect 276716 82288 276722 82300
rect 400214 82288 400220 82300
rect 400272 82288 400278 82340
rect 288158 82220 288164 82272
rect 288216 82260 288222 82272
rect 510614 82260 510620 82272
rect 288216 82232 510620 82260
rect 288216 82220 288222 82232
rect 510614 82220 510620 82232
rect 510672 82220 510678 82272
rect 293218 82152 293224 82204
rect 293276 82192 293282 82204
rect 546494 82192 546500 82204
rect 293276 82164 546500 82192
rect 293276 82152 293282 82164
rect 546494 82152 546500 82164
rect 546552 82152 546558 82204
rect 294782 82084 294788 82136
rect 294840 82124 294846 82136
rect 553394 82124 553400 82136
rect 294840 82096 553400 82124
rect 294840 82084 294846 82096
rect 553394 82084 553400 82096
rect 553452 82084 553458 82136
rect 301498 80928 301504 80980
rect 301556 80968 301562 80980
rect 404354 80968 404360 80980
rect 301556 80940 404360 80968
rect 301556 80928 301562 80940
rect 404354 80928 404360 80940
rect 404412 80928 404418 80980
rect 274266 80860 274272 80912
rect 274324 80900 274330 80912
rect 429194 80900 429200 80912
rect 274324 80872 429200 80900
rect 274324 80860 274330 80872
rect 429194 80860 429200 80872
rect 429252 80860 429258 80912
rect 274358 80792 274364 80844
rect 274416 80832 274422 80844
rect 431218 80832 431224 80844
rect 274416 80804 431224 80832
rect 274416 80792 274422 80804
rect 431218 80792 431224 80804
rect 431276 80792 431282 80844
rect 275738 80724 275744 80776
rect 275796 80764 275802 80776
rect 440326 80764 440332 80776
rect 275796 80736 440332 80764
rect 275796 80724 275802 80736
rect 440326 80724 440332 80736
rect 440384 80724 440390 80776
rect 297726 80656 297732 80708
rect 297784 80696 297790 80708
rect 571334 80696 571340 80708
rect 297784 80668 571340 80696
rect 297784 80656 297790 80668
rect 571334 80656 571340 80668
rect 571392 80656 571398 80708
rect 302878 79296 302884 79348
rect 302936 79336 302942 79348
rect 447134 79336 447140 79348
rect 302936 79308 447140 79336
rect 302936 79296 302942 79308
rect 447134 79296 447140 79308
rect 447192 79296 447198 79348
rect 309778 73108 309784 73160
rect 309836 73148 309842 73160
rect 579982 73148 579988 73160
rect 309836 73120 579988 73148
rect 309836 73108 309842 73120
rect 579982 73108 579988 73120
rect 580040 73108 580046 73160
rect 2774 71612 2780 71664
rect 2832 71652 2838 71664
rect 4798 71652 4804 71664
rect 2832 71624 4804 71652
rect 2832 71612 2838 71624
rect 4798 71612 4804 71624
rect 4856 71612 4862 71664
rect 454678 60664 454684 60716
rect 454736 60704 454742 60716
rect 580166 60704 580172 60716
rect 454736 60676 580172 60704
rect 454736 60664 454742 60676
rect 580166 60664 580172 60676
rect 580224 60664 580230 60716
rect 3050 59304 3056 59356
rect 3108 59344 3114 59356
rect 146938 59344 146944 59356
rect 3108 59316 146944 59344
rect 3108 59304 3114 59316
rect 146938 59304 146944 59316
rect 146996 59304 147002 59356
rect 3418 45500 3424 45552
rect 3476 45540 3482 45552
rect 148318 45540 148324 45552
rect 3476 45512 148324 45540
rect 3476 45500 3482 45512
rect 148318 45500 148324 45512
rect 148376 45500 148382 45552
rect 322198 37884 322204 37936
rect 322256 37924 322262 37936
rect 478874 37924 478880 37936
rect 322256 37896 478880 37924
rect 322256 37884 322262 37896
rect 478874 37884 478880 37896
rect 478932 37884 478938 37936
rect 312538 35164 312544 35216
rect 312596 35204 312602 35216
rect 425054 35204 425060 35216
rect 312596 35176 425060 35204
rect 312596 35164 312602 35176
rect 425054 35164 425060 35176
rect 425112 35164 425118 35216
rect 254854 33736 254860 33788
rect 254912 33776 254918 33788
rect 322934 33776 322940 33788
rect 254912 33748 322940 33776
rect 254912 33736 254918 33748
rect 322934 33736 322940 33748
rect 322992 33736 322998 33788
rect 323670 33736 323676 33788
rect 323728 33776 323734 33788
rect 456886 33776 456892 33788
rect 323728 33748 456892 33776
rect 323728 33736 323734 33748
rect 456886 33736 456892 33748
rect 456944 33736 456950 33788
rect 3142 33056 3148 33108
rect 3200 33096 3206 33108
rect 155218 33096 155224 33108
rect 3200 33068 155224 33096
rect 3200 33056 3206 33068
rect 155218 33056 155224 33068
rect 155276 33056 155282 33108
rect 305638 33056 305644 33108
rect 305696 33096 305702 33108
rect 580166 33096 580172 33108
rect 305696 33068 580172 33096
rect 305696 33056 305702 33068
rect 580166 33056 580172 33068
rect 580224 33056 580230 33108
rect 256234 31016 256240 31068
rect 256292 31056 256298 31068
rect 329834 31056 329840 31068
rect 256292 31028 329840 31056
rect 256292 31016 256298 31028
rect 329834 31016 329840 31028
rect 329892 31016 329898 31068
rect 253474 29588 253480 29640
rect 253532 29628 253538 29640
rect 311894 29628 311900 29640
rect 253532 29600 311900 29628
rect 253532 29588 253538 29600
rect 311894 29588 311900 29600
rect 311952 29588 311958 29640
rect 294874 28228 294880 28280
rect 294932 28268 294938 28280
rect 556246 28268 556252 28280
rect 294932 28240 556252 28268
rect 294932 28228 294938 28240
rect 556246 28228 556252 28240
rect 556304 28228 556310 28280
rect 33042 26868 33048 26920
rect 33100 26908 33106 26920
rect 202138 26908 202144 26920
rect 33100 26880 202144 26908
rect 33100 26868 33106 26880
rect 202138 26868 202144 26880
rect 202196 26868 202202 26920
rect 292022 26868 292028 26920
rect 292080 26908 292086 26920
rect 539686 26908 539692 26920
rect 292080 26880 539692 26908
rect 292080 26868 292086 26880
rect 539686 26868 539692 26880
rect 539744 26868 539750 26920
rect 296162 25508 296168 25560
rect 296220 25548 296226 25560
rect 564526 25548 564532 25560
rect 296220 25520 564532 25548
rect 296220 25508 296226 25520
rect 564526 25508 564532 25520
rect 564584 25508 564590 25560
rect 199930 24080 199936 24132
rect 199988 24120 199994 24132
rect 233602 24120 233608 24132
rect 199988 24092 233608 24120
rect 199988 24080 199994 24092
rect 233602 24080 233608 24092
rect 233660 24080 233666 24132
rect 282454 24080 282460 24132
rect 282512 24120 282518 24132
rect 481726 24120 481732 24132
rect 282512 24092 481732 24120
rect 282512 24080 282518 24092
rect 481726 24080 481732 24092
rect 481784 24080 481790 24132
rect 234062 23468 234068 23520
rect 234120 23508 234126 23520
rect 238294 23508 238300 23520
rect 234120 23480 238300 23508
rect 234120 23468 234126 23480
rect 238294 23468 238300 23480
rect 238352 23468 238358 23520
rect 233142 22720 233148 22772
rect 233200 22760 233206 22772
rect 239490 22760 239496 22772
rect 233200 22732 239496 22760
rect 233200 22720 233206 22732
rect 239490 22720 239496 22732
rect 239548 22720 239554 22772
rect 246666 22720 246672 22772
rect 246724 22760 246730 22772
rect 267734 22760 267740 22772
rect 246724 22732 267740 22760
rect 246724 22720 246730 22732
rect 267734 22720 267740 22732
rect 267792 22720 267798 22772
rect 293494 22720 293500 22772
rect 293552 22760 293558 22772
rect 548518 22760 548524 22772
rect 293552 22732 548524 22760
rect 293552 22720 293558 22732
rect 548518 22720 548524 22732
rect 548576 22720 548582 22772
rect 286502 21360 286508 21412
rect 286560 21400 286566 21412
rect 506566 21400 506572 21412
rect 286560 21372 506572 21400
rect 286560 21360 286566 21372
rect 506566 21360 506572 21372
rect 506624 21360 506630 21412
rect 3418 20612 3424 20664
rect 3476 20652 3482 20664
rect 144178 20652 144184 20664
rect 3476 20624 144184 20652
rect 3476 20612 3482 20624
rect 144178 20612 144184 20624
rect 144236 20612 144242 20664
rect 453298 20612 453304 20664
rect 453356 20652 453362 20664
rect 580166 20652 580172 20664
rect 453356 20624 580172 20652
rect 453356 20612 453362 20624
rect 580166 20612 580172 20624
rect 580224 20612 580230 20664
rect 252278 19932 252284 19984
rect 252336 19972 252342 19984
rect 300854 19972 300860 19984
rect 252336 19944 300860 19972
rect 252336 19932 252342 19944
rect 300854 19932 300860 19944
rect 300912 19932 300918 19984
rect 287882 18572 287888 18624
rect 287940 18612 287946 18624
rect 517514 18612 517520 18624
rect 287940 18584 517520 18612
rect 287940 18572 287946 18584
rect 517514 18572 517520 18584
rect 517572 18572 517578 18624
rect 262950 17212 262956 17264
rect 263008 17252 263014 17264
rect 284294 17252 284300 17264
rect 263008 17224 284300 17252
rect 263008 17212 263014 17224
rect 284294 17212 284300 17224
rect 284352 17212 284358 17264
rect 285214 17212 285220 17264
rect 285272 17252 285278 17264
rect 499574 17252 499580 17264
rect 285272 17224 499580 17252
rect 285272 17212 285278 17224
rect 499574 17212 499580 17224
rect 499632 17212 499638 17264
rect 258994 15988 259000 16040
rect 259052 16028 259058 16040
rect 340966 16028 340972 16040
rect 259052 16000 340972 16028
rect 259052 15988 259058 16000
rect 340966 15988 340972 16000
rect 341024 15988 341030 16040
rect 299106 15920 299112 15972
rect 299164 15960 299170 15972
rect 575106 15960 575112 15972
rect 299164 15932 575112 15960
rect 299164 15920 299170 15932
rect 575106 15920 575112 15932
rect 575164 15920 575170 15972
rect 245286 15852 245292 15904
rect 245344 15892 245350 15904
rect 253382 15892 253388 15904
rect 245344 15864 253388 15892
rect 245344 15852 245350 15864
rect 253382 15852 253388 15864
rect 253440 15852 253446 15904
rect 299014 15852 299020 15904
rect 299072 15892 299078 15904
rect 578602 15892 578608 15904
rect 299072 15864 578608 15892
rect 299072 15852 299078 15864
rect 578602 15852 578608 15864
rect 578660 15852 578666 15904
rect 289538 14492 289544 14544
rect 289596 14532 289602 14544
rect 521838 14532 521844 14544
rect 289596 14504 521844 14532
rect 289596 14492 289602 14504
rect 521838 14492 521844 14504
rect 521896 14492 521902 14544
rect 64782 14424 64788 14476
rect 64840 14464 64846 14476
rect 196618 14464 196624 14476
rect 64840 14436 196624 14464
rect 64840 14424 64846 14436
rect 196618 14424 196624 14436
rect 196676 14424 196682 14476
rect 289446 14424 289452 14476
rect 289504 14464 289510 14476
rect 525058 14464 525064 14476
rect 289504 14436 525064 14464
rect 289504 14424 289510 14436
rect 525058 14424 525064 14436
rect 525116 14424 525122 14476
rect 273070 13676 273076 13728
rect 273128 13716 273134 13728
rect 428366 13716 428372 13728
rect 273128 13688 428372 13716
rect 273128 13676 273134 13688
rect 428366 13676 428372 13688
rect 428424 13676 428430 13728
rect 274174 13608 274180 13660
rect 274232 13648 274238 13660
rect 432046 13648 432052 13660
rect 274232 13620 432052 13648
rect 274232 13608 274238 13620
rect 432046 13608 432052 13620
rect 432104 13608 432110 13660
rect 274450 13540 274456 13592
rect 274508 13580 274514 13592
rect 435082 13580 435088 13592
rect 274508 13552 435088 13580
rect 274508 13540 274514 13552
rect 435082 13540 435088 13552
rect 435140 13540 435146 13592
rect 275922 13472 275928 13524
rect 275980 13512 275986 13524
rect 439130 13512 439136 13524
rect 275980 13484 439136 13512
rect 275980 13472 275986 13484
rect 439130 13472 439136 13484
rect 439188 13472 439194 13524
rect 275830 13404 275836 13456
rect 275888 13444 275894 13456
rect 442626 13444 442632 13456
rect 275888 13416 442632 13444
rect 275888 13404 275894 13416
rect 442626 13404 442632 13416
rect 442684 13404 442690 13456
rect 277118 13336 277124 13388
rect 277176 13376 277182 13388
rect 445754 13376 445760 13388
rect 277176 13348 445760 13376
rect 277176 13336 277182 13348
rect 445754 13336 445760 13348
rect 445812 13336 445818 13388
rect 277210 13268 277216 13320
rect 277268 13308 277274 13320
rect 449802 13308 449808 13320
rect 277268 13280 449808 13308
rect 277268 13268 277274 13280
rect 449802 13268 449808 13280
rect 449860 13268 449866 13320
rect 276934 13200 276940 13252
rect 276992 13240 276998 13252
rect 453298 13240 453304 13252
rect 276992 13212 453304 13240
rect 276992 13200 276998 13212
rect 453298 13200 453304 13212
rect 453356 13200 453362 13252
rect 279970 13132 279976 13184
rect 280028 13172 280034 13184
rect 467098 13172 467104 13184
rect 280028 13144 467104 13172
rect 280028 13132 280034 13144
rect 467098 13132 467104 13144
rect 467156 13132 467162 13184
rect 119890 13064 119896 13116
rect 119948 13104 119954 13116
rect 219710 13104 219716 13116
rect 119948 13076 219716 13104
rect 119948 13064 119954 13076
rect 219710 13064 219716 13076
rect 219768 13064 219774 13116
rect 253290 13064 253296 13116
rect 253348 13104 253354 13116
rect 259454 13104 259460 13116
rect 253348 13076 259460 13104
rect 253348 13064 253354 13076
rect 259454 13064 259460 13076
rect 259512 13064 259518 13116
rect 281074 13064 281080 13116
rect 281132 13104 281138 13116
rect 470594 13104 470600 13116
rect 281132 13076 470600 13104
rect 281132 13064 281138 13076
rect 470594 13064 470600 13076
rect 470652 13064 470658 13116
rect 112806 12180 112812 12232
rect 112864 12220 112870 12232
rect 218882 12220 218888 12232
rect 112864 12192 218888 12220
rect 112864 12180 112870 12192
rect 218882 12180 218888 12192
rect 218940 12180 218946 12232
rect 110322 12112 110328 12164
rect 110380 12152 110386 12164
rect 218606 12152 218612 12164
rect 110380 12124 218612 12152
rect 110380 12112 110386 12124
rect 218606 12112 218612 12124
rect 218664 12112 218670 12164
rect 259086 12112 259092 12164
rect 259144 12152 259150 12164
rect 342898 12152 342904 12164
rect 259144 12124 342904 12152
rect 259144 12112 259150 12124
rect 342898 12112 342904 12124
rect 342956 12112 342962 12164
rect 106182 12044 106188 12096
rect 106240 12084 106246 12096
rect 218330 12084 218336 12096
rect 106240 12056 218336 12084
rect 106240 12044 106246 12056
rect 218330 12044 218336 12056
rect 218388 12044 218394 12096
rect 259178 12044 259184 12096
rect 259236 12084 259242 12096
rect 346946 12084 346952 12096
rect 259236 12056 346952 12084
rect 259236 12044 259242 12056
rect 346946 12044 346952 12056
rect 347004 12044 347010 12096
rect 103422 11976 103428 12028
rect 103480 12016 103486 12028
rect 216950 12016 216956 12028
rect 103480 11988 216956 12016
rect 103480 11976 103486 11988
rect 216950 11976 216956 11988
rect 217008 11976 217014 12028
rect 263502 11976 263508 12028
rect 263560 12016 263566 12028
rect 367738 12016 367744 12028
rect 263560 11988 367744 12016
rect 263560 11976 263566 11988
rect 367738 11976 367744 11988
rect 367796 11976 367802 12028
rect 99282 11908 99288 11960
rect 99340 11948 99346 11960
rect 216858 11948 216864 11960
rect 99340 11920 216864 11948
rect 99340 11908 99346 11920
rect 216858 11908 216864 11920
rect 216916 11908 216922 11960
rect 266170 11908 266176 11960
rect 266228 11948 266234 11960
rect 382366 11948 382372 11960
rect 266228 11920 382372 11948
rect 266228 11908 266234 11920
rect 382366 11908 382372 11920
rect 382424 11908 382430 11960
rect 31294 11840 31300 11892
rect 31352 11880 31358 11892
rect 204438 11880 204444 11892
rect 31352 11852 204444 11880
rect 31352 11840 31358 11852
rect 204438 11840 204444 11852
rect 204496 11840 204502 11892
rect 266078 11840 266084 11892
rect 266136 11880 266142 11892
rect 385586 11880 385592 11892
rect 266136 11852 385592 11880
rect 266136 11840 266142 11852
rect 385586 11840 385592 11852
rect 385644 11840 385650 11892
rect 28902 11772 28908 11824
rect 28960 11812 28966 11824
rect 204714 11812 204720 11824
rect 28960 11784 204720 11812
rect 28960 11772 28966 11784
rect 204714 11772 204720 11784
rect 204772 11772 204778 11824
rect 267458 11772 267464 11824
rect 267516 11812 267522 11824
rect 389450 11812 389456 11824
rect 267516 11784 389456 11812
rect 267516 11772 267522 11784
rect 389450 11772 389456 11784
rect 389508 11772 389514 11824
rect 23014 11704 23020 11756
rect 23072 11744 23078 11756
rect 203150 11744 203156 11756
rect 23072 11716 203156 11744
rect 23072 11704 23078 11716
rect 203150 11704 203156 11716
rect 203208 11704 203214 11756
rect 267366 11704 267372 11756
rect 267424 11744 267430 11756
rect 392578 11744 392584 11756
rect 267424 11716 392584 11744
rect 267424 11704 267430 11716
rect 392578 11704 392584 11716
rect 392636 11704 392642 11756
rect 423766 11704 423772 11756
rect 423824 11744 423830 11756
rect 424962 11744 424968 11756
rect 423824 11716 424968 11744
rect 423824 11704 423830 11716
rect 424962 11704 424968 11716
rect 425020 11704 425026 11756
rect 332686 11636 332692 11688
rect 332744 11676 332750 11688
rect 333882 11676 333888 11688
rect 332744 11648 333888 11676
rect 332744 11636 332750 11648
rect 333882 11636 333888 11648
rect 333940 11636 333946 11688
rect 374086 11636 374092 11688
rect 374144 11676 374150 11688
rect 375282 11676 375288 11688
rect 374144 11648 375288 11676
rect 374144 11636 374150 11648
rect 375282 11636 375288 11648
rect 375340 11636 375346 11688
rect 95142 10684 95148 10736
rect 95200 10724 95206 10736
rect 216214 10724 216220 10736
rect 95200 10696 216220 10724
rect 95200 10684 95206 10696
rect 216214 10684 216220 10696
rect 216272 10684 216278 10736
rect 92382 10616 92388 10668
rect 92440 10656 92446 10668
rect 215478 10656 215484 10668
rect 92440 10628 215484 10656
rect 92440 10616 92446 10628
rect 215478 10616 215484 10628
rect 215536 10616 215542 10668
rect 87966 10548 87972 10600
rect 88024 10588 88030 10600
rect 214282 10588 214288 10600
rect 88024 10560 214288 10588
rect 88024 10548 88030 10560
rect 214282 10548 214288 10560
rect 214340 10548 214346 10600
rect 81342 10480 81348 10532
rect 81400 10520 81406 10532
rect 212718 10520 212724 10532
rect 81400 10492 212724 10520
rect 81400 10480 81406 10492
rect 212718 10480 212724 10492
rect 212776 10480 212782 10532
rect 78582 10412 78588 10464
rect 78640 10452 78646 10464
rect 212902 10452 212908 10464
rect 78640 10424 212908 10452
rect 78640 10412 78646 10424
rect 212902 10412 212908 10424
rect 212960 10412 212966 10464
rect 74442 10344 74448 10396
rect 74500 10384 74506 10396
rect 213270 10384 213276 10396
rect 74500 10356 213276 10384
rect 74500 10344 74506 10356
rect 213270 10344 213276 10356
rect 213328 10344 213334 10396
rect 246758 10344 246764 10396
rect 246816 10384 246822 10396
rect 251910 10384 251916 10396
rect 246816 10356 251916 10384
rect 246816 10344 246822 10356
rect 251910 10344 251916 10356
rect 251968 10344 251974 10396
rect 60642 10276 60648 10328
rect 60700 10316 60706 10328
rect 210050 10316 210056 10328
rect 60700 10288 210056 10316
rect 60700 10276 60706 10288
rect 210050 10276 210056 10288
rect 210108 10276 210114 10328
rect 220446 10276 220452 10328
rect 220504 10316 220510 10328
rect 233970 10316 233976 10328
rect 220504 10288 233976 10316
rect 220504 10276 220510 10288
rect 233970 10276 233976 10288
rect 234028 10276 234034 10328
rect 250806 10276 250812 10328
rect 250864 10316 250870 10328
rect 298094 10316 298100 10328
rect 250864 10288 298100 10316
rect 250864 10276 250870 10288
rect 298094 10276 298100 10288
rect 298152 10276 298158 10328
rect 299198 10276 299204 10328
rect 299256 10316 299262 10328
rect 576946 10316 576952 10328
rect 299256 10288 576952 10316
rect 299256 10276 299262 10288
rect 576946 10276 576952 10288
rect 577004 10276 577010 10328
rect 111610 9392 111616 9444
rect 111668 9432 111674 9444
rect 218514 9432 218520 9444
rect 111668 9404 218520 9432
rect 111668 9392 111674 9404
rect 218514 9392 218520 9404
rect 218572 9392 218578 9444
rect 108114 9324 108120 9376
rect 108172 9364 108178 9376
rect 218146 9364 218152 9376
rect 108172 9336 218152 9364
rect 108172 9324 108178 9336
rect 218146 9324 218152 9336
rect 218204 9324 218210 9376
rect 104526 9256 104532 9308
rect 104584 9296 104590 9308
rect 217134 9296 217140 9308
rect 104584 9268 217140 9296
rect 104584 9256 104590 9268
rect 217134 9256 217140 9268
rect 217192 9256 217198 9308
rect 101030 9188 101036 9240
rect 101088 9228 101094 9240
rect 217226 9228 217232 9240
rect 101088 9200 217232 9228
rect 101088 9188 101094 9200
rect 217226 9188 217232 9200
rect 217284 9188 217290 9240
rect 97442 9120 97448 9172
rect 97500 9160 97506 9172
rect 216122 9160 216128 9172
rect 97500 9132 216128 9160
rect 97500 9120 97506 9132
rect 216122 9120 216128 9132
rect 216180 9120 216186 9172
rect 93946 9052 93952 9104
rect 94004 9092 94010 9104
rect 215662 9092 215668 9104
rect 94004 9064 215668 9092
rect 94004 9052 94010 9064
rect 215662 9052 215668 9064
rect 215720 9052 215726 9104
rect 281350 9052 281356 9104
rect 281408 9092 281414 9104
rect 469858 9092 469864 9104
rect 281408 9064 469864 9092
rect 281408 9052 281414 9064
rect 469858 9052 469864 9064
rect 469916 9052 469922 9104
rect 79686 8984 79692 9036
rect 79744 9024 79750 9036
rect 212626 9024 212632 9036
rect 79744 8996 212632 9024
rect 79744 8984 79750 8996
rect 212626 8984 212632 8996
rect 212684 8984 212690 9036
rect 226334 8984 226340 9036
rect 226392 9024 226398 9036
rect 233878 9024 233884 9036
rect 226392 8996 233884 9024
rect 226392 8984 226398 8996
rect 233878 8984 233884 8996
rect 233936 8984 233942 9036
rect 281166 8984 281172 9036
rect 281224 9024 281230 9036
rect 473446 9024 473452 9036
rect 281224 8996 473452 9024
rect 281224 8984 281230 8996
rect 473446 8984 473452 8996
rect 473504 8984 473510 9036
rect 76190 8916 76196 8968
rect 76248 8956 76254 8968
rect 212994 8956 213000 8968
rect 76248 8928 213000 8956
rect 76248 8916 76254 8928
rect 212994 8916 213000 8928
rect 213052 8916 213058 8968
rect 281258 8916 281264 8968
rect 281316 8956 281322 8968
rect 476942 8956 476948 8968
rect 281316 8928 476948 8956
rect 281316 8916 281322 8928
rect 476942 8916 476948 8928
rect 477000 8916 477006 8968
rect 222746 8304 222752 8356
rect 222804 8344 222810 8356
rect 231302 8344 231308 8356
rect 222804 8316 231308 8344
rect 222804 8304 222810 8316
rect 231302 8304 231308 8316
rect 231360 8304 231366 8356
rect 265894 8100 265900 8152
rect 265952 8140 265958 8152
rect 388254 8140 388260 8152
rect 265952 8112 388260 8140
rect 265952 8100 265958 8112
rect 388254 8100 388260 8112
rect 388312 8100 388318 8152
rect 267550 8032 267556 8084
rect 267608 8072 267614 8084
rect 391842 8072 391848 8084
rect 267608 8044 391848 8072
rect 267608 8032 267614 8044
rect 391842 8032 391848 8044
rect 391900 8032 391906 8084
rect 267182 7964 267188 8016
rect 267240 8004 267246 8016
rect 395246 8004 395252 8016
rect 267240 7976 395252 8004
rect 267240 7964 267246 7976
rect 395246 7964 395252 7976
rect 395304 7964 395310 8016
rect 268930 7896 268936 7948
rect 268988 7936 268994 7948
rect 398926 7936 398932 7948
rect 268988 7908 398932 7936
rect 268988 7896 268994 7908
rect 398926 7896 398932 7908
rect 398984 7896 398990 7948
rect 269022 7828 269028 7880
rect 269080 7868 269086 7880
rect 402514 7868 402520 7880
rect 269080 7840 402520 7868
rect 269080 7828 269086 7840
rect 402514 7828 402520 7840
rect 402572 7828 402578 7880
rect 270310 7760 270316 7812
rect 270368 7800 270374 7812
rect 406010 7800 406016 7812
rect 270368 7772 406016 7800
rect 270368 7760 270374 7772
rect 406010 7760 406016 7772
rect 406068 7760 406074 7812
rect 192018 7692 192024 7744
rect 192076 7732 192082 7744
rect 232590 7732 232596 7744
rect 192076 7704 232596 7732
rect 192076 7692 192082 7704
rect 232590 7692 232596 7704
rect 232648 7692 232654 7744
rect 270218 7692 270224 7744
rect 270276 7732 270282 7744
rect 409598 7732 409604 7744
rect 270276 7704 409604 7732
rect 270276 7692 270282 7704
rect 409598 7692 409604 7704
rect 409656 7692 409662 7744
rect 24210 7624 24216 7676
rect 24268 7664 24274 7676
rect 94498 7664 94504 7676
rect 24268 7636 94504 7664
rect 24268 7624 24274 7636
rect 94498 7624 94504 7636
rect 94556 7624 94562 7676
rect 145926 7624 145932 7676
rect 145984 7664 145990 7676
rect 224126 7664 224132 7676
rect 145984 7636 224132 7664
rect 145984 7624 145990 7636
rect 224126 7624 224132 7636
rect 224184 7624 224190 7676
rect 269942 7624 269948 7676
rect 270000 7664 270006 7676
rect 413094 7664 413100 7676
rect 270000 7636 413100 7664
rect 270000 7624 270006 7636
rect 413094 7624 413100 7636
rect 413152 7624 413158 7676
rect 43070 7556 43076 7608
rect 43128 7596 43134 7608
rect 188430 7596 188436 7608
rect 43128 7568 188436 7596
rect 43128 7556 43134 7568
rect 188430 7556 188436 7568
rect 188488 7556 188494 7608
rect 188522 7556 188528 7608
rect 188580 7596 188586 7608
rect 232222 7596 232228 7608
rect 188580 7568 232228 7596
rect 188580 7556 188586 7568
rect 232222 7556 232228 7568
rect 232280 7556 232286 7608
rect 253198 7556 253204 7608
rect 253256 7596 253262 7608
rect 266538 7596 266544 7608
rect 253256 7568 266544 7596
rect 253256 7556 253262 7568
rect 266538 7556 266544 7568
rect 266596 7556 266602 7608
rect 273162 7556 273168 7608
rect 273220 7596 273226 7608
rect 427262 7596 427268 7608
rect 273220 7568 427268 7596
rect 273220 7556 273226 7568
rect 427262 7556 427268 7568
rect 427320 7556 427326 7608
rect 99834 6876 99840 6928
rect 99892 6916 99898 6928
rect 104158 6916 104164 6928
rect 99892 6888 104164 6916
rect 99892 6876 99898 6888
rect 104158 6876 104164 6888
rect 104216 6876 104222 6928
rect 3418 6604 3424 6656
rect 3476 6644 3482 6656
rect 7558 6644 7564 6656
rect 3476 6616 7564 6644
rect 3476 6604 3482 6616
rect 7558 6604 7564 6616
rect 7616 6604 7622 6656
rect 215662 6536 215668 6588
rect 215720 6576 215726 6588
rect 236730 6576 236736 6588
rect 215720 6548 236736 6576
rect 215720 6536 215726 6548
rect 236730 6536 236736 6548
rect 236788 6536 236794 6588
rect 249242 6536 249248 6588
rect 249300 6576 249306 6588
rect 284478 6576 284484 6588
rect 249300 6548 284484 6576
rect 249300 6536 249306 6548
rect 284478 6536 284484 6548
rect 284536 6536 284542 6588
rect 342162 6576 342168 6588
rect 335326 6548 342168 6576
rect 205082 6468 205088 6520
rect 205140 6508 205146 6520
rect 234982 6508 234988 6520
rect 205140 6480 234988 6508
rect 205140 6468 205146 6480
rect 234982 6468 234988 6480
rect 235040 6468 235046 6520
rect 250898 6468 250904 6520
rect 250956 6508 250962 6520
rect 297266 6508 297272 6520
rect 250956 6480 297272 6508
rect 250956 6468 250962 6480
rect 297266 6468 297272 6480
rect 297324 6468 297330 6520
rect 194410 6400 194416 6452
rect 194468 6440 194474 6452
rect 232682 6440 232688 6452
rect 194468 6412 232688 6440
rect 194468 6400 194474 6412
rect 232682 6400 232688 6412
rect 232740 6400 232746 6452
rect 259362 6400 259368 6452
rect 259420 6440 259426 6452
rect 335326 6440 335354 6548
rect 342162 6536 342168 6548
rect 342220 6536 342226 6588
rect 345750 6508 345756 6520
rect 259420 6412 335354 6440
rect 340156 6480 345756 6508
rect 259420 6400 259426 6412
rect 190822 6332 190828 6384
rect 190880 6372 190886 6384
rect 232038 6372 232044 6384
rect 190880 6344 232044 6372
rect 190880 6332 190886 6344
rect 232038 6332 232044 6344
rect 232096 6332 232102 6384
rect 259270 6332 259276 6384
rect 259328 6372 259334 6384
rect 340156 6372 340184 6480
rect 345750 6468 345756 6480
rect 345808 6468 345814 6520
rect 418982 6508 418988 6520
rect 412606 6480 418988 6508
rect 341518 6400 341524 6452
rect 341576 6440 341582 6452
rect 379974 6440 379980 6452
rect 341576 6412 379980 6440
rect 341576 6400 341582 6412
rect 379974 6400 379980 6412
rect 380032 6400 380038 6452
rect 394234 6440 394240 6452
rect 383626 6412 394240 6440
rect 352834 6372 352840 6384
rect 259328 6344 340184 6372
rect 344986 6344 352840 6372
rect 259328 6332 259334 6344
rect 14734 6264 14740 6316
rect 14792 6304 14798 6316
rect 124858 6304 124864 6316
rect 14792 6276 124864 6304
rect 14792 6264 14798 6276
rect 124858 6264 124864 6276
rect 124916 6264 124922 6316
rect 187326 6264 187332 6316
rect 187384 6304 187390 6316
rect 232406 6304 232412 6316
rect 187384 6276 232412 6304
rect 187384 6264 187390 6276
rect 232406 6264 232412 6276
rect 232464 6264 232470 6316
rect 260650 6264 260656 6316
rect 260708 6304 260714 6316
rect 344986 6304 345014 6344
rect 352834 6332 352840 6344
rect 352892 6332 352898 6384
rect 260708 6276 345014 6304
rect 260708 6264 260714 6276
rect 352558 6264 352564 6316
rect 352616 6304 352622 6316
rect 383626 6304 383654 6412
rect 394234 6400 394240 6412
rect 394292 6400 394298 6452
rect 388438 6332 388444 6384
rect 388496 6372 388502 6384
rect 412606 6372 412634 6480
rect 418982 6468 418988 6480
rect 419040 6468 419046 6520
rect 422570 6440 422576 6452
rect 388496 6344 412634 6372
rect 416516 6412 422576 6440
rect 388496 6332 388502 6344
rect 352616 6276 383654 6304
rect 352616 6264 352622 6276
rect 393958 6264 393964 6316
rect 394016 6304 394022 6316
rect 416516 6304 416544 6412
rect 422570 6400 422576 6412
rect 422628 6400 422634 6452
rect 418798 6332 418804 6384
rect 418856 6372 418862 6384
rect 443822 6372 443828 6384
rect 418856 6344 443828 6372
rect 418856 6332 418862 6344
rect 443822 6332 443828 6344
rect 443880 6332 443886 6384
rect 394016 6276 416544 6304
rect 394016 6264 394022 6276
rect 71498 6196 71504 6248
rect 71556 6236 71562 6248
rect 71556 6208 204576 6236
rect 71556 6196 71562 6208
rect 62022 6128 62028 6180
rect 62080 6168 62086 6180
rect 204548 6168 204576 6208
rect 208578 6196 208584 6248
rect 208636 6236 208642 6248
rect 234798 6236 234804 6248
rect 208636 6208 234804 6236
rect 208636 6196 208642 6208
rect 234798 6196 234804 6208
rect 234856 6196 234862 6248
rect 249426 6196 249432 6248
rect 249484 6236 249490 6248
rect 287790 6236 287796 6248
rect 249484 6208 287796 6236
rect 249484 6196 249490 6208
rect 287790 6196 287796 6208
rect 287848 6196 287854 6248
rect 287974 6196 287980 6248
rect 288032 6236 288038 6248
rect 514754 6236 514760 6248
rect 288032 6208 514760 6236
rect 288032 6196 288038 6208
rect 514754 6196 514760 6208
rect 514812 6196 514818 6248
rect 209038 6168 209044 6180
rect 62080 6140 200114 6168
rect 204548 6140 209044 6168
rect 62080 6128 62086 6140
rect 200086 6100 200114 6140
rect 209038 6128 209044 6140
rect 209096 6128 209102 6180
rect 212166 6128 212172 6180
rect 212224 6168 212230 6180
rect 236270 6168 236276 6180
rect 212224 6140 236276 6168
rect 212224 6128 212230 6140
rect 236270 6128 236276 6140
rect 236328 6128 236334 6180
rect 249334 6128 249340 6180
rect 249392 6168 249398 6180
rect 291378 6168 291384 6180
rect 249392 6140 291384 6168
rect 249392 6128 249398 6140
rect 291378 6128 291384 6140
rect 291436 6128 291442 6180
rect 291930 6128 291936 6180
rect 291988 6168 291994 6180
rect 536006 6168 536012 6180
rect 291988 6140 536012 6168
rect 291988 6128 291994 6140
rect 536006 6128 536012 6140
rect 536064 6128 536070 6180
rect 210510 6100 210516 6112
rect 200086 6072 210516 6100
rect 210510 6060 210516 6072
rect 210568 6060 210574 6112
rect 124674 5516 124680 5568
rect 124732 5556 124738 5568
rect 126238 5556 126244 5568
rect 124732 5528 126244 5556
rect 124732 5516 124738 5528
rect 126238 5516 126244 5528
rect 126296 5516 126302 5568
rect 245470 5244 245476 5296
rect 245528 5284 245534 5296
rect 265342 5284 265348 5296
rect 245528 5256 265348 5284
rect 245528 5244 245534 5256
rect 265342 5244 265348 5256
rect 265400 5244 265406 5296
rect 304258 5244 304264 5296
rect 304316 5284 304322 5296
rect 358722 5284 358728 5296
rect 304316 5256 358728 5284
rect 304316 5244 304322 5256
rect 358722 5244 358728 5256
rect 358780 5244 358786 5296
rect 249702 5176 249708 5228
rect 249760 5216 249766 5228
rect 290182 5216 290188 5228
rect 249760 5188 290188 5216
rect 249760 5176 249766 5188
rect 290182 5176 290188 5188
rect 290240 5176 290246 5228
rect 309870 5176 309876 5228
rect 309928 5216 309934 5228
rect 372890 5216 372896 5228
rect 309928 5188 372896 5216
rect 309928 5176 309934 5188
rect 372890 5176 372896 5188
rect 372948 5176 372954 5228
rect 35986 5108 35992 5160
rect 36044 5148 36050 5160
rect 50338 5148 50344 5160
rect 36044 5120 50344 5148
rect 36044 5108 36050 5120
rect 50338 5108 50344 5120
rect 50396 5108 50402 5160
rect 58434 5108 58440 5160
rect 58492 5148 58498 5160
rect 58492 5120 64874 5148
rect 58492 5108 58498 5120
rect 39574 5040 39580 5092
rect 39632 5080 39638 5092
rect 58618 5080 58624 5092
rect 39632 5052 58624 5080
rect 39632 5040 39638 5052
rect 58618 5040 58624 5052
rect 58676 5040 58682 5092
rect 64846 5080 64874 5120
rect 131758 5108 131764 5160
rect 131816 5148 131822 5160
rect 222470 5148 222476 5160
rect 131816 5120 222476 5148
rect 131816 5108 131822 5120
rect 222470 5108 222476 5120
rect 222528 5108 222534 5160
rect 245378 5108 245384 5160
rect 245436 5148 245442 5160
rect 261754 5148 261760 5160
rect 245436 5120 261760 5148
rect 245436 5108 245442 5120
rect 261754 5108 261760 5120
rect 261812 5108 261818 5160
rect 262858 5108 262864 5160
rect 262916 5148 262922 5160
rect 355226 5148 355232 5160
rect 262916 5120 355232 5148
rect 262916 5108 262922 5120
rect 355226 5108 355232 5120
rect 355284 5108 355290 5160
rect 377398 5108 377404 5160
rect 377456 5148 377462 5160
rect 411806 5148 411812 5160
rect 377456 5120 411812 5148
rect 377456 5108 377462 5120
rect 411806 5108 411812 5120
rect 411864 5108 411870 5160
rect 411898 5108 411904 5160
rect 411956 5148 411962 5160
rect 436646 5148 436652 5160
rect 411956 5120 436652 5148
rect 411956 5108 411962 5120
rect 436646 5108 436652 5120
rect 436704 5108 436710 5160
rect 443638 5108 443644 5160
rect 443696 5148 443702 5160
rect 472250 5148 472256 5160
rect 443696 5120 472256 5148
rect 443696 5108 443702 5120
rect 472250 5108 472256 5120
rect 472308 5108 472314 5160
rect 209866 5080 209872 5092
rect 64846 5052 209872 5080
rect 209866 5040 209872 5052
rect 209924 5040 209930 5092
rect 246482 5040 246488 5092
rect 246540 5080 246546 5092
rect 268838 5080 268844 5092
rect 246540 5052 268844 5080
rect 246540 5040 246546 5052
rect 268838 5040 268844 5052
rect 268896 5040 268902 5092
rect 271782 5040 271788 5092
rect 271840 5080 271846 5092
rect 415486 5080 415492 5092
rect 271840 5052 415492 5080
rect 271840 5040 271846 5052
rect 415486 5040 415492 5052
rect 415544 5040 415550 5092
rect 436738 5040 436744 5092
rect 436796 5080 436802 5092
rect 465166 5080 465172 5092
rect 436796 5052 465172 5080
rect 436796 5040 436802 5052
rect 465166 5040 465172 5052
rect 465224 5040 465230 5092
rect 47854 4972 47860 5024
rect 47912 5012 47918 5024
rect 207842 5012 207848 5024
rect 47912 4984 207848 5012
rect 47912 4972 47918 4984
rect 207842 4972 207848 4984
rect 207900 4972 207906 5024
rect 221550 4972 221556 5024
rect 221608 5012 221614 5024
rect 237650 5012 237656 5024
rect 221608 4984 237656 5012
rect 221608 4972 221614 4984
rect 237650 4972 237656 4984
rect 237708 4972 237714 5024
rect 251818 4972 251824 5024
rect 251876 5012 251882 5024
rect 279510 5012 279516 5024
rect 251876 4984 279516 5012
rect 251876 4972 251882 4984
rect 279510 4972 279516 4984
rect 279568 4972 279574 5024
rect 286686 4972 286692 5024
rect 286744 5012 286750 5024
rect 504174 5012 504180 5024
rect 286744 4984 504180 5012
rect 286744 4972 286750 4984
rect 504174 4972 504180 4984
rect 504232 4972 504238 5024
rect 2866 4904 2872 4956
rect 2924 4944 2930 4956
rect 200482 4944 200488 4956
rect 2924 4916 200488 4944
rect 2924 4904 2930 4916
rect 200482 4904 200488 4916
rect 200540 4904 200546 4956
rect 218054 4904 218060 4956
rect 218112 4944 218118 4956
rect 236638 4944 236644 4956
rect 218112 4916 236644 4944
rect 218112 4904 218118 4916
rect 236638 4904 236644 4916
rect 236696 4904 236702 4956
rect 249518 4904 249524 4956
rect 249576 4944 249582 4956
rect 286594 4944 286600 4956
rect 249576 4916 286600 4944
rect 249576 4904 249582 4916
rect 286594 4904 286600 4916
rect 286652 4904 286658 4956
rect 289262 4904 289268 4956
rect 289320 4944 289326 4956
rect 519538 4944 519544 4956
rect 289320 4916 519544 4944
rect 289320 4904 289326 4916
rect 519538 4904 519544 4916
rect 519596 4904 519602 4956
rect 1670 4836 1676 4888
rect 1728 4876 1734 4888
rect 200390 4876 200396 4888
rect 1728 4848 200396 4876
rect 1728 4836 1734 4848
rect 200390 4836 200396 4848
rect 200448 4836 200454 4888
rect 214466 4836 214472 4888
rect 214524 4876 214530 4888
rect 236546 4876 236552 4888
rect 214524 4848 236552 4876
rect 214524 4836 214530 4848
rect 236546 4836 236552 4848
rect 236604 4836 236610 4888
rect 249610 4836 249616 4888
rect 249668 4876 249674 4888
rect 288986 4876 288992 4888
rect 249668 4848 288992 4876
rect 249668 4836 249674 4848
rect 288986 4836 288992 4848
rect 289044 4836 289050 4888
rect 289630 4836 289636 4888
rect 289688 4876 289694 4888
rect 523034 4876 523040 4888
rect 289688 4848 523040 4876
rect 289688 4836 289694 4848
rect 523034 4836 523040 4848
rect 523092 4836 523098 4888
rect 566 4768 572 4820
rect 624 4808 630 4820
rect 200574 4808 200580 4820
rect 624 4780 200580 4808
rect 624 4768 630 4780
rect 200574 4768 200580 4780
rect 200632 4768 200638 4820
rect 210970 4768 210976 4820
rect 211028 4808 211034 4820
rect 239030 4808 239036 4820
rect 211028 4780 239036 4808
rect 211028 4768 211034 4780
rect 239030 4768 239036 4780
rect 239088 4768 239094 4820
rect 250990 4768 250996 4820
rect 251048 4808 251054 4820
rect 293678 4808 293684 4820
rect 251048 4780 293684 4808
rect 251048 4768 251054 4780
rect 293678 4768 293684 4780
rect 293736 4768 293742 4820
rect 296254 4768 296260 4820
rect 296312 4808 296318 4820
rect 560846 4808 560852 4820
rect 296312 4780 560852 4808
rect 296312 4768 296318 4780
rect 560846 4768 560852 4780
rect 560904 4768 560910 4820
rect 74368 4168 74580 4196
rect 13538 4088 13544 4140
rect 13596 4128 13602 4140
rect 18598 4128 18604 4140
rect 13596 4100 18604 4128
rect 13596 4088 13602 4100
rect 18598 4088 18604 4100
rect 18656 4088 18662 4140
rect 67910 4088 67916 4140
rect 67968 4128 67974 4140
rect 74368 4128 74396 4168
rect 67968 4100 74396 4128
rect 74552 4128 74580 4168
rect 256988 4168 258488 4196
rect 97258 4128 97264 4140
rect 74552 4100 97264 4128
rect 67968 4088 67974 4100
rect 97258 4088 97264 4100
rect 97316 4088 97322 4140
rect 103330 4088 103336 4140
rect 103388 4128 103394 4140
rect 112438 4128 112444 4140
rect 103388 4100 112444 4128
rect 103388 4088 103394 4100
rect 112438 4088 112444 4100
rect 112496 4088 112502 4140
rect 129366 4088 129372 4140
rect 129424 4128 129430 4140
rect 221090 4128 221096 4140
rect 129424 4100 221096 4128
rect 129424 4088 129430 4100
rect 221090 4088 221096 4100
rect 221148 4088 221154 4140
rect 246298 4088 246304 4140
rect 246356 4128 246362 4140
rect 248782 4128 248788 4140
rect 246356 4100 248788 4128
rect 246356 4088 246362 4100
rect 248782 4088 248788 4100
rect 248840 4088 248846 4140
rect 252094 4088 252100 4140
rect 252152 4128 252158 4140
rect 256988 4128 257016 4168
rect 252152 4100 257016 4128
rect 252152 4088 252158 4100
rect 257062 4088 257068 4140
rect 257120 4128 257126 4140
rect 258350 4128 258356 4140
rect 257120 4100 258356 4128
rect 257120 4088 257126 4100
rect 258350 4088 258356 4100
rect 258408 4088 258414 4140
rect 12342 4020 12348 4072
rect 12400 4060 12406 4072
rect 17218 4060 17224 4072
rect 12400 4032 17224 4060
rect 12400 4020 12406 4032
rect 17218 4020 17224 4032
rect 17276 4020 17282 4072
rect 34790 4020 34796 4072
rect 34848 4060 34854 4072
rect 43438 4060 43444 4072
rect 34848 4032 43444 4060
rect 34848 4020 34854 4032
rect 43438 4020 43444 4032
rect 43496 4020 43502 4072
rect 50154 4020 50160 4072
rect 50212 4060 50218 4072
rect 79318 4060 79324 4072
rect 50212 4032 79324 4060
rect 50212 4020 50218 4032
rect 79318 4020 79324 4032
rect 79376 4020 79382 4072
rect 87414 4020 87420 4072
rect 87472 4060 87478 4072
rect 108298 4060 108304 4072
rect 87472 4032 108304 4060
rect 87472 4020 87478 4032
rect 108298 4020 108304 4032
rect 108356 4020 108362 4072
rect 117590 4020 117596 4072
rect 117648 4060 117654 4072
rect 217318 4060 217324 4072
rect 117648 4032 217324 4060
rect 117648 4020 117654 4032
rect 217318 4020 217324 4032
rect 217376 4020 217382 4072
rect 238110 4020 238116 4072
rect 238168 4060 238174 4072
rect 240594 4060 240600 4072
rect 238168 4032 240600 4060
rect 238168 4020 238174 4032
rect 240594 4020 240600 4032
rect 240652 4020 240658 4072
rect 243906 4020 243912 4072
rect 243964 4060 243970 4072
rect 254670 4060 254676 4072
rect 243964 4032 254676 4060
rect 243964 4020 243970 4032
rect 254670 4020 254676 4032
rect 254728 4020 254734 4072
rect 255958 4020 255964 4072
rect 256016 4060 256022 4072
rect 258074 4060 258080 4072
rect 256016 4032 258080 4060
rect 256016 4020 256022 4032
rect 258074 4020 258080 4032
rect 258132 4020 258138 4072
rect 258460 4060 258488 4168
rect 261478 4088 261484 4140
rect 261536 4128 261542 4140
rect 277118 4128 277124 4140
rect 261536 4100 277124 4128
rect 261536 4088 261542 4100
rect 277118 4088 277124 4100
rect 277176 4088 277182 4140
rect 278222 4088 278228 4140
rect 278280 4128 278286 4140
rect 284662 4128 284668 4140
rect 278280 4100 284668 4128
rect 278280 4088 278286 4100
rect 284662 4088 284668 4100
rect 284720 4088 284726 4140
rect 292574 4088 292580 4140
rect 292632 4128 292638 4140
rect 299566 4128 299572 4140
rect 292632 4100 299572 4128
rect 292632 4088 292638 4100
rect 299566 4088 299572 4100
rect 299624 4088 299630 4140
rect 363598 4088 363604 4140
rect 363656 4128 363662 4140
rect 364610 4128 364616 4140
rect 363656 4100 364616 4128
rect 363656 4088 363662 4100
rect 364610 4088 364616 4100
rect 364668 4088 364674 4140
rect 406378 4088 406384 4140
rect 406436 4128 406442 4140
rect 414290 4128 414296 4140
rect 406436 4100 414296 4128
rect 406436 4088 406442 4100
rect 414290 4088 414296 4100
rect 414348 4088 414354 4140
rect 471238 4088 471244 4140
rect 471296 4128 471302 4140
rect 475838 4128 475844 4140
rect 471296 4100 475844 4128
rect 471296 4088 471302 4100
rect 475838 4088 475844 4100
rect 475896 4088 475902 4140
rect 479518 4088 479524 4140
rect 479576 4128 479582 4140
rect 480530 4128 480536 4140
rect 479576 4100 480536 4128
rect 479576 4088 479582 4100
rect 480530 4088 480536 4100
rect 480588 4088 480594 4140
rect 566550 4088 566556 4140
rect 566608 4128 566614 4140
rect 568022 4128 568028 4140
rect 566608 4100 568028 4128
rect 566608 4088 566614 4100
rect 568022 4088 568028 4100
rect 568080 4088 568086 4140
rect 305546 4060 305552 4072
rect 258460 4032 305552 4060
rect 305546 4020 305552 4032
rect 305604 4020 305610 4072
rect 475378 4020 475384 4072
rect 475436 4060 475442 4072
rect 487614 4060 487620 4072
rect 475436 4032 487620 4060
rect 475436 4020 475442 4032
rect 487614 4020 487620 4032
rect 487672 4020 487678 4072
rect 20622 3952 20628 4004
rect 20680 3992 20686 4004
rect 20680 3964 35894 3992
rect 20680 3952 20686 3964
rect 21818 3816 21824 3868
rect 21876 3856 21882 3868
rect 29638 3856 29644 3868
rect 21876 3828 29644 3856
rect 21876 3816 21882 3828
rect 29638 3816 29644 3828
rect 29696 3816 29702 3868
rect 35866 3856 35894 3964
rect 37182 3952 37188 4004
rect 37240 3992 37246 4004
rect 47578 3992 47584 4004
rect 37240 3964 47584 3992
rect 37240 3952 37246 3964
rect 47578 3952 47584 3964
rect 47636 3952 47642 4004
rect 57330 3952 57336 4004
rect 57388 3992 57394 4004
rect 88978 3992 88984 4004
rect 57388 3964 88984 3992
rect 57388 3952 57394 3964
rect 88978 3952 88984 3964
rect 89036 3952 89042 4004
rect 96246 3952 96252 4004
rect 96304 3992 96310 4004
rect 105538 3992 105544 4004
rect 96304 3964 105544 3992
rect 96304 3952 96310 3964
rect 105538 3952 105544 3964
rect 105596 3952 105602 4004
rect 110506 3952 110512 4004
rect 110564 3992 110570 4004
rect 215938 3992 215944 4004
rect 110564 3964 215944 3992
rect 110564 3952 110570 3964
rect 215938 3952 215944 3964
rect 215996 3952 216002 4004
rect 225138 3952 225144 4004
rect 225196 3992 225202 4004
rect 234062 3992 234068 4004
rect 225196 3964 234068 3992
rect 225196 3952 225202 3964
rect 234062 3952 234068 3964
rect 234120 3952 234126 4004
rect 242434 3952 242440 4004
rect 242492 3992 242498 4004
rect 249978 3992 249984 4004
rect 242492 3964 249984 3992
rect 242492 3952 242498 3964
rect 249978 3952 249984 3964
rect 250036 3952 250042 4004
rect 252002 3952 252008 4004
rect 252060 3992 252066 4004
rect 307938 3992 307944 4004
rect 252060 3964 307944 3992
rect 252060 3952 252066 3964
rect 307938 3952 307944 3964
rect 307996 3952 308002 4004
rect 428458 3952 428464 4004
rect 428516 3992 428522 4004
rect 445018 3992 445024 4004
rect 428516 3964 445024 3992
rect 428516 3952 428522 3964
rect 445018 3952 445024 3964
rect 445076 3952 445082 4004
rect 472618 3952 472624 4004
rect 472676 3992 472682 4004
rect 491110 3992 491116 4004
rect 472676 3964 491116 3992
rect 472676 3952 472682 3964
rect 491110 3952 491116 3964
rect 491168 3952 491174 4004
rect 40678 3884 40684 3936
rect 40736 3924 40742 3936
rect 53098 3924 53104 3936
rect 40736 3896 53104 3924
rect 40736 3884 40742 3896
rect 53098 3884 53104 3896
rect 53156 3884 53162 3936
rect 54938 3884 54944 3936
rect 54996 3924 55002 3936
rect 61378 3924 61384 3936
rect 54996 3896 61384 3924
rect 54996 3884 55002 3896
rect 61378 3884 61384 3896
rect 61436 3884 61442 3936
rect 63218 3884 63224 3936
rect 63276 3924 63282 3936
rect 210234 3924 210240 3936
rect 63276 3896 210240 3924
rect 63276 3884 63282 3896
rect 210234 3884 210240 3896
rect 210292 3884 210298 3936
rect 223758 3884 223764 3936
rect 223816 3924 223822 3936
rect 228542 3924 228548 3936
rect 223816 3896 228548 3924
rect 223816 3884 223822 3896
rect 228542 3884 228548 3896
rect 228600 3884 228606 3936
rect 228726 3884 228732 3936
rect 228784 3924 228790 3936
rect 237926 3924 237932 3936
rect 228784 3896 237932 3924
rect 228784 3884 228790 3896
rect 237926 3884 237932 3896
rect 237984 3884 237990 3936
rect 260742 3884 260748 3936
rect 260800 3924 260806 3936
rect 349246 3924 349252 3936
rect 260800 3896 349252 3924
rect 260800 3884 260806 3896
rect 349246 3884 349252 3896
rect 349304 3884 349310 3936
rect 395338 3884 395344 3936
rect 395396 3924 395402 3936
rect 397730 3924 397736 3936
rect 395396 3896 397736 3924
rect 395396 3884 395402 3896
rect 397730 3884 397736 3896
rect 397788 3884 397794 3936
rect 425790 3884 425796 3936
rect 425848 3924 425854 3936
rect 450906 3924 450912 3936
rect 425848 3896 450912 3924
rect 425848 3884 425854 3896
rect 450906 3884 450912 3896
rect 450964 3884 450970 3936
rect 461578 3884 461584 3936
rect 461636 3924 461642 3936
rect 498194 3924 498200 3936
rect 461636 3896 498200 3924
rect 461636 3884 461642 3896
rect 498194 3884 498200 3896
rect 498252 3884 498258 3936
rect 39298 3856 39304 3868
rect 35866 3828 39304 3856
rect 39298 3816 39304 3828
rect 39356 3816 39362 3868
rect 52546 3816 52552 3868
rect 52604 3856 52610 3868
rect 208670 3856 208676 3868
rect 52604 3828 208676 3856
rect 52604 3816 52610 3828
rect 208670 3816 208676 3828
rect 208728 3816 208734 3868
rect 219250 3816 219256 3868
rect 219308 3856 219314 3868
rect 228358 3856 228364 3868
rect 219308 3828 228364 3856
rect 219308 3816 219314 3828
rect 228358 3816 228364 3828
rect 228416 3816 228422 3868
rect 244090 3816 244096 3868
rect 244148 3856 244154 3868
rect 255866 3856 255872 3868
rect 244148 3828 255872 3856
rect 244148 3816 244154 3828
rect 255866 3816 255872 3828
rect 255924 3816 255930 3868
rect 264882 3816 264888 3868
rect 264940 3856 264946 3868
rect 377674 3856 377680 3868
rect 264940 3828 377680 3856
rect 264940 3816 264946 3828
rect 377674 3816 377680 3828
rect 377732 3816 377738 3868
rect 392670 3816 392676 3868
rect 392728 3856 392734 3868
rect 408402 3856 408408 3868
rect 392728 3828 408408 3856
rect 392728 3816 392734 3828
rect 408402 3816 408408 3828
rect 408460 3816 408466 3868
rect 414658 3816 414664 3868
rect 414716 3856 414722 3868
rect 462774 3856 462780 3868
rect 414716 3828 462780 3856
rect 414716 3816 414722 3828
rect 462774 3816 462780 3828
rect 462832 3816 462838 3868
rect 468478 3816 468484 3868
rect 468536 3856 468542 3868
rect 494698 3856 494704 3868
rect 468536 3828 494704 3856
rect 468536 3816 468542 3828
rect 494698 3816 494704 3828
rect 494756 3816 494762 3868
rect 519630 3816 519636 3868
rect 519688 3856 519694 3868
rect 540790 3856 540796 3868
rect 519688 3828 540796 3856
rect 519688 3816 519694 3828
rect 540790 3816 540796 3828
rect 540848 3816 540854 3868
rect 547138 3816 547144 3868
rect 547196 3856 547202 3868
rect 552658 3856 552664 3868
rect 547196 3828 552664 3856
rect 547196 3816 547202 3828
rect 552658 3816 552664 3828
rect 552716 3816 552722 3868
rect 11146 3748 11152 3800
rect 11204 3788 11210 3800
rect 35158 3788 35164 3800
rect 11204 3760 35164 3788
rect 11204 3748 11210 3760
rect 35158 3748 35164 3760
rect 35216 3748 35222 3800
rect 44266 3748 44272 3800
rect 44324 3788 44330 3800
rect 207382 3788 207388 3800
rect 44324 3760 207388 3788
rect 44324 3748 44330 3760
rect 207382 3748 207388 3760
rect 207440 3748 207446 3800
rect 216858 3748 216864 3800
rect 216916 3788 216922 3800
rect 229738 3788 229744 3800
rect 216916 3760 229744 3788
rect 216916 3748 216922 3760
rect 229738 3748 229744 3760
rect 229796 3748 229802 3800
rect 245194 3748 245200 3800
rect 245252 3788 245258 3800
rect 262950 3788 262956 3800
rect 245252 3760 262956 3788
rect 245252 3748 245258 3760
rect 262950 3748 262956 3760
rect 263008 3748 263014 3800
rect 264238 3748 264244 3800
rect 264296 3788 264302 3800
rect 276014 3788 276020 3800
rect 264296 3760 276020 3788
rect 264296 3748 264302 3760
rect 276014 3748 276020 3760
rect 276072 3748 276078 3800
rect 278406 3748 278412 3800
rect 278464 3788 278470 3800
rect 454494 3788 454500 3800
rect 278464 3760 454500 3788
rect 278464 3748 278470 3760
rect 454494 3748 454500 3760
rect 454552 3748 454558 3800
rect 465718 3748 465724 3800
rect 465776 3788 465782 3800
rect 565630 3788 565636 3800
rect 465776 3760 565636 3788
rect 465776 3748 465782 3760
rect 565630 3748 565636 3760
rect 565688 3748 565694 3800
rect 16022 3680 16028 3732
rect 16080 3720 16086 3732
rect 16080 3692 16574 3720
rect 16080 3680 16086 3692
rect 7650 3612 7656 3664
rect 7708 3652 7714 3664
rect 16546 3652 16574 3692
rect 25314 3680 25320 3732
rect 25372 3720 25378 3732
rect 204622 3720 204628 3732
rect 25372 3692 204628 3720
rect 25372 3680 25378 3692
rect 204622 3680 204628 3692
rect 204680 3680 204686 3732
rect 213362 3680 213368 3732
rect 213420 3720 213426 3732
rect 228450 3720 228456 3732
rect 213420 3692 228456 3720
rect 213420 3680 213426 3692
rect 228450 3680 228456 3692
rect 228508 3680 228514 3732
rect 243998 3680 244004 3732
rect 244056 3720 244062 3732
rect 259454 3720 259460 3732
rect 244056 3692 259460 3720
rect 244056 3680 244062 3692
rect 259454 3680 259460 3692
rect 259512 3680 259518 3732
rect 260098 3680 260104 3732
rect 260156 3720 260162 3732
rect 278314 3720 278320 3732
rect 260156 3692 278320 3720
rect 260156 3680 260162 3692
rect 278314 3680 278320 3692
rect 278372 3680 278378 3732
rect 280062 3680 280068 3732
rect 280120 3720 280126 3732
rect 280120 3692 284616 3720
rect 280120 3680 280126 3692
rect 200022 3652 200028 3664
rect 7708 3624 15976 3652
rect 16546 3624 200028 3652
rect 7708 3612 7714 3624
rect 8754 3544 8760 3596
rect 8812 3584 8818 3596
rect 15838 3584 15844 3596
rect 8812 3556 15844 3584
rect 8812 3544 8818 3556
rect 15838 3544 15844 3556
rect 15896 3544 15902 3596
rect 15948 3584 15976 3624
rect 200022 3612 200028 3624
rect 200080 3612 200086 3664
rect 209774 3612 209780 3664
rect 209832 3652 209838 3664
rect 231210 3652 231216 3664
rect 209832 3624 231216 3652
rect 209832 3612 209838 3624
rect 231210 3612 231216 3624
rect 231268 3612 231274 3664
rect 242618 3612 242624 3664
rect 242676 3652 242682 3664
rect 251174 3652 251180 3664
rect 242676 3624 251180 3652
rect 242676 3612 242682 3624
rect 251174 3612 251180 3624
rect 251232 3612 251238 3664
rect 251910 3612 251916 3664
rect 251968 3652 251974 3664
rect 271230 3652 271236 3664
rect 251968 3624 271236 3652
rect 251968 3612 251974 3624
rect 271230 3612 271236 3624
rect 271288 3612 271294 3664
rect 280982 3612 280988 3664
rect 281040 3652 281046 3664
rect 284588 3652 284616 3692
rect 284662 3680 284668 3732
rect 284720 3720 284726 3732
rect 461578 3720 461584 3732
rect 284720 3692 461584 3720
rect 284720 3680 284726 3692
rect 461578 3680 461584 3692
rect 461636 3680 461642 3732
rect 467190 3680 467196 3732
rect 467248 3720 467254 3732
rect 573910 3720 573916 3732
rect 467248 3692 573916 3720
rect 467248 3680 467254 3692
rect 573910 3680 573916 3692
rect 573968 3680 573974 3732
rect 468662 3652 468668 3664
rect 281040 3624 284524 3652
rect 284588 3624 468668 3652
rect 281040 3612 281046 3624
rect 200390 3584 200396 3596
rect 15948 3556 200396 3584
rect 200390 3544 200396 3556
rect 200448 3544 200454 3596
rect 201770 3584 201776 3596
rect 200960 3556 201776 3584
rect 6454 3476 6460 3528
rect 6512 3516 6518 3528
rect 193122 3516 193128 3528
rect 6512 3488 193128 3516
rect 6512 3476 6518 3488
rect 193122 3476 193128 3488
rect 193180 3476 193186 3528
rect 193214 3476 193220 3528
rect 193272 3516 193278 3528
rect 194502 3516 194508 3528
rect 193272 3488 194508 3516
rect 193272 3476 193278 3488
rect 194502 3476 194508 3488
rect 194560 3476 194566 3528
rect 196802 3476 196808 3528
rect 196860 3516 196866 3528
rect 197262 3516 197268 3528
rect 196860 3488 197268 3516
rect 196860 3476 196866 3488
rect 197262 3476 197268 3488
rect 197320 3476 197326 3528
rect 197906 3476 197912 3528
rect 197964 3516 197970 3528
rect 198642 3516 198648 3528
rect 197964 3488 198648 3516
rect 197964 3476 197970 3488
rect 198642 3476 198648 3488
rect 198700 3476 198706 3528
rect 199102 3476 199108 3528
rect 199160 3516 199166 3528
rect 199930 3516 199936 3528
rect 199160 3488 199936 3516
rect 199160 3476 199166 3488
rect 199930 3476 199936 3488
rect 199988 3476 199994 3528
rect 200022 3476 200028 3528
rect 200080 3516 200086 3528
rect 200960 3516 200988 3556
rect 201770 3544 201776 3556
rect 201828 3544 201834 3596
rect 207382 3544 207388 3596
rect 207440 3584 207446 3596
rect 231118 3584 231124 3596
rect 207440 3556 231124 3584
rect 207440 3544 207446 3556
rect 231118 3544 231124 3556
rect 231176 3544 231182 3596
rect 246574 3544 246580 3596
rect 246632 3584 246638 3596
rect 271046 3584 271052 3596
rect 246632 3556 271052 3584
rect 246632 3544 246638 3556
rect 271046 3544 271052 3556
rect 271104 3544 271110 3596
rect 271138 3544 271144 3596
rect 271196 3584 271202 3596
rect 274818 3584 274824 3596
rect 271196 3556 274824 3584
rect 271196 3544 271202 3556
rect 274818 3544 274824 3556
rect 274876 3544 274882 3596
rect 281902 3544 281908 3596
rect 281960 3584 281966 3596
rect 284386 3584 284392 3596
rect 281960 3556 284392 3584
rect 281960 3544 281966 3556
rect 284386 3544 284392 3556
rect 284444 3544 284450 3596
rect 284496 3584 284524 3624
rect 468662 3612 468668 3624
rect 468720 3612 468726 3664
rect 475746 3652 475752 3664
rect 470566 3624 475752 3652
rect 470566 3584 470594 3624
rect 475746 3612 475752 3624
rect 475804 3612 475810 3664
rect 475838 3612 475844 3664
rect 475896 3652 475902 3664
rect 485222 3652 485228 3664
rect 475896 3624 485228 3652
rect 475896 3612 475902 3624
rect 485222 3612 485228 3624
rect 485280 3612 485286 3664
rect 485332 3624 488948 3652
rect 284496 3556 470594 3584
rect 472710 3544 472716 3596
rect 472768 3584 472774 3596
rect 474550 3584 474556 3596
rect 472768 3556 474556 3584
rect 472768 3544 472774 3556
rect 474550 3544 474556 3556
rect 474608 3544 474614 3596
rect 485038 3544 485044 3596
rect 485096 3584 485102 3596
rect 485332 3584 485360 3624
rect 485096 3556 485360 3584
rect 485096 3544 485102 3556
rect 486418 3544 486424 3596
rect 486476 3584 486482 3596
rect 488810 3584 488816 3596
rect 486476 3556 488816 3584
rect 486476 3544 486482 3556
rect 488810 3544 488816 3556
rect 488868 3544 488874 3596
rect 488920 3584 488948 3624
rect 489178 3612 489184 3664
rect 489236 3652 489242 3664
rect 515950 3652 515956 3664
rect 489236 3624 515956 3652
rect 489236 3612 489242 3624
rect 515950 3612 515956 3624
rect 516008 3612 516014 3664
rect 518158 3612 518164 3664
rect 518216 3652 518222 3664
rect 529106 3652 529112 3664
rect 518216 3624 529112 3652
rect 518216 3612 518222 3624
rect 529106 3612 529112 3624
rect 529164 3612 529170 3664
rect 529198 3612 529204 3664
rect 529256 3652 529262 3664
rect 531314 3652 531320 3664
rect 529256 3624 531320 3652
rect 529256 3612 529262 3624
rect 531314 3612 531320 3624
rect 531372 3612 531378 3664
rect 536098 3612 536104 3664
rect 536156 3652 536162 3664
rect 556154 3652 556160 3664
rect 536156 3624 556160 3652
rect 536156 3612 536162 3624
rect 556154 3612 556160 3624
rect 556212 3612 556218 3664
rect 547874 3584 547880 3596
rect 488920 3556 547880 3584
rect 547874 3544 547880 3556
rect 547932 3544 547938 3596
rect 560938 3544 560944 3596
rect 560996 3584 561002 3596
rect 563238 3584 563244 3596
rect 560996 3556 563244 3584
rect 560996 3544 561002 3556
rect 563238 3544 563244 3556
rect 563296 3544 563302 3596
rect 565078 3544 565084 3596
rect 565136 3584 565142 3596
rect 570322 3584 570328 3596
rect 565136 3556 570328 3584
rect 565136 3544 565142 3556
rect 570322 3544 570328 3556
rect 570380 3544 570386 3596
rect 200080 3488 200988 3516
rect 200080 3476 200086 3488
rect 201494 3476 201500 3528
rect 201552 3516 201558 3528
rect 223758 3516 223764 3528
rect 201552 3488 223764 3516
rect 201552 3476 201558 3488
rect 223758 3476 223764 3488
rect 223816 3476 223822 3528
rect 223942 3476 223948 3528
rect 224000 3516 224006 3528
rect 224862 3516 224868 3528
rect 224000 3488 224868 3516
rect 224000 3476 224006 3488
rect 224862 3476 224868 3488
rect 224920 3476 224926 3528
rect 229830 3476 229836 3528
rect 229888 3516 229894 3528
rect 230382 3516 230388 3528
rect 229888 3488 230388 3516
rect 229888 3476 229894 3488
rect 230382 3476 230388 3488
rect 230440 3476 230446 3528
rect 234614 3476 234620 3528
rect 234672 3516 234678 3528
rect 238202 3516 238208 3528
rect 234672 3488 238208 3516
rect 234672 3476 234678 3488
rect 238202 3476 238208 3488
rect 238260 3476 238266 3528
rect 242158 3476 242164 3528
rect 242216 3516 242222 3528
rect 242894 3516 242900 3528
rect 242216 3488 242900 3516
rect 242216 3476 242222 3488
rect 242894 3476 242900 3488
rect 242952 3476 242958 3528
rect 248046 3476 248052 3528
rect 248104 3516 248110 3528
rect 280706 3516 280712 3528
rect 248104 3488 280712 3516
rect 248104 3476 248110 3488
rect 280706 3476 280712 3488
rect 280764 3476 280770 3528
rect 282178 3476 282184 3528
rect 282236 3516 282242 3528
rect 283098 3516 283104 3528
rect 282236 3488 283104 3516
rect 282236 3476 282242 3488
rect 283098 3476 283104 3488
rect 283156 3476 283162 3528
rect 284294 3476 284300 3528
rect 284352 3516 284358 3528
rect 285398 3516 285404 3528
rect 284352 3488 285404 3516
rect 284352 3476 284358 3488
rect 285398 3476 285404 3488
rect 285456 3476 285462 3528
rect 300762 3476 300768 3528
rect 300820 3516 300826 3528
rect 302326 3516 302332 3528
rect 300820 3488 302332 3516
rect 300820 3476 300826 3488
rect 302326 3476 302332 3488
rect 302384 3476 302390 3528
rect 302436 3488 580120 3516
rect 4062 3408 4068 3460
rect 4120 3448 4126 3460
rect 200666 3448 200672 3460
rect 4120 3420 200672 3448
rect 4120 3408 4126 3420
rect 200666 3408 200672 3420
rect 200724 3408 200730 3460
rect 206186 3408 206192 3460
rect 206244 3448 206250 3460
rect 206244 3420 229094 3448
rect 206244 3408 206250 3420
rect 17034 3340 17040 3392
rect 17092 3380 17098 3392
rect 21358 3380 21364 3392
rect 17092 3352 21364 3380
rect 17092 3340 17098 3352
rect 21358 3340 21364 3352
rect 21416 3340 21422 3392
rect 27706 3340 27712 3392
rect 27764 3380 27770 3392
rect 28902 3380 28908 3392
rect 27764 3352 28908 3380
rect 27764 3340 27770 3352
rect 28902 3340 28908 3352
rect 28960 3340 28966 3392
rect 32398 3340 32404 3392
rect 32456 3380 32462 3392
rect 33042 3380 33048 3392
rect 32456 3352 33048 3380
rect 32456 3340 32462 3352
rect 33042 3340 33048 3352
rect 33100 3340 33106 3392
rect 33594 3340 33600 3392
rect 33652 3380 33658 3392
rect 40586 3380 40592 3392
rect 33652 3352 40592 3380
rect 33652 3340 33658 3352
rect 40586 3340 40592 3352
rect 40644 3340 40650 3392
rect 41874 3340 41880 3392
rect 41932 3380 41938 3392
rect 43530 3380 43536 3392
rect 41932 3352 43536 3380
rect 41932 3340 41938 3352
rect 43530 3340 43536 3352
rect 43588 3340 43594 3392
rect 51350 3340 51356 3392
rect 51408 3380 51414 3392
rect 54478 3380 54484 3392
rect 51408 3352 54484 3380
rect 51408 3340 51414 3352
rect 54478 3340 54484 3352
rect 54536 3340 54542 3392
rect 55186 3352 65472 3380
rect 19426 3272 19432 3324
rect 19484 3312 19490 3324
rect 25498 3312 25504 3324
rect 19484 3284 25504 3312
rect 19484 3272 19490 3284
rect 25498 3272 25504 3284
rect 25556 3272 25562 3324
rect 48958 3272 48964 3324
rect 49016 3312 49022 3324
rect 55186 3312 55214 3352
rect 49016 3284 55214 3312
rect 49016 3272 49022 3284
rect 56042 3272 56048 3324
rect 56100 3312 56106 3324
rect 57238 3312 57244 3324
rect 56100 3284 57244 3312
rect 56100 3272 56106 3284
rect 57238 3272 57244 3284
rect 57296 3272 57302 3324
rect 59630 3272 59636 3324
rect 59688 3312 59694 3324
rect 60642 3312 60648 3324
rect 59688 3284 60648 3312
rect 59688 3272 59694 3284
rect 60642 3272 60648 3284
rect 60700 3272 60706 3324
rect 60826 3272 60832 3324
rect 60884 3312 60890 3324
rect 65444 3312 65472 3352
rect 65518 3340 65524 3392
rect 65576 3380 65582 3392
rect 66162 3380 66168 3392
rect 65576 3352 66168 3380
rect 65576 3340 65582 3352
rect 66162 3340 66168 3352
rect 66220 3340 66226 3392
rect 69106 3340 69112 3392
rect 69164 3380 69170 3392
rect 70302 3380 70308 3392
rect 69164 3352 70308 3380
rect 69164 3340 69170 3352
rect 70302 3340 70308 3352
rect 70360 3340 70366 3392
rect 72602 3340 72608 3392
rect 72660 3380 72666 3392
rect 73062 3380 73068 3392
rect 72660 3352 73068 3380
rect 72660 3340 72666 3352
rect 73062 3340 73068 3352
rect 73120 3340 73126 3392
rect 73798 3340 73804 3392
rect 73856 3380 73862 3392
rect 74442 3380 74448 3392
rect 73856 3352 74448 3380
rect 73856 3340 73862 3352
rect 74442 3340 74448 3352
rect 74500 3340 74506 3392
rect 77386 3340 77392 3392
rect 77444 3380 77450 3392
rect 78582 3380 78588 3392
rect 77444 3352 78588 3380
rect 77444 3340 77450 3352
rect 78582 3340 78588 3352
rect 78640 3340 78646 3392
rect 78692 3352 98684 3380
rect 68278 3312 68284 3324
rect 60884 3284 65380 3312
rect 65444 3284 68284 3312
rect 60884 3272 60890 3284
rect 26510 3204 26516 3256
rect 26568 3244 26574 3256
rect 33778 3244 33784 3256
rect 26568 3216 33784 3244
rect 26568 3204 26574 3216
rect 33778 3204 33784 3216
rect 33836 3204 33842 3256
rect 64322 3204 64328 3256
rect 64380 3244 64386 3256
rect 64782 3244 64788 3256
rect 64380 3216 64788 3244
rect 64380 3204 64386 3216
rect 64782 3204 64788 3216
rect 64840 3204 64846 3256
rect 9950 3136 9956 3188
rect 10008 3176 10014 3188
rect 14458 3176 14464 3188
rect 10008 3148 14464 3176
rect 10008 3136 10014 3148
rect 14458 3136 14464 3148
rect 14516 3136 14522 3188
rect 18230 3136 18236 3188
rect 18288 3176 18294 3188
rect 22738 3176 22744 3188
rect 18288 3148 22744 3176
rect 18288 3136 18294 3148
rect 22738 3136 22744 3148
rect 22796 3136 22802 3188
rect 65352 3176 65380 3284
rect 68278 3272 68284 3284
rect 68336 3272 68342 3324
rect 66714 3204 66720 3256
rect 66772 3244 66778 3256
rect 75178 3244 75184 3256
rect 66772 3216 75184 3244
rect 66772 3204 66778 3216
rect 75178 3204 75184 3216
rect 75236 3204 75242 3256
rect 71038 3176 71044 3188
rect 65352 3148 71044 3176
rect 71038 3136 71044 3148
rect 71096 3136 71102 3188
rect 74994 3136 75000 3188
rect 75052 3176 75058 3188
rect 78692 3176 78720 3352
rect 98546 3312 98552 3324
rect 75052 3148 78720 3176
rect 78784 3284 98552 3312
rect 75052 3136 75058 3148
rect 28902 3068 28908 3120
rect 28960 3108 28966 3120
rect 32306 3108 32312 3120
rect 28960 3080 32312 3108
rect 28960 3068 28966 3080
rect 32306 3068 32312 3080
rect 32364 3068 32370 3120
rect 78582 3068 78588 3120
rect 78640 3108 78646 3120
rect 78784 3108 78812 3284
rect 98546 3272 98552 3284
rect 98604 3272 98610 3324
rect 98656 3312 98684 3352
rect 102226 3340 102232 3392
rect 102284 3380 102290 3392
rect 103422 3380 103428 3392
rect 102284 3352 103428 3380
rect 102284 3340 102290 3352
rect 103422 3340 103428 3352
rect 103480 3340 103486 3392
rect 105722 3340 105728 3392
rect 105780 3380 105786 3392
rect 106182 3380 106188 3392
rect 105780 3352 106188 3380
rect 105780 3340 105786 3352
rect 106182 3340 106188 3352
rect 106240 3340 106246 3392
rect 106918 3340 106924 3392
rect 106976 3380 106982 3392
rect 107562 3380 107568 3392
rect 106976 3352 107568 3380
rect 106976 3340 106982 3352
rect 107562 3340 107568 3352
rect 107620 3340 107626 3392
rect 109310 3340 109316 3392
rect 109368 3380 109374 3392
rect 110322 3380 110328 3392
rect 109368 3352 110328 3380
rect 109368 3340 109374 3352
rect 110322 3340 110328 3352
rect 110380 3340 110386 3392
rect 114002 3340 114008 3392
rect 114060 3380 114066 3392
rect 115198 3380 115204 3392
rect 114060 3352 115204 3380
rect 114060 3340 114066 3352
rect 115198 3340 115204 3352
rect 115256 3340 115262 3392
rect 116394 3340 116400 3392
rect 116452 3380 116458 3392
rect 117222 3380 117228 3392
rect 116452 3352 117228 3380
rect 116452 3340 116458 3352
rect 117222 3340 117228 3352
rect 117280 3340 117286 3392
rect 122282 3340 122288 3392
rect 122340 3380 122346 3392
rect 122742 3380 122748 3392
rect 122340 3352 122748 3380
rect 122340 3340 122346 3352
rect 122742 3340 122748 3352
rect 122800 3340 122806 3392
rect 123478 3340 123484 3392
rect 123536 3380 123542 3392
rect 124122 3380 124128 3392
rect 123536 3352 124128 3380
rect 123536 3340 123542 3352
rect 124122 3340 124128 3352
rect 124180 3340 124186 3392
rect 125870 3340 125876 3392
rect 125928 3380 125934 3392
rect 126882 3380 126888 3392
rect 125928 3352 126888 3380
rect 125928 3340 125934 3352
rect 126882 3340 126888 3352
rect 126940 3340 126946 3392
rect 130562 3340 130568 3392
rect 130620 3380 130626 3392
rect 131022 3380 131028 3392
rect 130620 3352 131028 3380
rect 130620 3340 130626 3352
rect 131022 3340 131028 3352
rect 131080 3340 131086 3392
rect 132954 3340 132960 3392
rect 133012 3380 133018 3392
rect 133782 3380 133788 3392
rect 133012 3352 133788 3380
rect 133012 3340 133018 3352
rect 133782 3340 133788 3352
rect 133840 3340 133846 3392
rect 134150 3340 134156 3392
rect 134208 3380 134214 3392
rect 135162 3380 135168 3392
rect 134208 3352 135168 3380
rect 134208 3340 134214 3352
rect 135162 3340 135168 3352
rect 135220 3340 135226 3392
rect 135254 3340 135260 3392
rect 135312 3380 135318 3392
rect 136542 3380 136548 3392
rect 135312 3352 136548 3380
rect 135312 3340 135318 3352
rect 136542 3340 136548 3352
rect 136600 3340 136606 3392
rect 138842 3340 138848 3392
rect 138900 3380 138906 3392
rect 139302 3380 139308 3392
rect 138900 3352 139308 3380
rect 138900 3340 138906 3352
rect 139302 3340 139308 3352
rect 139360 3340 139366 3392
rect 141234 3340 141240 3392
rect 141292 3380 141298 3392
rect 142062 3380 142068 3392
rect 141292 3352 142068 3380
rect 141292 3340 141298 3352
rect 142062 3340 142068 3352
rect 142120 3340 142126 3392
rect 142430 3340 142436 3392
rect 142488 3380 142494 3392
rect 143442 3380 143448 3392
rect 142488 3352 143448 3380
rect 142488 3340 142494 3352
rect 143442 3340 143448 3352
rect 143500 3340 143506 3392
rect 144730 3340 144736 3392
rect 144788 3380 144794 3392
rect 145558 3380 145564 3392
rect 144788 3352 145564 3380
rect 144788 3340 144794 3352
rect 145558 3340 145564 3352
rect 145616 3340 145622 3392
rect 147122 3340 147128 3392
rect 147180 3380 147186 3392
rect 147582 3380 147588 3392
rect 147180 3352 147588 3380
rect 147180 3340 147186 3352
rect 147582 3340 147588 3352
rect 147640 3340 147646 3392
rect 148318 3340 148324 3392
rect 148376 3380 148382 3392
rect 148962 3380 148968 3392
rect 148376 3352 148968 3380
rect 148376 3340 148382 3352
rect 148962 3340 148968 3352
rect 149020 3340 149026 3392
rect 149514 3340 149520 3392
rect 149572 3380 149578 3392
rect 150342 3380 150348 3392
rect 149572 3352 150348 3380
rect 149572 3340 149578 3352
rect 150342 3340 150348 3352
rect 150400 3340 150406 3392
rect 223850 3380 223856 3392
rect 150452 3352 223856 3380
rect 101398 3312 101404 3324
rect 98656 3284 101404 3312
rect 101398 3272 101404 3284
rect 101456 3272 101462 3324
rect 136450 3272 136456 3324
rect 136508 3312 136514 3324
rect 137278 3312 137284 3324
rect 136508 3284 137284 3312
rect 136508 3272 136514 3284
rect 137278 3272 137284 3284
rect 137336 3272 137342 3324
rect 140038 3272 140044 3324
rect 140096 3312 140102 3324
rect 150452 3312 150480 3352
rect 223850 3340 223856 3352
rect 223908 3340 223914 3392
rect 229066 3380 229094 3420
rect 232222 3408 232228 3460
rect 232280 3448 232286 3460
rect 233142 3448 233148 3460
rect 232280 3420 233148 3448
rect 232280 3408 232286 3420
rect 233142 3408 233148 3420
rect 233200 3408 233206 3460
rect 242710 3408 242716 3460
rect 242768 3448 242774 3460
rect 246390 3448 246396 3460
rect 242768 3420 246396 3448
rect 242768 3408 242774 3420
rect 246390 3408 246396 3420
rect 246448 3408 246454 3460
rect 250714 3408 250720 3460
rect 250772 3448 250778 3460
rect 294874 3448 294880 3460
rect 250772 3420 294880 3448
rect 250772 3408 250778 3420
rect 294874 3408 294880 3420
rect 294932 3408 294938 3460
rect 298922 3408 298928 3460
rect 298980 3448 298986 3460
rect 302436 3448 302464 3488
rect 580092 3448 580120 3488
rect 580258 3476 580264 3528
rect 580316 3516 580322 3528
rect 582190 3516 582196 3528
rect 580316 3488 582196 3516
rect 580316 3476 580322 3488
rect 582190 3476 582196 3488
rect 582248 3476 582254 3528
rect 580994 3448 581000 3460
rect 298980 3420 302464 3448
rect 306346 3420 567194 3448
rect 580092 3420 581000 3448
rect 298980 3408 298986 3420
rect 234890 3380 234896 3392
rect 229066 3352 234896 3380
rect 234890 3340 234896 3352
rect 234948 3340 234954 3392
rect 242802 3340 242808 3392
rect 242860 3380 242866 3392
rect 247586 3380 247592 3392
rect 242860 3352 247592 3380
rect 242860 3340 242866 3352
rect 247586 3340 247592 3352
rect 247644 3340 247650 3392
rect 257338 3340 257344 3392
rect 257396 3380 257402 3392
rect 270034 3380 270040 3392
rect 257396 3352 270040 3380
rect 257396 3340 257402 3352
rect 270034 3340 270040 3352
rect 270092 3340 270098 3392
rect 271046 3340 271052 3392
rect 271104 3380 271110 3392
rect 272426 3380 272432 3392
rect 271104 3352 272432 3380
rect 271104 3340 271110 3352
rect 272426 3340 272432 3352
rect 272484 3340 272490 3392
rect 296070 3340 296076 3392
rect 296128 3380 296134 3392
rect 299750 3380 299756 3392
rect 296128 3352 299756 3380
rect 296128 3340 296134 3352
rect 299750 3340 299756 3352
rect 299808 3340 299814 3392
rect 140096 3284 150480 3312
rect 140096 3272 140102 3284
rect 150618 3272 150624 3324
rect 150676 3312 150682 3324
rect 225322 3312 225328 3324
rect 150676 3284 225328 3312
rect 150676 3272 150682 3284
rect 225322 3272 225328 3284
rect 225380 3272 225386 3324
rect 233418 3272 233424 3324
rect 233476 3312 233482 3324
rect 239122 3312 239128 3324
rect 233476 3284 239128 3312
rect 233476 3272 233482 3284
rect 239122 3272 239128 3284
rect 239180 3272 239186 3324
rect 239306 3272 239312 3324
rect 239364 3312 239370 3324
rect 240318 3312 240324 3324
rect 239364 3284 240324 3312
rect 239364 3272 239370 3284
rect 240318 3272 240324 3284
rect 240376 3272 240382 3324
rect 253290 3272 253296 3324
rect 253348 3312 253354 3324
rect 260650 3312 260656 3324
rect 253348 3284 260656 3312
rect 253348 3272 253354 3284
rect 260650 3272 260656 3284
rect 260708 3272 260714 3324
rect 264330 3272 264336 3324
rect 264388 3312 264394 3324
rect 273622 3312 273628 3324
rect 264388 3284 273628 3312
rect 264388 3272 264394 3284
rect 273622 3272 273628 3284
rect 273680 3272 273686 3324
rect 80882 3204 80888 3256
rect 80940 3244 80946 3256
rect 81342 3244 81348 3256
rect 80940 3216 81348 3244
rect 80940 3204 80946 3216
rect 81342 3204 81348 3216
rect 81400 3204 81406 3256
rect 83274 3204 83280 3256
rect 83332 3244 83338 3256
rect 84102 3244 84108 3256
rect 83332 3216 84108 3244
rect 83332 3204 83338 3216
rect 84102 3204 84108 3216
rect 84160 3204 84166 3256
rect 84470 3204 84476 3256
rect 84528 3244 84534 3256
rect 87598 3244 87604 3256
rect 84528 3216 87604 3244
rect 84528 3204 84534 3216
rect 87598 3204 87604 3216
rect 87656 3204 87662 3256
rect 89162 3204 89168 3256
rect 89220 3244 89226 3256
rect 90358 3244 90364 3256
rect 89220 3216 90364 3244
rect 89220 3204 89226 3216
rect 90358 3204 90364 3216
rect 90416 3204 90422 3256
rect 91554 3204 91560 3256
rect 91612 3244 91618 3256
rect 92382 3244 92388 3256
rect 91612 3216 92388 3244
rect 91612 3204 91618 3216
rect 92382 3204 92388 3216
rect 92440 3204 92446 3256
rect 92750 3204 92756 3256
rect 92808 3244 92814 3256
rect 111058 3244 111064 3256
rect 92808 3216 111064 3244
rect 92808 3204 92814 3216
rect 111058 3204 111064 3216
rect 111116 3204 111122 3256
rect 115198 3204 115204 3256
rect 115256 3244 115262 3256
rect 116578 3244 116584 3256
rect 115256 3216 116584 3244
rect 115256 3204 115262 3216
rect 116578 3204 116584 3216
rect 116636 3204 116642 3256
rect 143534 3204 143540 3256
rect 143592 3244 143598 3256
rect 144822 3244 144828 3256
rect 143592 3216 144828 3244
rect 143592 3204 143598 3216
rect 144822 3204 144828 3216
rect 144880 3204 144886 3256
rect 154206 3204 154212 3256
rect 154264 3244 154270 3256
rect 155310 3244 155316 3256
rect 154264 3216 155316 3244
rect 154264 3204 154270 3216
rect 155310 3204 155316 3216
rect 155368 3204 155374 3256
rect 155402 3204 155408 3256
rect 155460 3244 155466 3256
rect 156598 3244 156604 3256
rect 155460 3216 156604 3244
rect 155460 3204 155466 3216
rect 156598 3204 156604 3216
rect 156656 3204 156662 3256
rect 158898 3204 158904 3256
rect 158956 3244 158962 3256
rect 160002 3244 160008 3256
rect 158956 3216 160008 3244
rect 158956 3204 158962 3216
rect 160002 3204 160008 3216
rect 160060 3204 160066 3256
rect 160094 3204 160100 3256
rect 160152 3244 160158 3256
rect 161198 3244 161204 3256
rect 160152 3216 161204 3244
rect 160152 3204 160158 3216
rect 161198 3204 161204 3216
rect 161256 3204 161262 3256
rect 163682 3204 163688 3256
rect 163740 3244 163746 3256
rect 164142 3244 164148 3256
rect 163740 3216 164148 3244
rect 163740 3204 163746 3216
rect 164142 3204 164148 3216
rect 164200 3204 164206 3256
rect 164878 3204 164884 3256
rect 164936 3244 164942 3256
rect 165522 3244 165528 3256
rect 164936 3216 165528 3244
rect 164936 3204 164942 3216
rect 165522 3204 165528 3216
rect 165580 3204 165586 3256
rect 166074 3204 166080 3256
rect 166132 3244 166138 3256
rect 166902 3244 166908 3256
rect 166132 3216 166908 3244
rect 166132 3204 166138 3216
rect 166902 3204 166908 3216
rect 166960 3204 166966 3256
rect 167178 3204 167184 3256
rect 167236 3244 167242 3256
rect 169018 3244 169024 3256
rect 167236 3216 169024 3244
rect 167236 3204 167242 3216
rect 169018 3204 169024 3216
rect 169076 3204 169082 3256
rect 173158 3204 173164 3256
rect 173216 3244 173222 3256
rect 173802 3244 173808 3256
rect 173216 3216 173808 3244
rect 173216 3204 173222 3216
rect 173802 3204 173808 3216
rect 173860 3204 173866 3256
rect 174262 3204 174268 3256
rect 174320 3244 174326 3256
rect 175182 3244 175188 3256
rect 174320 3216 175188 3244
rect 174320 3204 174326 3216
rect 175182 3204 175188 3216
rect 175240 3204 175246 3256
rect 175458 3204 175464 3256
rect 175516 3244 175522 3256
rect 176562 3244 176568 3256
rect 175516 3216 176568 3244
rect 175516 3204 175522 3216
rect 176562 3204 176568 3216
rect 176620 3204 176626 3256
rect 176654 3204 176660 3256
rect 176712 3244 176718 3256
rect 177942 3244 177948 3256
rect 176712 3216 177948 3244
rect 176712 3204 176718 3216
rect 177942 3204 177948 3216
rect 178000 3204 178006 3256
rect 180242 3204 180248 3256
rect 180300 3244 180306 3256
rect 180702 3244 180708 3256
rect 180300 3216 180708 3244
rect 180300 3204 180306 3216
rect 180702 3204 180708 3216
rect 180760 3204 180766 3256
rect 181438 3204 181444 3256
rect 181496 3244 181502 3256
rect 182082 3244 182088 3256
rect 181496 3216 182088 3244
rect 181496 3204 181502 3216
rect 182082 3204 182088 3216
rect 182140 3204 182146 3256
rect 182542 3204 182548 3256
rect 182600 3244 182606 3256
rect 183462 3244 183468 3256
rect 182600 3216 183468 3244
rect 182600 3204 182606 3216
rect 183462 3204 183468 3216
rect 183520 3204 183526 3256
rect 183738 3204 183744 3256
rect 183796 3244 183802 3256
rect 184842 3244 184848 3256
rect 183796 3216 184848 3244
rect 183796 3204 183802 3216
rect 184842 3204 184848 3216
rect 184900 3204 184906 3256
rect 186130 3204 186136 3256
rect 186188 3244 186194 3256
rect 186958 3244 186964 3256
rect 186188 3216 186964 3244
rect 186188 3204 186194 3216
rect 186958 3204 186964 3216
rect 187016 3204 187022 3256
rect 189718 3204 189724 3256
rect 189776 3244 189782 3256
rect 191098 3244 191104 3256
rect 189776 3216 191104 3244
rect 189776 3204 189782 3216
rect 191098 3204 191104 3216
rect 191156 3204 191162 3256
rect 193122 3204 193128 3256
rect 193180 3244 193186 3256
rect 200758 3244 200764 3256
rect 193180 3216 200764 3244
rect 193180 3204 193186 3216
rect 200758 3204 200764 3216
rect 200816 3204 200822 3256
rect 299290 3204 299296 3256
rect 299348 3244 299354 3256
rect 306346 3244 306374 3420
rect 307018 3340 307024 3392
rect 307076 3380 307082 3392
rect 309042 3380 309048 3392
rect 307076 3352 309048 3380
rect 307076 3340 307082 3352
rect 309042 3340 309048 3352
rect 309100 3340 309106 3392
rect 313918 3340 313924 3392
rect 313976 3380 313982 3392
rect 315022 3380 315028 3392
rect 313976 3352 315028 3380
rect 313976 3340 313982 3352
rect 315022 3340 315028 3352
rect 315080 3340 315086 3392
rect 316034 3340 316040 3392
rect 316092 3380 316098 3392
rect 317322 3380 317328 3392
rect 316092 3352 317328 3380
rect 316092 3340 316098 3352
rect 317322 3340 317328 3352
rect 317380 3340 317386 3392
rect 318150 3340 318156 3392
rect 318208 3380 318214 3392
rect 319714 3380 319720 3392
rect 318208 3352 319720 3380
rect 318208 3340 318214 3352
rect 319714 3340 319720 3352
rect 319772 3340 319778 3392
rect 323578 3340 323584 3392
rect 323636 3380 323642 3392
rect 325602 3380 325608 3392
rect 323636 3352 325608 3380
rect 323636 3340 323642 3352
rect 325602 3340 325608 3352
rect 325660 3340 325666 3392
rect 331858 3340 331864 3392
rect 331916 3380 331922 3392
rect 332686 3380 332692 3392
rect 331916 3352 332692 3380
rect 331916 3340 331922 3352
rect 332686 3340 332692 3352
rect 332744 3340 332750 3392
rect 335998 3340 336004 3392
rect 336056 3380 336062 3392
rect 337470 3380 337476 3392
rect 336056 3352 337476 3380
rect 336056 3340 336062 3352
rect 337470 3340 337476 3352
rect 337528 3340 337534 3392
rect 342990 3340 342996 3392
rect 343048 3380 343054 3392
rect 344554 3380 344560 3392
rect 343048 3352 344560 3380
rect 343048 3340 343054 3352
rect 344554 3340 344560 3352
rect 344612 3340 344618 3392
rect 345658 3340 345664 3392
rect 345716 3380 345722 3392
rect 348050 3380 348056 3392
rect 345716 3352 348056 3380
rect 345716 3340 345722 3352
rect 348050 3340 348056 3352
rect 348108 3340 348114 3392
rect 348418 3340 348424 3392
rect 348476 3380 348482 3392
rect 351638 3380 351644 3392
rect 348476 3352 351644 3380
rect 348476 3340 348482 3352
rect 351638 3340 351644 3352
rect 351696 3340 351702 3392
rect 364978 3340 364984 3392
rect 365036 3380 365042 3392
rect 367002 3380 367008 3392
rect 365036 3352 367008 3380
rect 365036 3340 365042 3352
rect 367002 3340 367008 3352
rect 367060 3340 367066 3392
rect 367830 3340 367836 3392
rect 367888 3380 367894 3392
rect 369394 3380 369400 3392
rect 367888 3352 369400 3380
rect 367888 3340 367894 3352
rect 369394 3340 369400 3352
rect 369452 3340 369458 3392
rect 382274 3340 382280 3392
rect 382332 3380 382338 3392
rect 383562 3380 383568 3392
rect 382332 3352 383568 3380
rect 382332 3340 382338 3352
rect 383562 3340 383568 3352
rect 383620 3340 383626 3392
rect 389818 3340 389824 3392
rect 389876 3380 389882 3392
rect 390646 3380 390652 3392
rect 389876 3352 390652 3380
rect 389876 3340 389882 3352
rect 390646 3340 390652 3352
rect 390704 3340 390710 3392
rect 398834 3340 398840 3392
rect 398892 3380 398898 3392
rect 400122 3380 400128 3392
rect 398892 3352 400128 3380
rect 398892 3340 398898 3352
rect 400122 3340 400128 3352
rect 400180 3340 400186 3392
rect 432598 3340 432604 3392
rect 432656 3380 432662 3392
rect 434438 3380 434444 3392
rect 432656 3352 434444 3380
rect 432656 3340 432662 3352
rect 434438 3340 434444 3352
rect 434496 3340 434502 3392
rect 435358 3340 435364 3392
rect 435416 3380 435422 3392
rect 437934 3380 437940 3392
rect 435416 3352 437940 3380
rect 435416 3340 435422 3352
rect 437934 3340 437940 3352
rect 437992 3340 437998 3392
rect 439498 3340 439504 3392
rect 439556 3380 439562 3392
rect 441522 3380 441528 3392
rect 439556 3352 441528 3380
rect 439556 3340 439562 3352
rect 441522 3340 441528 3352
rect 441580 3340 441586 3392
rect 454770 3340 454776 3392
rect 454828 3380 454834 3392
rect 455690 3380 455696 3392
rect 454828 3352 455696 3380
rect 454828 3340 454834 3352
rect 455690 3340 455696 3352
rect 455748 3340 455754 3392
rect 457438 3340 457444 3392
rect 457496 3380 457502 3392
rect 459186 3380 459192 3392
rect 457496 3352 459192 3380
rect 457496 3340 457502 3352
rect 459186 3340 459192 3352
rect 459244 3340 459250 3392
rect 490558 3340 490564 3392
rect 490616 3380 490622 3392
rect 492306 3380 492312 3392
rect 490616 3352 492312 3380
rect 490616 3340 490622 3352
rect 492306 3340 492312 3352
rect 492364 3340 492370 3392
rect 497458 3340 497464 3392
rect 497516 3380 497522 3392
rect 499390 3380 499396 3392
rect 497516 3352 499396 3380
rect 497516 3340 497522 3352
rect 499390 3340 499396 3352
rect 499448 3340 499454 3392
rect 502978 3340 502984 3392
rect 503036 3380 503042 3392
rect 505370 3380 505376 3392
rect 503036 3352 505376 3380
rect 503036 3340 503042 3352
rect 505370 3340 505376 3352
rect 505428 3340 505434 3392
rect 515398 3340 515404 3392
rect 515456 3380 515462 3392
rect 517146 3380 517152 3392
rect 515456 3352 517152 3380
rect 515456 3340 515462 3352
rect 517146 3340 517152 3352
rect 517204 3340 517210 3392
rect 522298 3340 522304 3392
rect 522356 3380 522362 3392
rect 524230 3380 524236 3392
rect 522356 3352 524236 3380
rect 522356 3340 522362 3352
rect 524230 3340 524236 3352
rect 524288 3340 524294 3392
rect 530578 3340 530584 3392
rect 530636 3380 530642 3392
rect 532510 3380 532516 3392
rect 530636 3352 532516 3380
rect 530636 3340 530642 3352
rect 532510 3340 532516 3352
rect 532568 3340 532574 3392
rect 540238 3340 540244 3392
rect 540296 3380 540302 3392
rect 541986 3380 541992 3392
rect 540296 3352 541992 3380
rect 540296 3340 540302 3352
rect 541986 3340 541992 3352
rect 542044 3340 542050 3392
rect 567166 3380 567194 3420
rect 580994 3408 581000 3420
rect 581052 3408 581058 3460
rect 583386 3380 583392 3392
rect 567166 3352 583392 3380
rect 583386 3340 583392 3352
rect 583444 3340 583450 3392
rect 347038 3272 347044 3324
rect 347096 3312 347102 3324
rect 350442 3312 350448 3324
rect 347096 3284 350448 3312
rect 347096 3272 347102 3284
rect 350442 3272 350448 3284
rect 350500 3272 350506 3324
rect 421558 3272 421564 3324
rect 421616 3312 421622 3324
rect 423766 3312 423772 3324
rect 421616 3284 423772 3312
rect 421616 3272 421622 3284
rect 423766 3272 423772 3284
rect 423824 3272 423830 3324
rect 431218 3272 431224 3324
rect 431276 3312 431282 3324
rect 433242 3312 433248 3324
rect 431276 3284 433248 3312
rect 431276 3272 431282 3284
rect 433242 3272 433248 3284
rect 433300 3272 433306 3324
rect 453390 3272 453396 3324
rect 453448 3312 453454 3324
rect 456886 3312 456892 3324
rect 453448 3284 456892 3312
rect 453448 3272 453454 3284
rect 456886 3272 456892 3284
rect 456944 3272 456950 3324
rect 529106 3272 529112 3324
rect 529164 3312 529170 3324
rect 534902 3312 534908 3324
rect 529164 3284 534908 3312
rect 529164 3272 529170 3284
rect 534902 3272 534908 3284
rect 534960 3272 534966 3324
rect 548518 3272 548524 3324
rect 548576 3312 548582 3324
rect 550266 3312 550272 3324
rect 548576 3284 550272 3312
rect 548576 3272 548582 3284
rect 550266 3272 550272 3284
rect 550324 3272 550330 3324
rect 299348 3216 306374 3244
rect 299348 3204 299354 3216
rect 382918 3204 382924 3256
rect 382976 3244 382982 3256
rect 384758 3244 384764 3256
rect 382976 3216 384764 3244
rect 382976 3204 382982 3216
rect 384758 3204 384764 3216
rect 384816 3204 384822 3256
rect 500310 3204 500316 3256
rect 500368 3244 500374 3256
rect 502978 3244 502984 3256
rect 500368 3216 502984 3244
rect 500368 3204 500374 3216
rect 502978 3204 502984 3216
rect 503036 3204 503042 3256
rect 556798 3204 556804 3256
rect 556856 3244 556862 3256
rect 559742 3244 559748 3256
rect 556856 3216 559748 3244
rect 556856 3204 556862 3216
rect 559742 3204 559748 3216
rect 559800 3204 559806 3256
rect 82078 3136 82084 3188
rect 82136 3176 82142 3188
rect 87414 3176 87420 3188
rect 82136 3148 87420 3176
rect 82136 3136 82142 3148
rect 87414 3136 87420 3148
rect 87472 3136 87478 3188
rect 98638 3136 98644 3188
rect 98696 3176 98702 3188
rect 99282 3176 99288 3188
rect 98696 3148 99288 3176
rect 98696 3136 98702 3148
rect 99282 3136 99288 3148
rect 99340 3136 99346 3188
rect 151814 3136 151820 3188
rect 151872 3176 151878 3188
rect 153102 3176 153108 3188
rect 151872 3148 153108 3176
rect 151872 3136 151878 3148
rect 153102 3136 153108 3148
rect 153160 3136 153166 3188
rect 157794 3136 157800 3188
rect 157852 3176 157858 3188
rect 159358 3176 159364 3188
rect 157852 3148 159364 3176
rect 157852 3136 157858 3148
rect 159358 3136 159364 3148
rect 159416 3136 159422 3188
rect 169570 3136 169576 3188
rect 169628 3176 169634 3188
rect 170398 3176 170404 3188
rect 169628 3148 170404 3176
rect 169628 3136 169634 3148
rect 170398 3136 170404 3148
rect 170456 3136 170462 3188
rect 231026 3136 231032 3188
rect 231084 3176 231090 3188
rect 238018 3176 238024 3188
rect 231084 3148 238024 3176
rect 231084 3136 231090 3148
rect 238018 3136 238024 3148
rect 238076 3136 238082 3188
rect 385678 3136 385684 3188
rect 385736 3176 385742 3188
rect 387150 3176 387156 3188
rect 385736 3148 387156 3176
rect 385736 3136 385742 3148
rect 387150 3136 387156 3148
rect 387208 3136 387214 3188
rect 413278 3136 413284 3188
rect 413336 3176 413342 3188
rect 416682 3176 416688 3188
rect 413336 3148 416688 3176
rect 413336 3136 413342 3148
rect 416682 3136 416688 3148
rect 416740 3136 416746 3188
rect 78640 3080 78812 3108
rect 78640 3068 78646 3080
rect 85666 3068 85672 3120
rect 85724 3108 85730 3120
rect 86862 3108 86868 3120
rect 85724 3080 86868 3108
rect 85724 3068 85730 3080
rect 86862 3068 86868 3080
rect 86920 3068 86926 3120
rect 90358 3068 90364 3120
rect 90416 3108 90422 3120
rect 93118 3108 93124 3120
rect 90416 3080 93124 3108
rect 90416 3068 90422 3080
rect 93118 3068 93124 3080
rect 93176 3068 93182 3120
rect 156598 3068 156604 3120
rect 156656 3108 156662 3120
rect 157978 3108 157984 3120
rect 156656 3080 157984 3108
rect 156656 3068 156662 3080
rect 157978 3068 157984 3080
rect 158036 3068 158042 3120
rect 168374 3068 168380 3120
rect 168432 3108 168438 3120
rect 169662 3108 169668 3120
rect 168432 3080 169668 3108
rect 168432 3068 168438 3080
rect 169662 3068 169668 3080
rect 169720 3068 169726 3120
rect 171962 3068 171968 3120
rect 172020 3108 172026 3120
rect 173066 3108 173072 3120
rect 172020 3080 173072 3108
rect 172020 3068 172026 3080
rect 173066 3068 173072 3080
rect 173124 3068 173130 3120
rect 324958 3068 324964 3120
rect 325016 3108 325022 3120
rect 326798 3108 326804 3120
rect 325016 3080 326804 3108
rect 325016 3068 325022 3080
rect 326798 3068 326804 3080
rect 326856 3068 326862 3120
rect 360838 3068 360844 3120
rect 360896 3108 360902 3120
rect 362310 3108 362316 3120
rect 360896 3080 362316 3108
rect 360896 3068 360902 3080
rect 362310 3068 362316 3080
rect 362368 3068 362374 3120
rect 237006 3000 237012 3052
rect 237064 3040 237070 3052
rect 241054 3040 241060 3052
rect 237064 3012 241060 3040
rect 237064 3000 237070 3012
rect 241054 3000 241060 3012
rect 241112 3000 241118 3052
rect 264146 3000 264152 3052
rect 264204 3040 264210 3052
rect 267826 3040 267832 3052
rect 264204 3012 267832 3040
rect 264204 3000 264210 3012
rect 267826 3000 267832 3012
rect 267884 3000 267890 3052
rect 511258 3000 511264 3052
rect 511316 3040 511322 3052
rect 513558 3040 513564 3052
rect 511316 3012 513564 3040
rect 511316 3000 511322 3012
rect 513558 3000 513564 3012
rect 513616 3000 513622 3052
rect 30098 2932 30104 2984
rect 30156 2972 30162 2984
rect 36538 2972 36544 2984
rect 30156 2944 36544 2972
rect 30156 2932 30162 2944
rect 36538 2932 36544 2944
rect 36596 2932 36602 2984
rect 126974 2932 126980 2984
rect 127032 2972 127038 2984
rect 128262 2972 128268 2984
rect 127032 2944 128268 2972
rect 127032 2932 127038 2944
rect 128262 2932 128268 2944
rect 128320 2932 128326 2984
rect 446398 2932 446404 2984
rect 446456 2972 446462 2984
rect 452102 2972 452108 2984
rect 446456 2944 452108 2972
rect 446456 2932 446462 2944
rect 452102 2932 452108 2944
rect 452160 2932 452166 2984
rect 464338 2932 464344 2984
rect 464396 2972 464402 2984
rect 466270 2972 466276 2984
rect 464396 2944 466276 2972
rect 464396 2932 464402 2944
rect 466270 2932 466276 2944
rect 466328 2932 466334 2984
rect 493318 2932 493324 2984
rect 493376 2972 493382 2984
rect 495894 2972 495900 2984
rect 493376 2944 495900 2972
rect 493376 2932 493382 2944
rect 495894 2932 495900 2944
rect 495952 2932 495958 2984
rect 504358 2932 504364 2984
rect 504416 2972 504422 2984
rect 510062 2972 510068 2984
rect 504416 2944 510068 2972
rect 504416 2932 504422 2944
rect 510062 2932 510068 2944
rect 510120 2932 510126 2984
rect 542998 2932 543004 2984
rect 543056 2972 543062 2984
rect 545482 2972 545488 2984
rect 543056 2944 545488 2972
rect 543056 2932 543062 2944
rect 545482 2932 545488 2944
rect 545540 2932 545546 2984
rect 70302 2864 70308 2916
rect 70360 2904 70366 2916
rect 76558 2904 76564 2916
rect 70360 2876 76564 2904
rect 70360 2864 70366 2876
rect 76558 2864 76564 2876
rect 76616 2864 76622 2916
rect 118786 2864 118792 2916
rect 118844 2904 118850 2916
rect 119982 2904 119988 2916
rect 118844 2876 119988 2904
rect 118844 2864 118850 2876
rect 119982 2864 119988 2876
rect 120040 2864 120046 2916
rect 184934 2864 184940 2916
rect 184992 2904 184998 2916
rect 188338 2904 188344 2916
rect 184992 2876 188344 2904
rect 184992 2864 184998 2876
rect 188338 2864 188344 2876
rect 188396 2864 188402 2916
rect 242526 2864 242532 2916
rect 242584 2904 242590 2916
rect 244090 2904 244096 2916
rect 242584 2876 244096 2904
rect 242584 2864 242590 2876
rect 244090 2864 244096 2876
rect 244148 2864 244154 2916
rect 369118 2864 369124 2916
rect 369176 2904 369182 2916
rect 371694 2904 371700 2916
rect 369176 2876 371700 2904
rect 369176 2864 369182 2876
rect 371694 2864 371700 2876
rect 371752 2864 371758 2916
rect 417510 2864 417516 2916
rect 417568 2904 417574 2916
rect 420178 2904 420184 2916
rect 417568 2876 420184 2904
rect 417568 2864 417574 2876
rect 420178 2864 420184 2876
rect 420236 2864 420242 2916
rect 525150 2864 525156 2916
rect 525208 2904 525214 2916
rect 527818 2904 527824 2916
rect 525208 2876 527824 2904
rect 525208 2864 525214 2876
rect 527818 2864 527824 2876
rect 527876 2864 527882 2916
<< via1 >>
rect 218980 700952 219032 701004
rect 252560 700952 252612 701004
rect 249616 700884 249668 700936
rect 348792 700884 348844 700936
rect 154120 700816 154172 700868
rect 255320 700816 255372 700868
rect 137836 700748 137888 700800
rect 255412 700748 255464 700800
rect 246948 700680 247000 700732
rect 413652 700680 413704 700732
rect 89168 700612 89220 700664
rect 258080 700612 258132 700664
rect 72976 700544 73028 700596
rect 258172 700544 258224 700596
rect 40500 700476 40552 700528
rect 41328 700476 41380 700528
rect 244188 700476 244240 700528
rect 478512 700476 478564 700528
rect 24308 700408 24360 700460
rect 260840 700408 260892 700460
rect 8116 700340 8168 700392
rect 259460 700340 259512 700392
rect 284944 700340 284996 700392
rect 332508 700340 332560 700392
rect 241428 700272 241480 700324
rect 543464 700272 543516 700324
rect 252468 700204 252520 700256
rect 283840 700204 283892 700256
rect 251088 700136 251140 700188
rect 267648 700136 267700 700188
rect 105452 699660 105504 699712
rect 106188 699660 106240 699712
rect 170312 699660 170364 699712
rect 171048 699660 171100 699712
rect 235172 699660 235224 699712
rect 240784 699660 240836 699712
rect 298744 699660 298796 699712
rect 300124 699660 300176 699712
rect 359464 699660 359516 699712
rect 364984 699660 365036 699712
rect 396724 699660 396776 699712
rect 397460 699660 397512 699712
rect 461584 699660 461636 699712
rect 462320 699660 462372 699712
rect 526444 699660 526496 699712
rect 527180 699660 527232 699712
rect 238668 696940 238720 696992
rect 580172 696940 580224 696992
rect 3424 683204 3476 683256
rect 262220 683204 262272 683256
rect 238576 683136 238628 683188
rect 580172 683136 580224 683188
rect 3424 670760 3476 670812
rect 263600 670760 263652 670812
rect 237288 670692 237340 670744
rect 580172 670692 580224 670744
rect 3424 656888 3476 656940
rect 262312 656888 262364 656940
rect 235908 643084 235960 643136
rect 580172 643084 580224 643136
rect 3424 632068 3476 632120
rect 264980 632068 265032 632120
rect 235816 630640 235868 630692
rect 580172 630640 580224 630692
rect 3148 618264 3200 618316
rect 266360 618264 266412 618316
rect 234528 616836 234580 616888
rect 580172 616836 580224 616888
rect 3240 605820 3292 605872
rect 265072 605820 265124 605872
rect 233148 590656 233200 590708
rect 579804 590656 579856 590708
rect 3332 579640 3384 579692
rect 266452 579640 266504 579692
rect 233056 576852 233108 576904
rect 580172 576852 580224 576904
rect 3424 565836 3476 565888
rect 269120 565836 269172 565888
rect 231768 563048 231820 563100
rect 579804 563048 579856 563100
rect 3424 553392 3476 553444
rect 267740 553392 267792 553444
rect 230388 536800 230440 536852
rect 580172 536800 580224 536852
rect 3424 527144 3476 527196
rect 269212 527144 269264 527196
rect 231676 524424 231728 524476
rect 580172 524424 580224 524476
rect 3424 514768 3476 514820
rect 271880 514768 271932 514820
rect 229008 510620 229060 510672
rect 580172 510620 580224 510672
rect 3056 500964 3108 501016
rect 270500 500964 270552 501016
rect 227628 484372 227680 484424
rect 580172 484372 580224 484424
rect 3424 474716 3476 474768
rect 271972 474716 272024 474768
rect 228916 470568 228968 470620
rect 579988 470568 580040 470620
rect 3240 462340 3292 462392
rect 273260 462340 273312 462392
rect 226248 456764 226300 456816
rect 580172 456764 580224 456816
rect 3148 448536 3200 448588
rect 273352 448536 273404 448588
rect 224868 430584 224920 430636
rect 580172 430584 580224 430636
rect 3424 422288 3476 422340
rect 274640 422288 274692 422340
rect 226156 418140 226208 418192
rect 580172 418140 580224 418192
rect 3148 409844 3200 409896
rect 276020 409844 276072 409896
rect 224776 404336 224828 404388
rect 580172 404336 580224 404388
rect 3424 397468 3476 397520
rect 276112 397468 276164 397520
rect 222016 378156 222068 378208
rect 580172 378156 580224 378208
rect 3424 371220 3476 371272
rect 277400 371220 277452 371272
rect 371608 368568 371660 368620
rect 376760 368568 376812 368620
rect 371700 368500 371752 368552
rect 381084 368500 381136 368552
rect 445208 368500 445260 368552
rect 452844 368500 452896 368552
rect 371608 367480 371660 367532
rect 374000 367480 374052 367532
rect 445668 367208 445720 367260
rect 452660 367208 452712 367260
rect 371516 367072 371568 367124
rect 380992 367072 381044 367124
rect 371608 365848 371660 365900
rect 378232 365848 378284 365900
rect 371240 365780 371292 365832
rect 375380 365780 375432 365832
rect 444932 365712 444984 365764
rect 448612 365712 448664 365764
rect 371240 364692 371292 364744
rect 374460 364692 374512 364744
rect 444932 364624 444984 364676
rect 449992 364624 450044 364676
rect 371608 364352 371660 364404
rect 378324 364352 378376 364404
rect 371608 363672 371660 363724
rect 375748 363672 375800 363724
rect 444564 363128 444616 363180
rect 447416 363128 447468 363180
rect 371424 362992 371476 363044
rect 377036 362992 377088 363044
rect 371700 362924 371752 362976
rect 378416 362924 378468 362976
rect 371424 361564 371476 361616
rect 376852 361564 376904 361616
rect 444932 361564 444984 361616
rect 450084 361564 450136 361616
rect 371608 360408 371660 360460
rect 375564 360408 375616 360460
rect 371700 360340 371752 360392
rect 374276 360340 374328 360392
rect 371516 360204 371568 360256
rect 375472 360204 375524 360256
rect 445668 360204 445720 360256
rect 449900 360204 449952 360256
rect 371884 359456 371936 359508
rect 379520 359456 379572 359508
rect 371332 358776 371384 358828
rect 383660 358776 383712 358828
rect 444472 358776 444524 358828
rect 447232 358776 447284 358828
rect 371424 357688 371476 357740
rect 375656 357688 375708 357740
rect 3148 357416 3200 357468
rect 278780 357416 278832 357468
rect 371516 357416 371568 357468
rect 382464 357416 382516 357468
rect 444932 357416 444984 357468
rect 448888 357416 448940 357468
rect 444564 356736 444616 356788
rect 448704 356736 448756 356788
rect 371332 356192 371384 356244
rect 378140 356192 378192 356244
rect 371240 356124 371292 356176
rect 381176 356124 381228 356176
rect 371424 356056 371476 356108
rect 382280 356056 382332 356108
rect 444380 355104 444432 355156
rect 446036 355104 446088 355156
rect 371240 354968 371292 355020
rect 372896 354968 372948 355020
rect 371700 354764 371752 354816
rect 376944 354764 376996 354816
rect 371516 354152 371568 354204
rect 374184 354152 374236 354204
rect 444472 353336 444524 353388
rect 447324 353336 447376 353388
rect 371700 353268 371752 353320
rect 374092 353268 374144 353320
rect 372068 352588 372120 352640
rect 377128 352588 377180 352640
rect 372252 352520 372304 352572
rect 379612 352520 379664 352572
rect 444380 351976 444432 352028
rect 447140 351976 447192 352028
rect 371608 348168 371660 348220
rect 374368 348168 374420 348220
rect 445208 345584 445260 345636
rect 450176 345584 450228 345636
rect 445668 345108 445720 345160
rect 452752 345108 452804 345160
rect 3332 345040 3384 345092
rect 278872 345040 278924 345092
rect 445668 343612 445720 343664
rect 454040 343612 454092 343664
rect 445668 342252 445720 342304
rect 451372 342252 451424 342304
rect 445116 340960 445168 341012
rect 448796 340960 448848 341012
rect 444748 340212 444800 340264
rect 446128 340212 446180 340264
rect 299940 337424 299992 337476
rect 438952 337424 439004 337476
rect 198556 337356 198608 337408
rect 366916 337356 366968 337408
rect 441252 336744 441304 336796
rect 441620 336744 441672 336796
rect 368940 335316 368992 335368
rect 369124 335316 369176 335368
rect 245568 327700 245620 327752
rect 396724 327700 396776 327752
rect 219348 324300 219400 324352
rect 580172 324300 580224 324352
rect 242716 323552 242768 323604
rect 461584 323552 461636 323604
rect 3424 318792 3476 318844
rect 280252 318792 280304 318844
rect 220636 311856 220688 311908
rect 580172 311856 580224 311908
rect 202788 305872 202840 305924
rect 252928 305872 252980 305924
rect 246856 305804 246908 305856
rect 359464 305804 359516 305856
rect 244280 305736 244332 305788
rect 429200 305736 429252 305788
rect 41328 305668 41380 305720
rect 259828 305668 259880 305720
rect 240048 305600 240100 305652
rect 526444 305600 526496 305652
rect 3240 304988 3292 305040
rect 282276 304988 282328 305040
rect 240784 304784 240836 304836
rect 252100 304784 252152 304836
rect 247776 304716 247828 304768
rect 284944 304716 284996 304768
rect 249524 304648 249576 304700
rect 298744 304648 298796 304700
rect 171048 304580 171100 304632
rect 254676 304580 254728 304632
rect 106188 304512 106240 304564
rect 257252 304512 257304 304564
rect 241704 304444 241756 304496
rect 494060 304444 494112 304496
rect 239128 304376 239180 304428
rect 558920 304376 558972 304428
rect 222752 304308 222804 304360
rect 580264 304308 580316 304360
rect 221004 304240 221056 304292
rect 580356 304240 580408 304292
rect 237380 303016 237432 303068
rect 238668 303016 238720 303068
rect 243452 303016 243504 303068
rect 244188 303016 244240 303068
rect 246028 303016 246080 303068
rect 246948 303016 247000 303068
rect 248604 303016 248656 303068
rect 249616 303016 249668 303068
rect 251180 303016 251232 303068
rect 252468 303016 252520 303068
rect 255320 303016 255372 303068
rect 256148 303016 256200 303068
rect 273260 303016 273312 303068
rect 274180 303016 274232 303068
rect 215024 302948 215076 303000
rect 316684 302948 316736 303000
rect 177396 302880 177448 302932
rect 287428 302880 287480 302932
rect 178684 302812 178736 302864
rect 298652 302812 298704 302864
rect 214104 302744 214156 302796
rect 447968 302744 448020 302796
rect 211528 302676 211580 302728
rect 446404 302676 446456 302728
rect 217600 302608 217652 302660
rect 464344 302608 464396 302660
rect 212448 302540 212500 302592
rect 461584 302540 461636 302592
rect 207204 302472 207256 302524
rect 457444 302472 457496 302524
rect 204628 302404 204680 302456
rect 454684 302404 454736 302456
rect 202052 302336 202104 302388
rect 453304 302336 453356 302388
rect 14464 302268 14516 302320
rect 292580 302268 292632 302320
rect 11704 302200 11756 302252
rect 290004 302200 290056 302252
rect 230480 302132 230532 302184
rect 231676 302132 231728 302184
rect 229652 302064 229704 302116
rect 230388 302064 230440 302116
rect 232228 302064 232280 302116
rect 233148 302064 233200 302116
rect 258080 302064 258132 302116
rect 259000 302064 259052 302116
rect 278780 302064 278832 302116
rect 279700 302064 279752 302116
rect 276020 301792 276072 301844
rect 277032 301792 277084 301844
rect 196624 301656 196676 301708
rect 281356 301656 281408 301708
rect 199384 301588 199436 301640
rect 285680 301588 285732 301640
rect 215852 301520 215904 301572
rect 304264 301520 304316 301572
rect 210700 301452 210752 301504
rect 301504 301452 301556 301504
rect 203800 301384 203852 301436
rect 309784 301384 309836 301436
rect 159364 301316 159416 301368
rect 288256 301316 288308 301368
rect 151084 301248 151136 301300
rect 291752 301248 291804 301300
rect 146944 301180 146996 301232
rect 295156 301180 295208 301232
rect 209872 301112 209924 301164
rect 465724 301112 465776 301164
rect 17224 301044 17276 301096
rect 283104 301044 283156 301096
rect 7564 300976 7616 301028
rect 296904 300976 296956 301028
rect 202972 300908 203024 300960
rect 582472 300908 582524 300960
rect 200396 300840 200448 300892
rect 582380 300840 582432 300892
rect 234804 300432 234856 300484
rect 235908 300432 235960 300484
rect 223672 300296 223724 300348
rect 224776 300296 224828 300348
rect 225328 300296 225380 300348
rect 226156 300296 226208 300348
rect 227904 300296 227956 300348
rect 228916 300296 228968 300348
rect 205548 300228 205600 300280
rect 307024 300228 307076 300280
rect 201224 300160 201276 300212
rect 305644 300160 305696 300212
rect 206376 300092 206428 300144
rect 313924 300092 313976 300144
rect 170404 300024 170456 300076
rect 290556 300024 290608 300076
rect 152464 299956 152516 300008
rect 288900 299956 288952 300008
rect 155224 299888 155276 299940
rect 295708 299888 295760 299940
rect 148324 299820 148376 299872
rect 294052 299820 294104 299872
rect 144184 299752 144236 299804
rect 297364 299752 297416 299804
rect 209320 299684 209372 299736
rect 443644 299684 443696 299736
rect 213552 299616 213604 299668
rect 450544 299616 450596 299668
rect 208308 299548 208360 299600
rect 449164 299548 449216 299600
rect 4804 299480 4856 299532
rect 293132 299480 293184 299532
rect 216680 299412 216732 299464
rect 220084 299412 220136 299464
rect 237196 299412 237248 299464
rect 199844 298460 199896 298512
rect 216680 299276 216732 299328
rect 217140 299276 217192 299328
rect 218060 299276 218112 299328
rect 218152 299276 218204 299328
rect 218704 299276 218756 299328
rect 218796 299276 218848 299328
rect 219900 299276 219952 299328
rect 220084 299276 220136 299328
rect 3516 298392 3568 298444
rect 3608 298324 3660 298376
rect 3424 298256 3476 298308
rect 237196 299276 237248 299328
rect 242164 299276 242216 299328
rect 242348 299276 242400 299328
rect 283564 299276 283616 299328
rect 284484 299276 284536 299328
rect 286508 299276 286560 299328
rect 299848 299276 299900 299328
rect 300124 299276 300176 299328
rect 434720 299072 434772 299124
rect 441712 299072 441764 299124
rect 318064 298460 318116 298512
rect 302792 298256 302844 298308
rect 322204 298256 322256 298308
rect 580172 298188 580224 298240
rect 580264 298120 580316 298172
rect 371240 298052 371292 298104
rect 381084 298052 381136 298104
rect 436100 297576 436152 297628
rect 441804 297576 441856 297628
rect 381084 297440 381136 297492
rect 382372 297440 382424 297492
rect 371240 297372 371292 297424
rect 379520 297372 379572 297424
rect 445668 296964 445720 297016
rect 447784 296964 447836 297016
rect 447784 296828 447836 296880
rect 452844 296828 452896 296880
rect 303068 296760 303120 296812
rect 369400 296760 369452 296812
rect 302884 296692 302936 296744
rect 369308 296692 369360 296744
rect 371240 296624 371292 296676
rect 376760 296624 376812 296676
rect 445668 295944 445720 295996
rect 452660 295944 452712 295996
rect 324964 295876 325016 295928
rect 371240 295876 371292 295928
rect 352564 295808 352616 295860
rect 369308 295808 369360 295860
rect 371240 295536 371292 295588
rect 373356 295536 373408 295588
rect 374000 295536 374052 295588
rect 376760 295400 376812 295452
rect 380900 295400 380952 295452
rect 370228 295332 370280 295384
rect 377404 295332 377456 295384
rect 380992 295332 381044 295384
rect 452660 295332 452712 295384
rect 454132 295332 454184 295384
rect 370136 295196 370188 295248
rect 378232 295196 378284 295248
rect 445668 295196 445720 295248
rect 448612 295196 448664 295248
rect 378232 294720 378284 294772
rect 381084 294720 381136 294772
rect 372344 294584 372396 294636
rect 372620 294584 372672 294636
rect 378232 294584 378284 294636
rect 448612 294040 448664 294092
rect 452660 294040 452712 294092
rect 180064 293972 180116 294024
rect 197912 293972 197964 294024
rect 302424 293972 302476 294024
rect 320824 293972 320876 294024
rect 371240 293972 371292 294024
rect 375380 293972 375432 294024
rect 445760 293972 445812 294024
rect 450268 293972 450320 294024
rect 2872 293904 2924 293956
rect 196624 293904 196676 293956
rect 371240 293224 371292 293276
rect 378324 293224 378376 293276
rect 371240 292884 371292 292936
rect 374460 292884 374512 292936
rect 374920 292884 374972 292936
rect 445668 292884 445720 292936
rect 446496 292884 446548 292936
rect 449992 292884 450044 292936
rect 378324 292544 378376 292596
rect 378508 292544 378560 292596
rect 371240 291864 371292 291916
rect 375748 291864 375800 291916
rect 378324 291864 378376 291916
rect 195244 291796 195296 291848
rect 198096 291796 198148 291848
rect 372344 291796 372396 291848
rect 373264 291796 373316 291848
rect 378416 291796 378468 291848
rect 302332 291184 302384 291236
rect 359464 291184 359516 291236
rect 371240 291184 371292 291236
rect 376024 291184 376076 291236
rect 377036 291184 377088 291236
rect 445668 291184 445720 291236
rect 447416 291184 447468 291236
rect 451280 291184 451332 291236
rect 448612 291116 448664 291168
rect 450084 291116 450136 291168
rect 445668 290572 445720 290624
rect 448612 290572 448664 290624
rect 372344 290504 372396 290556
rect 372804 290504 372856 290556
rect 376760 290504 376812 290556
rect 371240 290436 371292 290488
rect 376852 290436 376904 290488
rect 184204 289824 184256 289876
rect 197360 289824 197412 289876
rect 445668 289416 445720 289468
rect 445852 289416 445904 289468
rect 450084 289416 450136 289468
rect 371240 289008 371292 289060
rect 374276 289008 374328 289060
rect 375748 289008 375800 289060
rect 372344 288940 372396 288992
rect 374736 288940 374788 288992
rect 375472 288940 375524 288992
rect 372804 288532 372856 288584
rect 375564 288532 375616 288584
rect 371240 288328 371292 288380
rect 377128 288328 377180 288380
rect 383660 288328 383712 288380
rect 445668 288328 445720 288380
rect 447876 288328 447928 288380
rect 449900 288328 449952 288380
rect 445116 288056 445168 288108
rect 447232 288056 447284 288108
rect 448520 288056 448572 288108
rect 160100 287036 160152 287088
rect 197636 287036 197688 287088
rect 372344 287036 372396 287088
rect 382648 287036 382700 287088
rect 383568 287036 383620 287088
rect 371884 286560 371936 286612
rect 372344 286560 372396 286612
rect 371332 286424 371384 286476
rect 375656 286424 375708 286476
rect 371884 286356 371936 286408
rect 376116 286356 376168 286408
rect 382464 286356 382516 286408
rect 372528 286288 372580 286340
rect 379612 286288 379664 286340
rect 188344 285676 188396 285728
rect 197360 285676 197412 285728
rect 302792 285676 302844 285728
rect 353944 285676 353996 285728
rect 375656 285676 375708 285728
rect 380900 285676 380952 285728
rect 445668 285676 445720 285728
rect 448888 285676 448940 285728
rect 449900 285676 449952 285728
rect 371884 285608 371936 285660
rect 381176 285608 381228 285660
rect 371884 285064 371936 285116
rect 374644 285064 374696 285116
rect 378140 285064 378192 285116
rect 445668 284860 445720 284912
rect 446680 284860 446732 284912
rect 448704 284860 448756 284912
rect 381176 284384 381228 284436
rect 382556 284384 382608 284436
rect 371884 284316 371936 284368
rect 378140 284316 378192 284368
rect 382280 284316 382332 284368
rect 445484 283636 445536 283688
rect 446036 283636 446088 283688
rect 371884 283568 371936 283620
rect 376944 283568 376996 283620
rect 377220 283568 377272 283620
rect 371884 283160 371936 283212
rect 372896 283160 372948 283212
rect 375472 283160 375524 283212
rect 184296 282888 184348 282940
rect 197360 282888 197412 282940
rect 446036 282888 446088 282940
rect 448704 282888 448756 282940
rect 371884 282684 371936 282736
rect 374184 282684 374236 282736
rect 374552 282684 374604 282736
rect 445392 282480 445444 282532
rect 447232 282480 447284 282532
rect 371884 282140 371936 282192
rect 374092 282140 374144 282192
rect 374276 282140 374328 282192
rect 302424 281528 302476 281580
rect 356704 281528 356756 281580
rect 445116 281460 445168 281512
rect 446588 281460 446640 281512
rect 447140 281460 447192 281512
rect 444748 280576 444800 280628
rect 445944 280576 445996 280628
rect 447140 280576 447192 280628
rect 186964 280168 187016 280220
rect 197360 280168 197412 280220
rect 358084 280100 358136 280152
rect 360200 280100 360252 280152
rect 444564 280032 444616 280084
rect 444840 280032 444892 280084
rect 193956 278944 194008 278996
rect 197360 278944 197412 278996
rect 302608 278740 302660 278792
rect 358084 278740 358136 278792
rect 372160 278672 372212 278724
rect 372988 278672 373040 278724
rect 444380 278672 444432 278724
rect 445116 278672 445168 278724
rect 372344 277448 372396 277500
rect 374184 277448 374236 277500
rect 369124 277176 369176 277228
rect 369308 277176 369360 277228
rect 371608 276360 371660 276412
rect 372160 276360 372212 276412
rect 182824 276020 182876 276072
rect 197544 276020 197596 276072
rect 371608 276020 371660 276072
rect 374000 276020 374052 276072
rect 374368 276020 374420 276072
rect 196624 274864 196676 274916
rect 198372 274864 198424 274916
rect 445576 274592 445628 274644
rect 449256 274592 449308 274644
rect 452752 274592 452804 274644
rect 445668 273232 445720 273284
rect 450176 273232 450228 273284
rect 452936 273232 452988 273284
rect 371056 273164 371108 273216
rect 374368 273164 374420 273216
rect 445668 272484 445720 272536
rect 454040 272484 454092 272536
rect 181444 271872 181496 271924
rect 197360 271872 197412 271924
rect 371516 271464 371568 271516
rect 371516 271124 371568 271176
rect 371792 271124 371844 271176
rect 371976 271124 372028 271176
rect 358084 271056 358136 271108
rect 360660 271056 360712 271108
rect 445668 270580 445720 270632
rect 451372 270580 451424 270632
rect 178776 270512 178828 270564
rect 197360 270512 197412 270564
rect 302332 270444 302384 270496
rect 352564 270444 352616 270496
rect 445668 269084 445720 269136
rect 448796 269084 448848 269136
rect 452844 269084 452896 269136
rect 372160 268336 372212 268388
rect 372896 268336 372948 268388
rect 175924 267724 175976 267776
rect 197728 267724 197780 267776
rect 3240 267656 3292 267708
rect 17224 267656 17276 267708
rect 302424 267656 302476 267708
rect 324964 267656 325016 267708
rect 302516 266976 302568 267028
rect 370228 266976 370280 267028
rect 362868 266296 362920 266348
rect 435180 266296 435232 266348
rect 436008 266296 436060 266348
rect 441712 266296 441764 266348
rect 364892 266228 364944 266280
rect 437388 266228 437440 266280
rect 441804 266228 441856 266280
rect 302976 266160 303028 266212
rect 368940 266160 368992 266212
rect 369124 266160 369176 266212
rect 441344 266160 441396 266212
rect 441528 266160 441580 266212
rect 300124 266092 300176 266144
rect 366916 266092 366968 266144
rect 360936 265684 360988 265736
rect 431960 265684 432012 265736
rect 432604 265684 432656 265736
rect 300032 265616 300084 265668
rect 438860 265616 438912 265668
rect 174544 264936 174596 264988
rect 197360 264936 197412 264988
rect 360200 264936 360252 264988
rect 360936 264936 360988 264988
rect 180156 263576 180208 263628
rect 197912 263576 197964 263628
rect 196716 261808 196768 261860
rect 198648 261808 198700 261860
rect 302792 260788 302844 260840
rect 370136 260788 370188 260840
rect 195336 259496 195388 259548
rect 197728 259496 197780 259548
rect 464344 259360 464396 259412
rect 580172 259360 580224 259412
rect 191104 256708 191156 256760
rect 198096 256708 198148 256760
rect 302792 256708 302844 256760
rect 370872 256708 370924 256760
rect 188436 255280 188488 255332
rect 197360 255280 197412 255332
rect 187056 252560 187108 252612
rect 197360 252560 197412 252612
rect 171784 248412 171836 248464
rect 198188 248412 198240 248464
rect 302884 247664 302936 247716
rect 370504 247664 370556 247716
rect 304264 245556 304316 245608
rect 580172 245556 580224 245608
rect 171876 244264 171928 244316
rect 197360 244264 197412 244316
rect 192484 241544 192536 241596
rect 197728 241544 197780 241596
rect 370504 241476 370556 241528
rect 375380 241476 375432 241528
rect 303160 240728 303212 240780
rect 370320 240728 370372 240780
rect 171968 238756 172020 238808
rect 197360 238756 197412 238808
rect 184388 237396 184440 237448
rect 197360 237396 197412 237448
rect 303068 235220 303120 235272
rect 369216 235220 369268 235272
rect 172060 234608 172112 234660
rect 197544 234608 197596 234660
rect 191196 233384 191248 233436
rect 198188 233384 198240 233436
rect 447968 233180 448020 233232
rect 579988 233180 580040 233232
rect 369216 231684 369268 231736
rect 374920 231684 374972 231736
rect 177488 230460 177540 230512
rect 197636 230460 197688 230512
rect 302976 229712 303028 229764
rect 369400 229712 369452 229764
rect 177304 229100 177356 229152
rect 197360 229100 197412 229152
rect 369400 229100 369452 229152
rect 373264 229100 373316 229152
rect 303160 228352 303212 228404
rect 370228 228352 370280 228404
rect 436008 227740 436060 227792
rect 441896 227740 441948 227792
rect 316684 226992 316736 227044
rect 580264 226992 580316 227044
rect 437388 226244 437440 226296
rect 441712 226244 441764 226296
rect 303252 225632 303304 225684
rect 369952 225632 370004 225684
rect 302792 225564 302844 225616
rect 370136 225564 370188 225616
rect 371608 225564 371660 225616
rect 382372 225564 382424 225616
rect 445576 225564 445628 225616
rect 447784 225564 447836 225616
rect 454224 225564 454276 225616
rect 372712 225020 372764 225072
rect 371608 224952 371660 225004
rect 374460 224952 374512 225004
rect 379520 224952 379572 225004
rect 441804 224952 441856 225004
rect 302700 224340 302752 224392
rect 369860 224340 369912 224392
rect 302884 224272 302936 224324
rect 370044 224272 370096 224324
rect 302792 224204 302844 224256
rect 370320 224204 370372 224256
rect 372252 224204 372304 224256
rect 373356 224204 373408 224256
rect 377128 224204 377180 224256
rect 359556 224068 359608 224120
rect 376944 224136 376996 224188
rect 379612 224204 379664 224256
rect 359740 224000 359792 224052
rect 382464 224136 382516 224188
rect 382648 224136 382700 224188
rect 379520 224000 379572 224052
rect 380992 224000 381044 224052
rect 359648 223932 359700 223984
rect 383660 223932 383712 223984
rect 358912 223864 358964 223916
rect 372712 223864 372764 223916
rect 441804 223864 441856 223916
rect 452752 223864 452804 223916
rect 454132 223864 454184 223916
rect 372804 223796 372856 223848
rect 371608 223728 371660 223780
rect 379520 223728 379572 223780
rect 193864 223592 193916 223644
rect 198280 223592 198332 223644
rect 441712 223592 441764 223644
rect 441896 223592 441948 223644
rect 370872 223524 370924 223576
rect 371424 223524 371476 223576
rect 378232 223524 378284 223576
rect 380992 223524 381044 223576
rect 447508 223524 447560 223576
rect 450268 223524 450320 223576
rect 371608 223456 371660 223508
rect 377404 223456 377456 223508
rect 381176 223456 381228 223508
rect 445668 223116 445720 223168
rect 447508 223116 447560 223168
rect 371608 222640 371660 222692
rect 375564 222640 375616 222692
rect 381084 222640 381136 222692
rect 170496 222164 170548 222216
rect 197360 222164 197412 222216
rect 302792 222096 302844 222148
rect 358912 222096 358964 222148
rect 375380 222096 375432 222148
rect 378416 222096 378468 222148
rect 377036 222028 377088 222080
rect 378508 222028 378560 222080
rect 445668 221212 445720 221264
rect 451464 221212 451516 221264
rect 452660 221212 452712 221264
rect 370412 220872 370464 220924
rect 377036 220872 377088 220924
rect 374920 220736 374972 220788
rect 378324 220736 378376 220788
rect 445668 220736 445720 220788
rect 446496 220736 446548 220788
rect 448888 220736 448940 220788
rect 375656 220668 375708 220720
rect 378232 220668 378284 220720
rect 450176 219988 450228 220040
rect 451280 219988 451332 220040
rect 369860 219648 369912 219700
rect 375656 219648 375708 219700
rect 445668 219580 445720 219632
rect 450176 219580 450228 219632
rect 369860 219512 369912 219564
rect 370228 219512 370280 219564
rect 180248 219444 180300 219496
rect 197544 219444 197596 219496
rect 373264 219444 373316 219496
rect 374828 219444 374880 219496
rect 302792 219376 302844 219428
rect 359740 219376 359792 219428
rect 369860 219376 369912 219428
rect 376024 219376 376076 219428
rect 446128 218900 446180 218952
rect 448612 218900 448664 218952
rect 369952 218832 370004 218884
rect 373356 218832 373408 218884
rect 376760 218832 376812 218884
rect 370044 218696 370096 218748
rect 376852 218696 376904 218748
rect 445484 218424 445536 218476
rect 446128 218424 446180 218476
rect 196808 218152 196860 218204
rect 198464 218152 198516 218204
rect 376024 218016 376076 218068
rect 378232 218016 378284 218068
rect 370136 217948 370188 218000
rect 370412 217948 370464 218000
rect 374736 217948 374788 218000
rect 376852 217948 376904 218000
rect 445668 217336 445720 217388
rect 449992 217336 450044 217388
rect 370320 216928 370372 216980
rect 374920 216928 374972 216980
rect 375748 216928 375800 216980
rect 302792 216588 302844 216640
rect 359648 216588 359700 216640
rect 382648 216588 382700 216640
rect 383660 216588 383712 216640
rect 371608 216520 371660 216572
rect 382464 216520 382516 216572
rect 383752 216520 383804 216572
rect 372068 216384 372120 216436
rect 372804 216384 372856 216436
rect 375840 216384 375892 216436
rect 445668 216112 445720 216164
rect 447876 216112 447928 216164
rect 195428 215296 195480 215348
rect 197912 215296 197964 215348
rect 371608 215296 371660 215348
rect 382280 215296 382332 215348
rect 382648 215296 382700 215348
rect 447876 215296 447928 215348
rect 448796 215296 448848 215348
rect 3332 215228 3384 215280
rect 199384 215228 199436 215280
rect 445484 214752 445536 214804
rect 448520 214752 448572 214804
rect 450084 214752 450136 214804
rect 371608 214616 371660 214668
rect 376116 214616 376168 214668
rect 379612 214616 379664 214668
rect 371700 214548 371752 214600
rect 376944 214548 376996 214600
rect 191288 213936 191340 213988
rect 197360 213936 197412 213988
rect 302792 213868 302844 213920
rect 359556 213868 359608 213920
rect 445668 213868 445720 213920
rect 447324 213868 447376 213920
rect 449900 213868 449952 213920
rect 371700 213256 371752 213308
rect 374644 213256 374696 213308
rect 380900 213256 380952 213308
rect 371608 213188 371660 213240
rect 382556 213188 382608 213240
rect 371424 213052 371476 213104
rect 375748 213052 375800 213104
rect 380808 213052 380860 213104
rect 445668 212712 445720 212764
rect 446680 212712 446732 212764
rect 448612 212712 448664 212764
rect 446036 212440 446088 212492
rect 448704 212440 448756 212492
rect 373172 211964 373224 212016
rect 375472 211964 375524 212016
rect 371424 211828 371476 211880
rect 377220 211828 377272 211880
rect 370228 211760 370280 211812
rect 378140 211760 378192 211812
rect 445484 211556 445536 211608
rect 446036 211556 446088 211608
rect 188528 211148 188580 211200
rect 197728 211148 197780 211200
rect 373080 210604 373132 210656
rect 374552 210604 374604 210656
rect 445392 210468 445444 210520
rect 447232 210468 447284 210520
rect 445208 209176 445260 209228
rect 446588 209176 446640 209228
rect 187148 208360 187200 208412
rect 197360 208360 197412 208412
rect 446588 208360 446640 208412
rect 447416 208360 447468 208412
rect 444748 207884 444800 207936
rect 445944 207884 445996 207936
rect 447140 207884 447192 207936
rect 173164 207000 173216 207052
rect 197360 207000 197412 207052
rect 450544 206932 450596 206984
rect 579804 206932 579856 206984
rect 371608 206252 371660 206304
rect 374184 206252 374236 206304
rect 371700 205776 371752 205828
rect 372988 205776 373040 205828
rect 302332 205640 302384 205692
rect 359556 205640 359608 205692
rect 373816 205572 373868 205624
rect 374184 205572 374236 205624
rect 369124 205164 369176 205216
rect 369308 205164 369360 205216
rect 173256 204280 173308 204332
rect 197544 204280 197596 204332
rect 372068 204212 372120 204264
rect 374000 204212 374052 204264
rect 173348 202852 173400 202904
rect 197360 202852 197412 202904
rect 302792 202852 302844 202904
rect 359648 202852 359700 202904
rect 3056 202784 3108 202836
rect 177396 202784 177448 202836
rect 370136 202716 370188 202768
rect 374276 202716 374328 202768
rect 373172 202648 373224 202700
rect 375380 202648 375432 202700
rect 372620 202512 372672 202564
rect 373264 202512 373316 202564
rect 371608 201560 371660 201612
rect 374000 201560 374052 201612
rect 374368 201560 374420 201612
rect 445668 201492 445720 201544
rect 448520 201492 448572 201544
rect 452936 201492 452988 201544
rect 173440 200132 173492 200184
rect 197360 200132 197412 200184
rect 445668 200132 445720 200184
rect 449256 200132 449308 200184
rect 452660 200132 452712 200184
rect 445668 199452 445720 199504
rect 449900 199452 449952 199504
rect 454040 199452 454092 199504
rect 445668 198772 445720 198824
rect 451372 198772 451424 198824
rect 173532 198704 173584 198756
rect 197360 198704 197412 198756
rect 302516 198704 302568 198756
rect 359372 198704 359424 198756
rect 445668 197752 445720 197804
rect 447140 197752 447192 197804
rect 452844 197752 452896 197804
rect 302884 197208 302936 197260
rect 379612 197208 379664 197260
rect 302700 197140 302752 197192
rect 370320 197140 370372 197192
rect 359648 197072 359700 197124
rect 382464 197072 382516 197124
rect 359372 197004 359424 197056
rect 380900 197004 380952 197056
rect 359556 196936 359608 196988
rect 375748 196936 375800 196988
rect 302976 196664 303028 196716
rect 369860 196664 369912 196716
rect 303068 196596 303120 196648
rect 375380 196596 375432 196648
rect 369860 196052 369912 196104
rect 371148 196052 371200 196104
rect 173624 195984 173676 196036
rect 197360 195984 197412 196036
rect 322204 195916 322256 195968
rect 438768 195916 438820 195968
rect 302884 195236 302936 195288
rect 370504 195236 370556 195288
rect 302424 194488 302476 194540
rect 370964 194488 371016 194540
rect 372712 194488 372764 194540
rect 437388 194488 437440 194540
rect 441804 194488 441856 194540
rect 318064 194420 318116 194472
rect 366916 194420 366968 194472
rect 436008 194420 436060 194472
rect 441712 194420 441764 194472
rect 196900 194352 196952 194404
rect 198648 194352 198700 194404
rect 435180 193604 435232 193656
rect 436008 193604 436060 193656
rect 373080 193196 373132 193248
rect 374092 193196 374144 193248
rect 446404 193128 446456 193180
rect 580172 193128 580224 193180
rect 176016 191836 176068 191888
rect 197360 191836 197412 191888
rect 172428 190408 172480 190460
rect 188344 190408 188396 190460
rect 172428 188980 172480 189032
rect 184296 188980 184348 189032
rect 181536 187688 181588 187740
rect 197360 187688 197412 187740
rect 172428 187620 172480 187672
rect 186964 187620 187016 187672
rect 302700 187620 302752 187672
rect 374092 187620 374144 187672
rect 172428 186260 172480 186312
rect 193956 186260 194008 186312
rect 182916 184900 182968 184952
rect 197360 184900 197412 184952
rect 172336 184832 172388 184884
rect 196624 184832 196676 184884
rect 302792 184832 302844 184884
rect 370136 184832 370188 184884
rect 374276 184832 374328 184884
rect 172428 184764 172480 184816
rect 182824 184764 182876 184816
rect 172428 183472 172480 183524
rect 181444 183472 181496 183524
rect 178868 182792 178920 182844
rect 197544 182792 197596 182844
rect 172428 182044 172480 182096
rect 178776 182044 178828 182096
rect 172152 180820 172204 180872
rect 197360 180820 197412 180872
rect 172428 180548 172480 180600
rect 175924 180548 175976 180600
rect 461584 179324 461636 179376
rect 580172 179324 580224 179376
rect 172428 179188 172480 179240
rect 174544 179188 174596 179240
rect 191380 178032 191432 178084
rect 197544 178032 197596 178084
rect 172428 177964 172480 178016
rect 196716 177964 196768 178016
rect 172336 177896 172388 177948
rect 180156 177896 180208 177948
rect 180340 176672 180392 176724
rect 197360 176672 197412 176724
rect 172428 176604 172480 176656
rect 195336 176604 195388 176656
rect 171692 175176 171744 175228
rect 191104 175176 191156 175228
rect 302240 175176 302292 175228
rect 370872 175176 370924 175228
rect 369768 175108 369820 175160
rect 373816 175108 373868 175160
rect 446128 175176 446180 175228
rect 188344 173884 188396 173936
rect 197636 173884 197688 173936
rect 171508 173816 171560 173868
rect 188436 173816 188488 173868
rect 174544 172524 174596 172576
rect 197360 172524 197412 172576
rect 172428 172456 172480 172508
rect 187056 172456 187108 172508
rect 370136 172456 370188 172508
rect 371700 172456 371752 172508
rect 302792 171096 302844 171148
rect 370136 171096 370188 171148
rect 172428 171028 172480 171080
rect 198004 171028 198056 171080
rect 186964 169736 187016 169788
rect 197360 169736 197412 169788
rect 172428 169668 172480 169720
rect 198096 169668 198148 169720
rect 369676 169668 369728 169720
rect 374736 169668 374788 169720
rect 448704 169668 448756 169720
rect 369584 168308 369636 168360
rect 374644 168308 374696 168360
rect 450084 168308 450136 168360
rect 195336 167016 195388 167068
rect 197912 167016 197964 167068
rect 172428 166948 172480 167000
rect 192484 166948 192536 167000
rect 301504 166948 301556 167000
rect 580172 166948 580224 167000
rect 191104 166064 191156 166116
rect 198464 166064 198516 166116
rect 171784 164840 171836 164892
rect 191196 164840 191248 164892
rect 447416 164228 447468 164280
rect 3240 164160 3292 164212
rect 159364 164160 159416 164212
rect 172428 164160 172480 164212
rect 184388 164160 184440 164212
rect 370044 164160 370096 164212
rect 370504 164160 370556 164212
rect 370596 164160 370648 164212
rect 372988 164160 373040 164212
rect 449992 164160 450044 164212
rect 370228 162664 370280 162716
rect 371148 162664 371200 162716
rect 372068 162188 372120 162240
rect 444656 162188 444708 162240
rect 171784 162120 171836 162172
rect 191380 162120 191432 162172
rect 302700 162120 302752 162172
rect 370228 162120 370280 162172
rect 373264 162120 373316 162172
rect 447232 162120 447284 162172
rect 184296 161440 184348 161492
rect 197360 161440 197412 161492
rect 172244 161100 172296 161152
rect 177488 161100 177540 161152
rect 169208 160760 169260 160812
rect 180064 160760 180116 160812
rect 165160 160488 165212 160540
rect 195244 160692 195296 160744
rect 369860 160012 369912 160064
rect 446036 160080 446088 160132
rect 447324 160012 447376 160064
rect 369400 159944 369452 159996
rect 373908 159944 373960 159996
rect 180064 158720 180116 158772
rect 197360 158720 197412 158772
rect 162860 158652 162912 158704
rect 184204 158652 184256 158704
rect 166908 157972 166960 158024
rect 196624 157972 196676 158024
rect 371884 157972 371936 158024
rect 444472 157972 444524 158024
rect 177396 157360 177448 157412
rect 197360 157360 197412 157412
rect 369492 156612 369544 156664
rect 374552 156612 374604 156664
rect 444748 156612 444800 156664
rect 448612 156612 448664 156664
rect 436008 155864 436060 155916
rect 441712 155864 441764 155916
rect 188436 155184 188488 155236
rect 198188 155184 198240 155236
rect 372160 155184 372212 155236
rect 444564 155184 444616 155236
rect 171232 154504 171284 154556
rect 196808 154504 196860 154556
rect 302792 154504 302844 154556
rect 370044 154504 370096 154556
rect 370596 154504 370648 154556
rect 371700 154504 371752 154556
rect 382372 154504 382424 154556
rect 445668 154504 445720 154556
rect 454224 154504 454276 154556
rect 171600 153960 171652 154012
rect 180248 153960 180300 154012
rect 370136 153824 370188 153876
rect 444932 153824 444984 153876
rect 451464 153824 451516 153876
rect 437388 153552 437440 153604
rect 441896 153552 441948 153604
rect 371700 153348 371752 153400
rect 374460 153348 374512 153400
rect 172428 153144 172480 153196
rect 195428 153144 195480 153196
rect 302976 153144 303028 153196
rect 369768 153144 369820 153196
rect 371516 153144 371568 153196
rect 379520 153144 379572 153196
rect 443644 153144 443696 153196
rect 580172 153144 580224 153196
rect 172336 153076 172388 153128
rect 191288 153076 191340 153128
rect 302884 153076 302936 153128
rect 369676 153076 369728 153128
rect 371700 153076 371752 153128
rect 377128 153076 377180 153128
rect 302792 153008 302844 153060
rect 369584 153008 369636 153060
rect 369676 152736 369728 152788
rect 369952 152736 370004 152788
rect 302700 152464 302752 152516
rect 369216 152464 369268 152516
rect 369584 152464 369636 152516
rect 370320 152464 370372 152516
rect 359372 151988 359424 152040
rect 369308 151988 369360 152040
rect 359556 151920 359608 151972
rect 369124 151920 369176 151972
rect 369860 151920 369912 151972
rect 359004 151852 359056 151904
rect 369492 151852 369544 151904
rect 444840 151852 444892 151904
rect 452752 151852 452804 151904
rect 371700 151716 371752 151768
rect 381176 151716 381228 151768
rect 172336 151648 172388 151700
rect 187148 151648 187200 151700
rect 371516 151648 371568 151700
rect 380992 151648 381044 151700
rect 172428 151580 172480 151632
rect 188528 151580 188580 151632
rect 444840 151308 444892 151360
rect 447508 151308 447560 151360
rect 187056 151036 187108 151088
rect 198280 151036 198332 151088
rect 371700 151036 371752 151088
rect 375564 151036 375616 151088
rect 196716 150560 196768 150612
rect 198372 150560 198424 150612
rect 171876 150492 171928 150544
rect 173164 150492 173216 150544
rect 3424 150356 3476 150408
rect 11704 150356 11756 150408
rect 302792 150356 302844 150408
rect 359372 150356 359424 150408
rect 371700 150356 371752 150408
rect 378416 150356 378468 150408
rect 371516 150288 371568 150340
rect 377036 150288 377088 150340
rect 171508 150016 171560 150068
rect 173256 150016 173308 150068
rect 171692 149404 171744 149456
rect 173348 149404 173400 149456
rect 171692 148996 171744 149048
rect 173532 148996 173584 149048
rect 371700 148996 371752 149048
rect 378324 148996 378376 149048
rect 171876 148860 171928 148912
rect 173440 148860 173492 148912
rect 445300 148860 445352 148912
rect 448888 148860 448940 148912
rect 371700 148384 371752 148436
rect 374828 148384 374880 148436
rect 173164 148316 173216 148368
rect 198004 148316 198056 148368
rect 171692 148180 171744 148232
rect 173624 148180 173676 148232
rect 371700 148180 371752 148232
rect 375656 148180 375708 148232
rect 445576 148112 445628 148164
rect 450176 148112 450228 148164
rect 195244 147636 195296 147688
rect 198280 147636 198332 147688
rect 172428 147568 172480 147620
rect 196900 147568 196952 147620
rect 171876 147500 171928 147552
rect 176016 147500 176068 147552
rect 371240 147500 371292 147552
rect 378232 147500 378284 147552
rect 371240 146684 371292 146736
rect 373356 146684 373408 146736
rect 444840 146548 444892 146600
rect 446128 146548 446180 146600
rect 191196 146480 191248 146532
rect 197728 146480 197780 146532
rect 172336 146208 172388 146260
rect 182916 146208 182968 146260
rect 302792 146208 302844 146260
rect 359004 146208 359056 146260
rect 172428 146140 172480 146192
rect 181536 146140 181588 146192
rect 371516 146140 371568 146192
rect 376852 146140 376904 146192
rect 172244 146072 172296 146124
rect 178868 146072 178920 146124
rect 371700 146072 371752 146124
rect 376760 146072 376812 146124
rect 445484 146004 445536 146056
rect 449992 146004 450044 146056
rect 371700 145052 371752 145104
rect 374920 145052 374972 145104
rect 172428 144848 172480 144900
rect 188436 144848 188488 144900
rect 371516 144848 371568 144900
rect 383752 144848 383804 144900
rect 372068 144780 372120 144832
rect 382280 144780 382332 144832
rect 445116 144712 445168 144764
rect 448704 144712 448756 144764
rect 371700 144508 371752 144560
rect 375840 144508 375892 144560
rect 171692 144168 171744 144220
rect 188344 144168 188396 144220
rect 188528 143556 188580 143608
rect 197360 143556 197412 143608
rect 171876 143488 171928 143540
rect 180340 143488 180392 143540
rect 302792 143488 302844 143540
rect 359556 143488 359608 143540
rect 371240 143488 371292 143540
rect 379612 143488 379664 143540
rect 371700 143420 371752 143472
rect 376944 143420 376996 143472
rect 445116 143148 445168 143200
rect 450084 143148 450136 143200
rect 171784 142808 171836 142860
rect 186964 142808 187016 142860
rect 171508 142264 171560 142316
rect 174544 142264 174596 142316
rect 187148 142128 187200 142180
rect 197360 142128 197412 142180
rect 172428 142060 172480 142112
rect 195336 142060 195388 142112
rect 371516 142060 371568 142112
rect 382464 142060 382516 142112
rect 444380 142060 444432 142112
rect 444840 142060 444892 142112
rect 371240 141992 371292 142044
rect 380900 141992 380952 142044
rect 371700 141924 371752 141976
rect 375748 141924 375800 141976
rect 444380 141924 444432 141976
rect 447324 141924 447376 141976
rect 171692 141380 171744 141432
rect 191104 141380 191156 141432
rect 371700 140632 371752 140684
rect 378140 140632 378192 140684
rect 444380 140428 444432 140480
rect 446036 140428 446088 140480
rect 172336 140020 172388 140072
rect 198096 140020 198148 140072
rect 171692 139748 171744 139800
rect 173164 139748 173216 139800
rect 172428 139340 172480 139392
rect 184296 139340 184348 139392
rect 371516 139340 371568 139392
rect 374276 139340 374328 139392
rect 465724 139340 465776 139392
rect 580172 139340 580224 139392
rect 371700 139204 371752 139256
rect 375380 139204 375432 139256
rect 171600 139068 171652 139120
rect 180064 139068 180116 139120
rect 371700 138864 371752 138916
rect 374092 138864 374144 138916
rect 444380 138592 444432 138644
rect 447232 138592 447284 138644
rect 171508 138184 171560 138236
rect 177396 138184 177448 138236
rect 3240 137912 3292 137964
rect 152464 137912 152516 137964
rect 172060 137912 172112 137964
rect 187056 137912 187108 137964
rect 444380 137300 444432 137352
rect 447416 137300 447468 137352
rect 172428 137232 172480 137284
rect 196716 137232 196768 137284
rect 172520 136620 172572 136672
rect 197544 136620 197596 136672
rect 172244 136552 172296 136604
rect 195244 136552 195296 136604
rect 171692 136484 171744 136536
rect 191196 136484 191248 136536
rect 172336 135260 172388 135312
rect 198096 135260 198148 135312
rect 171232 135192 171284 135244
rect 198280 135192 198332 135244
rect 369216 135192 369268 135244
rect 369400 135192 369452 135244
rect 172428 135124 172480 135176
rect 188528 135124 188580 135176
rect 172244 135056 172296 135108
rect 187148 135056 187200 135108
rect 171140 132472 171192 132524
rect 197544 132472 197596 132524
rect 172428 131724 172480 131776
rect 197912 131724 197964 131776
rect 370228 130636 370280 130688
rect 373264 130636 373316 130688
rect 443920 130364 443972 130416
rect 448520 130364 448572 130416
rect 171876 130024 171928 130076
rect 179420 130024 179472 130076
rect 171508 129684 171560 129736
rect 197360 129684 197412 129736
rect 369860 129072 369912 129124
rect 374000 129072 374052 129124
rect 427820 129072 427872 129124
rect 370320 129004 370372 129056
rect 371424 129004 371476 129056
rect 430580 129004 430632 129056
rect 443644 128324 443696 128376
rect 452660 128324 452712 128376
rect 444380 128052 444432 128104
rect 449900 128052 449952 128104
rect 172520 127576 172572 127628
rect 198004 127576 198056 127628
rect 172336 126896 172388 126948
rect 197360 126896 197412 126948
rect 449164 126896 449216 126948
rect 580172 126896 580224 126948
rect 444380 126624 444432 126676
rect 447140 126624 447192 126676
rect 372436 126012 372488 126064
rect 443092 126012 443144 126064
rect 371792 125944 371844 125996
rect 443000 125944 443052 125996
rect 370412 125876 370464 125928
rect 371608 125876 371660 125928
rect 443644 125876 443696 125928
rect 172428 125740 172480 125792
rect 186964 125740 187016 125792
rect 172336 125672 172388 125724
rect 188344 125672 188396 125724
rect 172244 125604 172296 125656
rect 191104 125604 191156 125656
rect 179420 125536 179472 125588
rect 198556 125536 198608 125588
rect 370504 125468 370556 125520
rect 372620 125468 372672 125520
rect 441620 125468 441672 125520
rect 427820 125400 427872 125452
rect 444748 125400 444800 125452
rect 430580 125332 430632 125384
rect 444840 125332 444892 125384
rect 371332 125264 371384 125316
rect 441896 125264 441948 125316
rect 302792 125196 302844 125248
rect 370320 125196 370372 125248
rect 303068 125128 303120 125180
rect 369860 125128 369912 125180
rect 302884 125060 302936 125112
rect 370228 125060 370280 125112
rect 302976 124992 303028 125044
rect 369952 124992 370004 125044
rect 302608 124924 302660 124976
rect 370044 124924 370096 124976
rect 370780 124856 370832 124908
rect 441896 124856 441948 124908
rect 445852 124856 445904 124908
rect 172428 124312 172480 124364
rect 184204 124312 184256 124364
rect 171692 124244 171744 124296
rect 180064 124244 180116 124296
rect 172152 124176 172204 124228
rect 173164 124176 173216 124228
rect 302700 124108 302752 124160
rect 371240 124108 371292 124160
rect 302976 123564 303028 123616
rect 370412 123564 370464 123616
rect 302884 123428 302936 123480
rect 369952 123428 370004 123480
rect 160928 122952 160980 123004
rect 170496 122952 170548 123004
rect 162860 122884 162912 122936
rect 193864 122884 193916 122936
rect 164884 122816 164936 122868
rect 198740 122816 198792 122868
rect 166908 122748 166960 122800
rect 178684 122748 178736 122800
rect 320824 122748 320876 122800
rect 438860 122748 438912 122800
rect 168932 122680 168984 122732
rect 177304 122680 177356 122732
rect 359464 122680 359516 122732
rect 366916 122680 366968 122732
rect 437204 122680 437256 122732
rect 441804 122680 441856 122732
rect 435180 122612 435232 122664
rect 441712 122612 441764 122664
rect 172060 121388 172112 121440
rect 197544 121388 197596 121440
rect 302792 121388 302844 121440
rect 370136 121388 370188 121440
rect 188344 119348 188396 119400
rect 198004 119348 198056 119400
rect 171876 118600 171928 118652
rect 198096 118600 198148 118652
rect 302792 118600 302844 118652
rect 371792 118600 371844 118652
rect 171968 117240 172020 117292
rect 197544 117240 197596 117292
rect 171784 114452 171836 114504
rect 197360 114452 197412 114504
rect 313924 113092 313976 113144
rect 579804 113092 579856 113144
rect 3424 111732 3476 111784
rect 170404 111732 170456 111784
rect 191104 111732 191156 111784
rect 197360 111732 197412 111784
rect 302332 111732 302384 111784
rect 370596 111732 370648 111784
rect 302792 108944 302844 108996
rect 371332 108944 371384 108996
rect 186964 107584 187016 107636
rect 198556 107584 198608 107636
rect 184204 106224 184256 106276
rect 197544 106224 197596 106276
rect 180064 103436 180116 103488
rect 197912 103436 197964 103488
rect 173164 102076 173216 102128
rect 197544 102076 197596 102128
rect 302792 102076 302844 102128
rect 369860 102076 369912 102128
rect 457444 100648 457496 100700
rect 580172 100648 580224 100700
rect 196624 99356 196676 99408
rect 299480 99356 299532 99408
rect 112444 99288 112496 99340
rect 217600 99288 217652 99340
rect 278872 99288 278924 99340
rect 414664 99288 414716 99340
rect 98644 99220 98696 99272
rect 213368 99220 213420 99272
rect 240508 99220 240560 99272
rect 241060 99220 241112 99272
rect 271052 99220 271104 99272
rect 413284 99220 413336 99272
rect 97264 99152 97316 99204
rect 211528 99152 211580 99204
rect 271604 99152 271656 99204
rect 417424 99152 417476 99204
rect 88984 99084 89036 99136
rect 209780 99084 209832 99136
rect 272248 99084 272300 99136
rect 421564 99084 421616 99136
rect 93124 99016 93176 99068
rect 215392 99016 215444 99068
rect 273444 99016 273496 99068
rect 430580 99016 430632 99068
rect 87604 98948 87656 99000
rect 214380 98948 214432 99000
rect 274640 98948 274692 99000
rect 435364 98948 435416 99000
rect 71044 98880 71096 98932
rect 210332 98880 210384 98932
rect 275284 98880 275336 98932
rect 439504 98880 439556 98932
rect 43444 98812 43496 98864
rect 205916 98812 205968 98864
rect 276480 98812 276532 98864
rect 448520 98812 448572 98864
rect 22744 98744 22796 98796
rect 203064 98744 203116 98796
rect 283380 98744 283432 98796
rect 486424 98744 486476 98796
rect 33784 98676 33836 98728
rect 204536 98676 204588 98728
rect 290004 98676 290056 98728
rect 525064 98676 525116 98728
rect 21364 98608 21416 98660
rect 202880 98608 202932 98660
rect 297088 98608 297140 98660
rect 568580 98608 568632 98660
rect 259920 98540 259972 98592
rect 348424 98540 348476 98592
rect 259368 98472 259420 98524
rect 345664 98472 345716 98524
rect 258724 98404 258776 98456
rect 342904 98404 342956 98456
rect 211160 98268 211212 98320
rect 211436 98268 211488 98320
rect 211620 98268 211672 98320
rect 211988 98268 212040 98320
rect 216036 98268 216088 98320
rect 216404 98268 216456 98320
rect 238208 98268 238260 98320
rect 238484 98268 238536 98320
rect 274456 98064 274508 98116
rect 278228 98064 278280 98116
rect 278136 97996 278188 98048
rect 3424 97928 3476 97980
rect 14464 97928 14516 97980
rect 150348 97928 150400 97980
rect 225512 97928 225564 97980
rect 269028 97928 269080 97980
rect 282368 97928 282420 97980
rect 286784 97996 286836 98048
rect 286968 97996 287020 98048
rect 295984 97996 296036 98048
rect 296352 97996 296404 98048
rect 323676 97928 323728 97980
rect 126888 97860 126940 97912
rect 210884 97860 210936 97912
rect 231308 97860 231360 97912
rect 238024 97860 238076 97912
rect 246856 97860 246908 97912
rect 253204 97860 253256 97912
rect 272340 97860 272392 97912
rect 309876 97860 309928 97912
rect 124864 97792 124916 97844
rect 202512 97792 202564 97844
rect 202788 97792 202840 97844
rect 126244 97724 126296 97776
rect 210240 97724 210292 97776
rect 234528 97792 234580 97844
rect 247684 97792 247736 97844
rect 251824 97792 251876 97844
rect 272248 97792 272300 97844
rect 341524 97792 341576 97844
rect 210884 97724 210936 97776
rect 221464 97724 221516 97776
rect 245476 97724 245528 97776
rect 253020 97724 253072 97776
rect 259736 97724 259788 97776
rect 115204 97656 115256 97708
rect 219440 97656 219492 97708
rect 254124 97656 254176 97708
rect 111064 97588 111116 97640
rect 215760 97588 215812 97640
rect 241980 97588 242032 97640
rect 242716 97588 242768 97640
rect 247500 97588 247552 97640
rect 256792 97588 256844 97640
rect 256976 97656 257028 97708
rect 263140 97656 263192 97708
rect 267188 97724 267240 97776
rect 352564 97724 352616 97776
rect 347044 97656 347096 97708
rect 263876 97588 263928 97640
rect 264980 97588 265032 97640
rect 268200 97588 268252 97640
rect 270224 97588 270276 97640
rect 94504 97520 94556 97572
rect 204076 97520 204128 97572
rect 104164 97452 104216 97504
rect 217048 97520 217100 97572
rect 212540 97452 212592 97504
rect 225052 97520 225104 97572
rect 248696 97520 248748 97572
rect 263048 97520 263100 97572
rect 263692 97520 263744 97572
rect 272340 97520 272392 97572
rect 220176 97452 220228 97504
rect 229928 97452 229980 97504
rect 251088 97452 251140 97504
rect 263600 97452 263652 97504
rect 264796 97452 264848 97504
rect 272248 97452 272300 97504
rect 277952 97588 278004 97640
rect 369124 97588 369176 97640
rect 377404 97520 377456 97572
rect 278136 97452 278188 97504
rect 388444 97452 388496 97504
rect 213920 97384 213972 97436
rect 232964 97384 233016 97436
rect 243820 97384 243872 97436
rect 258264 97384 258316 97436
rect 262404 97384 262456 97436
rect 265072 97384 265124 97436
rect 265440 97384 265492 97436
rect 271052 97384 271104 97436
rect 58624 97316 58676 97368
rect 206744 97316 206796 97368
rect 208308 97316 208360 97368
rect 227536 97316 227588 97368
rect 227628 97316 227680 97368
rect 238760 97316 238812 97368
rect 263416 97316 263468 97368
rect 275652 97316 275704 97368
rect 25504 97248 25556 97300
rect 203340 97248 203392 97300
rect 204168 97248 204220 97300
rect 234712 97248 234764 97300
rect 253204 97248 253256 97300
rect 271144 97248 271196 97300
rect 191196 97180 191248 97232
rect 218244 97180 218296 97232
rect 243176 97180 243228 97232
rect 259460 97180 259512 97232
rect 265072 97180 265124 97232
rect 188436 97112 188488 97164
rect 207296 97112 207348 97164
rect 196624 97044 196676 97096
rect 210976 97112 211028 97164
rect 211160 97112 211212 97164
rect 222660 97112 222712 97164
rect 242992 97112 243044 97164
rect 250260 97112 250312 97164
rect 255964 97112 256016 97164
rect 256608 97112 256660 97164
rect 256792 97112 256844 97164
rect 260104 97112 260156 97164
rect 261208 97112 261260 97164
rect 268384 97180 268436 97232
rect 276572 97248 276624 97300
rect 276848 97316 276900 97368
rect 277216 97316 277268 97368
rect 278320 97384 278372 97436
rect 393964 97384 394016 97436
rect 277952 97316 278004 97368
rect 282644 97316 282696 97368
rect 283656 97316 283708 97368
rect 411904 97316 411956 97368
rect 283012 97248 283064 97300
rect 418804 97248 418856 97300
rect 271420 97180 271472 97232
rect 278136 97180 278188 97232
rect 278228 97180 278280 97232
rect 282184 97180 282236 97232
rect 210240 97044 210292 97096
rect 221280 97044 221332 97096
rect 241428 97044 241480 97096
rect 242164 97044 242216 97096
rect 242440 97044 242492 97096
rect 246304 97044 246356 97096
rect 199384 96976 199436 97028
rect 209136 96976 209188 97028
rect 204260 96908 204312 96960
rect 207756 96908 207808 96960
rect 223580 96908 223632 96960
rect 225236 96908 225288 96960
rect 244464 96908 244516 96960
rect 245292 96908 245344 96960
rect 245844 96908 245896 96960
rect 246488 96908 246540 96960
rect 247224 96908 247276 96960
rect 248236 96908 248288 96960
rect 203892 96840 203944 96892
rect 207940 96840 207992 96892
rect 237380 96840 237432 96892
rect 239220 96840 239272 96892
rect 241796 96840 241848 96892
rect 244372 96840 244424 96892
rect 245660 96840 245712 96892
rect 246672 96840 246724 96892
rect 249708 97044 249760 97096
rect 256148 97044 256200 97096
rect 256424 97044 256476 97096
rect 260564 97044 260616 97096
rect 262864 97044 262916 97096
rect 271236 97112 271288 97164
rect 278688 97112 278740 97164
rect 304264 97180 304316 97232
rect 287980 97112 288032 97164
rect 288256 97112 288308 97164
rect 288808 97112 288860 97164
rect 289728 97112 289780 97164
rect 292212 97112 292264 97164
rect 292488 97112 292540 97164
rect 296076 97112 296128 97164
rect 296352 97112 296404 97164
rect 296628 97112 296680 97164
rect 322204 97112 322256 97164
rect 274180 97044 274232 97096
rect 250444 96976 250496 97028
rect 251088 96976 251140 97028
rect 251456 96976 251508 97028
rect 252284 96976 252336 97028
rect 258172 96976 258224 97028
rect 259000 96976 259052 97028
rect 262772 96976 262824 97028
rect 263508 96976 263560 97028
rect 265624 96976 265676 97028
rect 266268 96976 266320 97028
rect 266452 96976 266504 97028
rect 267464 96976 267516 97028
rect 268660 96976 268712 97028
rect 269028 96976 269080 97028
rect 269212 96976 269264 97028
rect 270316 96976 270368 97028
rect 272064 96976 272116 97028
rect 278228 96976 278280 97028
rect 250076 96908 250128 96960
rect 250996 96908 251048 96960
rect 251916 96908 251968 96960
rect 252192 96908 252244 96960
rect 253112 96908 253164 96960
rect 253572 96908 253624 96960
rect 254860 96908 254912 96960
rect 255136 96908 255188 96960
rect 255504 96908 255556 96960
rect 256332 96908 256384 96960
rect 257620 96908 257672 96960
rect 257896 96908 257948 96960
rect 258540 96908 258592 96960
rect 259092 96908 259144 96960
rect 260196 96908 260248 96960
rect 260656 96908 260708 96960
rect 262956 96908 263008 96960
rect 263416 96908 263468 96960
rect 264428 96908 264480 96960
rect 264888 96908 264940 96960
rect 265808 96908 265860 96960
rect 266084 96908 266136 96960
rect 267004 96908 267056 96960
rect 267372 96908 267424 96960
rect 268016 96908 268068 96960
rect 268936 96908 268988 96960
rect 269672 96908 269724 96960
rect 270132 96908 270184 96960
rect 270868 96908 270920 96960
rect 271788 96908 271840 96960
rect 272432 96908 272484 96960
rect 272984 96908 273036 96960
rect 273260 96908 273312 96960
rect 273904 96908 273956 96960
rect 275652 96908 275704 96960
rect 275928 96908 275980 96960
rect 276296 96908 276348 96960
rect 279148 96976 279200 97028
rect 281172 96976 281224 97028
rect 280160 96908 280212 96960
rect 281356 96908 281408 96960
rect 281724 97044 281776 97096
rect 284300 97044 284352 97096
rect 286324 97044 286376 97096
rect 286692 97044 286744 97096
rect 286784 97044 286836 97096
rect 312544 97044 312596 97096
rect 282368 96976 282420 97028
rect 297640 96976 297692 97028
rect 298008 96976 298060 97028
rect 298100 96976 298152 97028
rect 299112 96976 299164 97028
rect 250720 96840 250772 96892
rect 250904 96840 250956 96892
rect 252008 96840 252060 96892
rect 252468 96840 252520 96892
rect 252652 96840 252704 96892
rect 253756 96840 253808 96892
rect 253940 96840 253992 96892
rect 255044 96840 255096 96892
rect 256700 96840 256752 96892
rect 257804 96840 257856 96892
rect 258908 96840 258960 96892
rect 259276 96840 259328 96892
rect 261576 96840 261628 96892
rect 261944 96840 261996 96892
rect 262588 96840 262640 96892
rect 263324 96840 263376 96892
rect 263784 96840 263836 96892
rect 264612 96840 264664 96892
rect 265900 96840 265952 96892
rect 266176 96840 266228 96892
rect 266820 96840 266872 96892
rect 267556 96840 267608 96892
rect 267832 96840 267884 96892
rect 268844 96840 268896 96892
rect 269948 96840 270000 96892
rect 270408 96840 270460 96892
rect 272892 96840 272944 96892
rect 273168 96840 273220 96892
rect 276664 96840 276716 96892
rect 277216 96840 277268 96892
rect 280896 96840 280948 96892
rect 281448 96840 281500 96892
rect 282184 96840 282236 96892
rect 283656 96840 283708 96892
rect 283840 96840 283892 96892
rect 284116 96840 284168 96892
rect 285128 96840 285180 96892
rect 285404 96840 285456 96892
rect 285772 96840 285824 96892
rect 286416 96840 286468 96892
rect 287152 96840 287204 96892
rect 288164 96840 288216 96892
rect 288624 96840 288676 96892
rect 289268 96840 289320 96892
rect 290556 96840 290608 96892
rect 290924 96840 290976 96892
rect 291384 96840 291436 96892
rect 291936 96840 291988 96892
rect 293040 96840 293092 96892
rect 293408 96840 293460 96892
rect 293500 96840 293552 96892
rect 293868 96840 293920 96892
rect 294604 96840 294656 96892
rect 295248 96840 295300 96892
rect 295432 96840 295484 96892
rect 296076 96840 296128 96892
rect 86868 96772 86920 96824
rect 236000 96772 236052 96824
rect 239036 96772 239088 96824
rect 244648 96772 244700 96824
rect 245384 96772 245436 96824
rect 246212 96772 246264 96824
rect 246764 96772 246816 96824
rect 248420 96772 248472 96824
rect 249248 96772 249300 96824
rect 249340 96772 249392 96824
rect 254492 96772 254544 96824
rect 255136 96772 255188 96824
rect 256056 96772 256108 96824
rect 256516 96772 256568 96824
rect 257344 96772 257396 96824
rect 257896 96772 257948 96824
rect 258356 96772 258408 96824
rect 259368 96772 259420 96824
rect 260472 96772 260524 96824
rect 260748 96772 260800 96824
rect 263968 96772 264020 96824
rect 264704 96772 264756 96824
rect 266636 96772 266688 96824
rect 267280 96772 267332 96824
rect 270684 96772 270736 96824
rect 271604 96772 271656 96824
rect 272616 96772 272668 96824
rect 214472 96704 214524 96756
rect 215944 96704 215996 96756
rect 218796 96704 218848 96756
rect 219440 96704 219492 96756
rect 223028 96704 223080 96756
rect 233884 96704 233936 96756
rect 238576 96704 238628 96756
rect 246028 96704 246080 96756
rect 246856 96704 246908 96756
rect 260932 96704 260984 96756
rect 261852 96704 261904 96756
rect 265164 96704 265216 96756
rect 266176 96704 266228 96756
rect 269856 96704 269908 96756
rect 270224 96704 270276 96756
rect 271880 96704 271932 96756
rect 272892 96704 272944 96756
rect 274916 96772 274968 96824
rect 275928 96772 275980 96824
rect 276112 96772 276164 96824
rect 277124 96772 277176 96824
rect 280344 96772 280396 96824
rect 281080 96772 281132 96824
rect 281172 96772 281224 96824
rect 282276 96772 282328 96824
rect 283564 96772 283616 96824
rect 284024 96772 284076 96824
rect 284576 96772 284628 96824
rect 285312 96772 285364 96824
rect 285956 96772 286008 96824
rect 286600 96772 286652 96824
rect 287888 96772 287940 96824
rect 288348 96772 288400 96824
rect 288992 96772 289044 96824
rect 289544 96772 289596 96824
rect 291844 96772 291896 96824
rect 292304 96772 292356 96824
rect 292580 96772 292632 96824
rect 293684 96772 293736 96824
rect 295616 96772 295668 96824
rect 296260 96772 296312 96824
rect 286784 96704 286836 96756
rect 289176 96704 289228 96756
rect 289636 96704 289688 96756
rect 290188 96704 290240 96756
rect 290832 96704 290884 96756
rect 291200 96704 291252 96756
rect 292120 96704 292172 96756
rect 294880 96704 294932 96756
rect 295064 96704 295116 96756
rect 295800 96704 295852 96756
rect 296536 96704 296588 96756
rect 198004 96636 198056 96688
rect 200856 96636 200908 96688
rect 202144 96636 202196 96688
rect 205548 96636 205600 96688
rect 209044 96636 209096 96688
rect 212172 96636 212224 96688
rect 217416 96636 217468 96688
rect 219992 96636 220044 96688
rect 222200 96636 222252 96688
rect 224040 96636 224092 96688
rect 233976 96636 234028 96688
rect 237564 96636 237616 96688
rect 238024 96636 238076 96688
rect 238944 96636 238996 96688
rect 240140 96636 240192 96688
rect 240968 96636 241020 96688
rect 242256 96636 242308 96688
rect 242808 96636 242860 96688
rect 248880 96636 248932 96688
rect 249524 96636 249576 96688
rect 259552 96636 259604 96688
rect 260748 96636 260800 96688
rect 261668 96636 261720 96688
rect 262128 96636 262180 96688
rect 264152 96636 264204 96688
rect 267004 96636 267056 96688
rect 269396 96636 269448 96688
rect 270408 96636 270460 96688
rect 274088 96636 274140 96688
rect 274548 96636 274600 96688
rect 275100 96636 275152 96688
rect 275744 96636 275796 96688
rect 276940 96636 276992 96688
rect 277308 96636 277360 96688
rect 277492 96636 277544 96688
rect 278320 96636 278372 96688
rect 278412 96636 278464 96688
rect 278688 96636 278740 96688
rect 280712 96636 280764 96688
rect 281172 96636 281224 96688
rect 281540 96636 281592 96688
rect 282828 96636 282880 96688
rect 282920 96636 282972 96688
rect 284116 96636 284168 96688
rect 284300 96636 284352 96688
rect 296628 96636 296680 96688
rect 296812 96772 296864 96824
rect 297640 96772 297692 96824
rect 298652 96908 298704 96960
rect 299020 96908 299072 96960
rect 298468 96840 298520 96892
rect 299204 96840 299256 96892
rect 298284 96772 298336 96824
rect 299388 96772 299440 96824
rect 301504 96704 301556 96756
rect 302884 96636 302936 96688
rect 176568 96568 176620 96620
rect 220176 96568 220228 96620
rect 254676 96568 254728 96620
rect 320180 96568 320232 96620
rect 161388 96500 161440 96552
rect 208308 96500 208360 96552
rect 257528 96500 257580 96552
rect 336004 96500 336056 96552
rect 183468 96432 183520 96484
rect 231124 96432 231176 96484
rect 271052 96432 271104 96484
rect 271236 96432 271288 96484
rect 284944 96432 284996 96484
rect 461584 96432 461636 96484
rect 179328 96364 179380 96416
rect 230480 96364 230532 96416
rect 284392 96364 284444 96416
rect 468484 96364 468536 96416
rect 173164 96296 173216 96348
rect 229284 96296 229336 96348
rect 231124 96296 231176 96348
rect 235356 96296 235408 96348
rect 283748 96296 283800 96348
rect 472624 96296 472676 96348
rect 169668 96228 169720 96280
rect 228732 96228 228784 96280
rect 281908 96228 281960 96280
rect 479524 96228 479576 96280
rect 165528 96160 165580 96212
rect 228088 96160 228140 96212
rect 283104 96160 283156 96212
rect 475384 96160 475436 96212
rect 133788 96092 133840 96144
rect 211160 96092 211212 96144
rect 282552 96092 282604 96144
rect 483020 96092 483072 96144
rect 131028 96024 131080 96076
rect 222292 96024 222344 96076
rect 285588 96024 285640 96076
rect 500960 96024 501012 96076
rect 54484 95956 54536 96008
rect 208676 95956 208728 96008
rect 245016 95956 245068 96008
rect 267832 95956 267884 96008
rect 286140 95956 286192 96008
rect 502984 95956 503036 96008
rect 17224 95888 17276 95940
rect 202052 95888 202104 95940
rect 228364 95888 228416 95940
rect 237472 95888 237524 95940
rect 248052 95888 248104 95940
rect 284392 95888 284444 95940
rect 294328 95888 294380 95940
rect 295064 95888 295116 95940
rect 295340 95888 295392 95940
rect 512000 95888 512052 95940
rect 186964 95820 187016 95872
rect 231768 95820 231820 95872
rect 253480 95820 253532 95872
rect 313280 95820 313332 95872
rect 191104 95752 191156 95804
rect 232320 95752 232372 95804
rect 251272 95752 251324 95804
rect 302332 95752 302384 95804
rect 197268 95684 197320 95736
rect 233516 95684 233568 95736
rect 251088 95684 251140 95736
rect 299664 95684 299716 95736
rect 200028 95616 200080 95668
rect 234160 95616 234212 95668
rect 263600 95616 263652 95668
rect 299480 95616 299532 95668
rect 194508 95548 194560 95600
rect 213920 95548 213972 95600
rect 249892 95548 249944 95600
rect 299572 95548 299624 95600
rect 287336 95480 287388 95532
rect 295340 95480 295392 95532
rect 235908 95276 235960 95328
rect 240232 95276 240284 95328
rect 210516 95208 210568 95260
rect 210700 95208 210752 95260
rect 238116 95208 238168 95260
rect 239404 95208 239456 95260
rect 171048 95140 171100 95192
rect 229100 95140 229152 95192
rect 261392 95140 261444 95192
rect 358820 95140 358872 95192
rect 162768 95072 162820 95124
rect 227720 95072 227772 95124
rect 295984 95072 296036 95124
rect 465724 95072 465776 95124
rect 147588 95004 147640 95056
rect 212540 95004 212592 95056
rect 293316 95004 293368 95056
rect 485044 95004 485096 95056
rect 159364 94936 159416 94988
rect 226892 94936 226944 94988
rect 288256 94936 288308 94988
rect 489184 94936 489236 94988
rect 155316 94868 155368 94920
rect 226248 94868 226300 94920
rect 286968 94868 287020 94920
rect 507860 94868 507912 94920
rect 144828 94800 144880 94852
rect 224500 94800 224552 94852
rect 230388 94800 230440 94852
rect 237380 94800 237432 94852
rect 292488 94800 292540 94852
rect 519544 94800 519596 94852
rect 137284 94732 137336 94784
rect 223304 94732 223356 94784
rect 290372 94732 290424 94784
rect 529940 94732 529992 94784
rect 128268 94664 128320 94716
rect 221648 94664 221700 94716
rect 234988 94664 235040 94716
rect 235172 94664 235224 94716
rect 291016 94664 291068 94716
rect 532700 94664 532752 94716
rect 121368 94596 121420 94648
rect 220636 94596 220688 94648
rect 232136 94596 232188 94648
rect 232412 94596 232464 94648
rect 101404 94528 101456 94580
rect 212816 94528 212868 94580
rect 212908 94528 212960 94580
rect 213092 94528 213144 94580
rect 216128 94528 216180 94580
rect 216496 94528 216548 94580
rect 216956 94528 217008 94580
rect 217324 94528 217376 94580
rect 218520 94528 218572 94580
rect 218888 94528 218940 94580
rect 219716 94528 219768 94580
rect 220360 94528 220412 94580
rect 220912 94528 220964 94580
rect 221556 94528 221608 94580
rect 228456 94528 228508 94580
rect 236368 94596 236420 94648
rect 291568 94596 291620 94648
rect 536840 94596 536892 94648
rect 234804 94528 234856 94580
rect 235448 94528 235500 94580
rect 236644 94528 236696 94580
rect 237104 94528 237156 94580
rect 239128 94528 239180 94580
rect 239680 94528 239732 94580
rect 240324 94528 240376 94580
rect 240692 94528 240744 94580
rect 278044 94528 278096 94580
rect 278412 94528 278464 94580
rect 292856 94528 292908 94580
rect 543740 94528 543792 94580
rect 29644 94460 29696 94512
rect 199844 94460 199896 94512
rect 200212 94460 200264 94512
rect 200580 94460 200632 94512
rect 201776 94460 201828 94512
rect 202604 94460 202656 94512
rect 204444 94460 204496 94512
rect 205180 94460 205232 94512
rect 212724 94460 212776 94512
rect 213276 94460 213328 94512
rect 217140 94460 217192 94512
rect 217692 94460 217744 94512
rect 221096 94460 221148 94512
rect 221924 94460 221976 94512
rect 232044 94460 232096 94512
rect 232412 94460 232464 94512
rect 241612 94460 241664 94512
rect 242532 94460 242584 94512
rect 243636 94460 243688 94512
rect 244096 94460 244148 94512
rect 247040 94460 247092 94512
rect 264244 94460 264296 94512
rect 278228 94460 278280 94512
rect 278596 94460 278648 94512
rect 297272 94460 297324 94512
rect 565084 94460 565136 94512
rect 173808 94392 173860 94444
rect 229468 94392 229520 94444
rect 255320 94392 255372 94444
rect 324412 94392 324464 94444
rect 188344 94324 188396 94376
rect 231492 94324 231544 94376
rect 252928 94324 252980 94376
rect 309140 94324 309192 94376
rect 200212 94256 200264 94308
rect 201132 94256 201184 94308
rect 198648 94188 198700 94240
rect 233700 94256 233752 94308
rect 252376 94256 252428 94308
rect 306380 94256 306432 94308
rect 212632 94188 212684 94240
rect 213460 94188 213512 94240
rect 218060 94188 218112 94240
rect 218336 94188 218388 94240
rect 263876 94188 263928 94240
rect 316040 94188 316092 94240
rect 199844 94120 199896 94172
rect 203708 94120 203760 94172
rect 212724 94120 212776 94172
rect 213644 94120 213696 94172
rect 251732 94120 251784 94172
rect 302240 94120 302292 94172
rect 170404 93780 170456 93832
rect 166908 93712 166960 93764
rect 228272 93712 228324 93764
rect 228548 93780 228600 93832
rect 234252 93780 234304 93832
rect 257712 93780 257764 93832
rect 338120 93780 338172 93832
rect 228824 93712 228876 93764
rect 262036 93712 262088 93764
rect 362960 93712 363012 93764
rect 160008 93644 160060 93696
rect 226984 93644 227036 93696
rect 266268 93644 266320 93696
rect 382924 93644 382976 93696
rect 153108 93576 153160 93628
rect 225788 93576 225840 93628
rect 270408 93576 270460 93628
rect 407212 93576 407264 93628
rect 145564 93508 145616 93560
rect 224592 93508 224644 93560
rect 277768 93508 277820 93560
rect 454776 93508 454828 93560
rect 142068 93440 142120 93492
rect 222200 93440 222252 93492
rect 293408 93440 293460 93492
rect 543004 93440 543056 93492
rect 136548 93372 136600 93424
rect 219440 93372 219492 93424
rect 295248 93372 295300 93424
rect 554780 93372 554832 93424
rect 135168 93304 135220 93356
rect 222752 93304 222804 93356
rect 295156 93304 295208 93356
rect 557540 93304 557592 93356
rect 61384 93236 61436 93288
rect 209228 93236 209280 93288
rect 296536 93236 296588 93288
rect 561680 93236 561732 93288
rect 36544 93168 36596 93220
rect 204996 93168 205048 93220
rect 246856 93168 246908 93220
rect 257344 93168 257396 93220
rect 298008 93168 298060 93220
rect 572812 93168 572864 93220
rect 15844 93100 15896 93152
rect 201592 93100 201644 93152
rect 243912 93100 243964 93152
rect 255964 93100 256016 93152
rect 299388 93100 299440 93152
rect 575480 93100 575532 93152
rect 177948 93032 178000 93084
rect 230020 93032 230072 93084
rect 257252 93032 257304 93084
rect 333980 93032 334032 93084
rect 180708 92964 180760 93016
rect 230756 92964 230808 93016
rect 256056 92964 256108 93016
rect 331220 92964 331272 93016
rect 184848 92896 184900 92948
rect 231400 92896 231452 92948
rect 256608 92896 256660 92948
rect 327080 92896 327132 92948
rect 195888 92828 195940 92880
rect 233148 92828 233200 92880
rect 229744 92556 229796 92608
rect 236828 92556 236880 92608
rect 231216 92488 231268 92540
rect 235632 92488 235684 92540
rect 175188 92420 175240 92472
rect 229652 92420 229704 92472
rect 238208 92420 238260 92472
rect 239864 92420 239916 92472
rect 263324 92420 263376 92472
rect 364984 92420 365036 92472
rect 169024 92352 169076 92404
rect 228640 92352 228692 92404
rect 263232 92352 263284 92404
rect 369860 92352 369912 92404
rect 164148 92284 164200 92336
rect 227996 92284 228048 92336
rect 264612 92284 264664 92336
rect 374000 92284 374052 92336
rect 156604 92216 156656 92268
rect 226524 92216 226576 92268
rect 268200 92216 268252 92268
rect 380900 92216 380952 92268
rect 148968 92148 149020 92200
rect 223580 92148 223632 92200
rect 265992 92148 266044 92200
rect 385684 92148 385736 92200
rect 137928 92080 137980 92132
rect 223396 92080 223448 92132
rect 267648 92080 267700 92132
rect 396080 92080 396132 92132
rect 128176 92012 128228 92064
rect 221740 92012 221792 92064
rect 275652 92012 275704 92064
rect 428464 92012 428516 92064
rect 84108 91944 84160 91996
rect 214196 91944 214248 91996
rect 250260 91944 250312 91996
rect 251272 91944 251324 91996
rect 274548 91944 274600 91996
rect 432604 91944 432656 91996
rect 70308 91876 70360 91928
rect 211712 91876 211764 91928
rect 276848 91876 276900 91928
rect 446404 91876 446456 91928
rect 66168 91808 66220 91860
rect 211436 91808 211488 91860
rect 279608 91808 279660 91860
rect 464344 91808 464396 91860
rect 45468 91740 45520 91792
rect 204260 91740 204312 91792
rect 224868 91740 224920 91792
rect 238484 91740 238536 91792
rect 246948 91740 247000 91792
rect 264336 91740 264388 91792
rect 289728 91740 289780 91792
rect 520280 91740 520332 91792
rect 182088 91672 182140 91724
rect 230848 91672 230900 91724
rect 260472 91672 260524 91724
rect 356060 91672 356112 91724
rect 254400 91604 254452 91656
rect 317420 91604 317472 91656
rect 177856 90992 177908 91044
rect 230204 90992 230256 91044
rect 260564 90992 260616 91044
rect 353300 90992 353352 91044
rect 161296 90924 161348 90976
rect 227168 90924 227220 90976
rect 271604 90924 271656 90976
rect 406384 90924 406436 90976
rect 153016 90856 153068 90908
rect 225972 90856 226024 90908
rect 278688 90856 278740 90908
rect 457444 90856 457496 90908
rect 143448 90788 143500 90840
rect 224132 90788 224184 90840
rect 282736 90788 282788 90840
rect 471244 90788 471296 90840
rect 139308 90720 139360 90772
rect 223764 90720 223816 90772
rect 282092 90720 282144 90772
rect 481640 90720 481692 90772
rect 116584 90652 116636 90704
rect 219624 90652 219676 90704
rect 283932 90652 283984 90704
rect 490564 90652 490616 90704
rect 105544 90584 105596 90636
rect 216036 90584 216088 90636
rect 285312 90584 285364 90636
rect 493324 90584 493376 90636
rect 86776 90516 86828 90568
rect 214656 90516 214708 90568
rect 286416 90516 286468 90568
rect 500224 90516 500276 90568
rect 73068 90448 73120 90500
rect 212264 90448 212316 90500
rect 287704 90448 287756 90500
rect 511264 90448 511316 90500
rect 68284 90380 68336 90432
rect 208216 90380 208268 90432
rect 290924 90380 290976 90432
rect 529204 90380 529256 90432
rect 18604 90312 18656 90364
rect 202236 90312 202288 90364
rect 248144 90312 248196 90364
rect 282184 90312 282236 90364
rect 296076 90312 296128 90364
rect 556804 90312 556856 90364
rect 254952 90244 255004 90296
rect 321560 90244 321612 90296
rect 253572 90176 253624 90228
rect 310520 90176 310572 90228
rect 252192 90108 252244 90160
rect 303620 90108 303672 90160
rect 267280 89632 267332 89684
rect 389824 89632 389876 89684
rect 268660 89564 268712 89616
rect 398840 89564 398892 89616
rect 297824 89496 297876 89548
rect 467104 89496 467156 89548
rect 157984 89428 158036 89480
rect 226616 89428 226668 89480
rect 281448 89428 281500 89480
rect 472716 89428 472768 89480
rect 122748 89360 122800 89412
rect 221556 89360 221608 89412
rect 285404 89360 285456 89412
rect 497464 89360 497516 89412
rect 119988 89292 120040 89344
rect 220268 89292 220320 89344
rect 286876 89292 286928 89344
rect 504364 89292 504416 89344
rect 108304 89224 108356 89276
rect 214104 89224 214156 89276
rect 286692 89224 286744 89276
rect 506480 89224 506532 89276
rect 53748 89156 53800 89208
rect 199384 89156 199436 89208
rect 292120 89156 292172 89208
rect 518164 89156 518216 89208
rect 47584 89088 47636 89140
rect 205824 89088 205876 89140
rect 288072 89088 288124 89140
rect 515404 89088 515456 89140
rect 43536 89020 43588 89072
rect 207204 89020 207256 89072
rect 289360 89020 289412 89072
rect 522304 89020 522356 89072
rect 40684 88952 40736 89004
rect 205732 88952 205784 89004
rect 293592 88952 293644 89004
rect 547972 88952 548024 89004
rect 257804 88884 257856 88936
rect 331864 88884 331916 88936
rect 256332 88816 256384 88868
rect 323584 88816 323636 88868
rect 256424 88272 256476 88324
rect 328460 88272 328512 88324
rect 257896 88204 257948 88256
rect 335360 88204 335412 88256
rect 261852 88136 261904 88188
rect 357440 88136 357492 88188
rect 263416 88068 263468 88120
rect 367744 88068 367796 88120
rect 124128 88000 124180 88052
rect 221188 88000 221240 88052
rect 270040 88000 270092 88052
rect 409880 88000 409932 88052
rect 117228 87932 117280 87984
rect 219808 87932 219860 87984
rect 272892 87932 272944 87984
rect 420920 87932 420972 87984
rect 75184 87864 75236 87916
rect 211252 87864 211304 87916
rect 294972 87864 295024 87916
rect 536104 87864 536156 87916
rect 57244 87796 57296 87848
rect 209412 87796 209464 87848
rect 292304 87796 292356 87848
rect 538220 87796 538272 87848
rect 53104 87728 53156 87780
rect 206836 87728 206888 87780
rect 292212 87728 292264 87780
rect 540244 87728 540296 87780
rect 46848 87660 46900 87712
rect 203524 87660 203576 87712
rect 295064 87660 295116 87712
rect 547144 87660 547196 87712
rect 14464 87592 14516 87644
rect 201684 87592 201736 87644
rect 296352 87592 296404 87644
rect 560944 87592 560996 87644
rect 253664 87524 253716 87576
rect 313924 87524 313976 87576
rect 307024 86912 307076 86964
rect 580172 86912 580224 86964
rect 257620 86844 257672 86896
rect 339500 86844 339552 86896
rect 261944 86776 261996 86828
rect 360200 86776 360252 86828
rect 261668 86708 261720 86760
rect 363604 86708 363656 86760
rect 264704 86640 264756 86692
rect 374092 86640 374144 86692
rect 268752 86572 268804 86624
rect 402980 86572 403032 86624
rect 107568 86504 107620 86556
rect 191196 86504 191248 86556
rect 271696 86504 271748 86556
rect 416780 86504 416832 86556
rect 90364 86436 90416 86488
rect 215116 86436 215168 86488
rect 277032 86436 277084 86488
rect 425704 86436 425756 86488
rect 79324 86368 79376 86420
rect 208860 86368 208912 86420
rect 278412 86368 278464 86420
rect 453396 86368 453448 86420
rect 76564 86300 76616 86352
rect 211620 86300 211672 86352
rect 297640 86300 297692 86352
rect 566464 86300 566516 86352
rect 35164 86232 35216 86284
rect 201868 86232 201920 86284
rect 248236 86232 248288 86284
rect 261484 86232 261536 86284
rect 296444 86232 296496 86284
rect 565820 86232 565872 86284
rect 255044 86164 255096 86216
rect 316132 86164 316184 86216
rect 3148 85484 3200 85536
rect 151084 85484 151136 85536
rect 253756 85416 253808 85468
rect 307024 85416 307076 85468
rect 263140 85348 263192 85400
rect 332692 85348 332744 85400
rect 267004 85280 267056 85332
rect 375380 85280 375432 85332
rect 264796 85212 264848 85264
rect 378140 85212 378192 85264
rect 272984 85144 273036 85196
rect 423772 85144 423824 85196
rect 278504 85076 278556 85128
rect 459560 85076 459612 85128
rect 282276 85008 282328 85060
rect 463700 85008 463752 85060
rect 284116 84940 284168 84992
rect 485780 84940 485832 84992
rect 284024 84872 284076 84924
rect 490012 84872 490064 84924
rect 5448 84804 5500 84856
rect 198004 84804 198056 84856
rect 290740 84804 290792 84856
rect 530584 84804 530636 84856
rect 255136 83988 255188 84040
rect 318064 83988 318116 84040
rect 256148 83920 256200 83972
rect 324964 83920 325016 83972
rect 261760 83852 261812 83904
rect 360844 83852 360896 83904
rect 268844 83784 268896 83836
rect 395344 83784 395396 83836
rect 282736 83716 282788 83768
rect 477500 83716 477552 83768
rect 283840 83648 283892 83700
rect 492680 83648 492732 83700
rect 285128 83580 285180 83632
rect 496820 83580 496872 83632
rect 290832 83512 290884 83564
rect 528560 83512 528612 83564
rect 293684 83444 293736 83496
rect 542360 83444 542412 83496
rect 271328 82492 271380 82544
rect 365812 82492 365864 82544
rect 271236 82424 271288 82476
rect 382280 82424 382332 82476
rect 270132 82356 270184 82408
rect 392584 82356 392636 82408
rect 276664 82288 276716 82340
rect 400220 82288 400272 82340
rect 288164 82220 288216 82272
rect 510620 82220 510672 82272
rect 293224 82152 293276 82204
rect 546500 82152 546552 82204
rect 294788 82084 294840 82136
rect 553400 82084 553452 82136
rect 301504 80928 301556 80980
rect 404360 80928 404412 80980
rect 274272 80860 274324 80912
rect 429200 80860 429252 80912
rect 274364 80792 274416 80844
rect 431224 80792 431276 80844
rect 275744 80724 275796 80776
rect 440332 80724 440384 80776
rect 297732 80656 297784 80708
rect 571340 80656 571392 80708
rect 302884 79296 302936 79348
rect 447140 79296 447192 79348
rect 309784 73108 309836 73160
rect 579988 73108 580040 73160
rect 2780 71612 2832 71664
rect 4804 71612 4856 71664
rect 454684 60664 454736 60716
rect 580172 60664 580224 60716
rect 3056 59304 3108 59356
rect 146944 59304 146996 59356
rect 3424 45500 3476 45552
rect 148324 45500 148376 45552
rect 322204 37884 322256 37936
rect 478880 37884 478932 37936
rect 312544 35164 312596 35216
rect 425060 35164 425112 35216
rect 254860 33736 254912 33788
rect 322940 33736 322992 33788
rect 323676 33736 323728 33788
rect 456892 33736 456944 33788
rect 3148 33056 3200 33108
rect 155224 33056 155276 33108
rect 305644 33056 305696 33108
rect 580172 33056 580224 33108
rect 256240 31016 256292 31068
rect 329840 31016 329892 31068
rect 253480 29588 253532 29640
rect 311900 29588 311952 29640
rect 294880 28228 294932 28280
rect 556252 28228 556304 28280
rect 33048 26868 33100 26920
rect 202144 26868 202196 26920
rect 292028 26868 292080 26920
rect 539692 26868 539744 26920
rect 296168 25508 296220 25560
rect 564532 25508 564584 25560
rect 199936 24080 199988 24132
rect 233608 24080 233660 24132
rect 282460 24080 282512 24132
rect 481732 24080 481784 24132
rect 234068 23468 234120 23520
rect 238300 23468 238352 23520
rect 233148 22720 233200 22772
rect 239496 22720 239548 22772
rect 246672 22720 246724 22772
rect 267740 22720 267792 22772
rect 293500 22720 293552 22772
rect 548524 22720 548576 22772
rect 286508 21360 286560 21412
rect 506572 21360 506624 21412
rect 3424 20612 3476 20664
rect 144184 20612 144236 20664
rect 453304 20612 453356 20664
rect 580172 20612 580224 20664
rect 252284 19932 252336 19984
rect 300860 19932 300912 19984
rect 287888 18572 287940 18624
rect 517520 18572 517572 18624
rect 262956 17212 263008 17264
rect 284300 17212 284352 17264
rect 285220 17212 285272 17264
rect 499580 17212 499632 17264
rect 259000 15988 259052 16040
rect 340972 15988 341024 16040
rect 299112 15920 299164 15972
rect 575112 15920 575164 15972
rect 245292 15852 245344 15904
rect 253388 15852 253440 15904
rect 299020 15852 299072 15904
rect 578608 15852 578660 15904
rect 289544 14492 289596 14544
rect 521844 14492 521896 14544
rect 64788 14424 64840 14476
rect 196624 14424 196676 14476
rect 289452 14424 289504 14476
rect 525064 14424 525116 14476
rect 273076 13676 273128 13728
rect 428372 13676 428424 13728
rect 274180 13608 274232 13660
rect 432052 13608 432104 13660
rect 274456 13540 274508 13592
rect 435088 13540 435140 13592
rect 275928 13472 275980 13524
rect 439136 13472 439188 13524
rect 275836 13404 275888 13456
rect 442632 13404 442684 13456
rect 277124 13336 277176 13388
rect 445760 13336 445812 13388
rect 277216 13268 277268 13320
rect 449808 13268 449860 13320
rect 276940 13200 276992 13252
rect 453304 13200 453356 13252
rect 279976 13132 280028 13184
rect 467104 13132 467156 13184
rect 119896 13064 119948 13116
rect 219716 13064 219768 13116
rect 253296 13064 253348 13116
rect 259460 13064 259512 13116
rect 281080 13064 281132 13116
rect 470600 13064 470652 13116
rect 112812 12180 112864 12232
rect 218888 12180 218940 12232
rect 110328 12112 110380 12164
rect 218612 12112 218664 12164
rect 259092 12112 259144 12164
rect 342904 12112 342956 12164
rect 106188 12044 106240 12096
rect 218336 12044 218388 12096
rect 259184 12044 259236 12096
rect 346952 12044 347004 12096
rect 103428 11976 103480 12028
rect 216956 11976 217008 12028
rect 263508 11976 263560 12028
rect 367744 11976 367796 12028
rect 99288 11908 99340 11960
rect 216864 11908 216916 11960
rect 266176 11908 266228 11960
rect 382372 11908 382424 11960
rect 31300 11840 31352 11892
rect 204444 11840 204496 11892
rect 266084 11840 266136 11892
rect 385592 11840 385644 11892
rect 28908 11772 28960 11824
rect 204720 11772 204772 11824
rect 267464 11772 267516 11824
rect 389456 11772 389508 11824
rect 23020 11704 23072 11756
rect 203156 11704 203208 11756
rect 267372 11704 267424 11756
rect 392584 11704 392636 11756
rect 423772 11704 423824 11756
rect 424968 11704 425020 11756
rect 332692 11636 332744 11688
rect 333888 11636 333940 11688
rect 374092 11636 374144 11688
rect 375288 11636 375340 11688
rect 95148 10684 95200 10736
rect 216220 10684 216272 10736
rect 92388 10616 92440 10668
rect 215484 10616 215536 10668
rect 87972 10548 88024 10600
rect 214288 10548 214340 10600
rect 81348 10480 81400 10532
rect 212724 10480 212776 10532
rect 78588 10412 78640 10464
rect 212908 10412 212960 10464
rect 74448 10344 74500 10396
rect 213276 10344 213328 10396
rect 246764 10344 246816 10396
rect 251916 10344 251968 10396
rect 60648 10276 60700 10328
rect 210056 10276 210108 10328
rect 220452 10276 220504 10328
rect 233976 10276 234028 10328
rect 250812 10276 250864 10328
rect 298100 10276 298152 10328
rect 299204 10276 299256 10328
rect 576952 10276 577004 10328
rect 111616 9392 111668 9444
rect 218520 9392 218572 9444
rect 108120 9324 108172 9376
rect 218152 9324 218204 9376
rect 104532 9256 104584 9308
rect 217140 9256 217192 9308
rect 101036 9188 101088 9240
rect 217232 9188 217284 9240
rect 97448 9120 97500 9172
rect 216128 9120 216180 9172
rect 93952 9052 94004 9104
rect 215668 9052 215720 9104
rect 281356 9052 281408 9104
rect 469864 9052 469916 9104
rect 79692 8984 79744 9036
rect 212632 8984 212684 9036
rect 226340 8984 226392 9036
rect 233884 8984 233936 9036
rect 281172 8984 281224 9036
rect 473452 8984 473504 9036
rect 76196 8916 76248 8968
rect 213000 8916 213052 8968
rect 281264 8916 281316 8968
rect 476948 8916 477000 8968
rect 222752 8304 222804 8356
rect 231308 8304 231360 8356
rect 265900 8100 265952 8152
rect 388260 8100 388312 8152
rect 267556 8032 267608 8084
rect 391848 8032 391900 8084
rect 267188 7964 267240 8016
rect 395252 7964 395304 8016
rect 268936 7896 268988 7948
rect 398932 7896 398984 7948
rect 269028 7828 269080 7880
rect 402520 7828 402572 7880
rect 270316 7760 270368 7812
rect 406016 7760 406068 7812
rect 192024 7692 192076 7744
rect 232596 7692 232648 7744
rect 270224 7692 270276 7744
rect 409604 7692 409656 7744
rect 24216 7624 24268 7676
rect 94504 7624 94556 7676
rect 145932 7624 145984 7676
rect 224132 7624 224184 7676
rect 269948 7624 270000 7676
rect 413100 7624 413152 7676
rect 43076 7556 43128 7608
rect 188436 7556 188488 7608
rect 188528 7556 188580 7608
rect 232228 7556 232280 7608
rect 253204 7556 253256 7608
rect 266544 7556 266596 7608
rect 273168 7556 273220 7608
rect 427268 7556 427320 7608
rect 99840 6876 99892 6928
rect 104164 6876 104216 6928
rect 3424 6604 3476 6656
rect 7564 6604 7616 6656
rect 215668 6536 215720 6588
rect 236736 6536 236788 6588
rect 249248 6536 249300 6588
rect 284484 6536 284536 6588
rect 205088 6468 205140 6520
rect 234988 6468 235040 6520
rect 250904 6468 250956 6520
rect 297272 6468 297324 6520
rect 194416 6400 194468 6452
rect 232688 6400 232740 6452
rect 259368 6400 259420 6452
rect 342168 6536 342220 6588
rect 190828 6332 190880 6384
rect 232044 6332 232096 6384
rect 259276 6332 259328 6384
rect 345756 6468 345808 6520
rect 341524 6400 341576 6452
rect 379980 6400 380032 6452
rect 14740 6264 14792 6316
rect 124864 6264 124916 6316
rect 187332 6264 187384 6316
rect 232412 6264 232464 6316
rect 260656 6264 260708 6316
rect 352840 6332 352892 6384
rect 352564 6264 352616 6316
rect 394240 6400 394292 6452
rect 388444 6332 388496 6384
rect 418988 6468 419040 6520
rect 393964 6264 394016 6316
rect 422576 6400 422628 6452
rect 418804 6332 418856 6384
rect 443828 6332 443880 6384
rect 71504 6196 71556 6248
rect 62028 6128 62080 6180
rect 208584 6196 208636 6248
rect 234804 6196 234856 6248
rect 249432 6196 249484 6248
rect 287796 6196 287848 6248
rect 287980 6196 288032 6248
rect 514760 6196 514812 6248
rect 209044 6128 209096 6180
rect 212172 6128 212224 6180
rect 236276 6128 236328 6180
rect 249340 6128 249392 6180
rect 291384 6128 291436 6180
rect 291936 6128 291988 6180
rect 536012 6128 536064 6180
rect 210516 6060 210568 6112
rect 124680 5516 124732 5568
rect 126244 5516 126296 5568
rect 245476 5244 245528 5296
rect 265348 5244 265400 5296
rect 304264 5244 304316 5296
rect 358728 5244 358780 5296
rect 249708 5176 249760 5228
rect 290188 5176 290240 5228
rect 309876 5176 309928 5228
rect 372896 5176 372948 5228
rect 35992 5108 36044 5160
rect 50344 5108 50396 5160
rect 58440 5108 58492 5160
rect 39580 5040 39632 5092
rect 58624 5040 58676 5092
rect 131764 5108 131816 5160
rect 222476 5108 222528 5160
rect 245384 5108 245436 5160
rect 261760 5108 261812 5160
rect 262864 5108 262916 5160
rect 355232 5108 355284 5160
rect 377404 5108 377456 5160
rect 411812 5108 411864 5160
rect 411904 5108 411956 5160
rect 436652 5108 436704 5160
rect 443644 5108 443696 5160
rect 472256 5108 472308 5160
rect 209872 5040 209924 5092
rect 246488 5040 246540 5092
rect 268844 5040 268896 5092
rect 271788 5040 271840 5092
rect 415492 5040 415544 5092
rect 436744 5040 436796 5092
rect 465172 5040 465224 5092
rect 47860 4972 47912 5024
rect 207848 4972 207900 5024
rect 221556 4972 221608 5024
rect 237656 4972 237708 5024
rect 251824 4972 251876 5024
rect 279516 4972 279568 5024
rect 286692 4972 286744 5024
rect 504180 4972 504232 5024
rect 2872 4904 2924 4956
rect 200488 4904 200540 4956
rect 218060 4904 218112 4956
rect 236644 4904 236696 4956
rect 249524 4904 249576 4956
rect 286600 4904 286652 4956
rect 289268 4904 289320 4956
rect 519544 4904 519596 4956
rect 1676 4836 1728 4888
rect 200396 4836 200448 4888
rect 214472 4836 214524 4888
rect 236552 4836 236604 4888
rect 249616 4836 249668 4888
rect 288992 4836 289044 4888
rect 289636 4836 289688 4888
rect 523040 4836 523092 4888
rect 572 4768 624 4820
rect 200580 4768 200632 4820
rect 210976 4768 211028 4820
rect 239036 4768 239088 4820
rect 250996 4768 251048 4820
rect 293684 4768 293736 4820
rect 296260 4768 296312 4820
rect 560852 4768 560904 4820
rect 13544 4088 13596 4140
rect 18604 4088 18656 4140
rect 67916 4088 67968 4140
rect 97264 4088 97316 4140
rect 103336 4088 103388 4140
rect 112444 4088 112496 4140
rect 129372 4088 129424 4140
rect 221096 4088 221148 4140
rect 246304 4088 246356 4140
rect 248788 4088 248840 4140
rect 252100 4088 252152 4140
rect 257068 4088 257120 4140
rect 258356 4088 258408 4140
rect 12348 4020 12400 4072
rect 17224 4020 17276 4072
rect 34796 4020 34848 4072
rect 43444 4020 43496 4072
rect 50160 4020 50212 4072
rect 79324 4020 79376 4072
rect 87420 4020 87472 4072
rect 108304 4020 108356 4072
rect 117596 4020 117648 4072
rect 217324 4020 217376 4072
rect 238116 4020 238168 4072
rect 240600 4020 240652 4072
rect 243912 4020 243964 4072
rect 254676 4020 254728 4072
rect 255964 4020 256016 4072
rect 258080 4020 258132 4072
rect 261484 4088 261536 4140
rect 277124 4088 277176 4140
rect 278228 4088 278280 4140
rect 284668 4088 284720 4140
rect 292580 4088 292632 4140
rect 299572 4088 299624 4140
rect 363604 4088 363656 4140
rect 364616 4088 364668 4140
rect 406384 4088 406436 4140
rect 414296 4088 414348 4140
rect 471244 4088 471296 4140
rect 475844 4088 475896 4140
rect 479524 4088 479576 4140
rect 480536 4088 480588 4140
rect 566556 4088 566608 4140
rect 568028 4088 568080 4140
rect 305552 4020 305604 4072
rect 475384 4020 475436 4072
rect 487620 4020 487672 4072
rect 20628 3952 20680 4004
rect 21824 3816 21876 3868
rect 29644 3816 29696 3868
rect 37188 3952 37240 4004
rect 47584 3952 47636 4004
rect 57336 3952 57388 4004
rect 88984 3952 89036 4004
rect 96252 3952 96304 4004
rect 105544 3952 105596 4004
rect 110512 3952 110564 4004
rect 215944 3952 215996 4004
rect 225144 3952 225196 4004
rect 234068 3952 234120 4004
rect 242440 3952 242492 4004
rect 249984 3952 250036 4004
rect 252008 3952 252060 4004
rect 307944 3952 307996 4004
rect 428464 3952 428516 4004
rect 445024 3952 445076 4004
rect 472624 3952 472676 4004
rect 491116 3952 491168 4004
rect 40684 3884 40736 3936
rect 53104 3884 53156 3936
rect 54944 3884 54996 3936
rect 61384 3884 61436 3936
rect 63224 3884 63276 3936
rect 210240 3884 210292 3936
rect 223764 3884 223816 3936
rect 228548 3884 228600 3936
rect 228732 3884 228784 3936
rect 237932 3884 237984 3936
rect 260748 3884 260800 3936
rect 349252 3884 349304 3936
rect 395344 3884 395396 3936
rect 397736 3884 397788 3936
rect 425796 3884 425848 3936
rect 450912 3884 450964 3936
rect 461584 3884 461636 3936
rect 498200 3884 498252 3936
rect 39304 3816 39356 3868
rect 52552 3816 52604 3868
rect 208676 3816 208728 3868
rect 219256 3816 219308 3868
rect 228364 3816 228416 3868
rect 244096 3816 244148 3868
rect 255872 3816 255924 3868
rect 264888 3816 264940 3868
rect 377680 3816 377732 3868
rect 392676 3816 392728 3868
rect 408408 3816 408460 3868
rect 414664 3816 414716 3868
rect 462780 3816 462832 3868
rect 468484 3816 468536 3868
rect 494704 3816 494756 3868
rect 519636 3816 519688 3868
rect 540796 3816 540848 3868
rect 547144 3816 547196 3868
rect 552664 3816 552716 3868
rect 11152 3748 11204 3800
rect 35164 3748 35216 3800
rect 44272 3748 44324 3800
rect 207388 3748 207440 3800
rect 216864 3748 216916 3800
rect 229744 3748 229796 3800
rect 245200 3748 245252 3800
rect 262956 3748 263008 3800
rect 264244 3748 264296 3800
rect 276020 3748 276072 3800
rect 278412 3748 278464 3800
rect 454500 3748 454552 3800
rect 465724 3748 465776 3800
rect 565636 3748 565688 3800
rect 16028 3680 16080 3732
rect 7656 3612 7708 3664
rect 25320 3680 25372 3732
rect 204628 3680 204680 3732
rect 213368 3680 213420 3732
rect 228456 3680 228508 3732
rect 244004 3680 244056 3732
rect 259460 3680 259512 3732
rect 260104 3680 260156 3732
rect 278320 3680 278372 3732
rect 280068 3680 280120 3732
rect 8760 3544 8812 3596
rect 15844 3544 15896 3596
rect 200028 3612 200080 3664
rect 209780 3612 209832 3664
rect 231216 3612 231268 3664
rect 242624 3612 242676 3664
rect 251180 3612 251232 3664
rect 251916 3612 251968 3664
rect 271236 3612 271288 3664
rect 280988 3612 281040 3664
rect 284668 3680 284720 3732
rect 461584 3680 461636 3732
rect 467196 3680 467248 3732
rect 573916 3680 573968 3732
rect 200396 3544 200448 3596
rect 6460 3476 6512 3528
rect 193128 3476 193180 3528
rect 193220 3476 193272 3528
rect 194508 3476 194560 3528
rect 196808 3476 196860 3528
rect 197268 3476 197320 3528
rect 197912 3476 197964 3528
rect 198648 3476 198700 3528
rect 199108 3476 199160 3528
rect 199936 3476 199988 3528
rect 200028 3476 200080 3528
rect 201776 3544 201828 3596
rect 207388 3544 207440 3596
rect 231124 3544 231176 3596
rect 246580 3544 246632 3596
rect 271052 3544 271104 3596
rect 271144 3544 271196 3596
rect 274824 3544 274876 3596
rect 281908 3544 281960 3596
rect 284392 3544 284444 3596
rect 468668 3612 468720 3664
rect 475752 3612 475804 3664
rect 475844 3612 475896 3664
rect 485228 3612 485280 3664
rect 472716 3544 472768 3596
rect 474556 3544 474608 3596
rect 485044 3544 485096 3596
rect 486424 3544 486476 3596
rect 488816 3544 488868 3596
rect 489184 3612 489236 3664
rect 515956 3612 516008 3664
rect 518164 3612 518216 3664
rect 529112 3612 529164 3664
rect 529204 3612 529256 3664
rect 531320 3612 531372 3664
rect 536104 3612 536156 3664
rect 556160 3612 556212 3664
rect 547880 3544 547932 3596
rect 560944 3544 560996 3596
rect 563244 3544 563296 3596
rect 565084 3544 565136 3596
rect 570328 3544 570380 3596
rect 201500 3476 201552 3528
rect 223764 3476 223816 3528
rect 223948 3476 224000 3528
rect 224868 3476 224920 3528
rect 229836 3476 229888 3528
rect 230388 3476 230440 3528
rect 234620 3476 234672 3528
rect 238208 3476 238260 3528
rect 242164 3476 242216 3528
rect 242900 3476 242952 3528
rect 248052 3476 248104 3528
rect 280712 3476 280764 3528
rect 282184 3476 282236 3528
rect 283104 3476 283156 3528
rect 284300 3476 284352 3528
rect 285404 3476 285456 3528
rect 300768 3476 300820 3528
rect 302332 3476 302384 3528
rect 4068 3408 4120 3460
rect 200672 3408 200724 3460
rect 206192 3408 206244 3460
rect 17040 3340 17092 3392
rect 21364 3340 21416 3392
rect 27712 3340 27764 3392
rect 28908 3340 28960 3392
rect 32404 3340 32456 3392
rect 33048 3340 33100 3392
rect 33600 3340 33652 3392
rect 40592 3340 40644 3392
rect 41880 3340 41932 3392
rect 43536 3340 43588 3392
rect 51356 3340 51408 3392
rect 54484 3340 54536 3392
rect 19432 3272 19484 3324
rect 25504 3272 25556 3324
rect 48964 3272 49016 3324
rect 56048 3272 56100 3324
rect 57244 3272 57296 3324
rect 59636 3272 59688 3324
rect 60648 3272 60700 3324
rect 60832 3272 60884 3324
rect 65524 3340 65576 3392
rect 66168 3340 66220 3392
rect 69112 3340 69164 3392
rect 70308 3340 70360 3392
rect 72608 3340 72660 3392
rect 73068 3340 73120 3392
rect 73804 3340 73856 3392
rect 74448 3340 74500 3392
rect 77392 3340 77444 3392
rect 78588 3340 78640 3392
rect 26516 3204 26568 3256
rect 33784 3204 33836 3256
rect 64328 3204 64380 3256
rect 64788 3204 64840 3256
rect 9956 3136 10008 3188
rect 14464 3136 14516 3188
rect 18236 3136 18288 3188
rect 22744 3136 22796 3188
rect 68284 3272 68336 3324
rect 66720 3204 66772 3256
rect 75184 3204 75236 3256
rect 71044 3136 71096 3188
rect 75000 3136 75052 3188
rect 28908 3068 28960 3120
rect 32312 3068 32364 3120
rect 78588 3068 78640 3120
rect 98552 3272 98604 3324
rect 102232 3340 102284 3392
rect 103428 3340 103480 3392
rect 105728 3340 105780 3392
rect 106188 3340 106240 3392
rect 106924 3340 106976 3392
rect 107568 3340 107620 3392
rect 109316 3340 109368 3392
rect 110328 3340 110380 3392
rect 114008 3340 114060 3392
rect 115204 3340 115256 3392
rect 116400 3340 116452 3392
rect 117228 3340 117280 3392
rect 122288 3340 122340 3392
rect 122748 3340 122800 3392
rect 123484 3340 123536 3392
rect 124128 3340 124180 3392
rect 125876 3340 125928 3392
rect 126888 3340 126940 3392
rect 130568 3340 130620 3392
rect 131028 3340 131080 3392
rect 132960 3340 133012 3392
rect 133788 3340 133840 3392
rect 134156 3340 134208 3392
rect 135168 3340 135220 3392
rect 135260 3340 135312 3392
rect 136548 3340 136600 3392
rect 138848 3340 138900 3392
rect 139308 3340 139360 3392
rect 141240 3340 141292 3392
rect 142068 3340 142120 3392
rect 142436 3340 142488 3392
rect 143448 3340 143500 3392
rect 144736 3340 144788 3392
rect 145564 3340 145616 3392
rect 147128 3340 147180 3392
rect 147588 3340 147640 3392
rect 148324 3340 148376 3392
rect 148968 3340 149020 3392
rect 149520 3340 149572 3392
rect 150348 3340 150400 3392
rect 101404 3272 101456 3324
rect 136456 3272 136508 3324
rect 137284 3272 137336 3324
rect 140044 3272 140096 3324
rect 223856 3340 223908 3392
rect 232228 3408 232280 3460
rect 233148 3408 233200 3460
rect 242716 3408 242768 3460
rect 246396 3408 246448 3460
rect 250720 3408 250772 3460
rect 294880 3408 294932 3460
rect 298928 3408 298980 3460
rect 580264 3476 580316 3528
rect 582196 3476 582248 3528
rect 234896 3340 234948 3392
rect 242808 3340 242860 3392
rect 247592 3340 247644 3392
rect 257344 3340 257396 3392
rect 270040 3340 270092 3392
rect 271052 3340 271104 3392
rect 272432 3340 272484 3392
rect 296076 3340 296128 3392
rect 299756 3340 299808 3392
rect 150624 3272 150676 3324
rect 225328 3272 225380 3324
rect 233424 3272 233476 3324
rect 239128 3272 239180 3324
rect 239312 3272 239364 3324
rect 240324 3272 240376 3324
rect 253296 3272 253348 3324
rect 260656 3272 260708 3324
rect 264336 3272 264388 3324
rect 273628 3272 273680 3324
rect 80888 3204 80940 3256
rect 81348 3204 81400 3256
rect 83280 3204 83332 3256
rect 84108 3204 84160 3256
rect 84476 3204 84528 3256
rect 87604 3204 87656 3256
rect 89168 3204 89220 3256
rect 90364 3204 90416 3256
rect 91560 3204 91612 3256
rect 92388 3204 92440 3256
rect 92756 3204 92808 3256
rect 111064 3204 111116 3256
rect 115204 3204 115256 3256
rect 116584 3204 116636 3256
rect 143540 3204 143592 3256
rect 144828 3204 144880 3256
rect 154212 3204 154264 3256
rect 155316 3204 155368 3256
rect 155408 3204 155460 3256
rect 156604 3204 156656 3256
rect 158904 3204 158956 3256
rect 160008 3204 160060 3256
rect 160100 3204 160152 3256
rect 161204 3204 161256 3256
rect 163688 3204 163740 3256
rect 164148 3204 164200 3256
rect 164884 3204 164936 3256
rect 165528 3204 165580 3256
rect 166080 3204 166132 3256
rect 166908 3204 166960 3256
rect 167184 3204 167236 3256
rect 169024 3204 169076 3256
rect 173164 3204 173216 3256
rect 173808 3204 173860 3256
rect 174268 3204 174320 3256
rect 175188 3204 175240 3256
rect 175464 3204 175516 3256
rect 176568 3204 176620 3256
rect 176660 3204 176712 3256
rect 177948 3204 178000 3256
rect 180248 3204 180300 3256
rect 180708 3204 180760 3256
rect 181444 3204 181496 3256
rect 182088 3204 182140 3256
rect 182548 3204 182600 3256
rect 183468 3204 183520 3256
rect 183744 3204 183796 3256
rect 184848 3204 184900 3256
rect 186136 3204 186188 3256
rect 186964 3204 187016 3256
rect 189724 3204 189776 3256
rect 191104 3204 191156 3256
rect 193128 3204 193180 3256
rect 200764 3204 200816 3256
rect 299296 3204 299348 3256
rect 307024 3340 307076 3392
rect 309048 3340 309100 3392
rect 313924 3340 313976 3392
rect 315028 3340 315080 3392
rect 316040 3340 316092 3392
rect 317328 3340 317380 3392
rect 318156 3340 318208 3392
rect 319720 3340 319772 3392
rect 323584 3340 323636 3392
rect 325608 3340 325660 3392
rect 331864 3340 331916 3392
rect 332692 3340 332744 3392
rect 336004 3340 336056 3392
rect 337476 3340 337528 3392
rect 342996 3340 343048 3392
rect 344560 3340 344612 3392
rect 345664 3340 345716 3392
rect 348056 3340 348108 3392
rect 348424 3340 348476 3392
rect 351644 3340 351696 3392
rect 364984 3340 365036 3392
rect 367008 3340 367060 3392
rect 367836 3340 367888 3392
rect 369400 3340 369452 3392
rect 382280 3340 382332 3392
rect 383568 3340 383620 3392
rect 389824 3340 389876 3392
rect 390652 3340 390704 3392
rect 398840 3340 398892 3392
rect 400128 3340 400180 3392
rect 432604 3340 432656 3392
rect 434444 3340 434496 3392
rect 435364 3340 435416 3392
rect 437940 3340 437992 3392
rect 439504 3340 439556 3392
rect 441528 3340 441580 3392
rect 454776 3340 454828 3392
rect 455696 3340 455748 3392
rect 457444 3340 457496 3392
rect 459192 3340 459244 3392
rect 490564 3340 490616 3392
rect 492312 3340 492364 3392
rect 497464 3340 497516 3392
rect 499396 3340 499448 3392
rect 502984 3340 503036 3392
rect 505376 3340 505428 3392
rect 515404 3340 515456 3392
rect 517152 3340 517204 3392
rect 522304 3340 522356 3392
rect 524236 3340 524288 3392
rect 530584 3340 530636 3392
rect 532516 3340 532568 3392
rect 540244 3340 540296 3392
rect 541992 3340 542044 3392
rect 581000 3408 581052 3460
rect 583392 3340 583444 3392
rect 347044 3272 347096 3324
rect 350448 3272 350500 3324
rect 421564 3272 421616 3324
rect 423772 3272 423824 3324
rect 431224 3272 431276 3324
rect 433248 3272 433300 3324
rect 453396 3272 453448 3324
rect 456892 3272 456944 3324
rect 529112 3272 529164 3324
rect 534908 3272 534960 3324
rect 548524 3272 548576 3324
rect 550272 3272 550324 3324
rect 382924 3204 382976 3256
rect 384764 3204 384816 3256
rect 500316 3204 500368 3256
rect 502984 3204 503036 3256
rect 556804 3204 556856 3256
rect 559748 3204 559800 3256
rect 82084 3136 82136 3188
rect 87420 3136 87472 3188
rect 98644 3136 98696 3188
rect 99288 3136 99340 3188
rect 151820 3136 151872 3188
rect 153108 3136 153160 3188
rect 157800 3136 157852 3188
rect 159364 3136 159416 3188
rect 169576 3136 169628 3188
rect 170404 3136 170456 3188
rect 231032 3136 231084 3188
rect 238024 3136 238076 3188
rect 385684 3136 385736 3188
rect 387156 3136 387208 3188
rect 413284 3136 413336 3188
rect 416688 3136 416740 3188
rect 85672 3068 85724 3120
rect 86868 3068 86920 3120
rect 90364 3068 90416 3120
rect 93124 3068 93176 3120
rect 156604 3068 156656 3120
rect 157984 3068 158036 3120
rect 168380 3068 168432 3120
rect 169668 3068 169720 3120
rect 171968 3068 172020 3120
rect 173072 3068 173124 3120
rect 324964 3068 325016 3120
rect 326804 3068 326856 3120
rect 360844 3068 360896 3120
rect 362316 3068 362368 3120
rect 237012 3000 237064 3052
rect 241060 3000 241112 3052
rect 264152 3000 264204 3052
rect 267832 3000 267884 3052
rect 511264 3000 511316 3052
rect 513564 3000 513616 3052
rect 30104 2932 30156 2984
rect 36544 2932 36596 2984
rect 126980 2932 127032 2984
rect 128268 2932 128320 2984
rect 446404 2932 446456 2984
rect 452108 2932 452160 2984
rect 464344 2932 464396 2984
rect 466276 2932 466328 2984
rect 493324 2932 493376 2984
rect 495900 2932 495952 2984
rect 504364 2932 504416 2984
rect 510068 2932 510120 2984
rect 543004 2932 543056 2984
rect 545488 2932 545540 2984
rect 70308 2864 70360 2916
rect 76564 2864 76616 2916
rect 118792 2864 118844 2916
rect 119988 2864 120040 2916
rect 184940 2864 184992 2916
rect 188344 2864 188396 2916
rect 242532 2864 242584 2916
rect 244096 2864 244148 2916
rect 369124 2864 369176 2916
rect 371700 2864 371752 2916
rect 417516 2864 417568 2916
rect 420184 2864 420236 2916
rect 525156 2864 525208 2916
rect 527824 2864 527876 2916
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429212 703582 429700 703610
rect 8128 700398 8156 703520
rect 24320 700466 24348 703520
rect 40512 700534 40540 703520
rect 72988 700602 73016 703520
rect 89180 700670 89208 703520
rect 89168 700664 89220 700670
rect 89168 700606 89220 700612
rect 72976 700596 73028 700602
rect 72976 700538 73028 700544
rect 40500 700528 40552 700534
rect 40500 700470 40552 700476
rect 41328 700528 41380 700534
rect 41328 700470 41380 700476
rect 24308 700460 24360 700466
rect 24308 700402 24360 700408
rect 8116 700392 8168 700398
rect 8116 700334 8168 700340
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 3436 683262 3464 684247
rect 3424 683256 3476 683262
rect 3424 683198 3476 683204
rect 3422 671256 3478 671265
rect 3422 671191 3478 671200
rect 3436 670818 3464 671191
rect 3424 670812 3476 670818
rect 3424 670754 3476 670760
rect 3422 658200 3478 658209
rect 3422 658135 3478 658144
rect 3436 656946 3464 658135
rect 3424 656940 3476 656946
rect 3424 656882 3476 656888
rect 3424 632120 3476 632126
rect 3422 632088 3424 632097
rect 3476 632088 3478 632097
rect 3422 632023 3478 632032
rect 3146 619168 3202 619177
rect 3146 619103 3202 619112
rect 3160 618322 3188 619103
rect 3148 618316 3200 618322
rect 3148 618258 3200 618264
rect 3238 606112 3294 606121
rect 3238 606047 3294 606056
rect 3252 605878 3280 606047
rect 3240 605872 3292 605878
rect 3240 605814 3292 605820
rect 3330 580000 3386 580009
rect 3330 579935 3386 579944
rect 3344 579698 3372 579935
rect 3332 579692 3384 579698
rect 3332 579634 3384 579640
rect 3422 566944 3478 566953
rect 3422 566879 3478 566888
rect 3436 565894 3464 566879
rect 3424 565888 3476 565894
rect 3424 565830 3476 565836
rect 3422 553888 3478 553897
rect 3422 553823 3478 553832
rect 3436 553450 3464 553823
rect 3424 553444 3476 553450
rect 3424 553386 3476 553392
rect 3422 527912 3478 527921
rect 3422 527847 3478 527856
rect 3436 527202 3464 527847
rect 3424 527196 3476 527202
rect 3424 527138 3476 527144
rect 3422 514856 3478 514865
rect 3422 514791 3424 514800
rect 3476 514791 3478 514800
rect 3424 514762 3476 514768
rect 3054 501800 3110 501809
rect 3054 501735 3110 501744
rect 3068 501022 3096 501735
rect 3056 501016 3108 501022
rect 3056 500958 3108 500964
rect 3422 475688 3478 475697
rect 3422 475623 3478 475632
rect 3436 474774 3464 475623
rect 3424 474768 3476 474774
rect 3424 474710 3476 474716
rect 3238 462632 3294 462641
rect 3238 462567 3294 462576
rect 3252 462398 3280 462567
rect 3240 462392 3292 462398
rect 3240 462334 3292 462340
rect 3146 449576 3202 449585
rect 3146 449511 3202 449520
rect 3160 448594 3188 449511
rect 3148 448588 3200 448594
rect 3148 448530 3200 448536
rect 3422 423600 3478 423609
rect 3422 423535 3478 423544
rect 3436 422346 3464 423535
rect 3424 422340 3476 422346
rect 3424 422282 3476 422288
rect 3146 410544 3202 410553
rect 3146 410479 3202 410488
rect 3160 409902 3188 410479
rect 3148 409896 3200 409902
rect 3148 409838 3200 409844
rect 3424 397520 3476 397526
rect 3422 397488 3424 397497
rect 3476 397488 3478 397497
rect 3422 397423 3478 397432
rect 3422 371376 3478 371385
rect 3422 371311 3478 371320
rect 3436 371278 3464 371311
rect 3424 371272 3476 371278
rect 3424 371214 3476 371220
rect 3146 358456 3202 358465
rect 3146 358391 3202 358400
rect 3160 357474 3188 358391
rect 3148 357468 3200 357474
rect 3148 357410 3200 357416
rect 3330 345400 3386 345409
rect 3330 345335 3386 345344
rect 3344 345098 3372 345335
rect 3332 345092 3384 345098
rect 3332 345034 3384 345040
rect 3422 319288 3478 319297
rect 3422 319223 3478 319232
rect 3436 318850 3464 319223
rect 3424 318844 3476 318850
rect 3424 318786 3476 318792
rect 3238 306232 3294 306241
rect 3238 306167 3294 306176
rect 3252 305046 3280 306167
rect 41340 305726 41368 700470
rect 105464 699718 105492 703520
rect 137848 700806 137876 703520
rect 154132 700874 154160 703520
rect 154120 700868 154172 700874
rect 154120 700810 154172 700816
rect 137836 700800 137888 700806
rect 137836 700742 137888 700748
rect 170324 699718 170352 703520
rect 105452 699712 105504 699718
rect 105452 699654 105504 699660
rect 106188 699712 106240 699718
rect 106188 699654 106240 699660
rect 170312 699712 170364 699718
rect 170312 699654 170364 699660
rect 171048 699712 171100 699718
rect 171048 699654 171100 699660
rect 41328 305720 41380 305726
rect 41328 305662 41380 305668
rect 3240 305040 3292 305046
rect 3240 304982 3292 304988
rect 106200 304570 106228 699654
rect 171060 304638 171088 699654
rect 198556 337408 198608 337414
rect 198556 337350 198608 337356
rect 171048 304632 171100 304638
rect 171048 304574 171100 304580
rect 106188 304564 106240 304570
rect 106188 304506 106240 304512
rect 177396 302932 177448 302938
rect 177396 302874 177448 302880
rect 14464 302320 14516 302326
rect 14464 302262 14516 302268
rect 11704 302252 11756 302258
rect 11704 302194 11756 302200
rect 7564 301028 7616 301034
rect 7564 300970 7616 300976
rect 4804 299532 4856 299538
rect 4804 299474 4856 299480
rect 3516 298444 3568 298450
rect 3516 298386 3568 298392
rect 3424 298308 3476 298314
rect 3424 298250 3476 298256
rect 2872 293956 2924 293962
rect 2872 293898 2924 293904
rect 2884 293185 2912 293898
rect 2870 293176 2926 293185
rect 2870 293111 2926 293120
rect 3240 267708 3292 267714
rect 3240 267650 3292 267656
rect 3252 267209 3280 267650
rect 3238 267200 3294 267209
rect 3238 267135 3294 267144
rect 3332 215280 3384 215286
rect 3332 215222 3384 215228
rect 3344 214985 3372 215222
rect 3330 214976 3386 214985
rect 3330 214911 3386 214920
rect 3056 202836 3108 202842
rect 3056 202778 3108 202784
rect 3068 201929 3096 202778
rect 3054 201920 3110 201929
rect 3054 201855 3110 201864
rect 3436 188873 3464 298250
rect 3528 241097 3556 298386
rect 3608 298376 3660 298382
rect 3608 298318 3660 298324
rect 3620 254153 3648 298318
rect 3606 254144 3662 254153
rect 3606 254079 3662 254088
rect 3514 241088 3570 241097
rect 3514 241023 3570 241032
rect 3422 188864 3478 188873
rect 3422 188799 3478 188808
rect 3240 164212 3292 164218
rect 3240 164154 3292 164160
rect 3252 162897 3280 164154
rect 3238 162888 3294 162897
rect 3238 162823 3294 162832
rect 3424 150408 3476 150414
rect 3424 150350 3476 150356
rect 3436 149841 3464 150350
rect 3422 149832 3478 149841
rect 3422 149767 3478 149776
rect 3240 137964 3292 137970
rect 3240 137906 3292 137912
rect 3252 136785 3280 137906
rect 3238 136776 3294 136785
rect 3238 136711 3294 136720
rect 3424 111784 3476 111790
rect 3424 111726 3476 111732
rect 3436 110673 3464 111726
rect 3422 110664 3478 110673
rect 3422 110599 3478 110608
rect 3424 97980 3476 97986
rect 3424 97922 3476 97928
rect 3436 97617 3464 97922
rect 3422 97608 3478 97617
rect 3422 97543 3478 97552
rect 3148 85536 3200 85542
rect 3148 85478 3200 85484
rect 3160 84697 3188 85478
rect 3146 84688 3202 84697
rect 3146 84623 3202 84632
rect 4816 71670 4844 299474
rect 5448 84856 5500 84862
rect 5448 84798 5500 84804
rect 2780 71664 2832 71670
rect 2778 71632 2780 71641
rect 4804 71664 4856 71670
rect 2832 71632 2834 71641
rect 4804 71606 4856 71612
rect 2778 71567 2834 71576
rect 3056 59356 3108 59362
rect 3056 59298 3108 59304
rect 3068 58585 3096 59298
rect 3054 58576 3110 58585
rect 3054 58511 3110 58520
rect 3424 45552 3476 45558
rect 3422 45520 3424 45529
rect 3476 45520 3478 45529
rect 3422 45455 3478 45464
rect 3148 33108 3200 33114
rect 3148 33050 3200 33056
rect 3160 32473 3188 33050
rect 3146 32464 3202 32473
rect 3146 32399 3202 32408
rect 3424 20664 3476 20670
rect 3424 20606 3476 20612
rect 3436 19417 3464 20606
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 5460 6914 5488 84798
rect 5276 6886 5488 6914
rect 3424 6656 3476 6662
rect 3424 6598 3476 6604
rect 3436 6497 3464 6598
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 2872 4956 2924 4962
rect 2872 4898 2924 4904
rect 1676 4888 1728 4894
rect 1676 4830 1728 4836
rect 572 4820 624 4826
rect 572 4762 624 4768
rect 584 480 612 4762
rect 1688 480 1716 4830
rect 2884 480 2912 4898
rect 4068 3460 4120 3466
rect 4068 3402 4120 3408
rect 4080 480 4108 3402
rect 5276 480 5304 6886
rect 7576 6662 7604 300970
rect 11716 150414 11744 302194
rect 11704 150408 11756 150414
rect 11704 150350 11756 150356
rect 14476 97986 14504 302262
rect 159364 301368 159416 301374
rect 159364 301310 159416 301316
rect 151084 301300 151136 301306
rect 151084 301242 151136 301248
rect 146944 301232 146996 301238
rect 146944 301174 146996 301180
rect 17224 301096 17276 301102
rect 17224 301038 17276 301044
rect 17236 267714 17264 301038
rect 144184 299804 144236 299810
rect 144184 299746 144236 299752
rect 17224 267708 17276 267714
rect 17224 267650 17276 267656
rect 112444 99340 112496 99346
rect 112444 99282 112496 99288
rect 98644 99272 98696 99278
rect 98644 99214 98696 99220
rect 97264 99204 97316 99210
rect 97264 99146 97316 99152
rect 88984 99136 89036 99142
rect 88984 99078 89036 99084
rect 87604 99000 87656 99006
rect 87604 98942 87656 98948
rect 71044 98932 71096 98938
rect 71044 98874 71096 98880
rect 43444 98864 43496 98870
rect 43444 98806 43496 98812
rect 22744 98796 22796 98802
rect 22744 98738 22796 98744
rect 21364 98660 21416 98666
rect 21364 98602 21416 98608
rect 14464 97980 14516 97986
rect 14464 97922 14516 97928
rect 17224 95940 17276 95946
rect 17224 95882 17276 95888
rect 15844 93152 15896 93158
rect 15844 93094 15896 93100
rect 14464 87644 14516 87650
rect 14464 87586 14516 87592
rect 7564 6656 7616 6662
rect 7564 6598 7616 6604
rect 13544 4140 13596 4146
rect 13544 4082 13596 4088
rect 12348 4072 12400 4078
rect 12348 4014 12400 4020
rect 11152 3800 11204 3806
rect 11152 3742 11204 3748
rect 7656 3664 7708 3670
rect 7656 3606 7708 3612
rect 6460 3528 6512 3534
rect 6460 3470 6512 3476
rect 6472 480 6500 3470
rect 7668 480 7696 3606
rect 8760 3596 8812 3602
rect 8760 3538 8812 3544
rect 8772 480 8800 3538
rect 9956 3188 10008 3194
rect 9956 3130 10008 3136
rect 9968 480 9996 3130
rect 11164 480 11192 3742
rect 12360 480 12388 4014
rect 13556 480 13584 4082
rect 14476 3194 14504 87586
rect 14740 6316 14792 6322
rect 14740 6258 14792 6264
rect 14464 3188 14516 3194
rect 14464 3130 14516 3136
rect 14752 480 14780 6258
rect 15856 3602 15884 93094
rect 17236 4078 17264 95882
rect 18604 90364 18656 90370
rect 18604 90306 18656 90312
rect 18616 4146 18644 90306
rect 18604 4140 18656 4146
rect 18604 4082 18656 4088
rect 17224 4072 17276 4078
rect 17224 4014 17276 4020
rect 20628 4004 20680 4010
rect 20628 3946 20680 3952
rect 16028 3732 16080 3738
rect 16028 3674 16080 3680
rect 15844 3596 15896 3602
rect 15844 3538 15896 3544
rect 16040 1850 16068 3674
rect 17040 3392 17092 3398
rect 17040 3334 17092 3340
rect 15948 1822 16068 1850
rect 15948 480 15976 1822
rect 17052 480 17080 3334
rect 19432 3324 19484 3330
rect 19432 3266 19484 3272
rect 18236 3188 18288 3194
rect 18236 3130 18288 3136
rect 18248 480 18276 3130
rect 19444 480 19472 3266
rect 20640 480 20668 3946
rect 21376 3398 21404 98602
rect 21824 3868 21876 3874
rect 21824 3810 21876 3816
rect 21364 3392 21416 3398
rect 21364 3334 21416 3340
rect 21836 480 21864 3810
rect 22756 3194 22784 98738
rect 33784 98728 33836 98734
rect 33784 98670 33836 98676
rect 25504 97300 25556 97306
rect 25504 97242 25556 97248
rect 23020 11756 23072 11762
rect 23020 11698 23072 11704
rect 22744 3188 22796 3194
rect 22744 3130 22796 3136
rect 23032 480 23060 11698
rect 24216 7676 24268 7682
rect 24216 7618 24268 7624
rect 24228 480 24256 7618
rect 25320 3732 25372 3738
rect 25320 3674 25372 3680
rect 25332 480 25360 3674
rect 25516 3330 25544 97242
rect 32402 97200 32458 97209
rect 32402 97135 32458 97144
rect 29644 94512 29696 94518
rect 29644 94454 29696 94460
rect 28908 11824 28960 11830
rect 28908 11766 28960 11772
rect 28920 3398 28948 11766
rect 29656 3874 29684 94454
rect 31300 11892 31352 11898
rect 31300 11834 31352 11840
rect 29644 3868 29696 3874
rect 29644 3810 29696 3816
rect 27712 3392 27764 3398
rect 27712 3334 27764 3340
rect 28908 3392 28960 3398
rect 28908 3334 28960 3340
rect 25504 3324 25556 3330
rect 25504 3266 25556 3272
rect 26516 3256 26568 3262
rect 26516 3198 26568 3204
rect 26528 480 26556 3198
rect 27724 480 27752 3334
rect 28908 3120 28960 3126
rect 28908 3062 28960 3068
rect 28920 480 28948 3062
rect 30104 2984 30156 2990
rect 30104 2926 30156 2932
rect 30116 480 30144 2926
rect 31312 480 31340 11834
rect 32416 6914 32444 97135
rect 33048 26920 33100 26926
rect 33048 26862 33100 26868
rect 32324 6886 32444 6914
rect 32324 3126 32352 6886
rect 33060 3398 33088 26862
rect 32404 3392 32456 3398
rect 32404 3334 32456 3340
rect 33048 3392 33100 3398
rect 33048 3334 33100 3340
rect 33600 3392 33652 3398
rect 33600 3334 33652 3340
rect 32312 3120 32364 3126
rect 32312 3062 32364 3068
rect 32416 480 32444 3334
rect 33612 480 33640 3334
rect 33796 3262 33824 98670
rect 39302 97472 39358 97481
rect 39302 97407 39358 97416
rect 38566 97336 38622 97345
rect 38566 97271 38622 97280
rect 36544 93220 36596 93226
rect 36544 93162 36596 93168
rect 35164 86284 35216 86290
rect 35164 86226 35216 86232
rect 34796 4072 34848 4078
rect 34796 4014 34848 4020
rect 33784 3256 33836 3262
rect 33784 3198 33836 3204
rect 34808 480 34836 4014
rect 35176 3806 35204 86226
rect 35992 5160 36044 5166
rect 35992 5102 36044 5108
rect 35164 3800 35216 3806
rect 35164 3742 35216 3748
rect 36004 480 36032 5102
rect 36556 2990 36584 93162
rect 38580 6914 38608 97271
rect 38396 6886 38608 6914
rect 37188 4004 37240 4010
rect 37188 3946 37240 3952
rect 36544 2984 36596 2990
rect 36544 2926 36596 2932
rect 37200 480 37228 3946
rect 38396 480 38424 6886
rect 39316 3874 39344 97407
rect 40684 89004 40736 89010
rect 40684 88946 40736 88952
rect 40696 6914 40724 88946
rect 43076 7608 43128 7614
rect 43076 7550 43128 7556
rect 40604 6886 40724 6914
rect 39580 5092 39632 5098
rect 39580 5034 39632 5040
rect 39304 3868 39356 3874
rect 39304 3810 39356 3816
rect 39592 480 39620 5034
rect 40604 3398 40632 6886
rect 40684 3936 40736 3942
rect 40684 3878 40736 3884
rect 40592 3392 40644 3398
rect 40592 3334 40644 3340
rect 40696 480 40724 3878
rect 41880 3392 41932 3398
rect 41880 3334 41932 3340
rect 41892 480 41920 3334
rect 43088 480 43116 7550
rect 43456 4078 43484 98806
rect 50342 97608 50398 97617
rect 50342 97543 50398 97552
rect 45468 91792 45520 91798
rect 45468 91734 45520 91740
rect 43536 89072 43588 89078
rect 43536 89014 43588 89020
rect 43444 4072 43496 4078
rect 43444 4014 43496 4020
rect 43548 3398 43576 89014
rect 44272 3800 44324 3806
rect 44272 3742 44324 3748
rect 43536 3392 43588 3398
rect 43536 3334 43588 3340
rect 44284 480 44312 3742
rect 45480 480 45508 91734
rect 47584 89140 47636 89146
rect 47584 89082 47636 89088
rect 46848 87712 46900 87718
rect 46848 87654 46900 87660
rect 46860 6914 46888 87654
rect 46676 6886 46888 6914
rect 46676 480 46704 6886
rect 47596 4010 47624 89082
rect 50356 5166 50384 97543
rect 58624 97368 58676 97374
rect 58624 97310 58676 97316
rect 54484 96008 54536 96014
rect 54484 95950 54536 95956
rect 53748 89208 53800 89214
rect 53748 89150 53800 89156
rect 53104 87780 53156 87786
rect 53104 87722 53156 87728
rect 50344 5160 50396 5166
rect 50344 5102 50396 5108
rect 47860 5024 47912 5030
rect 47860 4966 47912 4972
rect 47584 4004 47636 4010
rect 47584 3946 47636 3952
rect 47872 480 47900 4966
rect 50160 4072 50212 4078
rect 50160 4014 50212 4020
rect 48964 3324 49016 3330
rect 48964 3266 49016 3272
rect 48976 480 49004 3266
rect 50172 480 50200 4014
rect 53116 3942 53144 87722
rect 53104 3936 53156 3942
rect 53104 3878 53156 3884
rect 52552 3868 52604 3874
rect 52552 3810 52604 3816
rect 51356 3392 51408 3398
rect 51356 3334 51408 3340
rect 51368 480 51396 3334
rect 52564 480 52592 3810
rect 53760 480 53788 89150
rect 54496 3398 54524 95950
rect 57244 87848 57296 87854
rect 57244 87790 57296 87796
rect 54944 3936 54996 3942
rect 54944 3878 54996 3884
rect 54484 3392 54536 3398
rect 54484 3334 54536 3340
rect 54956 480 54984 3878
rect 57256 3330 57284 87790
rect 58440 5160 58492 5166
rect 58440 5102 58492 5108
rect 57336 4004 57388 4010
rect 57336 3946 57388 3952
rect 56048 3324 56100 3330
rect 56048 3266 56100 3272
rect 57244 3324 57296 3330
rect 57244 3266 57296 3272
rect 56060 480 56088 3266
rect 57348 1986 57376 3946
rect 57256 1958 57376 1986
rect 57256 480 57284 1958
rect 58452 480 58480 5102
rect 58636 5098 58664 97310
rect 61384 93288 61436 93294
rect 61384 93230 61436 93236
rect 60648 10328 60700 10334
rect 60648 10270 60700 10276
rect 58624 5092 58676 5098
rect 58624 5034 58676 5040
rect 60660 3330 60688 10270
rect 61396 3942 61424 93230
rect 70308 91928 70360 91934
rect 70308 91870 70360 91876
rect 66168 91860 66220 91866
rect 66168 91802 66220 91808
rect 64788 14476 64840 14482
rect 64788 14418 64840 14424
rect 62028 6180 62080 6186
rect 62028 6122 62080 6128
rect 61384 3936 61436 3942
rect 61384 3878 61436 3884
rect 59636 3324 59688 3330
rect 59636 3266 59688 3272
rect 60648 3324 60700 3330
rect 60648 3266 60700 3272
rect 60832 3324 60884 3330
rect 60832 3266 60884 3272
rect 59648 480 59676 3266
rect 60844 480 60872 3266
rect 62040 480 62068 6122
rect 63224 3936 63276 3942
rect 63224 3878 63276 3884
rect 63236 480 63264 3878
rect 64800 3262 64828 14418
rect 66180 3398 66208 91802
rect 68284 90432 68336 90438
rect 68284 90374 68336 90380
rect 67916 4140 67968 4146
rect 67916 4082 67968 4088
rect 65524 3392 65576 3398
rect 65524 3334 65576 3340
rect 66168 3392 66220 3398
rect 66168 3334 66220 3340
rect 64328 3256 64380 3262
rect 64328 3198 64380 3204
rect 64788 3256 64840 3262
rect 64788 3198 64840 3204
rect 64340 480 64368 3198
rect 65536 480 65564 3334
rect 66720 3256 66772 3262
rect 66720 3198 66772 3204
rect 66732 480 66760 3198
rect 67928 480 67956 4082
rect 68296 3330 68324 90374
rect 70320 3398 70348 91870
rect 69112 3392 69164 3398
rect 69112 3334 69164 3340
rect 70308 3392 70360 3398
rect 70308 3334 70360 3340
rect 68284 3324 68336 3330
rect 68284 3266 68336 3272
rect 69124 480 69152 3334
rect 71056 3194 71084 98874
rect 86868 96824 86920 96830
rect 86868 96766 86920 96772
rect 84108 91996 84160 92002
rect 84108 91938 84160 91944
rect 73068 90500 73120 90506
rect 73068 90442 73120 90448
rect 71504 6248 71556 6254
rect 71504 6190 71556 6196
rect 71044 3188 71096 3194
rect 71044 3130 71096 3136
rect 70308 2916 70360 2922
rect 70308 2858 70360 2864
rect 70320 480 70348 2858
rect 71516 480 71544 6190
rect 73080 3398 73108 90442
rect 75184 87916 75236 87922
rect 75184 87858 75236 87864
rect 74448 10396 74500 10402
rect 74448 10338 74500 10344
rect 74460 3398 74488 10338
rect 72608 3392 72660 3398
rect 72608 3334 72660 3340
rect 73068 3392 73120 3398
rect 73068 3334 73120 3340
rect 73804 3392 73856 3398
rect 73804 3334 73856 3340
rect 74448 3392 74500 3398
rect 74448 3334 74500 3340
rect 72620 480 72648 3334
rect 73816 480 73844 3334
rect 75196 3262 75224 87858
rect 79324 86420 79376 86426
rect 79324 86362 79376 86368
rect 76564 86352 76616 86358
rect 76564 86294 76616 86300
rect 76196 8968 76248 8974
rect 76196 8910 76248 8916
rect 75184 3256 75236 3262
rect 75184 3198 75236 3204
rect 75000 3188 75052 3194
rect 75000 3130 75052 3136
rect 75012 480 75040 3130
rect 76208 480 76236 8910
rect 76576 2922 76604 86294
rect 78588 10464 78640 10470
rect 78588 10406 78640 10412
rect 78600 3398 78628 10406
rect 79336 4078 79364 86362
rect 81348 10532 81400 10538
rect 81348 10474 81400 10480
rect 79692 9036 79744 9042
rect 79692 8978 79744 8984
rect 79324 4072 79376 4078
rect 79324 4014 79376 4020
rect 77392 3392 77444 3398
rect 77392 3334 77444 3340
rect 78588 3392 78640 3398
rect 78588 3334 78640 3340
rect 76564 2916 76616 2922
rect 76564 2858 76616 2864
rect 77404 480 77432 3334
rect 78588 3120 78640 3126
rect 78588 3062 78640 3068
rect 78600 480 78628 3062
rect 79704 480 79732 8978
rect 81360 3262 81388 10474
rect 84120 3262 84148 91938
rect 86776 90568 86828 90574
rect 86776 90510 86828 90516
rect 80888 3256 80940 3262
rect 80888 3198 80940 3204
rect 81348 3256 81400 3262
rect 81348 3198 81400 3204
rect 83280 3256 83332 3262
rect 83280 3198 83332 3204
rect 84108 3256 84160 3262
rect 84108 3198 84160 3204
rect 84476 3256 84528 3262
rect 84476 3198 84528 3204
rect 80900 480 80928 3198
rect 82084 3188 82136 3194
rect 82084 3130 82136 3136
rect 82096 480 82124 3130
rect 83292 480 83320 3198
rect 84488 480 84516 3198
rect 85672 3120 85724 3126
rect 85672 3062 85724 3068
rect 85684 480 85712 3062
rect 86788 2938 86816 90510
rect 86880 3126 86908 96766
rect 87420 4072 87472 4078
rect 87420 4014 87472 4020
rect 87432 3194 87460 4014
rect 87616 3262 87644 98942
rect 87972 10600 88024 10606
rect 87972 10542 88024 10548
rect 87604 3256 87656 3262
rect 87604 3198 87656 3204
rect 87420 3188 87472 3194
rect 87420 3130 87472 3136
rect 86868 3120 86920 3126
rect 86868 3062 86920 3068
rect 86788 2910 86908 2938
rect 86880 480 86908 2910
rect 87984 480 88012 10542
rect 88996 4010 89024 99078
rect 93124 99068 93176 99074
rect 93124 99010 93176 99016
rect 90364 86488 90416 86494
rect 90364 86430 90416 86436
rect 88984 4004 89036 4010
rect 88984 3946 89036 3952
rect 90376 3262 90404 86430
rect 92388 10668 92440 10674
rect 92388 10610 92440 10616
rect 92400 3262 92428 10610
rect 89168 3256 89220 3262
rect 89168 3198 89220 3204
rect 90364 3256 90416 3262
rect 90364 3198 90416 3204
rect 91560 3256 91612 3262
rect 91560 3198 91612 3204
rect 92388 3256 92440 3262
rect 92388 3198 92440 3204
rect 92756 3256 92808 3262
rect 92756 3198 92808 3204
rect 89180 480 89208 3198
rect 90364 3120 90416 3126
rect 90364 3062 90416 3068
rect 90376 480 90404 3062
rect 91572 480 91600 3198
rect 92768 480 92796 3198
rect 93136 3126 93164 99010
rect 94504 97572 94556 97578
rect 94504 97514 94556 97520
rect 93952 9104 94004 9110
rect 93952 9046 94004 9052
rect 93124 3120 93176 3126
rect 93124 3062 93176 3068
rect 93964 480 93992 9046
rect 94516 7682 94544 97514
rect 95148 10736 95200 10742
rect 95148 10678 95200 10684
rect 94504 7676 94556 7682
rect 94504 7618 94556 7624
rect 95160 480 95188 10678
rect 97276 4146 97304 99146
rect 97448 9172 97500 9178
rect 97448 9114 97500 9120
rect 97264 4140 97316 4146
rect 97264 4082 97316 4088
rect 96252 4004 96304 4010
rect 96252 3946 96304 3952
rect 96264 480 96292 3946
rect 97460 480 97488 9114
rect 98656 6914 98684 99214
rect 111064 97640 111116 97646
rect 111064 97582 111116 97588
rect 104164 97504 104216 97510
rect 104164 97446 104216 97452
rect 101404 94580 101456 94586
rect 101404 94522 101456 94528
rect 99288 11960 99340 11966
rect 99288 11902 99340 11908
rect 98564 6886 98684 6914
rect 98564 3330 98592 6886
rect 98552 3324 98604 3330
rect 98552 3266 98604 3272
rect 99300 3194 99328 11902
rect 101036 9240 101088 9246
rect 101036 9182 101088 9188
rect 99840 6928 99892 6934
rect 99840 6870 99892 6876
rect 98644 3188 98696 3194
rect 98644 3130 98696 3136
rect 99288 3188 99340 3194
rect 99288 3130 99340 3136
rect 98656 480 98684 3130
rect 99852 480 99880 6870
rect 101048 480 101076 9182
rect 101416 3330 101444 94522
rect 103428 12028 103480 12034
rect 103428 11970 103480 11976
rect 103336 4140 103388 4146
rect 103336 4082 103388 4088
rect 102232 3392 102284 3398
rect 102232 3334 102284 3340
rect 101404 3324 101456 3330
rect 101404 3266 101456 3272
rect 102244 480 102272 3334
rect 103348 480 103376 4082
rect 103440 3398 103468 11970
rect 104176 6934 104204 97446
rect 105544 90636 105596 90642
rect 105544 90578 105596 90584
rect 104532 9308 104584 9314
rect 104532 9250 104584 9256
rect 104164 6928 104216 6934
rect 104164 6870 104216 6876
rect 103428 3392 103480 3398
rect 103428 3334 103480 3340
rect 104544 480 104572 9250
rect 105556 4010 105584 90578
rect 108304 89276 108356 89282
rect 108304 89218 108356 89224
rect 107568 86556 107620 86562
rect 107568 86498 107620 86504
rect 106188 12096 106240 12102
rect 106188 12038 106240 12044
rect 105544 4004 105596 4010
rect 105544 3946 105596 3952
rect 106200 3398 106228 12038
rect 107580 3398 107608 86498
rect 108120 9376 108172 9382
rect 108120 9318 108172 9324
rect 105728 3392 105780 3398
rect 105728 3334 105780 3340
rect 106188 3392 106240 3398
rect 106188 3334 106240 3340
rect 106924 3392 106976 3398
rect 106924 3334 106976 3340
rect 107568 3392 107620 3398
rect 107568 3334 107620 3340
rect 105740 480 105768 3334
rect 106936 480 106964 3334
rect 108132 480 108160 9318
rect 108316 4078 108344 89218
rect 110328 12164 110380 12170
rect 110328 12106 110380 12112
rect 108304 4072 108356 4078
rect 108304 4014 108356 4020
rect 110340 3398 110368 12106
rect 110512 4004 110564 4010
rect 110512 3946 110564 3952
rect 109316 3392 109368 3398
rect 109316 3334 109368 3340
rect 110328 3392 110380 3398
rect 110328 3334 110380 3340
rect 109328 480 109356 3334
rect 110524 480 110552 3946
rect 111076 3262 111104 97582
rect 111616 9444 111668 9450
rect 111616 9386 111668 9392
rect 111064 3256 111116 3262
rect 111064 3198 111116 3204
rect 111628 480 111656 9386
rect 112456 4146 112484 99282
rect 126888 97912 126940 97918
rect 126888 97854 126940 97860
rect 124864 97844 124916 97850
rect 124864 97786 124916 97792
rect 115204 97708 115256 97714
rect 115204 97650 115256 97656
rect 112812 12232 112864 12238
rect 112812 12174 112864 12180
rect 112444 4140 112496 4146
rect 112444 4082 112496 4088
rect 112824 480 112852 12174
rect 115216 3398 115244 97650
rect 121368 94648 121420 94654
rect 121368 94590 121420 94596
rect 116584 90704 116636 90710
rect 116584 90646 116636 90652
rect 114008 3392 114060 3398
rect 114008 3334 114060 3340
rect 115204 3392 115256 3398
rect 115204 3334 115256 3340
rect 116400 3392 116452 3398
rect 116400 3334 116452 3340
rect 114020 480 114048 3334
rect 115204 3256 115256 3262
rect 115204 3198 115256 3204
rect 115216 480 115244 3198
rect 116412 480 116440 3334
rect 116596 3262 116624 90646
rect 119988 89344 120040 89350
rect 119988 89286 120040 89292
rect 117228 87984 117280 87990
rect 117228 87926 117280 87932
rect 117240 3398 117268 87926
rect 119896 13116 119948 13122
rect 119896 13058 119948 13064
rect 117596 4072 117648 4078
rect 117596 4014 117648 4020
rect 117228 3392 117280 3398
rect 117228 3334 117280 3340
rect 116584 3256 116636 3262
rect 116584 3198 116636 3204
rect 117608 480 117636 4014
rect 118792 2916 118844 2922
rect 118792 2858 118844 2864
rect 118804 480 118832 2858
rect 119908 480 119936 13058
rect 120000 2922 120028 89286
rect 121380 6914 121408 94590
rect 122748 89412 122800 89418
rect 122748 89354 122800 89360
rect 121104 6886 121408 6914
rect 119988 2916 120040 2922
rect 119988 2858 120040 2864
rect 121104 480 121132 6886
rect 122760 3398 122788 89354
rect 124128 88052 124180 88058
rect 124128 87994 124180 88000
rect 124140 3398 124168 87994
rect 124876 6322 124904 97786
rect 126244 97776 126296 97782
rect 126244 97718 126296 97724
rect 124864 6316 124916 6322
rect 124864 6258 124916 6264
rect 126256 5574 126284 97718
rect 124680 5568 124732 5574
rect 124680 5510 124732 5516
rect 126244 5568 126296 5574
rect 126244 5510 126296 5516
rect 122288 3392 122340 3398
rect 122288 3334 122340 3340
rect 122748 3392 122800 3398
rect 122748 3334 122800 3340
rect 123484 3392 123536 3398
rect 123484 3334 123536 3340
rect 124128 3392 124180 3398
rect 124128 3334 124180 3340
rect 122300 480 122328 3334
rect 123496 480 123524 3334
rect 124692 480 124720 5510
rect 126900 3398 126928 97854
rect 133788 96144 133840 96150
rect 133788 96086 133840 96092
rect 131028 96076 131080 96082
rect 131028 96018 131080 96024
rect 128268 94716 128320 94722
rect 128268 94658 128320 94664
rect 128176 92064 128228 92070
rect 128176 92006 128228 92012
rect 125876 3392 125928 3398
rect 125876 3334 125928 3340
rect 126888 3392 126940 3398
rect 126888 3334 126940 3340
rect 125888 480 125916 3334
rect 126980 2984 127032 2990
rect 126980 2926 127032 2932
rect 126992 480 127020 2926
rect 128188 480 128216 92006
rect 128280 2990 128308 94658
rect 129372 4140 129424 4146
rect 129372 4082 129424 4088
rect 128268 2984 128320 2990
rect 128268 2926 128320 2932
rect 129384 480 129412 4082
rect 131040 3398 131068 96018
rect 131764 5160 131816 5166
rect 131764 5102 131816 5108
rect 130568 3392 130620 3398
rect 130568 3334 130620 3340
rect 131028 3392 131080 3398
rect 131028 3334 131080 3340
rect 130580 480 130608 3334
rect 131776 480 131804 5102
rect 133800 3398 133828 96086
rect 137284 94784 137336 94790
rect 137284 94726 137336 94732
rect 136548 93424 136600 93430
rect 136548 93366 136600 93372
rect 135168 93356 135220 93362
rect 135168 93298 135220 93304
rect 135180 3398 135208 93298
rect 136560 3398 136588 93366
rect 132960 3392 133012 3398
rect 132960 3334 133012 3340
rect 133788 3392 133840 3398
rect 133788 3334 133840 3340
rect 134156 3392 134208 3398
rect 134156 3334 134208 3340
rect 135168 3392 135220 3398
rect 135168 3334 135220 3340
rect 135260 3392 135312 3398
rect 135260 3334 135312 3340
rect 136548 3392 136600 3398
rect 136548 3334 136600 3340
rect 132972 480 133000 3334
rect 134168 480 134196 3334
rect 135272 480 135300 3334
rect 137296 3330 137324 94726
rect 142068 93492 142120 93498
rect 142068 93434 142120 93440
rect 137928 92132 137980 92138
rect 137928 92074 137980 92080
rect 137940 6914 137968 92074
rect 139308 90772 139360 90778
rect 139308 90714 139360 90720
rect 137664 6886 137968 6914
rect 136456 3324 136508 3330
rect 136456 3266 136508 3272
rect 137284 3324 137336 3330
rect 137284 3266 137336 3272
rect 136468 480 136496 3266
rect 137664 480 137692 6886
rect 139320 3398 139348 90714
rect 142080 3398 142108 93434
rect 143448 90840 143500 90846
rect 143448 90782 143500 90788
rect 143460 3398 143488 90782
rect 144196 20670 144224 299746
rect 144828 94852 144880 94858
rect 144828 94794 144880 94800
rect 144184 20664 144236 20670
rect 144184 20606 144236 20612
rect 138848 3392 138900 3398
rect 138848 3334 138900 3340
rect 139308 3392 139360 3398
rect 139308 3334 139360 3340
rect 141240 3392 141292 3398
rect 141240 3334 141292 3340
rect 142068 3392 142120 3398
rect 142068 3334 142120 3340
rect 142436 3392 142488 3398
rect 142436 3334 142488 3340
rect 143448 3392 143500 3398
rect 143448 3334 143500 3340
rect 144736 3392 144788 3398
rect 144736 3334 144788 3340
rect 138860 480 138888 3334
rect 140044 3324 140096 3330
rect 140044 3266 140096 3272
rect 140056 480 140084 3266
rect 141252 480 141280 3334
rect 142448 480 142476 3334
rect 143540 3256 143592 3262
rect 143540 3198 143592 3204
rect 143552 480 143580 3198
rect 144748 480 144776 3334
rect 144840 3262 144868 94794
rect 145564 93560 145616 93566
rect 145564 93502 145616 93508
rect 145576 3398 145604 93502
rect 146956 59362 146984 301174
rect 148324 299872 148376 299878
rect 148324 299814 148376 299820
rect 147588 95056 147640 95062
rect 147588 94998 147640 95004
rect 146944 59356 146996 59362
rect 146944 59298 146996 59304
rect 145932 7676 145984 7682
rect 145932 7618 145984 7624
rect 145564 3392 145616 3398
rect 145564 3334 145616 3340
rect 144828 3256 144880 3262
rect 144828 3198 144880 3204
rect 145944 480 145972 7618
rect 147600 3398 147628 94998
rect 148336 45558 148364 299814
rect 150348 97980 150400 97986
rect 150348 97922 150400 97928
rect 148968 92200 149020 92206
rect 148968 92142 149020 92148
rect 148324 45552 148376 45558
rect 148324 45494 148376 45500
rect 148980 3398 149008 92142
rect 150360 3398 150388 97922
rect 151096 85542 151124 301242
rect 152464 300008 152516 300014
rect 152464 299950 152516 299956
rect 152476 137970 152504 299950
rect 155224 299940 155276 299946
rect 155224 299882 155276 299888
rect 152464 137964 152516 137970
rect 152464 137906 152516 137912
rect 153108 93628 153160 93634
rect 153108 93570 153160 93576
rect 153016 90908 153068 90914
rect 153016 90850 153068 90856
rect 151084 85536 151136 85542
rect 151084 85478 151136 85484
rect 147128 3392 147180 3398
rect 147128 3334 147180 3340
rect 147588 3392 147640 3398
rect 147588 3334 147640 3340
rect 148324 3392 148376 3398
rect 148324 3334 148376 3340
rect 148968 3392 149020 3398
rect 148968 3334 149020 3340
rect 149520 3392 149572 3398
rect 149520 3334 149572 3340
rect 150348 3392 150400 3398
rect 150348 3334 150400 3340
rect 147140 480 147168 3334
rect 148336 480 148364 3334
rect 149532 480 149560 3334
rect 150624 3324 150676 3330
rect 150624 3266 150676 3272
rect 150636 480 150664 3266
rect 151820 3188 151872 3194
rect 151820 3130 151872 3136
rect 151832 480 151860 3130
rect 153028 480 153056 90850
rect 153120 3194 153148 93570
rect 155236 33114 155264 299882
rect 159376 164218 159404 301310
rect 170404 300076 170456 300082
rect 170404 300018 170456 300024
rect 160100 287088 160152 287094
rect 160100 287030 160152 287036
rect 160112 171134 160140 287030
rect 160112 171106 160600 171134
rect 159364 164212 159416 164218
rect 159364 164154 159416 164160
rect 160572 160698 160600 171106
rect 169208 160812 169260 160818
rect 169208 160754 169260 160760
rect 169220 160698 169248 160754
rect 160572 160670 160954 160698
rect 168958 160670 169248 160698
rect 165160 160540 165212 160546
rect 165160 160482 165212 160488
rect 165172 160426 165200 160482
rect 164910 160398 165200 160426
rect 162872 158710 162900 160004
rect 162860 158704 162912 158710
rect 162860 158646 162912 158652
rect 166920 158030 166948 160004
rect 166908 158024 166960 158030
rect 166908 157966 166960 157972
rect 160940 123010 160968 124100
rect 160928 123004 160980 123010
rect 160928 122946 160980 122952
rect 162872 122942 162900 124100
rect 162860 122936 162912 122942
rect 162860 122878 162912 122884
rect 164896 122874 164924 124100
rect 164884 122868 164936 122874
rect 164884 122810 164936 122816
rect 166920 122806 166948 124100
rect 166908 122800 166960 122806
rect 166908 122742 166960 122748
rect 168944 122738 168972 124100
rect 168932 122732 168984 122738
rect 168932 122674 168984 122680
rect 170416 111790 170444 300018
rect 175924 267776 175976 267782
rect 175924 267718 175976 267724
rect 174544 264988 174596 264994
rect 174544 264930 174596 264936
rect 171784 248464 171836 248470
rect 171784 248406 171836 248412
rect 170496 222216 170548 222222
rect 170496 222158 170548 222164
rect 170508 123010 170536 222158
rect 171692 175228 171744 175234
rect 171692 175170 171744 175176
rect 171704 174865 171732 175170
rect 171690 174856 171746 174865
rect 171690 174791 171746 174800
rect 171508 173868 171560 173874
rect 171508 173810 171560 173816
rect 171520 173641 171548 173810
rect 171506 173632 171562 173641
rect 171506 173567 171562 173576
rect 171796 170513 171824 248406
rect 171876 244316 171928 244322
rect 171876 244258 171928 244264
rect 171782 170504 171838 170513
rect 171782 170439 171838 170448
rect 171888 168201 171916 244258
rect 171968 238808 172020 238814
rect 171968 238750 172020 238756
rect 171874 168192 171930 168201
rect 171874 168127 171930 168136
rect 171784 164892 171836 164898
rect 171784 164834 171836 164840
rect 171796 162353 171824 164834
rect 171980 164529 172008 238750
rect 172060 234660 172112 234666
rect 172060 234602 172112 234608
rect 171966 164520 172022 164529
rect 171966 164455 172022 164464
rect 172072 163577 172100 234602
rect 173164 207052 173216 207058
rect 173164 206994 173216 207000
rect 172428 190460 172480 190466
rect 172428 190402 172480 190408
rect 172440 189961 172468 190402
rect 172426 189952 172482 189961
rect 172426 189887 172482 189896
rect 172428 189032 172480 189038
rect 172428 188974 172480 188980
rect 172440 188737 172468 188974
rect 172426 188728 172482 188737
rect 172426 188663 172482 188672
rect 172428 187672 172480 187678
rect 172428 187614 172480 187620
rect 172440 187377 172468 187614
rect 172426 187368 172482 187377
rect 172426 187303 172482 187312
rect 172428 186312 172480 186318
rect 172428 186254 172480 186260
rect 172440 186153 172468 186254
rect 172426 186144 172482 186153
rect 172426 186079 172482 186088
rect 172336 184884 172388 184890
rect 172336 184826 172388 184832
rect 172348 184385 172376 184826
rect 172428 184816 172480 184822
rect 172426 184784 172428 184793
rect 172480 184784 172482 184793
rect 172426 184719 172482 184728
rect 172334 184376 172390 184385
rect 172334 184311 172390 184320
rect 172428 183524 172480 183530
rect 172428 183466 172480 183472
rect 172440 183025 172468 183466
rect 172426 183016 172482 183025
rect 172426 182951 172482 182960
rect 172428 182096 172480 182102
rect 172428 182038 172480 182044
rect 172440 181801 172468 182038
rect 172426 181792 172482 181801
rect 172426 181727 172482 181736
rect 172152 180872 172204 180878
rect 172152 180814 172204 180820
rect 172058 163568 172114 163577
rect 172058 163503 172114 163512
rect 171782 162344 171838 162353
rect 171782 162279 171838 162288
rect 171784 162172 171836 162178
rect 171784 162114 171836 162120
rect 171232 154556 171284 154562
rect 171232 154498 171284 154504
rect 171244 153241 171272 154498
rect 171600 154012 171652 154018
rect 171600 153954 171652 153960
rect 171612 153785 171640 153954
rect 171598 153776 171654 153785
rect 171598 153711 171654 153720
rect 171230 153232 171286 153241
rect 171230 153167 171286 153176
rect 171508 150068 171560 150074
rect 171508 150010 171560 150016
rect 171520 149977 171548 150010
rect 171506 149968 171562 149977
rect 171506 149903 171562 149912
rect 171692 149456 171744 149462
rect 171690 149424 171692 149433
rect 171744 149424 171746 149433
rect 171690 149359 171746 149368
rect 171692 149048 171744 149054
rect 171692 148990 171744 148996
rect 171704 148345 171732 148990
rect 171690 148336 171746 148345
rect 171690 148271 171746 148280
rect 171692 148232 171744 148238
rect 171692 148174 171744 148180
rect 171704 147801 171732 148174
rect 171690 147792 171746 147801
rect 171690 147727 171746 147736
rect 171692 144220 171744 144226
rect 171692 144162 171744 144168
rect 171704 142497 171732 144162
rect 171796 143585 171824 162114
rect 171876 150544 171928 150550
rect 171874 150512 171876 150521
rect 171928 150512 171930 150521
rect 171874 150447 171930 150456
rect 171876 148912 171928 148918
rect 171874 148880 171876 148889
rect 171928 148880 171930 148889
rect 171874 148815 171930 148824
rect 171876 147552 171928 147558
rect 171876 147494 171928 147500
rect 171888 146713 171916 147494
rect 171874 146704 171930 146713
rect 171874 146639 171930 146648
rect 172164 144129 172192 180814
rect 172428 180600 172480 180606
rect 172426 180568 172428 180577
rect 172480 180568 172482 180577
rect 172426 180503 172482 180512
rect 172428 179240 172480 179246
rect 172426 179208 172428 179217
rect 172480 179208 172482 179217
rect 172426 179143 172482 179152
rect 172428 178016 172480 178022
rect 172334 177984 172390 177993
rect 172428 177958 172480 177964
rect 172334 177919 172336 177928
rect 172388 177919 172390 177928
rect 172336 177890 172388 177896
rect 172440 177449 172468 177958
rect 172426 177440 172482 177449
rect 172426 177375 172482 177384
rect 172428 176656 172480 176662
rect 172428 176598 172480 176604
rect 172440 176089 172468 176598
rect 172426 176080 172482 176089
rect 172426 176015 172482 176024
rect 172428 172508 172480 172514
rect 172428 172450 172480 172456
rect 172440 172417 172468 172450
rect 172426 172408 172482 172417
rect 172426 172343 172482 172352
rect 172428 171080 172480 171086
rect 172426 171048 172428 171057
rect 172480 171048 172482 171057
rect 172426 170983 172482 170992
rect 172428 169720 172480 169726
rect 172428 169662 172480 169668
rect 172440 169153 172468 169662
rect 172426 169144 172482 169153
rect 172426 169079 172482 169088
rect 172428 167000 172480 167006
rect 172428 166942 172480 166948
rect 172440 166705 172468 166942
rect 172426 166696 172482 166705
rect 172426 166631 172482 166640
rect 172428 164212 172480 164218
rect 172428 164154 172480 164160
rect 172440 164121 172468 164154
rect 172426 164112 172482 164121
rect 172426 164047 172482 164056
rect 172244 161152 172296 161158
rect 172244 161094 172296 161100
rect 172256 160993 172284 161094
rect 172242 160984 172298 160993
rect 172242 160919 172298 160928
rect 172428 153196 172480 153202
rect 172428 153138 172480 153144
rect 172336 153128 172388 153134
rect 172336 153070 172388 153076
rect 172348 152153 172376 153070
rect 172440 152697 172468 153138
rect 172426 152688 172482 152697
rect 172426 152623 172482 152632
rect 172334 152144 172390 152153
rect 172334 152079 172390 152088
rect 172336 151700 172388 151706
rect 172336 151642 172388 151648
rect 172348 151065 172376 151642
rect 172428 151632 172480 151638
rect 172426 151600 172428 151609
rect 172480 151600 172482 151609
rect 172426 151535 172482 151544
rect 172334 151056 172390 151065
rect 172334 150991 172390 151000
rect 173176 150550 173204 206994
rect 173256 204332 173308 204338
rect 173256 204274 173308 204280
rect 173164 150544 173216 150550
rect 173164 150486 173216 150492
rect 173268 150074 173296 204274
rect 173348 202904 173400 202910
rect 173348 202846 173400 202852
rect 173256 150068 173308 150074
rect 173256 150010 173308 150016
rect 173360 149462 173388 202846
rect 173440 200184 173492 200190
rect 173440 200126 173492 200132
rect 173348 149456 173400 149462
rect 173348 149398 173400 149404
rect 173452 148918 173480 200126
rect 173532 198756 173584 198762
rect 173532 198698 173584 198704
rect 173544 149054 173572 198698
rect 173624 196036 173676 196042
rect 173624 195978 173676 195984
rect 173532 149048 173584 149054
rect 173532 148990 173584 148996
rect 173440 148912 173492 148918
rect 173440 148854 173492 148860
rect 173164 148368 173216 148374
rect 173164 148310 173216 148316
rect 172428 147620 172480 147626
rect 172428 147562 172480 147568
rect 172440 147257 172468 147562
rect 172426 147248 172482 147257
rect 172426 147183 172482 147192
rect 172336 146260 172388 146266
rect 172336 146202 172388 146208
rect 172242 146160 172298 146169
rect 172242 146095 172244 146104
rect 172296 146095 172298 146104
rect 172244 146066 172296 146072
rect 172348 145081 172376 146202
rect 172428 146192 172480 146198
rect 172428 146134 172480 146140
rect 172440 145625 172468 146134
rect 172426 145616 172482 145625
rect 172426 145551 172482 145560
rect 172334 145072 172390 145081
rect 172334 145007 172390 145016
rect 172428 144900 172480 144906
rect 172428 144842 172480 144848
rect 172440 144537 172468 144842
rect 172426 144528 172482 144537
rect 172426 144463 172482 144472
rect 172150 144120 172206 144129
rect 172150 144055 172206 144064
rect 171782 143576 171838 143585
rect 171782 143511 171838 143520
rect 171876 143540 171928 143546
rect 171876 143482 171928 143488
rect 171888 143041 171916 143482
rect 171874 143032 171930 143041
rect 171874 142967 171930 142976
rect 171784 142860 171836 142866
rect 171784 142802 171836 142808
rect 171690 142488 171746 142497
rect 171690 142423 171746 142432
rect 171508 142316 171560 142322
rect 171508 142258 171560 142264
rect 171520 141953 171548 142258
rect 171506 141944 171562 141953
rect 171506 141879 171562 141888
rect 171692 141432 171744 141438
rect 171796 141409 171824 142802
rect 172428 142112 172480 142118
rect 172428 142054 172480 142060
rect 171692 141374 171744 141380
rect 171782 141400 171838 141409
rect 171704 140321 171732 141374
rect 171782 141335 171838 141344
rect 172440 140865 172468 142054
rect 172426 140856 172482 140865
rect 172426 140791 172482 140800
rect 171690 140312 171746 140321
rect 171690 140247 171746 140256
rect 172336 140072 172388 140078
rect 172336 140014 172388 140020
rect 171692 139800 171744 139806
rect 171690 139768 171692 139777
rect 171744 139768 171746 139777
rect 171690 139703 171746 139712
rect 171600 139120 171652 139126
rect 171600 139062 171652 139068
rect 171612 138689 171640 139062
rect 171598 138680 171654 138689
rect 171598 138615 171654 138624
rect 171508 138236 171560 138242
rect 171508 138178 171560 138184
rect 171520 138145 171548 138178
rect 171506 138136 171562 138145
rect 171506 138071 171562 138080
rect 172060 137964 172112 137970
rect 172060 137906 172112 137912
rect 172072 137601 172100 137906
rect 172058 137592 172114 137601
rect 172058 137527 172114 137536
rect 172348 137057 172376 140014
rect 173176 139806 173204 148310
rect 173636 148238 173664 195978
rect 174556 179246 174584 264930
rect 175936 180606 175964 267718
rect 177304 229152 177356 229158
rect 177304 229094 177356 229100
rect 176016 191888 176068 191894
rect 176016 191830 176068 191836
rect 175924 180600 175976 180606
rect 175924 180542 175976 180548
rect 174544 179240 174596 179246
rect 174544 179182 174596 179188
rect 174544 172576 174596 172582
rect 174544 172518 174596 172524
rect 173624 148232 173676 148238
rect 173624 148174 173676 148180
rect 174556 142322 174584 172518
rect 176028 147558 176056 191830
rect 176016 147552 176068 147558
rect 176016 147494 176068 147500
rect 174544 142316 174596 142322
rect 174544 142258 174596 142264
rect 173164 139800 173216 139806
rect 173164 139742 173216 139748
rect 172428 139392 172480 139398
rect 172428 139334 172480 139340
rect 172440 139233 172468 139334
rect 172426 139224 172482 139233
rect 172426 139159 172482 139168
rect 172428 137284 172480 137290
rect 172428 137226 172480 137232
rect 172334 137048 172390 137057
rect 172334 136983 172390 136992
rect 172244 136604 172296 136610
rect 172244 136546 172296 136552
rect 171692 136536 171744 136542
rect 171692 136478 171744 136484
rect 171704 135425 171732 136478
rect 172256 135969 172284 136546
rect 172440 136513 172468 137226
rect 172520 136672 172572 136678
rect 172520 136614 172572 136620
rect 172426 136504 172482 136513
rect 172426 136439 172482 136448
rect 172242 135960 172298 135969
rect 172242 135895 172298 135904
rect 171690 135416 171746 135425
rect 171690 135351 171746 135360
rect 172336 135312 172388 135318
rect 172336 135254 172388 135260
rect 171232 135244 171284 135250
rect 171232 135186 171284 135192
rect 171244 133929 171272 135186
rect 172244 135108 172296 135114
rect 172244 135050 172296 135056
rect 172256 134337 172284 135050
rect 172242 134328 172298 134337
rect 172242 134263 172298 134272
rect 171230 133920 171286 133929
rect 171230 133855 171286 133864
rect 172348 132841 172376 135254
rect 172428 135176 172480 135182
rect 172428 135118 172480 135124
rect 172440 134881 172468 135118
rect 172426 134872 172482 134881
rect 172426 134807 172482 134816
rect 172426 133376 172482 133385
rect 172532 133362 172560 136614
rect 172482 133334 172560 133362
rect 172426 133311 172482 133320
rect 172334 132832 172390 132841
rect 172334 132767 172390 132776
rect 171140 132524 171192 132530
rect 171140 132466 171192 132472
rect 171152 132297 171180 132466
rect 171138 132288 171194 132297
rect 171138 132223 171194 132232
rect 172428 131776 172480 131782
rect 172426 131744 172428 131753
rect 172480 131744 172482 131753
rect 172426 131679 172482 131688
rect 171506 131200 171562 131209
rect 171506 131135 171562 131144
rect 171520 129742 171548 131135
rect 172334 130656 172390 130665
rect 172334 130591 172390 130600
rect 171874 130112 171930 130121
rect 171874 130047 171876 130056
rect 171928 130047 171930 130056
rect 171876 130018 171928 130024
rect 171508 129736 171560 129742
rect 171508 129678 171560 129684
rect 172058 129024 172114 129033
rect 172058 128959 172114 128968
rect 171874 128480 171930 128489
rect 171874 128415 171930 128424
rect 171782 127392 171838 127401
rect 171782 127327 171838 127336
rect 171690 124672 171746 124681
rect 171690 124607 171746 124616
rect 171704 124302 171732 124607
rect 171692 124296 171744 124302
rect 171692 124238 171744 124244
rect 170496 123004 170548 123010
rect 170496 122946 170548 122952
rect 171796 114510 171824 127327
rect 171888 118658 171916 128415
rect 171966 127936 172022 127945
rect 171966 127871 172022 127880
rect 171876 118652 171928 118658
rect 171876 118594 171928 118600
rect 171980 117298 172008 127871
rect 172072 121446 172100 128959
rect 172348 126954 172376 130591
rect 172426 129568 172482 129577
rect 172482 129526 172560 129554
rect 172426 129503 172482 129512
rect 172532 127634 172560 129526
rect 172520 127628 172572 127634
rect 172520 127570 172572 127576
rect 172336 126948 172388 126954
rect 172336 126890 172388 126896
rect 172242 126848 172298 126857
rect 172242 126783 172298 126792
rect 172256 125662 172284 126783
rect 172334 126304 172390 126313
rect 172334 126239 172390 126248
rect 172348 125730 172376 126239
rect 172428 125792 172480 125798
rect 172426 125760 172428 125769
rect 172480 125760 172482 125769
rect 172336 125724 172388 125730
rect 172426 125695 172482 125704
rect 172336 125666 172388 125672
rect 172244 125656 172296 125662
rect 172244 125598 172296 125604
rect 172426 125216 172482 125225
rect 172426 125151 172482 125160
rect 172440 124370 172468 125151
rect 172428 124364 172480 124370
rect 172428 124306 172480 124312
rect 172150 124264 172206 124273
rect 172150 124199 172152 124208
rect 172204 124199 172206 124208
rect 173164 124228 173216 124234
rect 172152 124170 172204 124176
rect 173164 124170 173216 124176
rect 172060 121440 172112 121446
rect 172060 121382 172112 121388
rect 171968 117292 172020 117298
rect 171968 117234 172020 117240
rect 171784 114504 171836 114510
rect 171784 114446 171836 114452
rect 170404 111784 170456 111790
rect 170404 111726 170456 111732
rect 173176 102134 173204 124170
rect 177316 122738 177344 229094
rect 177408 202842 177436 302874
rect 178684 302864 178736 302870
rect 178684 302806 178736 302812
rect 177488 230512 177540 230518
rect 177488 230454 177540 230460
rect 177396 202836 177448 202842
rect 177396 202778 177448 202784
rect 177500 161158 177528 230454
rect 177488 161152 177540 161158
rect 177488 161094 177540 161100
rect 177396 157412 177448 157418
rect 177396 157354 177448 157360
rect 177408 138242 177436 157354
rect 177396 138236 177448 138242
rect 177396 138178 177448 138184
rect 178696 122806 178724 302806
rect 196624 301708 196676 301714
rect 196624 301650 196676 301656
rect 180064 294024 180116 294030
rect 180064 293966 180116 293972
rect 178776 270564 178828 270570
rect 178776 270506 178828 270512
rect 178788 182102 178816 270506
rect 178868 182844 178920 182850
rect 178868 182786 178920 182792
rect 178776 182096 178828 182102
rect 178776 182038 178828 182044
rect 178880 146130 178908 182786
rect 180076 160818 180104 293966
rect 196636 293962 196664 301650
rect 198568 298897 198596 337350
rect 202800 305930 202828 703520
rect 218992 701010 219020 703520
rect 218980 701004 219032 701010
rect 218980 700946 219032 700952
rect 235184 699718 235212 703520
rect 252560 701004 252612 701010
rect 252560 700946 252612 700952
rect 249616 700936 249668 700942
rect 249616 700878 249668 700884
rect 246948 700732 247000 700738
rect 246948 700674 247000 700680
rect 244188 700528 244240 700534
rect 244188 700470 244240 700476
rect 241428 700324 241480 700330
rect 241428 700266 241480 700272
rect 235172 699712 235224 699718
rect 235172 699654 235224 699660
rect 240784 699712 240836 699718
rect 240784 699654 240836 699660
rect 238668 696992 238720 696998
rect 238668 696934 238720 696940
rect 238576 683188 238628 683194
rect 238576 683130 238628 683136
rect 237288 670744 237340 670750
rect 237288 670686 237340 670692
rect 235908 643136 235960 643142
rect 235908 643078 235960 643084
rect 235816 630692 235868 630698
rect 235816 630634 235868 630640
rect 234528 616888 234580 616894
rect 234528 616830 234580 616836
rect 233148 590708 233200 590714
rect 233148 590650 233200 590656
rect 233056 576904 233108 576910
rect 233056 576846 233108 576852
rect 231768 563100 231820 563106
rect 231768 563042 231820 563048
rect 230388 536852 230440 536858
rect 230388 536794 230440 536800
rect 229008 510672 229060 510678
rect 229008 510614 229060 510620
rect 227628 484424 227680 484430
rect 227628 484366 227680 484372
rect 226248 456816 226300 456822
rect 226248 456758 226300 456764
rect 224868 430636 224920 430642
rect 224868 430578 224920 430584
rect 224776 404388 224828 404394
rect 224776 404330 224828 404336
rect 222016 378208 222068 378214
rect 222016 378150 222068 378156
rect 219348 324352 219400 324358
rect 219348 324294 219400 324300
rect 202788 305924 202840 305930
rect 202788 305866 202840 305872
rect 215024 303000 215076 303006
rect 215024 302942 215076 302948
rect 214104 302796 214156 302802
rect 214104 302738 214156 302744
rect 211528 302728 211580 302734
rect 211528 302670 211580 302676
rect 207204 302524 207256 302530
rect 207204 302466 207256 302472
rect 204628 302456 204680 302462
rect 204628 302398 204680 302404
rect 202052 302388 202104 302394
rect 202052 302330 202104 302336
rect 199384 301640 199436 301646
rect 199384 301582 199436 301588
rect 198554 298888 198610 298897
rect 198554 298823 198610 298832
rect 197910 294536 197966 294545
rect 197910 294471 197966 294480
rect 197924 294030 197952 294471
rect 197912 294024 197964 294030
rect 197912 293966 197964 293972
rect 196624 293956 196676 293962
rect 196624 293898 196676 293904
rect 198094 292360 198150 292369
rect 198094 292295 198150 292304
rect 198108 291854 198136 292295
rect 195244 291848 195296 291854
rect 195244 291790 195296 291796
rect 198096 291848 198148 291854
rect 198096 291790 198148 291796
rect 184204 289876 184256 289882
rect 184204 289818 184256 289824
rect 182824 276072 182876 276078
rect 182824 276014 182876 276020
rect 181444 271924 181496 271930
rect 181444 271866 181496 271872
rect 180156 263628 180208 263634
rect 180156 263570 180208 263576
rect 180168 177954 180196 263570
rect 180248 219496 180300 219502
rect 180248 219438 180300 219444
rect 180156 177948 180208 177954
rect 180156 177890 180208 177896
rect 180064 160812 180116 160818
rect 180064 160754 180116 160760
rect 180064 158772 180116 158778
rect 180064 158714 180116 158720
rect 178868 146124 178920 146130
rect 178868 146066 178920 146072
rect 180076 139126 180104 158714
rect 180260 154018 180288 219438
rect 181456 183530 181484 271866
rect 181536 187740 181588 187746
rect 181536 187682 181588 187688
rect 181444 183524 181496 183530
rect 181444 183466 181496 183472
rect 180340 176724 180392 176730
rect 180340 176666 180392 176672
rect 180248 154012 180300 154018
rect 180248 153954 180300 153960
rect 180352 143546 180380 176666
rect 181548 146198 181576 187682
rect 182836 184822 182864 276014
rect 182916 184952 182968 184958
rect 182916 184894 182968 184900
rect 182824 184816 182876 184822
rect 182824 184758 182876 184764
rect 182928 146266 182956 184894
rect 184216 158710 184244 289818
rect 188344 285728 188396 285734
rect 188344 285670 188396 285676
rect 184296 282940 184348 282946
rect 184296 282882 184348 282888
rect 184308 189038 184336 282882
rect 186964 280220 187016 280226
rect 186964 280162 187016 280168
rect 184388 237448 184440 237454
rect 184388 237390 184440 237396
rect 184296 189032 184348 189038
rect 184296 188974 184348 188980
rect 184400 164218 184428 237390
rect 186976 187678 187004 280162
rect 187056 252612 187108 252618
rect 187056 252554 187108 252560
rect 186964 187672 187016 187678
rect 186964 187614 187016 187620
rect 187068 172514 187096 252554
rect 187148 208412 187200 208418
rect 187148 208354 187200 208360
rect 187056 172508 187108 172514
rect 187056 172450 187108 172456
rect 186964 169788 187016 169794
rect 186964 169730 187016 169736
rect 184388 164212 184440 164218
rect 184388 164154 184440 164160
rect 184296 161492 184348 161498
rect 184296 161434 184348 161440
rect 184204 158704 184256 158710
rect 184204 158646 184256 158652
rect 182916 146260 182968 146266
rect 182916 146202 182968 146208
rect 181536 146192 181588 146198
rect 181536 146134 181588 146140
rect 180340 143540 180392 143546
rect 180340 143482 180392 143488
rect 184308 139398 184336 161434
rect 186976 142866 187004 169730
rect 187160 151706 187188 208354
rect 188356 190466 188384 285670
rect 193956 278996 194008 279002
rect 193956 278938 194008 278944
rect 191104 256760 191156 256766
rect 191104 256702 191156 256708
rect 188436 255332 188488 255338
rect 188436 255274 188488 255280
rect 188344 190460 188396 190466
rect 188344 190402 188396 190408
rect 188344 173936 188396 173942
rect 188344 173878 188396 173884
rect 187148 151700 187200 151706
rect 187148 151642 187200 151648
rect 187056 151088 187108 151094
rect 187056 151030 187108 151036
rect 186964 142860 187016 142866
rect 186964 142802 187016 142808
rect 184296 139392 184348 139398
rect 184296 139334 184348 139340
rect 180064 139120 180116 139126
rect 180064 139062 180116 139068
rect 187068 137970 187096 151030
rect 188356 144226 188384 173878
rect 188448 173874 188476 255274
rect 188528 211200 188580 211206
rect 188528 211142 188580 211148
rect 188436 173868 188488 173874
rect 188436 173810 188488 173816
rect 188436 155236 188488 155242
rect 188436 155178 188488 155184
rect 188448 144906 188476 155178
rect 188540 151638 188568 211142
rect 191116 175234 191144 256702
rect 192484 241596 192536 241602
rect 192484 241538 192536 241544
rect 191196 233436 191248 233442
rect 191196 233378 191248 233384
rect 191104 175228 191156 175234
rect 191104 175170 191156 175176
rect 191104 166116 191156 166122
rect 191104 166058 191156 166064
rect 188528 151632 188580 151638
rect 188528 151574 188580 151580
rect 188436 144900 188488 144906
rect 188436 144842 188488 144848
rect 188344 144220 188396 144226
rect 188344 144162 188396 144168
rect 188528 143608 188580 143614
rect 188528 143550 188580 143556
rect 187148 142180 187200 142186
rect 187148 142122 187200 142128
rect 187056 137964 187108 137970
rect 187056 137906 187108 137912
rect 187160 135114 187188 142122
rect 188540 135182 188568 143550
rect 191116 141438 191144 166058
rect 191208 164898 191236 233378
rect 191288 213988 191340 213994
rect 191288 213930 191340 213936
rect 191196 164892 191248 164898
rect 191196 164834 191248 164840
rect 191300 153134 191328 213930
rect 191380 178084 191432 178090
rect 191380 178026 191432 178032
rect 191392 162178 191420 178026
rect 192496 167006 192524 241538
rect 193864 223644 193916 223650
rect 193864 223586 193916 223592
rect 192484 167000 192536 167006
rect 192484 166942 192536 166948
rect 191380 162172 191432 162178
rect 191380 162114 191432 162120
rect 191288 153128 191340 153134
rect 191288 153070 191340 153076
rect 191196 146532 191248 146538
rect 191196 146474 191248 146480
rect 191104 141432 191156 141438
rect 191104 141374 191156 141380
rect 191208 136542 191236 146474
rect 191196 136536 191248 136542
rect 191196 136478 191248 136484
rect 188528 135176 188580 135182
rect 188528 135118 188580 135124
rect 187148 135108 187200 135114
rect 187148 135050 187200 135056
rect 179420 130076 179472 130082
rect 179420 130018 179472 130024
rect 179432 125594 179460 130018
rect 186964 125792 187016 125798
rect 186964 125734 187016 125740
rect 179420 125588 179472 125594
rect 179420 125530 179472 125536
rect 184204 124364 184256 124370
rect 184204 124306 184256 124312
rect 180064 124296 180116 124302
rect 180064 124238 180116 124244
rect 178684 122800 178736 122806
rect 178684 122742 178736 122748
rect 177304 122732 177356 122738
rect 177304 122674 177356 122680
rect 180076 103494 180104 124238
rect 184216 106282 184244 124306
rect 186976 107642 187004 125734
rect 188344 125724 188396 125730
rect 188344 125666 188396 125672
rect 188356 119406 188384 125666
rect 191104 125656 191156 125662
rect 191104 125598 191156 125604
rect 188344 119400 188396 119406
rect 188344 119342 188396 119348
rect 191116 111790 191144 125598
rect 193876 122942 193904 223586
rect 193968 186318 193996 278938
rect 193956 186312 194008 186318
rect 193956 186254 194008 186260
rect 195256 160750 195284 291790
rect 197358 290184 197414 290193
rect 197358 290119 197414 290128
rect 197372 289882 197400 290119
rect 197360 289876 197412 289882
rect 197360 289818 197412 289824
rect 197634 288008 197690 288017
rect 197634 287943 197690 287952
rect 197648 287094 197676 287943
rect 197636 287088 197688 287094
rect 197636 287030 197688 287036
rect 197358 285832 197414 285841
rect 197358 285767 197414 285776
rect 197372 285734 197400 285767
rect 197360 285728 197412 285734
rect 197360 285670 197412 285676
rect 197358 283656 197414 283665
rect 197358 283591 197414 283600
rect 197372 282946 197400 283591
rect 197360 282940 197412 282946
rect 197360 282882 197412 282888
rect 197358 281480 197414 281489
rect 197358 281415 197414 281424
rect 197372 280226 197400 281415
rect 197360 280220 197412 280226
rect 197360 280162 197412 280168
rect 197358 279304 197414 279313
rect 197358 279239 197414 279248
rect 197372 279002 197400 279239
rect 197360 278996 197412 279002
rect 197360 278938 197412 278944
rect 197542 277128 197598 277137
rect 197542 277063 197598 277072
rect 197556 276078 197584 277063
rect 197544 276072 197596 276078
rect 197544 276014 197596 276020
rect 198370 274952 198426 274961
rect 196624 274916 196676 274922
rect 198370 274887 198372 274896
rect 196624 274858 196676 274864
rect 198424 274887 198426 274896
rect 198372 274858 198424 274864
rect 195336 259548 195388 259554
rect 195336 259490 195388 259496
rect 195348 176662 195376 259490
rect 195428 215348 195480 215354
rect 195428 215290 195480 215296
rect 195336 176656 195388 176662
rect 195336 176598 195388 176604
rect 195336 167068 195388 167074
rect 195336 167010 195388 167016
rect 195244 160744 195296 160750
rect 195244 160686 195296 160692
rect 195244 147688 195296 147694
rect 195244 147630 195296 147636
rect 195256 136610 195284 147630
rect 195348 142118 195376 167010
rect 195440 153202 195468 215290
rect 196636 184890 196664 274858
rect 197358 272776 197414 272785
rect 197358 272711 197414 272720
rect 197372 271930 197400 272711
rect 197360 271924 197412 271930
rect 197360 271866 197412 271872
rect 197358 270600 197414 270609
rect 197358 270535 197360 270544
rect 197412 270535 197414 270544
rect 197360 270506 197412 270512
rect 197726 268424 197782 268433
rect 197726 268359 197782 268368
rect 197740 267782 197768 268359
rect 197728 267776 197780 267782
rect 197728 267718 197780 267724
rect 197358 266248 197414 266257
rect 197358 266183 197414 266192
rect 197372 264994 197400 266183
rect 197360 264988 197412 264994
rect 197360 264930 197412 264936
rect 197910 264072 197966 264081
rect 197910 264007 197966 264016
rect 197924 263634 197952 264007
rect 197912 263628 197964 263634
rect 197912 263570 197964 263576
rect 198646 261896 198702 261905
rect 196716 261860 196768 261866
rect 198646 261831 198648 261840
rect 196716 261802 196768 261808
rect 198700 261831 198702 261840
rect 198648 261802 198700 261808
rect 196624 184884 196676 184890
rect 196624 184826 196676 184832
rect 196728 178022 196756 261802
rect 197726 259720 197782 259729
rect 197726 259655 197782 259664
rect 197740 259554 197768 259655
rect 197728 259548 197780 259554
rect 197728 259490 197780 259496
rect 198094 257544 198150 257553
rect 198094 257479 198150 257488
rect 198108 256766 198136 257479
rect 198096 256760 198148 256766
rect 198096 256702 198148 256708
rect 197358 255368 197414 255377
rect 197358 255303 197360 255312
rect 197412 255303 197414 255312
rect 197360 255274 197412 255280
rect 197358 253192 197414 253201
rect 197358 253127 197414 253136
rect 197372 252618 197400 253127
rect 197360 252612 197412 252618
rect 197360 252554 197412 252560
rect 198002 251016 198058 251025
rect 198002 250951 198058 250960
rect 197358 244488 197414 244497
rect 197358 244423 197414 244432
rect 197372 244322 197400 244423
rect 197360 244316 197412 244322
rect 197360 244258 197412 244264
rect 197726 242312 197782 242321
rect 197726 242247 197782 242256
rect 197740 241602 197768 242247
rect 197728 241596 197780 241602
rect 197728 241538 197780 241544
rect 197358 240136 197414 240145
rect 197358 240071 197414 240080
rect 197372 238814 197400 240071
rect 197360 238808 197412 238814
rect 197360 238750 197412 238756
rect 197358 237960 197414 237969
rect 197358 237895 197414 237904
rect 197372 237454 197400 237895
rect 197360 237448 197412 237454
rect 197360 237390 197412 237396
rect 197542 235784 197598 235793
rect 197542 235719 197598 235728
rect 197556 234666 197584 235719
rect 197544 234660 197596 234666
rect 197544 234602 197596 234608
rect 197634 231432 197690 231441
rect 197634 231367 197690 231376
rect 197648 230518 197676 231367
rect 197636 230512 197688 230518
rect 197636 230454 197688 230460
rect 197358 229256 197414 229265
rect 197358 229191 197414 229200
rect 197372 229158 197400 229191
rect 197360 229152 197412 229158
rect 197360 229094 197412 229100
rect 197358 222728 197414 222737
rect 197358 222663 197414 222672
rect 197372 222222 197400 222663
rect 197360 222216 197412 222222
rect 197360 222158 197412 222164
rect 197542 220552 197598 220561
rect 197542 220487 197598 220496
rect 197556 219502 197584 220487
rect 197544 219496 197596 219502
rect 197544 219438 197596 219444
rect 196808 218204 196860 218210
rect 196808 218146 196860 218152
rect 196716 178016 196768 178022
rect 196716 177958 196768 177964
rect 196624 158024 196676 158030
rect 196624 157966 196676 157972
rect 195428 153196 195480 153202
rect 195428 153138 195480 153144
rect 195336 142112 195388 142118
rect 195336 142054 195388 142060
rect 195244 136604 195296 136610
rect 195244 136546 195296 136552
rect 193864 122936 193916 122942
rect 193864 122878 193916 122884
rect 191104 111784 191156 111790
rect 191104 111726 191156 111732
rect 186964 107636 187016 107642
rect 186964 107578 187016 107584
rect 184204 106276 184256 106282
rect 184204 106218 184256 106224
rect 180064 103488 180116 103494
rect 180064 103430 180116 103436
rect 173164 102128 173216 102134
rect 173164 102070 173216 102076
rect 196636 99414 196664 157966
rect 196820 154562 196848 218146
rect 197910 216200 197966 216209
rect 197910 216135 197966 216144
rect 197924 215354 197952 216135
rect 197912 215348 197964 215354
rect 197912 215290 197964 215296
rect 197358 214024 197414 214033
rect 197358 213959 197360 213968
rect 197412 213959 197414 213968
rect 197360 213930 197412 213936
rect 197726 211848 197782 211857
rect 197726 211783 197782 211792
rect 197740 211206 197768 211783
rect 197728 211200 197780 211206
rect 197728 211142 197780 211148
rect 197358 209672 197414 209681
rect 197358 209607 197414 209616
rect 197372 208418 197400 209607
rect 197360 208412 197412 208418
rect 197360 208354 197412 208360
rect 197358 207496 197414 207505
rect 197358 207431 197414 207440
rect 197372 207058 197400 207431
rect 197360 207052 197412 207058
rect 197360 206994 197412 207000
rect 197542 205320 197598 205329
rect 197542 205255 197598 205264
rect 197556 204338 197584 205255
rect 197544 204332 197596 204338
rect 197544 204274 197596 204280
rect 197358 203144 197414 203153
rect 197358 203079 197414 203088
rect 197372 202910 197400 203079
rect 197360 202904 197412 202910
rect 197360 202846 197412 202852
rect 197358 200968 197414 200977
rect 197358 200903 197414 200912
rect 197372 200190 197400 200903
rect 197360 200184 197412 200190
rect 197360 200126 197412 200132
rect 197358 198792 197414 198801
rect 197358 198727 197360 198736
rect 197412 198727 197414 198736
rect 197360 198698 197412 198704
rect 197358 196616 197414 196625
rect 197358 196551 197414 196560
rect 197372 196042 197400 196551
rect 197360 196036 197412 196042
rect 197360 195978 197412 195984
rect 196900 194404 196952 194410
rect 196900 194346 196952 194352
rect 196808 154556 196860 154562
rect 196808 154498 196860 154504
rect 196716 150612 196768 150618
rect 196716 150554 196768 150560
rect 196728 137290 196756 150554
rect 196912 147626 196940 194346
rect 197358 192264 197414 192273
rect 197358 192199 197414 192208
rect 197372 191894 197400 192199
rect 197360 191888 197412 191894
rect 197360 191830 197412 191836
rect 197542 190088 197598 190097
rect 197542 190023 197598 190032
rect 197358 187912 197414 187921
rect 197358 187847 197414 187856
rect 197372 187746 197400 187847
rect 197360 187740 197412 187746
rect 197360 187682 197412 187688
rect 197358 185736 197414 185745
rect 197358 185671 197414 185680
rect 197372 184958 197400 185671
rect 197360 184952 197412 184958
rect 197360 184894 197412 184900
rect 197556 182850 197584 190023
rect 197544 182844 197596 182850
rect 197544 182786 197596 182792
rect 197358 181384 197414 181393
rect 197358 181319 197414 181328
rect 197372 180878 197400 181319
rect 197360 180872 197412 180878
rect 197360 180814 197412 180820
rect 197542 179208 197598 179217
rect 197542 179143 197598 179152
rect 197556 178090 197584 179143
rect 197544 178084 197596 178090
rect 197544 178026 197596 178032
rect 197358 177032 197414 177041
rect 197358 176967 197414 176976
rect 197372 176730 197400 176967
rect 197360 176724 197412 176730
rect 197360 176666 197412 176672
rect 197634 174856 197690 174865
rect 197634 174791 197690 174800
rect 197648 173942 197676 174791
rect 197636 173936 197688 173942
rect 197636 173878 197688 173884
rect 197358 172680 197414 172689
rect 197358 172615 197414 172624
rect 197372 172582 197400 172615
rect 197360 172576 197412 172582
rect 197360 172518 197412 172524
rect 198016 171086 198044 250951
rect 198186 248840 198242 248849
rect 198186 248775 198242 248784
rect 198200 248470 198228 248775
rect 198188 248464 198240 248470
rect 198188 248406 198240 248412
rect 198094 246664 198150 246673
rect 198094 246599 198150 246608
rect 198004 171080 198056 171086
rect 198004 171022 198056 171028
rect 197358 170504 197414 170513
rect 197358 170439 197414 170448
rect 197372 169794 197400 170439
rect 197360 169788 197412 169794
rect 197360 169730 197412 169736
rect 198108 169726 198136 246599
rect 198186 233608 198242 233617
rect 198186 233543 198242 233552
rect 198200 233442 198228 233543
rect 198188 233436 198240 233442
rect 198188 233378 198240 233384
rect 198738 227080 198794 227089
rect 198738 227015 198794 227024
rect 198278 224904 198334 224913
rect 198278 224839 198334 224848
rect 198292 223650 198320 224839
rect 198280 223644 198332 223650
rect 198280 223586 198332 223592
rect 198462 218376 198518 218385
rect 198462 218311 198518 218320
rect 198476 218210 198504 218311
rect 198464 218204 198516 218210
rect 198464 218146 198516 218152
rect 198646 194440 198702 194449
rect 198646 194375 198648 194384
rect 198700 194375 198702 194384
rect 198648 194346 198700 194352
rect 198186 183560 198242 183569
rect 198186 183495 198242 183504
rect 198096 169720 198148 169726
rect 198096 169662 198148 169668
rect 197910 168328 197966 168337
rect 197910 168263 197966 168272
rect 197924 167074 197952 168263
rect 197912 167068 197964 167074
rect 197912 167010 197964 167016
rect 198002 163976 198058 163985
rect 198002 163911 198058 163920
rect 197358 161800 197414 161809
rect 197358 161735 197414 161744
rect 197372 161498 197400 161735
rect 197360 161492 197412 161498
rect 197360 161434 197412 161440
rect 197358 159624 197414 159633
rect 197358 159559 197414 159568
rect 197372 158778 197400 159559
rect 197360 158772 197412 158778
rect 197360 158714 197412 158720
rect 197358 157448 197414 157457
rect 197358 157383 197360 157392
rect 197412 157383 197414 157392
rect 197360 157354 197412 157360
rect 198016 148374 198044 163911
rect 198200 155242 198228 183495
rect 198462 166152 198518 166161
rect 198462 166087 198464 166096
rect 198516 166087 198518 166096
rect 198464 166058 198516 166064
rect 198278 155272 198334 155281
rect 198188 155236 198240 155242
rect 198278 155207 198334 155216
rect 198188 155178 198240 155184
rect 198094 153096 198150 153105
rect 198094 153031 198150 153040
rect 198004 148368 198056 148374
rect 198004 148310 198056 148316
rect 196900 147620 196952 147626
rect 196900 147562 196952 147568
rect 197726 146568 197782 146577
rect 197726 146503 197728 146512
rect 197780 146503 197782 146512
rect 197728 146474 197780 146480
rect 197358 144392 197414 144401
rect 197358 144327 197414 144336
rect 197372 143614 197400 144327
rect 197360 143608 197412 143614
rect 197360 143550 197412 143556
rect 197358 142216 197414 142225
rect 197358 142151 197360 142160
rect 197412 142151 197414 142160
rect 197360 142122 197412 142128
rect 198108 140078 198136 153031
rect 198292 151094 198320 155207
rect 198280 151088 198332 151094
rect 198280 151030 198332 151036
rect 198370 150920 198426 150929
rect 198370 150855 198426 150864
rect 198384 150618 198412 150855
rect 198372 150612 198424 150618
rect 198372 150554 198424 150560
rect 198278 148744 198334 148753
rect 198278 148679 198334 148688
rect 198292 147694 198320 148679
rect 198280 147688 198332 147694
rect 198280 147630 198332 147636
rect 198096 140072 198148 140078
rect 198096 140014 198148 140020
rect 198278 140040 198334 140049
rect 198278 139975 198334 139984
rect 197542 137864 197598 137873
rect 197542 137799 197598 137808
rect 196716 137284 196768 137290
rect 196716 137226 196768 137232
rect 197556 136678 197584 137799
rect 197544 136672 197596 136678
rect 197544 136614 197596 136620
rect 198094 135688 198150 135697
rect 198094 135623 198150 135632
rect 198108 135318 198136 135623
rect 198096 135312 198148 135318
rect 198096 135254 198148 135260
rect 198292 135250 198320 139975
rect 198280 135244 198332 135250
rect 198280 135186 198332 135192
rect 197542 133512 197598 133521
rect 197542 133447 197598 133456
rect 197556 132530 197584 133447
rect 197544 132524 197596 132530
rect 197544 132466 197596 132472
rect 197912 131776 197964 131782
rect 197912 131718 197964 131724
rect 197924 131345 197952 131718
rect 197910 131336 197966 131345
rect 197910 131271 197966 131280
rect 197360 129736 197412 129742
rect 197360 129678 197412 129684
rect 197372 129169 197400 129678
rect 197358 129160 197414 129169
rect 197358 129095 197414 129104
rect 198004 127628 198056 127634
rect 198004 127570 198056 127576
rect 197358 126984 197414 126993
rect 197358 126919 197360 126928
rect 197412 126919 197414 126928
rect 197360 126890 197412 126896
rect 198016 122641 198044 127570
rect 198556 125588 198608 125594
rect 198556 125530 198608 125536
rect 198568 124817 198596 125530
rect 198554 124808 198610 124817
rect 198554 124743 198610 124752
rect 198752 122874 198780 227015
rect 199396 215286 199424 301582
rect 200396 300892 200448 300898
rect 200396 300834 200448 300840
rect 200408 299948 200436 300834
rect 201224 300212 201276 300218
rect 201224 300154 201276 300160
rect 201236 299948 201264 300154
rect 202064 299948 202092 302330
rect 203800 301436 203852 301442
rect 203800 301378 203852 301384
rect 202972 300960 203024 300966
rect 202972 300902 203024 300908
rect 202984 299948 203012 300902
rect 203812 299948 203840 301378
rect 204640 299948 204668 302398
rect 205548 300280 205600 300286
rect 205548 300222 205600 300228
rect 205560 299948 205588 300222
rect 206376 300144 206428 300150
rect 206376 300086 206428 300092
rect 206388 299948 206416 300086
rect 207216 299948 207244 302466
rect 210700 301504 210752 301510
rect 210700 301446 210752 301452
rect 209872 301164 209924 301170
rect 209872 301106 209924 301112
rect 209884 299948 209912 301106
rect 210712 299948 210740 301446
rect 211540 299948 211568 302670
rect 212448 302592 212500 302598
rect 212448 302534 212500 302540
rect 212460 299948 212488 302534
rect 214116 299948 214144 302738
rect 215036 299948 215064 302942
rect 217600 302660 217652 302666
rect 217600 302602 217652 302608
rect 215852 301572 215904 301578
rect 215852 301514 215904 301520
rect 215864 299948 215892 301514
rect 217612 299948 217640 302602
rect 219360 299948 219388 324294
rect 220636 311908 220688 311914
rect 220636 311850 220688 311856
rect 220648 299962 220676 311850
rect 221004 304292 221056 304298
rect 221004 304234 221056 304240
rect 220202 299934 220676 299962
rect 221016 299948 221044 304234
rect 222028 299962 222056 378150
rect 222752 304360 222804 304366
rect 222752 304302 222804 304308
rect 221950 299934 222056 299962
rect 222764 299948 222792 304302
rect 224788 300354 224816 404330
rect 223672 300348 223724 300354
rect 223672 300290 223724 300296
rect 224776 300348 224828 300354
rect 224776 300290 224828 300296
rect 223684 299948 223712 300290
rect 224880 299962 224908 430578
rect 226156 418192 226208 418198
rect 226156 418134 226208 418140
rect 226168 300354 226196 418134
rect 225328 300348 225380 300354
rect 225328 300290 225380 300296
rect 226156 300348 226208 300354
rect 226156 300290 226208 300296
rect 224526 299934 224908 299962
rect 225340 299948 225368 300290
rect 226260 299948 226288 456758
rect 227640 306374 227668 484366
rect 228916 470620 228968 470626
rect 228916 470562 228968 470568
rect 227456 306346 227668 306374
rect 227456 299962 227484 306346
rect 228928 300354 228956 470562
rect 227904 300348 227956 300354
rect 227904 300290 227956 300296
rect 228916 300348 228968 300354
rect 228916 300290 228968 300296
rect 227102 299934 227484 299962
rect 227916 299948 227944 300290
rect 229020 299962 229048 510614
rect 230400 302122 230428 536794
rect 231676 524476 231728 524482
rect 231676 524418 231728 524424
rect 231688 302190 231716 524418
rect 230480 302184 230532 302190
rect 230480 302126 230532 302132
rect 231676 302184 231728 302190
rect 231676 302126 231728 302132
rect 229652 302116 229704 302122
rect 229652 302058 229704 302064
rect 230388 302116 230440 302122
rect 230388 302058 230440 302064
rect 228850 299934 229048 299962
rect 229664 299948 229692 302058
rect 230492 299948 230520 302126
rect 231780 299962 231808 563042
rect 232228 302116 232280 302122
rect 232228 302058 232280 302064
rect 231426 299934 231808 299962
rect 232240 299948 232268 302058
rect 233068 299962 233096 576846
rect 233160 302122 233188 590650
rect 234540 306374 234568 616830
rect 234448 306346 234568 306374
rect 233148 302116 233200 302122
rect 233148 302058 233200 302064
rect 234448 299962 234476 306346
rect 234804 300484 234856 300490
rect 234804 300426 234856 300432
rect 233068 299934 233174 299962
rect 234002 299934 234476 299962
rect 234816 299948 234844 300426
rect 235828 299962 235856 630634
rect 235920 300490 235948 643078
rect 237300 306374 237328 670686
rect 237024 306346 237328 306374
rect 235908 300484 235960 300490
rect 235908 300426 235960 300432
rect 237024 299962 237052 306346
rect 237380 303068 237432 303074
rect 237380 303010 237432 303016
rect 235750 299934 235856 299962
rect 236578 299934 237052 299962
rect 237392 299948 237420 303010
rect 238588 299962 238616 683130
rect 238680 303074 238708 696934
rect 240048 305652 240100 305658
rect 240048 305594 240100 305600
rect 239128 304428 239180 304434
rect 239128 304370 239180 304376
rect 238668 303068 238720 303074
rect 238668 303010 238720 303016
rect 238326 299934 238616 299962
rect 239140 299948 239168 304370
rect 240060 299948 240088 305594
rect 240796 304842 240824 699654
rect 241440 306374 241468 700266
rect 242716 323604 242768 323610
rect 242716 323546 242768 323552
rect 241256 306346 241468 306374
rect 240784 304836 240836 304842
rect 240784 304778 240836 304784
rect 241256 299962 241284 306346
rect 241704 304496 241756 304502
rect 241704 304438 241756 304444
rect 240902 299934 241284 299962
rect 241716 299948 241744 304438
rect 242728 299962 242756 323546
rect 244200 303074 244228 700470
rect 245568 327752 245620 327758
rect 245568 327694 245620 327700
rect 244280 305788 244332 305794
rect 244280 305730 244332 305736
rect 243452 303068 243504 303074
rect 243452 303010 243504 303016
rect 244188 303068 244240 303074
rect 244188 303010 244240 303016
rect 242650 299934 242756 299962
rect 243464 299948 243492 303010
rect 244292 299948 244320 305730
rect 245580 299962 245608 327694
rect 246856 305856 246908 305862
rect 246856 305798 246908 305804
rect 246028 303068 246080 303074
rect 246028 303010 246080 303016
rect 245226 299934 245608 299962
rect 246040 299948 246068 303010
rect 246868 299962 246896 305798
rect 246960 303074 246988 700674
rect 247776 304768 247828 304774
rect 247776 304710 247828 304716
rect 246948 303068 247000 303074
rect 246948 303010 247000 303016
rect 246868 299934 246974 299962
rect 247788 299948 247816 304710
rect 249524 304700 249576 304706
rect 249524 304642 249576 304648
rect 248604 303068 248656 303074
rect 248604 303010 248656 303016
rect 248616 299948 248644 303010
rect 249536 299948 249564 304642
rect 249628 303074 249656 700878
rect 252468 700256 252520 700262
rect 252468 700198 252520 700204
rect 251088 700188 251140 700194
rect 251088 700130 251140 700136
rect 251100 306374 251128 700130
rect 250824 306346 251128 306374
rect 249616 303068 249668 303074
rect 249616 303010 249668 303016
rect 250824 299962 250852 306346
rect 252100 304836 252152 304842
rect 252100 304778 252152 304784
rect 251180 303068 251232 303074
rect 251180 303010 251232 303016
rect 250378 299934 250852 299962
rect 251192 299948 251220 303010
rect 252112 299948 252140 304778
rect 252480 303074 252508 700198
rect 252572 325694 252600 700946
rect 255320 700868 255372 700874
rect 255320 700810 255372 700816
rect 252572 325666 253336 325694
rect 252928 305924 252980 305930
rect 252928 305866 252980 305872
rect 252468 303068 252520 303074
rect 252468 303010 252520 303016
rect 252940 299948 252968 305866
rect 253308 299962 253336 325666
rect 254676 304632 254728 304638
rect 254676 304574 254728 304580
rect 253308 299934 253782 299962
rect 254688 299948 254716 304574
rect 255332 303074 255360 700810
rect 255412 700800 255464 700806
rect 255412 700742 255464 700748
rect 255320 303068 255372 303074
rect 255320 303010 255372 303016
rect 255424 299962 255452 700742
rect 258080 700664 258132 700670
rect 258080 700606 258132 700612
rect 257252 304564 257304 304570
rect 257252 304506 257304 304512
rect 256148 303068 256200 303074
rect 256148 303010 256200 303016
rect 256160 299962 256188 303010
rect 255424 299934 255530 299962
rect 256160 299934 256450 299962
rect 257264 299948 257292 304506
rect 258092 302122 258120 700606
rect 258172 700596 258224 700602
rect 258172 700538 258224 700544
rect 258080 302116 258132 302122
rect 258080 302058 258132 302064
rect 258184 299962 258212 700538
rect 260840 700460 260892 700466
rect 260840 700402 260892 700408
rect 259460 700392 259512 700398
rect 259460 700334 259512 700340
rect 259472 325694 259500 700334
rect 260852 325694 260880 700402
rect 267660 700194 267688 703520
rect 283852 700262 283880 703520
rect 284944 700392 284996 700398
rect 284944 700334 284996 700340
rect 283840 700256 283892 700262
rect 283840 700198 283892 700204
rect 267648 700188 267700 700194
rect 267648 700130 267700 700136
rect 262220 683256 262272 683262
rect 262220 683198 262272 683204
rect 259472 325666 260328 325694
rect 260852 325666 261248 325694
rect 259828 305720 259880 305726
rect 259828 305662 259880 305668
rect 259000 302116 259052 302122
rect 259000 302058 259052 302064
rect 258106 299934 258212 299962
rect 259012 299948 259040 302058
rect 259840 299948 259868 305662
rect 260300 299962 260328 325666
rect 261220 299962 261248 325666
rect 262232 299962 262260 683198
rect 263600 670812 263652 670818
rect 263600 670754 263652 670760
rect 262312 656940 262364 656946
rect 262312 656882 262364 656888
rect 262324 325694 262352 656882
rect 263612 325694 263640 670754
rect 264980 632120 265032 632126
rect 264980 632062 265032 632068
rect 262324 325666 262904 325694
rect 263612 325666 263824 325694
rect 262876 299962 262904 325666
rect 263796 299962 263824 325666
rect 260300 299934 260682 299962
rect 261220 299934 261602 299962
rect 262232 299934 262430 299962
rect 262876 299934 263350 299962
rect 263796 299934 264178 299962
rect 264992 299948 265020 632062
rect 266360 618316 266412 618322
rect 266360 618258 266412 618264
rect 265072 605872 265124 605878
rect 265072 605814 265124 605820
rect 265084 325694 265112 605814
rect 265084 325666 265480 325694
rect 265452 299962 265480 325666
rect 266372 299962 266400 618258
rect 266452 579692 266504 579698
rect 266452 579634 266504 579640
rect 266464 325694 266492 579634
rect 269120 565888 269172 565894
rect 269120 565830 269172 565836
rect 267740 553444 267792 553450
rect 267740 553386 267792 553392
rect 267752 325694 267780 553386
rect 266464 325666 267136 325694
rect 267752 325666 268056 325694
rect 267108 299962 267136 325666
rect 268028 299962 268056 325666
rect 269132 299962 269160 565830
rect 269212 527196 269264 527202
rect 269212 527138 269264 527144
rect 269224 325694 269252 527138
rect 271880 514820 271932 514826
rect 271880 514762 271932 514768
rect 270500 501016 270552 501022
rect 270500 500958 270552 500964
rect 270512 325694 270540 500958
rect 269224 325666 269896 325694
rect 270512 325666 270632 325694
rect 269868 299962 269896 325666
rect 270604 299962 270632 325666
rect 265452 299934 265926 299962
rect 266372 299934 266754 299962
rect 267108 299934 267582 299962
rect 268028 299934 268502 299962
rect 269132 299934 269330 299962
rect 269868 299934 270250 299962
rect 270604 299934 271078 299962
rect 271892 299948 271920 514762
rect 271972 474768 272024 474774
rect 271972 474710 272024 474716
rect 271984 325694 272012 474710
rect 273260 462392 273312 462398
rect 273260 462334 273312 462340
rect 271984 325666 272472 325694
rect 272444 299962 272472 325666
rect 273272 303074 273300 462334
rect 273352 448588 273404 448594
rect 273352 448530 273404 448536
rect 273260 303068 273312 303074
rect 273260 303010 273312 303016
rect 273364 299962 273392 448530
rect 274640 422340 274692 422346
rect 274640 422282 274692 422288
rect 274652 325694 274680 422282
rect 276020 409896 276072 409902
rect 276020 409838 276072 409844
rect 274652 325666 275048 325694
rect 274180 303068 274232 303074
rect 274180 303010 274232 303016
rect 274192 299962 274220 303010
rect 275020 299962 275048 325666
rect 276032 301850 276060 409838
rect 276112 397520 276164 397526
rect 276112 397462 276164 397468
rect 276020 301844 276072 301850
rect 276020 301786 276072 301792
rect 276124 299962 276152 397462
rect 277400 371272 277452 371278
rect 277400 371214 277452 371220
rect 277412 325694 277440 371214
rect 278780 357468 278832 357474
rect 278780 357410 278832 357416
rect 277412 325666 277624 325694
rect 277032 301844 277084 301850
rect 277032 301786 277084 301792
rect 272444 299934 272826 299962
rect 273364 299934 273654 299962
rect 274192 299934 274482 299962
rect 275020 299934 275402 299962
rect 276124 299934 276230 299962
rect 277044 299948 277072 301786
rect 277596 299962 277624 325666
rect 278792 302122 278820 357410
rect 278872 345092 278924 345098
rect 278872 345034 278924 345040
rect 278780 302116 278832 302122
rect 278780 302058 278832 302064
rect 278884 299962 278912 345034
rect 280252 318844 280304 318850
rect 280252 318786 280304 318792
rect 279700 302116 279752 302122
rect 279700 302058 279752 302064
rect 277596 299934 277978 299962
rect 278806 299934 278912 299962
rect 279712 299948 279740 302058
rect 280264 299962 280292 318786
rect 282276 305040 282328 305046
rect 282276 304982 282328 304988
rect 281356 301708 281408 301714
rect 281356 301650 281408 301656
rect 280264 299934 280554 299962
rect 281368 299948 281396 301650
rect 282288 299948 282316 304982
rect 284956 304774 284984 700334
rect 300136 699718 300164 703520
rect 332520 700398 332548 703520
rect 348804 700942 348832 703520
rect 348792 700936 348844 700942
rect 348792 700878 348844 700884
rect 332508 700392 332560 700398
rect 332508 700334 332560 700340
rect 364996 699718 365024 703520
rect 397472 699718 397500 703520
rect 413664 700738 413692 703520
rect 413652 700732 413704 700738
rect 413652 700674 413704 700680
rect 298744 699712 298796 699718
rect 298744 699654 298796 699660
rect 300124 699712 300176 699718
rect 300124 699654 300176 699660
rect 359464 699712 359516 699718
rect 359464 699654 359516 699660
rect 364984 699712 365036 699718
rect 364984 699654 365036 699660
rect 396724 699712 396776 699718
rect 396724 699654 396776 699660
rect 397460 699712 397512 699718
rect 397460 699654 397512 699660
rect 284944 304768 284996 304774
rect 284944 304710 284996 304716
rect 298756 304706 298784 699654
rect 299940 337476 299992 337482
rect 299940 337418 299992 337424
rect 298744 304700 298796 304706
rect 298744 304642 298796 304648
rect 287428 302932 287480 302938
rect 287428 302874 287480 302880
rect 285680 301640 285732 301646
rect 285680 301582 285732 301588
rect 283104 301096 283156 301102
rect 283104 301038 283156 301044
rect 283116 299948 283144 301038
rect 285692 299948 285720 301582
rect 287440 299948 287468 302874
rect 298652 302864 298704 302870
rect 298652 302806 298704 302812
rect 292580 302320 292632 302326
rect 292580 302262 292632 302268
rect 290004 302252 290056 302258
rect 290004 302194 290056 302200
rect 288256 301368 288308 301374
rect 288256 301310 288308 301316
rect 288268 299948 288296 301310
rect 288900 300008 288952 300014
rect 288952 299956 289202 299962
rect 288900 299950 289202 299956
rect 288912 299934 289202 299950
rect 290016 299948 290044 302194
rect 291752 301300 291804 301306
rect 291752 301242 291804 301248
rect 290556 300076 290608 300082
rect 290556 300018 290608 300024
rect 290568 299962 290596 300018
rect 290568 299934 290858 299962
rect 291764 299948 291792 301242
rect 292592 299948 292620 302262
rect 295156 301232 295208 301238
rect 295156 301174 295208 301180
rect 295168 299948 295196 301174
rect 296904 301028 296956 301034
rect 296904 300970 296956 300976
rect 295720 299946 296102 299962
rect 296916 299948 296944 300970
rect 298664 299948 298692 302806
rect 295708 299940 296102 299946
rect 295760 299934 296102 299940
rect 295708 299882 295760 299888
rect 294052 299872 294104 299878
rect 294104 299820 294354 299826
rect 294052 299814 294354 299820
rect 294064 299798 294354 299814
rect 297376 299810 297758 299826
rect 297364 299804 297758 299810
rect 297416 299798 297758 299804
rect 297364 299746 297416 299752
rect 209320 299736 209372 299742
rect 208978 299684 209320 299690
rect 208978 299678 209372 299684
rect 208978 299662 209360 299678
rect 213302 299674 213592 299690
rect 213302 299668 213604 299674
rect 213302 299662 213552 299668
rect 213552 299610 213604 299616
rect 208308 299600 208360 299606
rect 208150 299548 208308 299554
rect 217046 299568 217102 299577
rect 208150 299542 208360 299548
rect 208150 299526 208348 299542
rect 216798 299526 217046 299554
rect 217046 299503 217102 299512
rect 218058 299568 218114 299577
rect 218114 299526 218192 299554
rect 293144 299538 293526 299554
rect 218058 299503 218114 299512
rect 216680 299464 216732 299470
rect 216680 299406 216732 299412
rect 218058 299432 218114 299441
rect 216692 299334 216720 299406
rect 218058 299367 218114 299376
rect 218072 299334 218100 299367
rect 218164 299334 218192 299526
rect 293132 299532 293526 299538
rect 293184 299526 293526 299532
rect 293132 299474 293184 299480
rect 220084 299464 220136 299470
rect 218794 299432 218850 299441
rect 220084 299406 220136 299412
rect 237196 299464 237248 299470
rect 237196 299406 237248 299412
rect 218794 299367 218850 299376
rect 218808 299334 218836 299367
rect 220096 299334 220124 299406
rect 237208 299334 237236 299406
rect 216680 299328 216732 299334
rect 217140 299328 217192 299334
rect 216680 299270 216732 299276
rect 217138 299296 217140 299305
rect 218060 299328 218112 299334
rect 217192 299296 217194 299305
rect 218060 299270 218112 299276
rect 218152 299328 218204 299334
rect 218704 299328 218756 299334
rect 218152 299270 218204 299276
rect 218454 299276 218704 299282
rect 218454 299270 218756 299276
rect 218796 299328 218848 299334
rect 219900 299328 219952 299334
rect 218796 299270 218848 299276
rect 219898 299296 219900 299305
rect 220084 299328 220136 299334
rect 219952 299296 219954 299305
rect 218454 299254 218744 299270
rect 217138 299231 217194 299240
rect 220084 299270 220136 299276
rect 237196 299328 237248 299334
rect 237196 299270 237248 299276
rect 242164 299328 242216 299334
rect 242348 299328 242400 299334
rect 242216 299288 242348 299316
rect 242164 299270 242216 299276
rect 242348 299270 242400 299276
rect 283564 299328 283616 299334
rect 284484 299328 284536 299334
rect 283616 299276 283958 299282
rect 283564 299270 283958 299276
rect 286508 299328 286560 299334
rect 284536 299276 284878 299282
rect 284484 299270 284878 299276
rect 299848 299328 299900 299334
rect 286560 299276 286626 299282
rect 286508 299270 286626 299276
rect 283576 299254 283958 299270
rect 284496 299254 284878 299270
rect 286520 299254 286626 299270
rect 299506 299276 299848 299282
rect 299506 299270 299900 299276
rect 299506 299254 299888 299270
rect 219898 299231 219954 299240
rect 199844 298512 199896 298518
rect 199844 298454 199896 298460
rect 199856 296721 199884 298454
rect 199842 296712 199898 296721
rect 199842 296647 199898 296656
rect 199384 215280 199436 215286
rect 199384 215222 199436 215228
rect 198740 122868 198792 122874
rect 198740 122810 198792 122816
rect 198002 122632 198058 122641
rect 198002 122567 198058 122576
rect 197544 121440 197596 121446
rect 197544 121382 197596 121388
rect 197556 120465 197584 121382
rect 197542 120456 197598 120465
rect 197542 120391 197598 120400
rect 198004 119400 198056 119406
rect 198004 119342 198056 119348
rect 197544 117292 197596 117298
rect 197544 117234 197596 117240
rect 197556 116113 197584 117234
rect 197542 116104 197598 116113
rect 197542 116039 197598 116048
rect 197360 114504 197412 114510
rect 197360 114446 197412 114452
rect 197372 113937 197400 114446
rect 197358 113928 197414 113937
rect 197358 113863 197414 113872
rect 197360 111784 197412 111790
rect 197358 111752 197360 111761
rect 197412 111752 197414 111761
rect 197358 111687 197414 111696
rect 198016 109585 198044 119342
rect 198096 118652 198148 118658
rect 198096 118594 198148 118600
rect 198108 118289 198136 118594
rect 198094 118280 198150 118289
rect 198094 118215 198150 118224
rect 198002 109576 198058 109585
rect 198002 109511 198058 109520
rect 198556 107636 198608 107642
rect 198556 107578 198608 107584
rect 198568 107409 198596 107578
rect 198554 107400 198610 107409
rect 198554 107335 198610 107344
rect 197544 106276 197596 106282
rect 197544 106218 197596 106224
rect 197556 105233 197584 106218
rect 197542 105224 197598 105233
rect 197542 105159 197598 105168
rect 197912 103488 197964 103494
rect 197912 103430 197964 103436
rect 197924 103057 197952 103430
rect 197910 103048 197966 103057
rect 197910 102983 197966 102992
rect 197544 102128 197596 102134
rect 197544 102070 197596 102076
rect 197556 101017 197584 102070
rect 197542 101008 197598 101017
rect 197542 100943 197598 100952
rect 299952 100722 299980 337418
rect 359476 305862 359504 699654
rect 371698 369744 371754 369753
rect 371698 369679 371754 369688
rect 371606 368656 371662 368665
rect 371606 368591 371608 368600
rect 371660 368591 371662 368600
rect 371608 368562 371660 368568
rect 371712 368558 371740 369679
rect 371882 369200 371938 369209
rect 371882 369135 371938 369144
rect 371700 368552 371752 368558
rect 371700 368494 371752 368500
rect 371606 368112 371662 368121
rect 371606 368047 371662 368056
rect 371514 367568 371570 367577
rect 371620 367538 371648 368047
rect 371514 367503 371570 367512
rect 371608 367532 371660 367538
rect 371528 367130 371556 367503
rect 371608 367474 371660 367480
rect 371516 367124 371568 367130
rect 371516 367066 371568 367072
rect 371606 367024 371662 367033
rect 371606 366959 371662 366968
rect 371238 365936 371294 365945
rect 371620 365906 371648 366959
rect 371238 365871 371294 365880
rect 371608 365900 371660 365906
rect 371252 365838 371280 365871
rect 371608 365842 371660 365848
rect 371240 365832 371292 365838
rect 371240 365774 371292 365780
rect 371606 365392 371662 365401
rect 371606 365327 371662 365336
rect 371238 364848 371294 364857
rect 371238 364783 371294 364792
rect 371252 364750 371280 364783
rect 371240 364744 371292 364750
rect 371240 364686 371292 364692
rect 371620 364410 371648 365327
rect 371608 364404 371660 364410
rect 371608 364346 371660 364352
rect 371698 364304 371754 364313
rect 371698 364239 371754 364248
rect 371606 363760 371662 363769
rect 371606 363695 371608 363704
rect 371660 363695 371662 363704
rect 371608 363666 371660 363672
rect 371422 363216 371478 363225
rect 371422 363151 371478 363160
rect 371436 363050 371464 363151
rect 371424 363044 371476 363050
rect 371424 362986 371476 362992
rect 371712 362982 371740 364239
rect 371700 362976 371752 362982
rect 371700 362918 371752 362924
rect 371422 362128 371478 362137
rect 371422 362063 371478 362072
rect 371436 361622 371464 362063
rect 371424 361616 371476 361622
rect 371424 361558 371476 361564
rect 371514 361584 371570 361593
rect 371514 361519 371570 361528
rect 371528 360262 371556 361519
rect 371698 361040 371754 361049
rect 371698 360975 371754 360984
rect 371606 360496 371662 360505
rect 371606 360431 371608 360440
rect 371660 360431 371662 360440
rect 371608 360402 371660 360408
rect 371712 360398 371740 360975
rect 371700 360392 371752 360398
rect 371700 360334 371752 360340
rect 371516 360256 371568 360262
rect 371516 360198 371568 360204
rect 371330 360088 371386 360097
rect 371330 360023 371386 360032
rect 371344 358834 371372 360023
rect 371896 359514 371924 369135
rect 376760 368620 376812 368626
rect 376760 368562 376812 368568
rect 374000 367532 374052 367538
rect 374000 367474 374052 367480
rect 372526 366480 372582 366489
rect 372582 366438 372660 366466
rect 372526 366415 372582 366424
rect 372066 359544 372122 359553
rect 371884 359508 371936 359514
rect 372066 359479 372122 359488
rect 371884 359450 371936 359456
rect 371332 358828 371384 358834
rect 371332 358770 371384 358776
rect 371514 358456 371570 358465
rect 371514 358391 371570 358400
rect 371422 357912 371478 357921
rect 371422 357847 371478 357856
rect 371436 357746 371464 357847
rect 371424 357740 371476 357746
rect 371424 357682 371476 357688
rect 371528 357474 371556 358391
rect 371516 357468 371568 357474
rect 371516 357410 371568 357416
rect 371238 357368 371294 357377
rect 371238 357303 371294 357312
rect 371252 356182 371280 357303
rect 371330 356824 371386 356833
rect 371330 356759 371386 356768
rect 371344 356250 371372 356759
rect 371422 356280 371478 356289
rect 371332 356244 371384 356250
rect 371422 356215 371478 356224
rect 371332 356186 371384 356192
rect 371240 356176 371292 356182
rect 371240 356118 371292 356124
rect 371436 356114 371464 356215
rect 371424 356108 371476 356114
rect 371424 356050 371476 356056
rect 371698 355736 371754 355745
rect 371698 355671 371754 355680
rect 371238 355192 371294 355201
rect 371238 355127 371294 355136
rect 371252 355026 371280 355127
rect 371240 355020 371292 355026
rect 371240 354962 371292 354968
rect 371712 354822 371740 355671
rect 371700 354816 371752 354822
rect 371700 354758 371752 354764
rect 371514 354648 371570 354657
rect 371514 354583 371570 354592
rect 371528 354210 371556 354583
rect 371516 354204 371568 354210
rect 371516 354146 371568 354152
rect 371698 354104 371754 354113
rect 371698 354039 371754 354048
rect 371712 353326 371740 354039
rect 371700 353320 371752 353326
rect 371700 353262 371752 353268
rect 372080 352646 372108 359479
rect 372250 359000 372306 359009
rect 372250 358935 372306 358944
rect 372068 352640 372120 352646
rect 372068 352582 372120 352588
rect 372264 352578 372292 358935
rect 372252 352572 372304 352578
rect 372252 352514 372304 352520
rect 371330 351928 371386 351937
rect 371330 351863 371386 351872
rect 370318 349344 370374 349353
rect 370318 349279 370374 349288
rect 369306 348528 369362 348537
rect 369306 348463 369362 348472
rect 369320 345014 369348 348463
rect 370042 346896 370098 346905
rect 370042 346831 370098 346840
rect 369950 345264 370006 345273
rect 369950 345199 370006 345208
rect 369044 344986 369348 345014
rect 360212 340054 360962 340082
rect 359464 305856 359516 305862
rect 359464 305798 359516 305804
rect 316684 303000 316736 303006
rect 316684 302942 316736 302948
rect 304264 301572 304316 301578
rect 304264 301514 304316 301520
rect 301504 301504 301556 301510
rect 301504 301446 301556 301452
rect 300124 299328 300176 299334
rect 300124 299270 300176 299276
rect 300136 266150 300164 299270
rect 300124 266144 300176 266150
rect 300124 266086 300176 266092
rect 300032 265668 300084 265674
rect 300032 265610 300084 265616
rect 299874 100694 299980 100722
rect 300044 100178 300072 265610
rect 301516 167006 301544 301446
rect 302790 298344 302846 298353
rect 302790 298279 302792 298288
rect 302844 298279 302846 298288
rect 302792 298250 302844 298256
rect 303068 296812 303120 296818
rect 303068 296754 303120 296760
rect 302884 296744 302936 296750
rect 302884 296686 302936 296692
rect 302422 295216 302478 295225
rect 302422 295151 302478 295160
rect 302436 294030 302464 295151
rect 302424 294024 302476 294030
rect 302424 293966 302476 293972
rect 302330 291952 302386 291961
rect 302330 291887 302386 291896
rect 302344 291242 302372 291887
rect 302332 291236 302384 291242
rect 302332 291178 302384 291184
rect 302792 285728 302844 285734
rect 302790 285696 302792 285705
rect 302844 285696 302846 285705
rect 302790 285631 302846 285640
rect 302422 282432 302478 282441
rect 302422 282367 302478 282376
rect 302436 281586 302464 282367
rect 302424 281580 302476 281586
rect 302424 281522 302476 281528
rect 302606 279304 302662 279313
rect 302606 279239 302662 279248
rect 302620 278798 302648 279239
rect 302608 278792 302660 278798
rect 302608 278734 302660 278740
rect 302896 272921 302924 296686
rect 302974 288824 303030 288833
rect 302974 288759 303030 288768
rect 302882 272912 302938 272921
rect 302882 272847 302938 272856
rect 302332 270496 302384 270502
rect 302332 270438 302384 270444
rect 302344 269793 302372 270438
rect 302330 269784 302386 269793
rect 302330 269719 302386 269728
rect 302424 267708 302476 267714
rect 302424 267650 302476 267656
rect 302436 266665 302464 267650
rect 302516 267028 302568 267034
rect 302516 266970 302568 266976
rect 302422 266656 302478 266665
rect 302422 266591 302478 266600
rect 302528 263401 302556 266970
rect 302988 266218 303016 288759
rect 303080 276185 303108 296754
rect 303066 276176 303122 276185
rect 303066 276111 303122 276120
rect 302976 266212 303028 266218
rect 302976 266154 303028 266160
rect 302514 263392 302570 263401
rect 302514 263327 302570 263336
rect 302792 260840 302844 260846
rect 302792 260782 302844 260788
rect 302804 260273 302832 260782
rect 302790 260264 302846 260273
rect 302790 260199 302846 260208
rect 302790 257136 302846 257145
rect 302790 257071 302846 257080
rect 302804 256766 302832 257071
rect 302792 256760 302844 256766
rect 302792 256702 302844 256708
rect 302882 253872 302938 253881
rect 302882 253807 302938 253816
rect 302896 247722 302924 253807
rect 303158 250744 303214 250753
rect 303158 250679 303214 250688
rect 302884 247716 302936 247722
rect 302884 247658 302936 247664
rect 303066 247616 303122 247625
rect 303066 247551 303122 247560
rect 302974 244352 303030 244361
rect 302974 244287 303030 244296
rect 302790 241224 302846 241233
rect 302790 241159 302846 241168
rect 302804 229094 302832 241159
rect 302882 231704 302938 231713
rect 302882 231639 302938 231648
rect 302712 229066 302832 229094
rect 302712 224398 302740 229066
rect 302790 228440 302846 228449
rect 302790 228375 302846 228384
rect 302804 225622 302832 228375
rect 302792 225616 302844 225622
rect 302792 225558 302844 225564
rect 302790 225312 302846 225321
rect 302790 225247 302846 225256
rect 302700 224392 302752 224398
rect 302700 224334 302752 224340
rect 302804 224262 302832 225247
rect 302896 224330 302924 231639
rect 302988 229770 303016 244287
rect 303080 235278 303108 247551
rect 303172 240786 303200 250679
rect 304276 245614 304304 301514
rect 309784 301436 309836 301442
rect 309784 301378 309836 301384
rect 307024 300280 307076 300286
rect 307024 300222 307076 300228
rect 305644 300212 305696 300218
rect 305644 300154 305696 300160
rect 304264 245608 304316 245614
rect 304264 245550 304316 245556
rect 303160 240780 303212 240786
rect 303160 240722 303212 240728
rect 303158 238096 303214 238105
rect 303158 238031 303214 238040
rect 303068 235272 303120 235278
rect 303068 235214 303120 235220
rect 302976 229764 303028 229770
rect 302976 229706 303028 229712
rect 303172 228410 303200 238031
rect 303250 234832 303306 234841
rect 303250 234767 303306 234776
rect 303160 228404 303212 228410
rect 303160 228346 303212 228352
rect 303264 225690 303292 234767
rect 303252 225684 303304 225690
rect 303252 225626 303304 225632
rect 302884 224324 302936 224330
rect 302884 224266 302936 224272
rect 302792 224256 302844 224262
rect 302792 224198 302844 224204
rect 302790 222184 302846 222193
rect 302790 222119 302792 222128
rect 302844 222119 302846 222128
rect 302792 222090 302844 222096
rect 302792 219428 302844 219434
rect 302792 219370 302844 219376
rect 302804 218929 302832 219370
rect 302790 218920 302846 218929
rect 302790 218855 302846 218864
rect 302792 216640 302844 216646
rect 302792 216582 302844 216588
rect 302804 215801 302832 216582
rect 302790 215792 302846 215801
rect 302790 215727 302846 215736
rect 302792 213920 302844 213926
rect 302792 213862 302844 213868
rect 302804 212673 302832 213862
rect 302790 212664 302846 212673
rect 302790 212599 302846 212608
rect 302882 209400 302938 209409
rect 302882 209335 302938 209344
rect 302330 206272 302386 206281
rect 302330 206207 302386 206216
rect 302344 205698 302372 206207
rect 302332 205692 302384 205698
rect 302332 205634 302384 205640
rect 302790 203144 302846 203153
rect 302790 203079 302846 203088
rect 302804 202910 302832 203079
rect 302792 202904 302844 202910
rect 302792 202846 302844 202852
rect 302514 199880 302570 199889
rect 302514 199815 302570 199824
rect 302528 198762 302556 199815
rect 302516 198756 302568 198762
rect 302516 198698 302568 198704
rect 302896 197266 302924 209335
rect 302884 197260 302936 197266
rect 302884 197202 302936 197208
rect 302700 197192 302752 197198
rect 302700 197134 302752 197140
rect 302712 196761 302740 197134
rect 302698 196752 302754 196761
rect 302698 196687 302754 196696
rect 302976 196716 303028 196722
rect 302976 196658 303028 196664
rect 302884 195288 302936 195294
rect 302884 195230 302936 195236
rect 302424 194540 302476 194546
rect 302424 194482 302476 194488
rect 302436 193633 302464 194482
rect 302422 193624 302478 193633
rect 302422 193559 302478 193568
rect 302700 187672 302752 187678
rect 302700 187614 302752 187620
rect 302712 187241 302740 187614
rect 302698 187232 302754 187241
rect 302698 187167 302754 187176
rect 302792 184884 302844 184890
rect 302792 184826 302844 184832
rect 302804 184113 302832 184826
rect 302790 184104 302846 184113
rect 302790 184039 302846 184048
rect 302896 177721 302924 195230
rect 302988 180849 303016 196658
rect 303068 196648 303120 196654
rect 303068 196590 303120 196596
rect 303080 190369 303108 196590
rect 303066 190360 303122 190369
rect 303066 190295 303122 190304
rect 302974 180840 303030 180849
rect 302974 180775 303030 180784
rect 302882 177712 302938 177721
rect 302882 177647 302938 177656
rect 302240 175228 302292 175234
rect 302240 175170 302292 175176
rect 302252 174593 302280 175170
rect 302238 174584 302294 174593
rect 302238 174519 302294 174528
rect 302790 171320 302846 171329
rect 302790 171255 302846 171264
rect 302804 171154 302832 171255
rect 302792 171148 302844 171154
rect 302792 171090 302844 171096
rect 302698 168192 302754 168201
rect 302698 168127 302754 168136
rect 301504 167000 301556 167006
rect 301504 166942 301556 166948
rect 302606 164928 302662 164937
rect 302606 164863 302662 164872
rect 302620 161474 302648 164863
rect 302712 162178 302740 168127
rect 302700 162172 302752 162178
rect 302700 162114 302752 162120
rect 302974 161800 303030 161809
rect 302974 161735 303030 161744
rect 302620 161446 302740 161474
rect 302712 152522 302740 161446
rect 302790 158672 302846 158681
rect 302790 158607 302846 158616
rect 302804 154562 302832 158607
rect 302882 155408 302938 155417
rect 302882 155343 302938 155352
rect 302792 154556 302844 154562
rect 302792 154498 302844 154504
rect 302896 153134 302924 155343
rect 302988 153202 303016 161735
rect 302976 153196 303028 153202
rect 302976 153138 303028 153144
rect 302884 153128 302936 153134
rect 302884 153070 302936 153076
rect 302792 153060 302844 153066
rect 302792 153002 302844 153008
rect 302700 152516 302752 152522
rect 302700 152458 302752 152464
rect 302804 152289 302832 153002
rect 302790 152280 302846 152289
rect 302790 152215 302846 152224
rect 302792 150408 302844 150414
rect 302792 150350 302844 150356
rect 302804 149161 302832 150350
rect 302790 149152 302846 149161
rect 302790 149087 302846 149096
rect 302792 146260 302844 146266
rect 302792 146202 302844 146208
rect 302804 145897 302832 146202
rect 302790 145888 302846 145897
rect 302790 145823 302846 145832
rect 302792 143540 302844 143546
rect 302792 143482 302844 143488
rect 302804 142769 302832 143482
rect 302790 142760 302846 142769
rect 302790 142695 302846 142704
rect 302882 139632 302938 139641
rect 302882 139567 302938 139576
rect 302790 130112 302846 130121
rect 302790 130047 302846 130056
rect 302606 126848 302662 126857
rect 302606 126783 302662 126792
rect 302620 124982 302648 126783
rect 302804 125254 302832 130047
rect 302792 125248 302844 125254
rect 302792 125190 302844 125196
rect 302896 125118 302924 139567
rect 302974 136368 303030 136377
rect 302974 136303 303030 136312
rect 302884 125112 302936 125118
rect 302884 125054 302936 125060
rect 302988 125050 303016 136303
rect 303066 133240 303122 133249
rect 303066 133175 303122 133184
rect 303080 125186 303108 133175
rect 303068 125180 303120 125186
rect 303068 125122 303120 125128
rect 302976 125044 303028 125050
rect 302976 124986 303028 124992
rect 302608 124976 302660 124982
rect 302608 124918 302660 124924
rect 302700 124160 302752 124166
rect 302700 124102 302752 124108
rect 302712 123729 302740 124102
rect 302698 123720 302754 123729
rect 302698 123655 302754 123664
rect 302976 123616 303028 123622
rect 302976 123558 303028 123564
rect 302884 123480 302936 123486
rect 302884 123422 302936 123428
rect 302792 121440 302844 121446
rect 302792 121382 302844 121388
rect 302804 120601 302832 121382
rect 302790 120592 302846 120601
rect 302790 120527 302846 120536
rect 302792 118652 302844 118658
rect 302792 118594 302844 118600
rect 302804 117337 302832 118594
rect 302790 117328 302846 117337
rect 302790 117263 302846 117272
rect 302332 111784 302384 111790
rect 302332 111726 302384 111732
rect 302344 111081 302372 111726
rect 302330 111072 302386 111081
rect 302330 111007 302386 111016
rect 302792 108996 302844 109002
rect 302792 108938 302844 108944
rect 302804 107817 302832 108938
rect 302790 107808 302846 107817
rect 302790 107743 302846 107752
rect 302896 104689 302924 123422
rect 302988 114209 303016 123558
rect 302974 114200 303030 114209
rect 302974 114135 303030 114144
rect 302882 104680 302938 104689
rect 302882 104615 302938 104624
rect 302792 102128 302844 102134
rect 302792 102070 302844 102076
rect 302804 101561 302832 102070
rect 302790 101552 302846 101561
rect 302790 101487 302846 101496
rect 299952 100150 300072 100178
rect 200146 100014 200252 100042
rect 200330 100014 200436 100042
rect 196624 99408 196676 99414
rect 196624 99350 196676 99356
rect 191196 97232 191248 97238
rect 191196 97174 191248 97180
rect 188436 97164 188488 97170
rect 188436 97106 188488 97112
rect 176568 96620 176620 96626
rect 176568 96562 176620 96568
rect 161388 96552 161440 96558
rect 161388 96494 161440 96500
rect 159364 94988 159416 94994
rect 159364 94930 159416 94936
rect 155316 94920 155368 94926
rect 155316 94862 155368 94868
rect 155224 33108 155276 33114
rect 155224 33050 155276 33056
rect 155328 3262 155356 94862
rect 156604 92268 156656 92274
rect 156604 92210 156656 92216
rect 156616 3262 156644 92210
rect 157984 89480 158036 89486
rect 157984 89422 158036 89428
rect 154212 3256 154264 3262
rect 154212 3198 154264 3204
rect 155316 3256 155368 3262
rect 155316 3198 155368 3204
rect 155408 3256 155460 3262
rect 155408 3198 155460 3204
rect 156604 3256 156656 3262
rect 156604 3198 156656 3204
rect 153108 3188 153160 3194
rect 153108 3130 153160 3136
rect 154224 480 154252 3198
rect 155420 480 155448 3198
rect 157800 3188 157852 3194
rect 157800 3130 157852 3136
rect 156604 3120 156656 3126
rect 156604 3062 156656 3068
rect 156616 480 156644 3062
rect 157812 480 157840 3130
rect 157996 3126 158024 89422
rect 158904 3256 158956 3262
rect 158904 3198 158956 3204
rect 157984 3120 158036 3126
rect 157984 3062 158036 3068
rect 158916 480 158944 3198
rect 159376 3194 159404 94930
rect 160008 93696 160060 93702
rect 160008 93638 160060 93644
rect 160020 3262 160048 93638
rect 161296 90976 161348 90982
rect 161296 90918 161348 90924
rect 161308 16574 161336 90918
rect 161216 16546 161336 16574
rect 161216 3262 161244 16546
rect 161400 6914 161428 96494
rect 173164 96348 173216 96354
rect 173164 96290 173216 96296
rect 169668 96280 169720 96286
rect 169668 96222 169720 96228
rect 165528 96212 165580 96218
rect 165528 96154 165580 96160
rect 162768 95124 162820 95130
rect 162768 95066 162820 95072
rect 162780 6914 162808 95066
rect 164148 92336 164200 92342
rect 164148 92278 164200 92284
rect 161308 6886 161428 6914
rect 162504 6886 162808 6914
rect 160008 3256 160060 3262
rect 160008 3198 160060 3204
rect 160100 3256 160152 3262
rect 160100 3198 160152 3204
rect 161204 3256 161256 3262
rect 161204 3198 161256 3204
rect 159364 3188 159416 3194
rect 159364 3130 159416 3136
rect 160112 480 160140 3198
rect 161308 480 161336 6886
rect 162504 480 162532 6886
rect 164160 3262 164188 92278
rect 165540 3262 165568 96154
rect 166908 93764 166960 93770
rect 166908 93706 166960 93712
rect 166920 3262 166948 93706
rect 169024 92404 169076 92410
rect 169024 92346 169076 92352
rect 169036 3262 169064 92346
rect 163688 3256 163740 3262
rect 163688 3198 163740 3204
rect 164148 3256 164200 3262
rect 164148 3198 164200 3204
rect 164884 3256 164936 3262
rect 164884 3198 164936 3204
rect 165528 3256 165580 3262
rect 165528 3198 165580 3204
rect 166080 3256 166132 3262
rect 166080 3198 166132 3204
rect 166908 3256 166960 3262
rect 166908 3198 166960 3204
rect 167184 3256 167236 3262
rect 167184 3198 167236 3204
rect 169024 3256 169076 3262
rect 169024 3198 169076 3204
rect 163700 480 163728 3198
rect 164896 480 164924 3198
rect 166092 480 166120 3198
rect 167196 480 167224 3198
rect 169576 3188 169628 3194
rect 169576 3130 169628 3136
rect 168380 3120 168432 3126
rect 168380 3062 168432 3068
rect 168392 480 168420 3062
rect 169588 480 169616 3130
rect 169680 3126 169708 96222
rect 171048 95192 171100 95198
rect 171048 95134 171100 95140
rect 170404 93832 170456 93838
rect 170404 93774 170456 93780
rect 170416 3194 170444 93774
rect 171060 6914 171088 95134
rect 173176 6914 173204 96290
rect 173808 94444 173860 94450
rect 173808 94386 173860 94392
rect 170784 6886 171088 6914
rect 173084 6886 173204 6914
rect 170404 3188 170456 3194
rect 170404 3130 170456 3136
rect 169668 3120 169720 3126
rect 169668 3062 169720 3068
rect 170784 480 170812 6886
rect 173084 3126 173112 6886
rect 173820 3262 173848 94386
rect 175188 92472 175240 92478
rect 175188 92414 175240 92420
rect 175200 3262 175228 92414
rect 176580 3262 176608 96562
rect 183468 96484 183520 96490
rect 183468 96426 183520 96432
rect 179328 96416 179380 96422
rect 179328 96358 179380 96364
rect 177948 93084 178000 93090
rect 177948 93026 178000 93032
rect 177856 91044 177908 91050
rect 177856 90986 177908 90992
rect 173164 3256 173216 3262
rect 173164 3198 173216 3204
rect 173808 3256 173860 3262
rect 173808 3198 173860 3204
rect 174268 3256 174320 3262
rect 174268 3198 174320 3204
rect 175188 3256 175240 3262
rect 175188 3198 175240 3204
rect 175464 3256 175516 3262
rect 175464 3198 175516 3204
rect 176568 3256 176620 3262
rect 176568 3198 176620 3204
rect 176660 3256 176712 3262
rect 176660 3198 176712 3204
rect 171968 3120 172020 3126
rect 171968 3062 172020 3068
rect 173072 3120 173124 3126
rect 173072 3062 173124 3068
rect 171980 480 172008 3062
rect 173176 480 173204 3198
rect 174280 480 174308 3198
rect 175476 480 175504 3198
rect 176672 480 176700 3198
rect 177868 480 177896 90986
rect 177960 3262 177988 93026
rect 179340 6914 179368 96358
rect 180708 93016 180760 93022
rect 180708 92958 180760 92964
rect 179064 6886 179368 6914
rect 177948 3256 178000 3262
rect 177948 3198 178000 3204
rect 179064 480 179092 6886
rect 180720 3262 180748 92958
rect 182088 91724 182140 91730
rect 182088 91666 182140 91672
rect 182100 3262 182128 91666
rect 183480 3262 183508 96426
rect 186964 95872 187016 95878
rect 186964 95814 187016 95820
rect 184848 92948 184900 92954
rect 184848 92890 184900 92896
rect 184860 3262 184888 92890
rect 186976 3262 187004 95814
rect 188344 94376 188396 94382
rect 188344 94318 188396 94324
rect 187332 6316 187384 6322
rect 187332 6258 187384 6264
rect 180248 3256 180300 3262
rect 180248 3198 180300 3204
rect 180708 3256 180760 3262
rect 180708 3198 180760 3204
rect 181444 3256 181496 3262
rect 181444 3198 181496 3204
rect 182088 3256 182140 3262
rect 182088 3198 182140 3204
rect 182548 3256 182600 3262
rect 182548 3198 182600 3204
rect 183468 3256 183520 3262
rect 183468 3198 183520 3204
rect 183744 3256 183796 3262
rect 183744 3198 183796 3204
rect 184848 3256 184900 3262
rect 184848 3198 184900 3204
rect 186136 3256 186188 3262
rect 186136 3198 186188 3204
rect 186964 3256 187016 3262
rect 186964 3198 187016 3204
rect 180260 480 180288 3198
rect 181456 480 181484 3198
rect 182560 480 182588 3198
rect 183756 480 183784 3198
rect 184940 2916 184992 2922
rect 184940 2858 184992 2864
rect 184952 480 184980 2858
rect 186148 480 186176 3198
rect 187344 480 187372 6258
rect 188356 2922 188384 94318
rect 188448 7614 188476 97106
rect 191104 95804 191156 95810
rect 191104 95746 191156 95752
rect 188436 7608 188488 7614
rect 188436 7550 188488 7556
rect 188528 7608 188580 7614
rect 188528 7550 188580 7556
rect 188344 2916 188396 2922
rect 188344 2858 188396 2864
rect 188540 480 188568 7550
rect 190828 6384 190880 6390
rect 190828 6326 190880 6332
rect 189724 3256 189776 3262
rect 189724 3198 189776 3204
rect 189736 480 189764 3198
rect 190840 480 190868 6326
rect 191116 3262 191144 95746
rect 191208 86562 191236 97174
rect 196624 97096 196676 97102
rect 196624 97038 196676 97044
rect 194508 95600 194560 95606
rect 194508 95542 194560 95548
rect 191196 86556 191248 86562
rect 191196 86498 191248 86504
rect 192024 7744 192076 7750
rect 192024 7686 192076 7692
rect 191104 3256 191156 3262
rect 191104 3198 191156 3204
rect 192036 480 192064 7686
rect 194416 6452 194468 6458
rect 194416 6394 194468 6400
rect 193128 3528 193180 3534
rect 193128 3470 193180 3476
rect 193220 3528 193272 3534
rect 193220 3470 193272 3476
rect 193140 3262 193168 3470
rect 193128 3256 193180 3262
rect 193128 3198 193180 3204
rect 193232 480 193260 3470
rect 194428 480 194456 6394
rect 194520 3534 194548 95542
rect 195888 92880 195940 92886
rect 195888 92822 195940 92828
rect 195900 6914 195928 92822
rect 196636 14482 196664 97038
rect 199384 97028 199436 97034
rect 199384 96970 199436 96976
rect 198004 96688 198056 96694
rect 198004 96630 198056 96636
rect 197268 95736 197320 95742
rect 197268 95678 197320 95684
rect 196624 14476 196676 14482
rect 196624 14418 196676 14424
rect 195624 6886 195928 6914
rect 194508 3528 194560 3534
rect 194508 3470 194560 3476
rect 195624 480 195652 6886
rect 197280 3534 197308 95678
rect 198016 84862 198044 96630
rect 198648 94240 198700 94246
rect 198648 94182 198700 94188
rect 198004 84856 198056 84862
rect 198004 84798 198056 84804
rect 198660 3534 198688 94182
rect 199396 89214 199424 96970
rect 200028 95668 200080 95674
rect 200028 95610 200080 95616
rect 199844 94512 199896 94518
rect 199844 94454 199896 94460
rect 199856 94178 199884 94454
rect 199844 94172 199896 94178
rect 199844 94114 199896 94120
rect 199384 89208 199436 89214
rect 199384 89150 199436 89156
rect 199936 24132 199988 24138
rect 199936 24074 199988 24080
rect 199948 3534 199976 24074
rect 200040 4026 200068 95610
rect 200224 94518 200252 100014
rect 200212 94512 200264 94518
rect 200212 94454 200264 94460
rect 200212 94308 200264 94314
rect 200212 94250 200264 94256
rect 200224 16574 200252 94250
rect 200224 16546 200344 16574
rect 200316 4706 200344 16546
rect 200408 4894 200436 100014
rect 200500 4962 200528 100028
rect 200580 94512 200632 94518
rect 200580 94454 200632 94460
rect 200488 4956 200540 4962
rect 200488 4898 200540 4904
rect 200396 4888 200448 4894
rect 200396 4830 200448 4836
rect 200592 4826 200620 94454
rect 200580 4820 200632 4826
rect 200580 4762 200632 4768
rect 200316 4678 200436 4706
rect 200040 3998 200344 4026
rect 200028 3664 200080 3670
rect 200028 3606 200080 3612
rect 200040 3534 200068 3606
rect 196808 3528 196860 3534
rect 196808 3470 196860 3476
rect 197268 3528 197320 3534
rect 197268 3470 197320 3476
rect 197912 3528 197964 3534
rect 197912 3470 197964 3476
rect 198648 3528 198700 3534
rect 198648 3470 198700 3476
rect 199108 3528 199160 3534
rect 199108 3470 199160 3476
rect 199936 3528 199988 3534
rect 199936 3470 199988 3476
rect 200028 3528 200080 3534
rect 200028 3470 200080 3476
rect 196820 480 196848 3470
rect 197924 480 197952 3470
rect 199120 480 199148 3470
rect 200316 480 200344 3998
rect 200408 3602 200436 4678
rect 200396 3596 200448 3602
rect 200396 3538 200448 3544
rect 200684 3466 200712 100028
rect 200868 96694 200896 100028
rect 200960 100014 201066 100042
rect 201144 100014 201342 100042
rect 201526 100014 201632 100042
rect 200856 96688 200908 96694
rect 200856 96630 200908 96636
rect 200960 84194 200988 100014
rect 201144 94314 201172 100014
rect 201132 94308 201184 94314
rect 201132 94250 201184 94256
rect 201604 93158 201632 100014
rect 201592 93152 201644 93158
rect 201592 93094 201644 93100
rect 201696 87650 201724 100028
rect 201776 94512 201828 94518
rect 201776 94454 201828 94460
rect 201684 87644 201736 87650
rect 201684 87586 201736 87592
rect 200776 84166 200988 84194
rect 200672 3460 200724 3466
rect 200672 3402 200724 3408
rect 200776 3262 200804 84166
rect 201788 3602 201816 94454
rect 201880 86290 201908 100028
rect 202064 95946 202092 100028
rect 202156 100014 202354 100042
rect 202156 99374 202184 100014
rect 202156 99346 202276 99374
rect 202144 96688 202196 96694
rect 202144 96630 202196 96636
rect 202052 95940 202104 95946
rect 202052 95882 202104 95888
rect 201868 86284 201920 86290
rect 201868 86226 201920 86232
rect 202156 26926 202184 96630
rect 202248 90370 202276 99346
rect 202524 97850 202552 100028
rect 202616 100014 202722 100042
rect 202512 97844 202564 97850
rect 202512 97786 202564 97792
rect 202616 94518 202644 100014
rect 202892 98666 202920 100028
rect 203076 98802 203104 100028
rect 203064 98796 203116 98802
rect 203064 98738 203116 98744
rect 202880 98660 202932 98666
rect 202880 98602 202932 98608
rect 202788 97844 202840 97850
rect 202788 97786 202840 97792
rect 202604 94512 202656 94518
rect 202604 94454 202656 94460
rect 202236 90364 202288 90370
rect 202236 90306 202288 90312
rect 202144 26920 202196 26926
rect 202144 26862 202196 26868
rect 202800 6914 202828 97786
rect 203352 97306 203380 100028
rect 203536 97481 203564 100028
rect 203522 97472 203578 97481
rect 203522 97407 203578 97416
rect 203340 97300 203392 97306
rect 203340 97242 203392 97248
rect 203720 94178 203748 100028
rect 203812 100014 203918 100042
rect 203708 94172 203760 94178
rect 203708 94114 203760 94120
rect 203812 94058 203840 100014
rect 204088 97578 204116 100028
rect 204378 100014 204484 100042
rect 204076 97572 204128 97578
rect 204076 97514 204128 97520
rect 204168 97300 204220 97306
rect 204168 97242 204220 97248
rect 203892 96892 203944 96898
rect 203892 96834 203944 96840
rect 203168 94030 203840 94058
rect 203168 11762 203196 94030
rect 203904 89714 203932 96834
rect 203536 89686 203932 89714
rect 203536 87718 203564 89686
rect 203524 87712 203576 87718
rect 203524 87654 203576 87660
rect 203156 11756 203208 11762
rect 203156 11698 203208 11704
rect 204180 6914 204208 97242
rect 204260 96960 204312 96966
rect 204260 96902 204312 96908
rect 204272 91798 204300 96902
rect 204456 96098 204484 100014
rect 204548 98734 204576 100028
rect 204536 98728 204588 98734
rect 204536 98670 204588 98676
rect 204456 96070 204576 96098
rect 204444 94512 204496 94518
rect 204444 94454 204496 94460
rect 204260 91792 204312 91798
rect 204260 91734 204312 91740
rect 204456 11898 204484 94454
rect 204548 89714 204576 96070
rect 204548 89686 204668 89714
rect 204444 11892 204496 11898
rect 204444 11834 204496 11840
rect 202708 6886 202828 6914
rect 203904 6886 204208 6914
rect 201776 3596 201828 3602
rect 201776 3538 201828 3544
rect 201500 3528 201552 3534
rect 201500 3470 201552 3476
rect 200764 3256 200816 3262
rect 200764 3198 200816 3204
rect 201512 480 201540 3470
rect 202708 480 202736 6886
rect 203904 480 203932 6886
rect 204640 3738 204668 89686
rect 204732 11830 204760 100028
rect 204916 97209 204944 100028
rect 205008 100014 205114 100042
rect 205192 100014 205298 100042
rect 204902 97200 204958 97209
rect 204902 97135 204958 97144
rect 205008 93226 205036 100014
rect 205192 94518 205220 100014
rect 205560 96694 205588 100028
rect 205548 96688 205600 96694
rect 205548 96630 205600 96636
rect 205180 94512 205232 94518
rect 205180 94454 205232 94460
rect 204996 93220 205048 93226
rect 204996 93162 205048 93168
rect 205744 89010 205772 100028
rect 205928 98870 205956 100028
rect 205916 98864 205968 98870
rect 205916 98806 205968 98812
rect 206112 97617 206140 100028
rect 206204 100014 206310 100042
rect 206098 97608 206154 97617
rect 206098 97543 206154 97552
rect 206204 89714 206232 100014
rect 206572 97345 206600 100028
rect 206756 97374 206784 100028
rect 206848 100014 206954 100042
rect 207138 100014 207244 100042
rect 206744 97368 206796 97374
rect 206558 97336 206614 97345
rect 206744 97310 206796 97316
rect 206558 97271 206614 97280
rect 205836 89686 206232 89714
rect 205836 89146 205864 89686
rect 205824 89140 205876 89146
rect 205824 89082 205876 89088
rect 205732 89004 205784 89010
rect 205732 88946 205784 88952
rect 206848 87786 206876 100014
rect 207216 89078 207244 100014
rect 207308 97170 207336 100028
rect 207400 100014 207598 100042
rect 207296 97164 207348 97170
rect 207296 97106 207348 97112
rect 207204 89072 207256 89078
rect 207204 89014 207256 89020
rect 206836 87780 206888 87786
rect 206836 87722 206888 87728
rect 204720 11824 204772 11830
rect 204720 11766 204772 11772
rect 205088 6520 205140 6526
rect 205088 6462 205140 6468
rect 204628 3732 204680 3738
rect 204628 3674 204680 3680
rect 205100 480 205128 6462
rect 207400 3806 207428 100014
rect 207768 96966 207796 100028
rect 207756 96960 207808 96966
rect 207756 96902 207808 96908
rect 207952 96898 207980 100028
rect 208044 100014 208150 100042
rect 208228 100014 208334 100042
rect 207940 96892 207992 96898
rect 207940 96834 207992 96840
rect 208044 84194 208072 100014
rect 208228 90438 208256 100014
rect 208308 97368 208360 97374
rect 208308 97310 208360 97316
rect 208320 96558 208348 97310
rect 208308 96552 208360 96558
rect 208308 96494 208360 96500
rect 208216 90432 208268 90438
rect 208216 90374 208268 90380
rect 208596 89714 208624 100028
rect 208688 100014 208794 100042
rect 208688 96014 208716 100014
rect 208676 96008 208728 96014
rect 208676 95950 208728 95956
rect 208596 89686 208900 89714
rect 208872 86426 208900 89686
rect 208860 86420 208912 86426
rect 208860 86362 208912 86368
rect 208964 84194 208992 100028
rect 209148 97034 209176 100028
rect 209240 100014 209346 100042
rect 209424 100014 209622 100042
rect 209136 97028 209188 97034
rect 209136 96970 209188 96976
rect 209044 96688 209096 96694
rect 209044 96630 209096 96636
rect 207860 84166 208072 84194
rect 208688 84166 208992 84194
rect 207860 5030 207888 84166
rect 208584 6248 208636 6254
rect 208584 6190 208636 6196
rect 207848 5024 207900 5030
rect 207848 4966 207900 4972
rect 207388 3800 207440 3806
rect 207388 3742 207440 3748
rect 207388 3596 207440 3602
rect 207388 3538 207440 3544
rect 206192 3460 206244 3466
rect 206192 3402 206244 3408
rect 206204 480 206232 3402
rect 207400 480 207428 3538
rect 208596 480 208624 6190
rect 208688 3874 208716 84166
rect 209056 6186 209084 96630
rect 209240 93294 209268 100014
rect 209228 93288 209280 93294
rect 209228 93230 209280 93236
rect 209424 87854 209452 100014
rect 209792 99142 209820 100028
rect 209884 100014 209990 100042
rect 210068 100014 210174 100042
rect 209780 99136 209832 99142
rect 209780 99078 209832 99084
rect 209412 87848 209464 87854
rect 209412 87790 209464 87796
rect 209044 6180 209096 6186
rect 209044 6122 209096 6128
rect 209884 5098 209912 100014
rect 210068 10334 210096 100014
rect 210344 98938 210372 100028
rect 210332 98932 210384 98938
rect 210332 98874 210384 98880
rect 210240 97776 210292 97782
rect 210240 97718 210292 97724
rect 210252 97102 210280 97718
rect 210240 97096 210292 97102
rect 210240 97038 210292 97044
rect 210528 95266 210556 100028
rect 210620 100014 210818 100042
rect 210516 95260 210568 95266
rect 210516 95202 210568 95208
rect 210620 91780 210648 100014
rect 210884 97912 210936 97918
rect 210884 97854 210936 97860
rect 210896 97782 210924 97854
rect 210884 97776 210936 97782
rect 210884 97718 210936 97724
rect 210988 97170 211016 100028
rect 211172 98326 211200 100028
rect 211264 100014 211370 100042
rect 211160 98320 211212 98326
rect 211160 98262 211212 98268
rect 210976 97164 211028 97170
rect 210976 97106 211028 97112
rect 211160 97164 211212 97170
rect 211160 97106 211212 97112
rect 211172 96150 211200 97106
rect 211160 96144 211212 96150
rect 211160 96086 211212 96092
rect 210700 95260 210752 95266
rect 210700 95202 210752 95208
rect 210252 91752 210648 91780
rect 210056 10328 210108 10334
rect 210056 10270 210108 10276
rect 209872 5092 209924 5098
rect 209872 5034 209924 5040
rect 210252 3942 210280 91752
rect 210712 86954 210740 95202
rect 211264 87922 211292 100014
rect 211540 99210 211568 100028
rect 211724 100014 211830 100042
rect 211528 99204 211580 99210
rect 211528 99146 211580 99152
rect 211436 98320 211488 98326
rect 211436 98262 211488 98268
rect 211620 98320 211672 98326
rect 211620 98262 211672 98268
rect 211448 91866 211476 98262
rect 211436 91860 211488 91866
rect 211436 91802 211488 91808
rect 211252 87916 211304 87922
rect 211252 87858 211304 87864
rect 210528 86926 210740 86954
rect 210528 6118 210556 86926
rect 211632 86358 211660 98262
rect 211724 91934 211752 100014
rect 212000 98326 212028 100028
rect 211988 98320 212040 98326
rect 211988 98262 212040 98268
rect 212184 96694 212212 100028
rect 212276 100014 212382 100042
rect 212566 100014 212764 100042
rect 212172 96688 212224 96694
rect 212172 96630 212224 96636
rect 211712 91928 211764 91934
rect 211712 91870 211764 91876
rect 212276 90506 212304 100014
rect 212540 97504 212592 97510
rect 212540 97446 212592 97452
rect 212552 95062 212580 97446
rect 212540 95056 212592 95062
rect 212540 94998 212592 95004
rect 212736 94518 212764 100014
rect 212828 94586 212856 100028
rect 212816 94580 212868 94586
rect 212816 94522 212868 94528
rect 212908 94580 212960 94586
rect 212908 94522 212960 94528
rect 212724 94512 212776 94518
rect 212724 94454 212776 94460
rect 212632 94240 212684 94246
rect 212632 94182 212684 94188
rect 212264 90500 212316 90506
rect 212264 90442 212316 90448
rect 211620 86352 211672 86358
rect 211620 86294 211672 86300
rect 212644 9042 212672 94182
rect 212724 94172 212776 94178
rect 212724 94114 212776 94120
rect 212736 10538 212764 94114
rect 212724 10532 212776 10538
rect 212724 10474 212776 10480
rect 212920 10470 212948 94522
rect 212908 10464 212960 10470
rect 212908 10406 212960 10412
rect 212632 9036 212684 9042
rect 212632 8978 212684 8984
rect 213012 8974 213040 100028
rect 213104 100014 213210 100042
rect 213104 94586 213132 100014
rect 213380 99278 213408 100028
rect 213472 100014 213578 100042
rect 213656 100014 213854 100042
rect 214038 100014 214144 100042
rect 213368 99272 213420 99278
rect 213368 99214 213420 99220
rect 213092 94580 213144 94586
rect 213092 94522 213144 94528
rect 213276 94512 213328 94518
rect 213276 94454 213328 94460
rect 213288 10402 213316 94454
rect 213472 94246 213500 100014
rect 213460 94240 213512 94246
rect 213460 94182 213512 94188
rect 213656 94178 213684 100014
rect 213920 97436 213972 97442
rect 213920 97378 213972 97384
rect 213932 95606 213960 97378
rect 213920 95600 213972 95606
rect 213920 95542 213972 95548
rect 213644 94172 213696 94178
rect 213644 94114 213696 94120
rect 214116 89282 214144 100014
rect 214208 92002 214236 100028
rect 214392 99006 214420 100028
rect 214484 100014 214590 100042
rect 214668 100014 214774 100042
rect 214852 100014 215050 100042
rect 215128 100014 215234 100042
rect 214380 99000 214432 99006
rect 214380 98942 214432 98948
rect 214484 96762 214512 100014
rect 214472 96756 214524 96762
rect 214472 96698 214524 96704
rect 214196 91996 214248 92002
rect 214196 91938 214248 91944
rect 214668 90574 214696 100014
rect 214656 90568 214708 90574
rect 214656 90510 214708 90516
rect 214852 89714 214880 100014
rect 214300 89686 214880 89714
rect 214104 89276 214156 89282
rect 214104 89218 214156 89224
rect 214300 10606 214328 89686
rect 215128 86494 215156 100014
rect 215404 99074 215432 100028
rect 215496 100014 215602 100042
rect 215392 99068 215444 99074
rect 215392 99010 215444 99016
rect 215116 86488 215168 86494
rect 215116 86430 215168 86436
rect 215496 10674 215524 100014
rect 215772 97646 215800 100028
rect 215864 100014 216062 100042
rect 216246 100014 216352 100042
rect 215760 97640 215812 97646
rect 215760 97582 215812 97588
rect 215864 89714 215892 100014
rect 216036 98320 216088 98326
rect 216036 98262 216088 98268
rect 215944 96756 215996 96762
rect 215944 96698 215996 96704
rect 215680 89686 215892 89714
rect 215484 10668 215536 10674
rect 215484 10610 215536 10616
rect 214288 10600 214340 10606
rect 214288 10542 214340 10548
rect 213276 10396 213328 10402
rect 213276 10338 213328 10344
rect 215680 9110 215708 89686
rect 215668 9104 215720 9110
rect 215668 9046 215720 9052
rect 213000 8968 213052 8974
rect 213000 8910 213052 8916
rect 215668 6588 215720 6594
rect 215668 6530 215720 6536
rect 212172 6180 212224 6186
rect 212172 6122 212224 6128
rect 210516 6112 210568 6118
rect 210516 6054 210568 6060
rect 210976 4820 211028 4826
rect 210976 4762 211028 4768
rect 210240 3936 210292 3942
rect 210240 3878 210292 3884
rect 208676 3868 208728 3874
rect 208676 3810 208728 3816
rect 209780 3664 209832 3670
rect 209780 3606 209832 3612
rect 209792 480 209820 3606
rect 210988 480 211016 4762
rect 212184 480 212212 6122
rect 214472 4888 214524 4894
rect 214472 4830 214524 4836
rect 213368 3732 213420 3738
rect 213368 3674 213420 3680
rect 213380 480 213408 3674
rect 214484 480 214512 4830
rect 215680 480 215708 6530
rect 215956 4010 215984 96698
rect 216048 90642 216076 98262
rect 216128 94580 216180 94586
rect 216128 94522 216180 94528
rect 216036 90636 216088 90642
rect 216036 90578 216088 90584
rect 216140 9178 216168 94522
rect 216324 89714 216352 100014
rect 216416 98326 216444 100028
rect 216508 100014 216614 100042
rect 216798 100014 216904 100042
rect 216404 98320 216456 98326
rect 216404 98262 216456 98268
rect 216508 94586 216536 100014
rect 216496 94580 216548 94586
rect 216496 94522 216548 94528
rect 216232 89686 216352 89714
rect 216232 10742 216260 89686
rect 216876 11966 216904 100014
rect 217060 97578 217088 100028
rect 217048 97572 217100 97578
rect 217048 97514 217100 97520
rect 216956 94580 217008 94586
rect 216956 94522 217008 94528
rect 216968 12034 216996 94522
rect 217140 94512 217192 94518
rect 217140 94454 217192 94460
rect 216956 12028 217008 12034
rect 216956 11970 217008 11976
rect 216864 11960 216916 11966
rect 216864 11902 216916 11908
rect 216220 10736 216272 10742
rect 216220 10678 216272 10684
rect 217152 9314 217180 94454
rect 217140 9308 217192 9314
rect 217140 9250 217192 9256
rect 217244 9246 217272 100028
rect 217336 100014 217442 100042
rect 217336 94586 217364 100014
rect 217612 99346 217640 100028
rect 217704 100014 217810 100042
rect 217600 99340 217652 99346
rect 217600 99282 217652 99288
rect 217416 96688 217468 96694
rect 217416 96630 217468 96636
rect 217324 94580 217376 94586
rect 217324 94522 217376 94528
rect 217428 84194 217456 96630
rect 217704 94518 217732 100014
rect 217692 94512 217744 94518
rect 217692 94454 217744 94460
rect 218072 94246 218100 100028
rect 218256 97238 218284 100028
rect 218348 100014 218454 100042
rect 218638 100014 218744 100042
rect 218244 97232 218296 97238
rect 218244 97174 218296 97180
rect 218348 94602 218376 100014
rect 218164 94574 218376 94602
rect 218520 94580 218572 94586
rect 218060 94240 218112 94246
rect 218060 94182 218112 94188
rect 217336 84166 217456 84194
rect 217232 9240 217284 9246
rect 217232 9182 217284 9188
rect 216128 9172 216180 9178
rect 216128 9114 216180 9120
rect 217336 4078 217364 84166
rect 218164 9382 218192 94574
rect 218520 94522 218572 94528
rect 218336 94240 218388 94246
rect 218336 94182 218388 94188
rect 218348 12102 218376 94182
rect 218336 12096 218388 12102
rect 218336 12038 218388 12044
rect 218532 9450 218560 94522
rect 218716 84194 218744 100014
rect 218808 96762 218836 100028
rect 218900 100014 219098 100042
rect 219176 100014 219282 100042
rect 218796 96756 218848 96762
rect 218796 96698 218848 96704
rect 218900 94586 218928 100014
rect 218888 94580 218940 94586
rect 218888 94522 218940 94528
rect 219176 84194 219204 100014
rect 219452 97714 219480 100028
rect 219440 97708 219492 97714
rect 219440 97650 219492 97656
rect 219440 96756 219492 96762
rect 219440 96698 219492 96704
rect 219452 93430 219480 96698
rect 219440 93424 219492 93430
rect 219440 93366 219492 93372
rect 219636 90710 219664 100028
rect 219716 94580 219768 94586
rect 219716 94522 219768 94528
rect 219624 90704 219676 90710
rect 219624 90646 219676 90652
rect 218624 84166 218744 84194
rect 218900 84166 219204 84194
rect 218624 12170 218652 84166
rect 218900 12238 218928 84166
rect 219728 13122 219756 94522
rect 219820 87990 219848 100028
rect 220004 96694 220032 100028
rect 220176 97504 220228 97510
rect 220176 97446 220228 97452
rect 219992 96688 220044 96694
rect 219992 96630 220044 96636
rect 220188 96626 220216 97446
rect 220176 96620 220228 96626
rect 220176 96562 220228 96568
rect 220280 89350 220308 100028
rect 220372 100014 220478 100042
rect 220372 94586 220400 100014
rect 220648 94654 220676 100028
rect 220846 100014 220952 100042
rect 221030 100014 221228 100042
rect 220636 94648 220688 94654
rect 220636 94590 220688 94596
rect 220924 94586 220952 100014
rect 220360 94580 220412 94586
rect 220360 94522 220412 94528
rect 220912 94580 220964 94586
rect 220912 94522 220964 94528
rect 221096 94512 221148 94518
rect 221096 94454 221148 94460
rect 220268 89344 220320 89350
rect 220268 89286 220320 89292
rect 219808 87984 219860 87990
rect 219808 87926 219860 87932
rect 219716 13116 219768 13122
rect 219716 13058 219768 13064
rect 218888 12232 218940 12238
rect 218888 12174 218940 12180
rect 218612 12164 218664 12170
rect 218612 12106 218664 12112
rect 220452 10328 220504 10334
rect 220452 10270 220504 10276
rect 218520 9444 218572 9450
rect 218520 9386 218572 9392
rect 218152 9376 218204 9382
rect 218152 9318 218204 9324
rect 218060 4956 218112 4962
rect 218060 4898 218112 4904
rect 217324 4072 217376 4078
rect 217324 4014 217376 4020
rect 215944 4004 215996 4010
rect 215944 3946 215996 3952
rect 216864 3800 216916 3806
rect 216864 3742 216916 3748
rect 216876 480 216904 3742
rect 218072 480 218100 4898
rect 219256 3868 219308 3874
rect 219256 3810 219308 3816
rect 219268 480 219296 3810
rect 220464 480 220492 10270
rect 221108 4146 221136 94454
rect 221200 88058 221228 100014
rect 221292 97102 221320 100028
rect 221476 97782 221504 100028
rect 221464 97776 221516 97782
rect 221464 97718 221516 97724
rect 221280 97096 221332 97102
rect 221280 97038 221332 97044
rect 221660 94722 221688 100028
rect 221752 100014 221858 100042
rect 221936 100014 222042 100042
rect 221648 94716 221700 94722
rect 221648 94658 221700 94664
rect 221556 94580 221608 94586
rect 221556 94522 221608 94528
rect 221568 89418 221596 94522
rect 221752 92070 221780 100014
rect 221936 94518 221964 100014
rect 222200 96688 222252 96694
rect 222200 96630 222252 96636
rect 221924 94512 221976 94518
rect 221924 94454 221976 94460
rect 222212 93498 222240 96630
rect 222304 96082 222332 100028
rect 222292 96076 222344 96082
rect 222292 96018 222344 96024
rect 222200 93492 222252 93498
rect 222200 93434 222252 93440
rect 221740 92064 221792 92070
rect 221740 92006 221792 92012
rect 221556 89412 221608 89418
rect 221556 89354 221608 89360
rect 221188 88052 221240 88058
rect 221188 87994 221240 88000
rect 222488 5166 222516 100028
rect 222672 97170 222700 100028
rect 222764 100014 222870 100042
rect 222660 97164 222712 97170
rect 222660 97106 222712 97112
rect 222764 93362 222792 100014
rect 223040 96762 223068 100028
rect 223028 96756 223080 96762
rect 223028 96698 223080 96704
rect 223316 94790 223344 100028
rect 223408 100014 223514 100042
rect 223698 100014 223804 100042
rect 223304 94784 223356 94790
rect 223304 94726 223356 94732
rect 222752 93356 222804 93362
rect 222752 93298 222804 93304
rect 223408 92138 223436 100014
rect 223580 96960 223632 96966
rect 223580 96902 223632 96908
rect 223592 92206 223620 96902
rect 223580 92200 223632 92206
rect 223580 92142 223632 92148
rect 223396 92132 223448 92138
rect 223396 92074 223448 92080
rect 223776 90778 223804 100014
rect 223764 90772 223816 90778
rect 223764 90714 223816 90720
rect 222752 8356 222804 8362
rect 222752 8298 222804 8304
rect 222476 5160 222528 5166
rect 222476 5102 222528 5108
rect 221556 5024 221608 5030
rect 221556 4966 221608 4972
rect 221096 4140 221148 4146
rect 221096 4082 221148 4088
rect 221568 480 221596 4966
rect 222764 480 222792 8298
rect 223764 3936 223816 3942
rect 223764 3878 223816 3884
rect 223776 3534 223804 3878
rect 223764 3528 223816 3534
rect 223764 3470 223816 3476
rect 223868 3398 223896 100028
rect 224052 96694 224080 100028
rect 224144 100014 224250 100042
rect 224040 96688 224092 96694
rect 224040 96630 224092 96636
rect 224144 90846 224172 100014
rect 224512 94858 224540 100028
rect 224604 100014 224710 100042
rect 224788 100014 224894 100042
rect 224500 94852 224552 94858
rect 224500 94794 224552 94800
rect 224604 93566 224632 100014
rect 224592 93560 224644 93566
rect 224592 93502 224644 93508
rect 224132 90840 224184 90846
rect 224132 90782 224184 90788
rect 224788 89714 224816 100014
rect 225064 97578 225092 100028
rect 225052 97572 225104 97578
rect 225052 97514 225104 97520
rect 225248 96966 225276 100028
rect 225524 97986 225552 100028
rect 225616 100014 225722 100042
rect 225800 100014 225906 100042
rect 225984 100014 226090 100042
rect 225512 97980 225564 97986
rect 225512 97922 225564 97928
rect 225236 96960 225288 96966
rect 225236 96902 225288 96908
rect 224868 91792 224920 91798
rect 224868 91734 224920 91740
rect 224144 89686 224816 89714
rect 224144 7682 224172 89686
rect 224132 7676 224184 7682
rect 224132 7618 224184 7624
rect 224880 3534 224908 91734
rect 225616 89714 225644 100014
rect 225800 93634 225828 100014
rect 225788 93628 225840 93634
rect 225788 93570 225840 93576
rect 225984 90914 226012 100014
rect 226260 94926 226288 100028
rect 226248 94920 226300 94926
rect 226248 94862 226300 94868
rect 226536 92274 226564 100028
rect 226628 100014 226734 100042
rect 226524 92268 226576 92274
rect 226524 92210 226576 92216
rect 225972 90908 226024 90914
rect 225972 90850 226024 90856
rect 225340 89686 225644 89714
rect 225144 4004 225196 4010
rect 225144 3946 225196 3952
rect 223948 3528 224000 3534
rect 223948 3470 224000 3476
rect 224868 3528 224920 3534
rect 224868 3470 224920 3476
rect 223856 3392 223908 3398
rect 223856 3334 223908 3340
rect 223960 480 223988 3470
rect 225156 480 225184 3946
rect 225340 3330 225368 89686
rect 226628 89486 226656 100014
rect 226904 94994 226932 100028
rect 226996 100014 227102 100042
rect 227180 100014 227286 100042
rect 226892 94988 226944 94994
rect 226892 94930 226944 94936
rect 226996 93702 227024 100014
rect 226984 93696 227036 93702
rect 226984 93638 227036 93644
rect 227180 90982 227208 100014
rect 227548 97374 227576 100028
rect 227536 97368 227588 97374
rect 227536 97310 227588 97316
rect 227628 97368 227680 97374
rect 227628 97310 227680 97316
rect 227168 90976 227220 90982
rect 227168 90918 227220 90924
rect 226616 89480 226668 89486
rect 226616 89422 226668 89428
rect 226340 9036 226392 9042
rect 226340 8978 226392 8984
rect 225328 3324 225380 3330
rect 225328 3266 225380 3272
rect 226352 480 226380 8978
rect 227640 6914 227668 97310
rect 227732 95130 227760 100028
rect 227930 100014 228036 100042
rect 227720 95124 227772 95130
rect 227720 95066 227772 95072
rect 228008 92342 228036 100014
rect 228100 96218 228128 100028
rect 228088 96212 228140 96218
rect 228088 96154 228140 96160
rect 228284 93770 228312 100028
rect 228376 100014 228574 100042
rect 228376 99374 228404 100014
rect 228376 99346 228680 99374
rect 228364 95940 228416 95946
rect 228364 95882 228416 95888
rect 228272 93764 228324 93770
rect 228272 93706 228324 93712
rect 227996 92336 228048 92342
rect 227996 92278 228048 92284
rect 227548 6886 227668 6914
rect 227548 480 227576 6886
rect 228376 3874 228404 95882
rect 228456 94580 228508 94586
rect 228456 94522 228508 94528
rect 228364 3868 228416 3874
rect 228364 3810 228416 3816
rect 228468 3738 228496 94522
rect 228548 93832 228600 93838
rect 228548 93774 228600 93780
rect 228560 3942 228588 93774
rect 228652 92410 228680 99346
rect 228744 96286 228772 100028
rect 228836 100014 228942 100042
rect 228732 96280 228784 96286
rect 228732 96222 228784 96228
rect 228836 93770 228864 100014
rect 229112 95198 229140 100028
rect 229296 96354 229324 100028
rect 229284 96348 229336 96354
rect 229284 96290 229336 96296
rect 229100 95192 229152 95198
rect 229100 95134 229152 95140
rect 229480 94450 229508 100028
rect 229664 100014 229770 100042
rect 229468 94444 229520 94450
rect 229468 94386 229520 94392
rect 228824 93764 228876 93770
rect 228824 93706 228876 93712
rect 229664 92478 229692 100014
rect 229940 97510 229968 100028
rect 230032 100014 230138 100042
rect 230216 100014 230322 100042
rect 229928 97504 229980 97510
rect 229928 97446 229980 97452
rect 230032 93090 230060 100014
rect 230020 93084 230072 93090
rect 230020 93026 230072 93032
rect 229744 92608 229796 92614
rect 229744 92550 229796 92556
rect 229652 92472 229704 92478
rect 229652 92414 229704 92420
rect 228640 92404 228692 92410
rect 228640 92346 228692 92352
rect 228548 3936 228600 3942
rect 228548 3878 228600 3884
rect 228732 3936 228784 3942
rect 228732 3878 228784 3884
rect 228456 3732 228508 3738
rect 228456 3674 228508 3680
rect 228744 480 228772 3878
rect 229756 3806 229784 92550
rect 230216 91050 230244 100014
rect 230492 96422 230520 100028
rect 230480 96416 230532 96422
rect 230480 96358 230532 96364
rect 230388 94852 230440 94858
rect 230388 94794 230440 94800
rect 230204 91044 230256 91050
rect 230204 90986 230256 90992
rect 229744 3800 229796 3806
rect 229744 3742 229796 3748
rect 230400 3534 230428 94794
rect 230768 93022 230796 100028
rect 230860 100014 230966 100042
rect 230756 93016 230808 93022
rect 230756 92958 230808 92964
rect 230860 91730 230888 100014
rect 231136 96490 231164 100028
rect 231334 100014 231440 100042
rect 231308 97912 231360 97918
rect 231308 97854 231360 97860
rect 231124 96484 231176 96490
rect 231124 96426 231176 96432
rect 231124 96348 231176 96354
rect 231124 96290 231176 96296
rect 230848 91724 230900 91730
rect 230848 91666 230900 91672
rect 231136 3602 231164 96290
rect 231216 92540 231268 92546
rect 231216 92482 231268 92488
rect 231228 3670 231256 92482
rect 231320 8362 231348 97854
rect 231412 92954 231440 100014
rect 231504 94382 231532 100028
rect 231780 95878 231808 100028
rect 231978 100014 232084 100042
rect 232162 100014 232268 100042
rect 231768 95872 231820 95878
rect 231768 95814 231820 95820
rect 232056 94518 232084 100014
rect 232240 95146 232268 100014
rect 232332 95810 232360 100028
rect 232424 100014 232530 100042
rect 232608 100014 232806 100042
rect 232320 95804 232372 95810
rect 232320 95746 232372 95752
rect 232240 95118 232360 95146
rect 232136 94648 232188 94654
rect 232136 94590 232188 94596
rect 232044 94512 232096 94518
rect 232044 94454 232096 94460
rect 231492 94376 231544 94382
rect 231492 94318 231544 94324
rect 231400 92948 231452 92954
rect 231400 92890 231452 92896
rect 232148 84194 232176 94590
rect 232332 86954 232360 95118
rect 232424 94654 232452 100014
rect 232412 94648 232464 94654
rect 232412 94590 232464 94596
rect 232412 94512 232464 94518
rect 232412 94454 232464 94460
rect 232056 84166 232176 84194
rect 232240 86926 232360 86954
rect 231308 8356 231360 8362
rect 231308 8298 231360 8304
rect 232056 6390 232084 84166
rect 232240 7614 232268 86926
rect 232228 7608 232280 7614
rect 232228 7550 232280 7556
rect 232044 6384 232096 6390
rect 232044 6326 232096 6332
rect 232424 6322 232452 94454
rect 232608 7750 232636 100014
rect 232976 97442 233004 100028
rect 233068 100014 233174 100042
rect 232964 97436 233016 97442
rect 232964 97378 233016 97384
rect 233068 84194 233096 100014
rect 233344 99374 233372 100028
rect 233252 99346 233372 99374
rect 233252 96642 233280 99346
rect 233160 96614 233280 96642
rect 233160 92886 233188 96614
rect 233528 95742 233556 100028
rect 233516 95736 233568 95742
rect 233516 95678 233568 95684
rect 233712 94314 233740 100028
rect 233804 100014 234002 100042
rect 233700 94308 233752 94314
rect 233700 94250 233752 94256
rect 233148 92880 233200 92886
rect 233148 92822 233200 92828
rect 233804 89714 233832 100014
rect 233884 96756 233936 96762
rect 233884 96698 233936 96704
rect 232700 84166 233096 84194
rect 233620 89686 233832 89714
rect 232596 7744 232648 7750
rect 232596 7686 232648 7692
rect 232700 6458 232728 84166
rect 233620 24138 233648 89686
rect 233608 24132 233660 24138
rect 233608 24074 233660 24080
rect 233148 22772 233200 22778
rect 233148 22714 233200 22720
rect 232688 6452 232740 6458
rect 232688 6394 232740 6400
rect 232412 6316 232464 6322
rect 232412 6258 232464 6264
rect 231216 3664 231268 3670
rect 231216 3606 231268 3612
rect 231124 3596 231176 3602
rect 231124 3538 231176 3544
rect 229836 3528 229888 3534
rect 229836 3470 229888 3476
rect 230388 3528 230440 3534
rect 230388 3470 230440 3476
rect 229848 480 229876 3470
rect 233160 3466 233188 22714
rect 233896 9042 233924 96698
rect 233976 96688 234028 96694
rect 233976 96630 234028 96636
rect 233988 10334 234016 96630
rect 234172 95674 234200 100028
rect 234264 100014 234370 100042
rect 234160 95668 234212 95674
rect 234160 95610 234212 95616
rect 234264 93838 234292 100014
rect 234540 97850 234568 100028
rect 234528 97844 234580 97850
rect 234528 97786 234580 97792
rect 234724 97306 234752 100028
rect 234712 97300 234764 97306
rect 234712 97242 234764 97248
rect 235000 94722 235028 100028
rect 235092 100014 235198 100042
rect 234988 94716 235040 94722
rect 234988 94658 235040 94664
rect 234804 94580 234856 94586
rect 234804 94522 234856 94528
rect 234252 93832 234304 93838
rect 234252 93774 234304 93780
rect 234068 23520 234120 23526
rect 234068 23462 234120 23468
rect 233976 10328 234028 10334
rect 233976 10270 234028 10276
rect 233884 9036 233936 9042
rect 233884 8978 233936 8984
rect 234080 4010 234108 23462
rect 234816 6254 234844 94522
rect 235092 91780 235120 100014
rect 235368 96354 235396 100028
rect 235460 100014 235566 100042
rect 235644 100014 235750 100042
rect 235356 96348 235408 96354
rect 235356 96290 235408 96296
rect 235172 94716 235224 94722
rect 235172 94658 235224 94664
rect 234908 91752 235120 91780
rect 234804 6248 234856 6254
rect 234804 6190 234856 6196
rect 234068 4004 234120 4010
rect 234068 3946 234120 3952
rect 234620 3528 234672 3534
rect 234620 3470 234672 3476
rect 232228 3460 232280 3466
rect 232228 3402 232280 3408
rect 233148 3460 233200 3466
rect 233148 3402 233200 3408
rect 231032 3188 231084 3194
rect 231032 3130 231084 3136
rect 231044 480 231072 3130
rect 232240 480 232268 3402
rect 233424 3324 233476 3330
rect 233424 3266 233476 3272
rect 233436 480 233464 3266
rect 234632 480 234660 3470
rect 234908 3398 234936 91752
rect 235184 86954 235212 94658
rect 235460 94586 235488 100014
rect 235448 94580 235500 94586
rect 235448 94522 235500 94528
rect 235644 92546 235672 100014
rect 236012 96830 236040 100028
rect 236210 100014 236316 100042
rect 236000 96824 236052 96830
rect 236000 96766 236052 96772
rect 235908 95328 235960 95334
rect 235908 95270 235960 95276
rect 235632 92540 235684 92546
rect 235632 92482 235684 92488
rect 235000 86926 235212 86954
rect 235000 6526 235028 86926
rect 235920 6914 235948 95270
rect 235828 6886 235948 6914
rect 234988 6520 235040 6526
rect 234988 6462 235040 6468
rect 234896 3392 234948 3398
rect 234896 3334 234948 3340
rect 235828 480 235856 6886
rect 236288 6186 236316 100014
rect 236380 94654 236408 100028
rect 236368 94648 236420 94654
rect 236368 94590 236420 94596
rect 236276 6180 236328 6186
rect 236276 6122 236328 6128
rect 236564 4894 236592 100028
rect 236644 94580 236696 94586
rect 236644 94522 236696 94528
rect 236656 4962 236684 94522
rect 236748 6594 236776 100028
rect 236840 100014 237038 100042
rect 237116 100014 237222 100042
rect 237406 100014 237512 100042
rect 236840 92614 236868 100014
rect 237116 94586 237144 100014
rect 237380 96892 237432 96898
rect 237380 96834 237432 96840
rect 237392 94858 237420 96834
rect 237484 95946 237512 100014
rect 237576 96694 237604 100028
rect 237668 100014 237774 100042
rect 237564 96688 237616 96694
rect 237564 96630 237616 96636
rect 237472 95940 237524 95946
rect 237472 95882 237524 95888
rect 237380 94852 237432 94858
rect 237380 94794 237432 94800
rect 237104 94580 237156 94586
rect 237104 94522 237156 94528
rect 236828 92608 236880 92614
rect 236828 92550 236880 92556
rect 236736 6588 236788 6594
rect 236736 6530 236788 6536
rect 237668 5030 237696 100014
rect 238036 97918 238064 100028
rect 238220 98326 238248 100028
rect 238312 100014 238418 100042
rect 238208 98320 238260 98326
rect 238208 98262 238260 98268
rect 238024 97912 238076 97918
rect 238024 97854 238076 97860
rect 238024 96688 238076 96694
rect 238024 96630 238076 96636
rect 238036 6914 238064 96630
rect 238116 95260 238168 95266
rect 238116 95202 238168 95208
rect 237944 6886 238064 6914
rect 237656 5024 237708 5030
rect 237656 4966 237708 4972
rect 236644 4956 236696 4962
rect 236644 4898 236696 4904
rect 236552 4888 236604 4894
rect 236552 4830 236604 4836
rect 237944 3942 237972 6886
rect 238128 4162 238156 95202
rect 238208 92472 238260 92478
rect 238208 92414 238260 92420
rect 238036 4134 238156 4162
rect 237932 3936 237984 3942
rect 237932 3878 237984 3884
rect 238036 3194 238064 4134
rect 238116 4072 238168 4078
rect 238116 4014 238168 4020
rect 238024 3188 238076 3194
rect 238024 3130 238076 3136
rect 237012 3052 237064 3058
rect 237012 2994 237064 3000
rect 237024 480 237052 2994
rect 238128 480 238156 4014
rect 238220 3534 238248 92414
rect 238312 23526 238340 100014
rect 238484 98320 238536 98326
rect 238484 98262 238536 98268
rect 238496 91798 238524 98262
rect 238588 96762 238616 100028
rect 238772 97374 238800 100028
rect 238760 97368 238812 97374
rect 238760 97310 238812 97316
rect 238576 96756 238628 96762
rect 238576 96698 238628 96704
rect 238956 96694 238984 100028
rect 239232 96898 239260 100028
rect 239220 96892 239272 96898
rect 239220 96834 239272 96840
rect 239036 96824 239088 96830
rect 239036 96766 239088 96772
rect 238944 96688 238996 96694
rect 238944 96630 238996 96636
rect 238484 91792 238536 91798
rect 238484 91734 238536 91740
rect 238300 23520 238352 23526
rect 238300 23462 238352 23468
rect 239048 4826 239076 96766
rect 239416 95266 239444 100028
rect 239508 100014 239614 100042
rect 239692 100014 239798 100042
rect 239876 100014 239982 100042
rect 239404 95260 239456 95266
rect 239404 95202 239456 95208
rect 239128 94580 239180 94586
rect 239128 94522 239180 94528
rect 239036 4820 239088 4826
rect 239036 4762 239088 4768
rect 238208 3528 238260 3534
rect 238208 3470 238260 3476
rect 239140 3330 239168 94522
rect 239508 22778 239536 100014
rect 239692 94586 239720 100014
rect 239680 94580 239732 94586
rect 239680 94522 239732 94528
rect 239876 92478 239904 100014
rect 240140 96688 240192 96694
rect 240140 96630 240192 96636
rect 239864 92472 239916 92478
rect 239864 92414 239916 92420
rect 239496 22772 239548 22778
rect 239496 22714 239548 22720
rect 239128 3324 239180 3330
rect 239128 3266 239180 3272
rect 239312 3324 239364 3330
rect 239312 3266 239364 3272
rect 239324 480 239352 3266
rect 240152 490 240180 96630
rect 240244 95334 240272 100028
rect 240442 100014 240548 100042
rect 240520 99278 240548 100014
rect 240508 99272 240560 99278
rect 240508 99214 240560 99220
rect 240232 95328 240284 95334
rect 240232 95270 240284 95276
rect 240324 94580 240376 94586
rect 240324 94522 240376 94528
rect 240336 3330 240364 94522
rect 240612 4078 240640 100028
rect 240704 100014 240810 100042
rect 240704 94586 240732 100014
rect 240980 96694 241008 100028
rect 241270 100014 241376 100042
rect 241060 99272 241112 99278
rect 241060 99214 241112 99220
rect 240968 96688 241020 96694
rect 240968 96630 241020 96636
rect 240692 94580 240744 94586
rect 240692 94522 240744 94528
rect 240600 4072 240652 4078
rect 240600 4014 240652 4020
rect 240324 3324 240376 3330
rect 240324 3266 240376 3272
rect 241072 3058 241100 99214
rect 241348 89714 241376 100014
rect 241440 97102 241468 100028
rect 241428 97096 241480 97102
rect 241428 97038 241480 97044
rect 241624 94518 241652 100028
rect 241808 96898 241836 100028
rect 241992 97646 242020 100028
rect 241980 97640 242032 97646
rect 241980 97582 242032 97588
rect 242164 97096 242216 97102
rect 242164 97038 242216 97044
rect 241796 96892 241848 96898
rect 241796 96834 241848 96840
rect 241612 94512 241664 94518
rect 241612 94454 241664 94460
rect 241348 89686 241468 89714
rect 241440 3482 241468 89686
rect 242176 3534 242204 97038
rect 242268 96694 242296 100028
rect 242452 97102 242480 100028
rect 242544 100014 242650 100042
rect 242728 100014 242834 100042
rect 242440 97096 242492 97102
rect 242440 97038 242492 97044
rect 242256 96688 242308 96694
rect 242256 96630 242308 96636
rect 242544 94602 242572 100014
rect 242728 99374 242756 100014
rect 242452 94574 242572 94602
rect 242636 99346 242756 99374
rect 242452 4010 242480 94574
rect 242532 94512 242584 94518
rect 242532 94454 242584 94460
rect 242440 4004 242492 4010
rect 242440 3946 242492 3952
rect 242164 3528 242216 3534
rect 241440 3454 241744 3482
rect 242164 3470 242216 3476
rect 241060 3052 241112 3058
rect 241060 2994 241112 3000
rect 240336 598 240548 626
rect 240336 490 240364 598
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240152 462 240364 490
rect 240520 480 240548 598
rect 241716 480 241744 3454
rect 242544 2922 242572 94454
rect 242636 3670 242664 99346
rect 242716 97640 242768 97646
rect 242716 97582 242768 97588
rect 242624 3664 242676 3670
rect 242624 3606 242676 3612
rect 242728 3466 242756 97582
rect 243004 97170 243032 100028
rect 243188 97238 243216 100028
rect 243478 100014 243584 100042
rect 243176 97232 243228 97238
rect 243176 97174 243228 97180
rect 242992 97164 243044 97170
rect 242992 97106 243044 97112
rect 242808 96688 242860 96694
rect 242808 96630 242860 96636
rect 242716 3460 242768 3466
rect 242716 3402 242768 3408
rect 242820 3398 242848 96630
rect 243556 89714 243584 100014
rect 243648 94518 243676 100028
rect 243832 97442 243860 100028
rect 243924 100014 244030 100042
rect 243820 97436 243872 97442
rect 243820 97378 243872 97384
rect 243636 94512 243688 94518
rect 243636 94454 243688 94460
rect 243924 93158 243952 100014
rect 244200 94602 244228 100028
rect 244476 96966 244504 100028
rect 244464 96960 244516 96966
rect 244464 96902 244516 96908
rect 244372 96892 244424 96898
rect 244372 96834 244424 96840
rect 244016 94574 244228 94602
rect 243912 93152 243964 93158
rect 243912 93094 243964 93100
rect 243556 89686 243952 89714
rect 243924 4078 243952 89686
rect 243912 4072 243964 4078
rect 243912 4014 243964 4020
rect 244016 3738 244044 94574
rect 244096 94512 244148 94518
rect 244096 94454 244148 94460
rect 244108 3874 244136 94454
rect 244384 16574 244412 96834
rect 244660 96830 244688 100028
rect 244858 100014 244964 100042
rect 244648 96824 244700 96830
rect 244648 96766 244700 96772
rect 244936 93854 244964 100014
rect 245028 96014 245056 100028
rect 245226 100014 245424 100042
rect 245292 96960 245344 96966
rect 245292 96902 245344 96908
rect 245396 96914 245424 100014
rect 245488 97782 245516 100028
rect 245476 97776 245528 97782
rect 245476 97718 245528 97724
rect 245016 96008 245068 96014
rect 245016 95950 245068 95956
rect 244936 93826 245240 93854
rect 244384 16546 245148 16574
rect 244096 3868 244148 3874
rect 244096 3810 244148 3816
rect 244004 3732 244056 3738
rect 244004 3674 244056 3680
rect 242900 3528 242952 3534
rect 242900 3470 242952 3476
rect 245120 3482 245148 16546
rect 245212 3806 245240 93826
rect 245304 15910 245332 96902
rect 245396 96886 245516 96914
rect 245672 96898 245700 100028
rect 245856 96966 245884 100028
rect 245844 96960 245896 96966
rect 245844 96902 245896 96908
rect 245384 96824 245436 96830
rect 245384 96766 245436 96772
rect 245292 15904 245344 15910
rect 245292 15846 245344 15852
rect 245396 5166 245424 96766
rect 245488 5302 245516 96886
rect 245660 96892 245712 96898
rect 245660 96834 245712 96840
rect 246040 96762 246068 100028
rect 246224 96830 246252 100028
rect 246514 100014 246620 100042
rect 246698 100014 246804 100042
rect 246304 97096 246356 97102
rect 246304 97038 246356 97044
rect 246212 96824 246264 96830
rect 246212 96766 246264 96772
rect 246028 96756 246080 96762
rect 246028 96698 246080 96704
rect 245476 5296 245528 5302
rect 245476 5238 245528 5244
rect 245384 5160 245436 5166
rect 245384 5102 245436 5108
rect 246316 4146 246344 97038
rect 246488 96960 246540 96966
rect 246488 96902 246540 96908
rect 246500 5098 246528 96902
rect 246488 5092 246540 5098
rect 246488 5034 246540 5040
rect 246304 4140 246356 4146
rect 246304 4082 246356 4088
rect 245200 3800 245252 3806
rect 245200 3742 245252 3748
rect 246592 3602 246620 100014
rect 246776 96914 246804 100014
rect 246868 97918 246896 100028
rect 246856 97912 246908 97918
rect 246856 97854 246908 97860
rect 246672 96892 246724 96898
rect 246776 96886 246988 96914
rect 246672 96834 246724 96840
rect 246684 22778 246712 96834
rect 246764 96824 246816 96830
rect 246764 96766 246816 96772
rect 246672 22772 246724 22778
rect 246672 22714 246724 22720
rect 246776 10402 246804 96766
rect 246856 96756 246908 96762
rect 246856 96698 246908 96704
rect 246868 93226 246896 96698
rect 246856 93220 246908 93226
rect 246856 93162 246908 93168
rect 246960 91798 246988 96886
rect 247052 94518 247080 100028
rect 247236 96966 247264 100028
rect 247512 97646 247540 100028
rect 247696 97850 247724 100028
rect 247894 100014 248000 100042
rect 247684 97844 247736 97850
rect 247684 97786 247736 97792
rect 247500 97640 247552 97646
rect 247500 97582 247552 97588
rect 247224 96960 247276 96966
rect 247224 96902 247276 96908
rect 247040 94512 247092 94518
rect 247040 94454 247092 94460
rect 247972 93854 248000 100014
rect 248064 95946 248092 100028
rect 248156 100014 248262 100042
rect 248052 95940 248104 95946
rect 248052 95882 248104 95888
rect 247972 93826 248092 93854
rect 246948 91792 247000 91798
rect 246948 91734 247000 91740
rect 246764 10396 246816 10402
rect 246764 10338 246816 10344
rect 246580 3596 246632 3602
rect 246580 3538 246632 3544
rect 248064 3534 248092 93826
rect 248156 90370 248184 100014
rect 248236 96960 248288 96966
rect 248236 96902 248288 96908
rect 248144 90364 248196 90370
rect 248144 90306 248196 90312
rect 248248 86290 248276 96902
rect 248432 96830 248460 100028
rect 248708 97578 248736 100028
rect 248696 97572 248748 97578
rect 248696 97514 248748 97520
rect 248420 96824 248472 96830
rect 248420 96766 248472 96772
rect 248892 96694 248920 100028
rect 249090 100014 249196 100042
rect 249274 100014 249380 100042
rect 249458 100014 249656 100042
rect 249168 96948 249196 100014
rect 249352 97050 249380 100014
rect 249352 97022 249564 97050
rect 249168 96920 249472 96948
rect 249248 96824 249300 96830
rect 249248 96766 249300 96772
rect 249340 96824 249392 96830
rect 249340 96766 249392 96772
rect 248880 96688 248932 96694
rect 248880 96630 248932 96636
rect 248236 86284 248288 86290
rect 248236 86226 248288 86232
rect 249260 6594 249288 96766
rect 249248 6588 249300 6594
rect 249248 6530 249300 6536
rect 249352 6186 249380 96766
rect 249444 6254 249472 96920
rect 249536 96778 249564 97022
rect 249628 96948 249656 100014
rect 249720 97102 249748 100028
rect 249708 97096 249760 97102
rect 249708 97038 249760 97044
rect 249628 96920 249748 96948
rect 249536 96750 249656 96778
rect 249524 96688 249576 96694
rect 249524 96630 249576 96636
rect 249432 6248 249484 6254
rect 249432 6190 249484 6196
rect 249340 6180 249392 6186
rect 249340 6122 249392 6128
rect 249536 4962 249564 96630
rect 249524 4956 249576 4962
rect 249524 4898 249576 4904
rect 249628 4894 249656 96750
rect 249720 5234 249748 96920
rect 249904 95606 249932 100028
rect 250088 96966 250116 100028
rect 250286 100014 250392 100042
rect 250260 97164 250312 97170
rect 250260 97106 250312 97112
rect 250076 96960 250128 96966
rect 250076 96902 250128 96908
rect 249892 95600 249944 95606
rect 249892 95542 249944 95548
rect 250272 92002 250300 97106
rect 250364 96778 250392 100014
rect 250456 97034 250484 100028
rect 250444 97028 250496 97034
rect 250444 96970 250496 96976
rect 250732 96898 250760 100028
rect 250824 100014 250930 100042
rect 250720 96892 250772 96898
rect 250720 96834 250772 96840
rect 250364 96750 250760 96778
rect 250260 91996 250312 92002
rect 250260 91938 250312 91944
rect 249708 5228 249760 5234
rect 249708 5170 249760 5176
rect 249616 4888 249668 4894
rect 249616 4830 249668 4836
rect 248788 4140 248840 4146
rect 248788 4082 248840 4088
rect 248052 3528 248104 3534
rect 242808 3392 242860 3398
rect 242808 3334 242860 3340
rect 242532 2916 242584 2922
rect 242532 2858 242584 2864
rect 242912 480 242940 3470
rect 245120 3454 245240 3482
rect 248052 3470 248104 3476
rect 244096 2916 244148 2922
rect 244096 2858 244148 2864
rect 244108 480 244136 2858
rect 245212 480 245240 3454
rect 246396 3460 246448 3466
rect 246396 3402 246448 3408
rect 246408 480 246436 3402
rect 247592 3392 247644 3398
rect 247592 3334 247644 3340
rect 247604 480 247632 3334
rect 248800 480 248828 4082
rect 249984 4004 250036 4010
rect 249984 3946 250036 3952
rect 249996 480 250024 3946
rect 250732 3466 250760 96750
rect 250824 10334 250852 100014
rect 251100 97510 251128 100028
rect 251088 97504 251140 97510
rect 251088 97446 251140 97452
rect 251088 97028 251140 97034
rect 251088 96970 251140 96976
rect 250996 96960 251048 96966
rect 250996 96902 251048 96908
rect 250904 96892 250956 96898
rect 250904 96834 250956 96840
rect 250812 10328 250864 10334
rect 250812 10270 250864 10276
rect 250916 6526 250944 96834
rect 250904 6520 250956 6526
rect 250904 6462 250956 6468
rect 251008 4826 251036 96902
rect 251100 95742 251128 96970
rect 251284 95810 251312 100028
rect 251468 97034 251496 100028
rect 251456 97028 251508 97034
rect 251456 96970 251508 96976
rect 251272 95804 251324 95810
rect 251272 95746 251324 95752
rect 251088 95736 251140 95742
rect 251088 95678 251140 95684
rect 251744 94178 251772 100028
rect 251824 97844 251876 97850
rect 251824 97786 251876 97792
rect 251732 94172 251784 94178
rect 251732 94114 251784 94120
rect 251272 91996 251324 92002
rect 251272 91938 251324 91944
rect 251284 16574 251312 91938
rect 251284 16546 251772 16574
rect 250996 4820 251048 4826
rect 250996 4762 251048 4768
rect 251180 3664 251232 3670
rect 251180 3606 251232 3612
rect 250720 3460 250772 3466
rect 250720 3402 250772 3408
rect 251192 480 251220 3606
rect 251744 3482 251772 16546
rect 251836 5030 251864 97786
rect 251928 96966 251956 100028
rect 251916 96960 251968 96966
rect 251916 96902 251968 96908
rect 252008 96892 252060 96898
rect 252008 96834 252060 96840
rect 251916 10396 251968 10402
rect 251916 10338 251968 10344
rect 251824 5024 251876 5030
rect 251824 4966 251876 4972
rect 251928 3670 251956 10338
rect 252020 4010 252048 96834
rect 252112 4146 252140 100028
rect 252310 100014 252416 100042
rect 252284 97028 252336 97034
rect 252284 96970 252336 96976
rect 252192 96960 252244 96966
rect 252192 96902 252244 96908
rect 252204 90166 252232 96902
rect 252192 90160 252244 90166
rect 252192 90102 252244 90108
rect 252296 19990 252324 96970
rect 252388 94314 252416 100014
rect 252480 96898 252508 100028
rect 252664 96898 252692 100028
rect 252468 96892 252520 96898
rect 252468 96834 252520 96840
rect 252652 96892 252704 96898
rect 252652 96834 252704 96840
rect 252940 94382 252968 100028
rect 253020 97776 253072 97782
rect 253020 97718 253072 97724
rect 252928 94376 252980 94382
rect 252928 94318 252980 94324
rect 252376 94308 252428 94314
rect 252376 94250 252428 94256
rect 253032 93854 253060 97718
rect 253124 96966 253152 100028
rect 253322 100014 253428 100042
rect 253204 97912 253256 97918
rect 253204 97854 253256 97860
rect 253216 97306 253244 97854
rect 253204 97300 253256 97306
rect 253204 97242 253256 97248
rect 253112 96960 253164 96966
rect 253112 96902 253164 96908
rect 253400 93854 253428 100014
rect 253492 95878 253520 100028
rect 253572 96960 253624 96966
rect 253572 96902 253624 96908
rect 253480 95872 253532 95878
rect 253480 95814 253532 95820
rect 253032 93826 253244 93854
rect 253400 93826 253520 93854
rect 252284 19984 252336 19990
rect 252284 19926 252336 19932
rect 253216 7614 253244 93826
rect 253492 29646 253520 93826
rect 253584 90234 253612 96902
rect 253572 90228 253624 90234
rect 253572 90170 253624 90176
rect 253676 87582 253704 100028
rect 253952 96898 253980 100028
rect 254136 97714 254164 100028
rect 254334 100014 254440 100042
rect 254124 97708 254176 97714
rect 254124 97650 254176 97656
rect 253756 96892 253808 96898
rect 253756 96834 253808 96840
rect 253940 96892 253992 96898
rect 253940 96834 253992 96840
rect 253664 87576 253716 87582
rect 253664 87518 253716 87524
rect 253768 85474 253796 96834
rect 254412 91662 254440 100014
rect 254504 96830 254532 100028
rect 254492 96824 254544 96830
rect 254492 96766 254544 96772
rect 254688 96626 254716 100028
rect 254860 96960 254912 96966
rect 254860 96902 254912 96908
rect 254676 96620 254728 96626
rect 254676 96562 254728 96568
rect 254400 91656 254452 91662
rect 254400 91598 254452 91604
rect 253756 85468 253808 85474
rect 253756 85410 253808 85416
rect 254872 33794 254900 96902
rect 254964 90302 254992 100028
rect 255148 96966 255176 100028
rect 255136 96960 255188 96966
rect 255136 96902 255188 96908
rect 255044 96892 255096 96898
rect 255044 96834 255096 96840
rect 254952 90296 255004 90302
rect 254952 90238 255004 90244
rect 255056 86222 255084 96834
rect 255136 96824 255188 96830
rect 255136 96766 255188 96772
rect 255044 86216 255096 86222
rect 255044 86158 255096 86164
rect 255148 84046 255176 96766
rect 255332 94450 255360 100028
rect 255516 96966 255544 100028
rect 255714 100014 255912 100042
rect 255504 96960 255556 96966
rect 255884 96948 255912 100014
rect 255976 97170 256004 100028
rect 255964 97164 256016 97170
rect 255964 97106 256016 97112
rect 256160 97102 256188 100028
rect 256252 100014 256358 100042
rect 256148 97096 256200 97102
rect 256148 97038 256200 97044
rect 255884 96920 256188 96948
rect 255504 96902 255556 96908
rect 256056 96824 256108 96830
rect 256056 96766 256108 96772
rect 255320 94444 255372 94450
rect 255320 94386 255372 94392
rect 255964 93152 256016 93158
rect 255964 93094 256016 93100
rect 255136 84040 255188 84046
rect 255136 83982 255188 83988
rect 254860 33788 254912 33794
rect 254860 33730 254912 33736
rect 253480 29640 253532 29646
rect 253480 29582 253532 29588
rect 253388 15904 253440 15910
rect 253388 15846 253440 15852
rect 253296 13116 253348 13122
rect 253296 13058 253348 13064
rect 253204 7608 253256 7614
rect 253204 7550 253256 7556
rect 253308 7426 253336 13058
rect 253216 7398 253336 7426
rect 252100 4140 252152 4146
rect 252100 4082 252152 4088
rect 252008 4004 252060 4010
rect 252008 3946 252060 3952
rect 251916 3664 251968 3670
rect 251916 3606 251968 3612
rect 251744 3454 252416 3482
rect 252388 480 252416 3454
rect 253216 3210 253244 7398
rect 253400 6914 253428 15846
rect 253308 6886 253428 6914
rect 253308 3330 253336 6886
rect 255976 4078 256004 93094
rect 256068 93022 256096 96766
rect 256056 93016 256108 93022
rect 256056 92958 256108 92964
rect 256160 83978 256188 96920
rect 256148 83972 256200 83978
rect 256148 83914 256200 83920
rect 256252 31074 256280 100014
rect 256424 97096 256476 97102
rect 256424 97038 256476 97044
rect 256332 96960 256384 96966
rect 256332 96902 256384 96908
rect 256344 88874 256372 96902
rect 256332 88868 256384 88874
rect 256332 88810 256384 88816
rect 256436 88330 256464 97038
rect 256528 96830 256556 100028
rect 256608 97164 256660 97170
rect 256608 97106 256660 97112
rect 256516 96824 256568 96830
rect 256516 96766 256568 96772
rect 256620 92954 256648 97106
rect 256712 96898 256740 100028
rect 256988 97714 257016 100028
rect 257186 100014 257292 100042
rect 256976 97708 257028 97714
rect 256976 97650 257028 97656
rect 256792 97640 256844 97646
rect 256792 97582 256844 97588
rect 256804 97170 256832 97582
rect 256792 97164 256844 97170
rect 256792 97106 256844 97112
rect 256700 96892 256752 96898
rect 256700 96834 256752 96840
rect 257264 93090 257292 100014
rect 257356 96830 257384 100028
rect 257344 96824 257396 96830
rect 257344 96766 257396 96772
rect 257540 96558 257568 100028
rect 257620 96960 257672 96966
rect 257620 96902 257672 96908
rect 257528 96552 257580 96558
rect 257528 96494 257580 96500
rect 257344 93220 257396 93226
rect 257344 93162 257396 93168
rect 257252 93084 257304 93090
rect 257252 93026 257304 93032
rect 256608 92948 256660 92954
rect 256608 92890 256660 92896
rect 256424 88324 256476 88330
rect 256424 88266 256476 88272
rect 256240 31068 256292 31074
rect 256240 31010 256292 31016
rect 257068 4140 257120 4146
rect 257068 4082 257120 4088
rect 254676 4072 254728 4078
rect 254676 4014 254728 4020
rect 255964 4072 256016 4078
rect 255964 4014 256016 4020
rect 253296 3324 253348 3330
rect 253296 3266 253348 3272
rect 253216 3182 253520 3210
rect 253492 480 253520 3182
rect 254688 480 254716 4014
rect 255872 3868 255924 3874
rect 255872 3810 255924 3816
rect 255884 480 255912 3810
rect 257080 480 257108 4082
rect 257356 3398 257384 93162
rect 257632 86902 257660 96902
rect 257724 93838 257752 100028
rect 257908 96966 257936 100028
rect 258184 97034 258212 100028
rect 258264 97436 258316 97442
rect 258264 97378 258316 97384
rect 258172 97028 258224 97034
rect 258172 96970 258224 96976
rect 257896 96960 257948 96966
rect 257896 96902 257948 96908
rect 257804 96892 257856 96898
rect 257804 96834 257856 96840
rect 257712 93832 257764 93838
rect 257712 93774 257764 93780
rect 257816 88942 257844 96834
rect 257896 96824 257948 96830
rect 257896 96766 257948 96772
rect 257804 88936 257856 88942
rect 257804 88878 257856 88884
rect 257908 88262 257936 96766
rect 258276 93854 258304 97378
rect 258368 96830 258396 100028
rect 258552 96966 258580 100028
rect 258736 98462 258764 100028
rect 258724 98456 258776 98462
rect 258724 98398 258776 98404
rect 258540 96960 258592 96966
rect 258540 96902 258592 96908
rect 258920 96898 258948 100028
rect 259000 97028 259052 97034
rect 259000 96970 259052 96976
rect 258908 96892 258960 96898
rect 258908 96834 258960 96840
rect 258356 96824 258408 96830
rect 258356 96766 258408 96772
rect 258276 93826 258396 93854
rect 257896 88256 257948 88262
rect 257896 88198 257948 88204
rect 257620 86896 257672 86902
rect 257620 86838 257672 86844
rect 258368 4146 258396 93826
rect 259012 16046 259040 96970
rect 259092 96960 259144 96966
rect 259092 96902 259144 96908
rect 259000 16040 259052 16046
rect 259000 15982 259052 15988
rect 259104 12170 259132 96902
rect 259092 12164 259144 12170
rect 259092 12106 259144 12112
rect 259196 12102 259224 100028
rect 259380 98530 259408 100028
rect 259368 98524 259420 98530
rect 259368 98466 259420 98472
rect 259460 97232 259512 97238
rect 259460 97174 259512 97180
rect 259276 96892 259328 96898
rect 259276 96834 259328 96840
rect 259184 12096 259236 12102
rect 259184 12038 259236 12044
rect 259288 6390 259316 96834
rect 259368 96824 259420 96830
rect 259368 96766 259420 96772
rect 259380 6458 259408 96766
rect 259472 13122 259500 97174
rect 259564 96694 259592 100028
rect 259748 97782 259776 100028
rect 259932 98598 259960 100028
rect 259920 98592 259972 98598
rect 259920 98534 259972 98540
rect 259736 97776 259788 97782
rect 259736 97718 259788 97724
rect 260104 97164 260156 97170
rect 260104 97106 260156 97112
rect 259552 96688 259604 96694
rect 259552 96630 259604 96636
rect 259460 13116 259512 13122
rect 259460 13058 259512 13064
rect 259368 6452 259420 6458
rect 259368 6394 259420 6400
rect 259276 6384 259328 6390
rect 259276 6326 259328 6332
rect 258356 4140 258408 4146
rect 258356 4082 258408 4088
rect 258080 4072 258132 4078
rect 258080 4014 258132 4020
rect 257344 3392 257396 3398
rect 257344 3334 257396 3340
rect 258092 2122 258120 4014
rect 260116 3738 260144 97106
rect 260208 96966 260236 100028
rect 260406 100014 260512 100042
rect 260196 96960 260248 96966
rect 260484 96948 260512 100014
rect 260576 97102 260604 100028
rect 260564 97096 260616 97102
rect 260564 97038 260616 97044
rect 260656 96960 260708 96966
rect 260484 96920 260604 96948
rect 260196 96902 260248 96908
rect 260472 96824 260524 96830
rect 260472 96766 260524 96772
rect 260484 91730 260512 96766
rect 260472 91724 260524 91730
rect 260472 91666 260524 91672
rect 260576 91050 260604 96920
rect 260656 96902 260708 96908
rect 260564 91044 260616 91050
rect 260564 90986 260616 90992
rect 260668 6322 260696 96902
rect 260760 96830 260788 100028
rect 260748 96824 260800 96830
rect 260748 96766 260800 96772
rect 260944 96762 260972 100028
rect 261220 97170 261248 100028
rect 261208 97164 261260 97170
rect 261208 97106 261260 97112
rect 260932 96756 260984 96762
rect 260932 96698 260984 96704
rect 260748 96688 260800 96694
rect 260748 96630 260800 96636
rect 260656 6316 260708 6322
rect 260656 6258 260708 6264
rect 260760 3942 260788 96630
rect 261404 95198 261432 100028
rect 261588 96898 261616 100028
rect 261576 96892 261628 96898
rect 261576 96834 261628 96840
rect 261668 96688 261720 96694
rect 261668 96630 261720 96636
rect 261392 95192 261444 95198
rect 261392 95134 261444 95140
rect 261680 86766 261708 96630
rect 261668 86760 261720 86766
rect 261668 86702 261720 86708
rect 261484 86284 261536 86290
rect 261484 86226 261536 86232
rect 261496 4146 261524 86226
rect 261772 83910 261800 100028
rect 261970 100014 262076 100042
rect 261944 96892 261996 96898
rect 261944 96834 261996 96840
rect 261852 96756 261904 96762
rect 261852 96698 261904 96704
rect 261864 88194 261892 96698
rect 261852 88188 261904 88194
rect 261852 88130 261904 88136
rect 261956 86834 261984 96834
rect 262048 93770 262076 100014
rect 262140 96694 262168 100028
rect 262416 97442 262444 100028
rect 262404 97436 262456 97442
rect 262404 97378 262456 97384
rect 262600 96898 262628 100028
rect 262784 97034 262812 100028
rect 262864 97096 262916 97102
rect 262864 97038 262916 97044
rect 262772 97028 262824 97034
rect 262772 96970 262824 96976
rect 262588 96892 262640 96898
rect 262588 96834 262640 96840
rect 262128 96688 262180 96694
rect 262128 96630 262180 96636
rect 262036 93764 262088 93770
rect 262036 93706 262088 93712
rect 261944 86828 261996 86834
rect 261944 86770 261996 86776
rect 261760 83904 261812 83910
rect 261760 83846 261812 83852
rect 262876 5166 262904 97038
rect 262968 96966 262996 100028
rect 263166 100014 263272 100042
rect 263140 97708 263192 97714
rect 263140 97650 263192 97656
rect 263048 97572 263100 97578
rect 263048 97514 263100 97520
rect 262956 96960 263008 96966
rect 262956 96902 263008 96908
rect 263060 96812 263088 97514
rect 262968 96784 263088 96812
rect 262968 17270 262996 96784
rect 263152 85406 263180 97650
rect 263244 92410 263272 100014
rect 263428 97374 263456 100028
rect 263626 100014 263732 100042
rect 263704 97578 263732 100014
rect 263692 97572 263744 97578
rect 263692 97514 263744 97520
rect 263600 97504 263652 97510
rect 263600 97446 263652 97452
rect 263416 97368 263468 97374
rect 263416 97310 263468 97316
rect 263508 97028 263560 97034
rect 263508 96970 263560 96976
rect 263416 96960 263468 96966
rect 263416 96902 263468 96908
rect 263324 96892 263376 96898
rect 263324 96834 263376 96840
rect 263336 92478 263364 96834
rect 263324 92472 263376 92478
rect 263324 92414 263376 92420
rect 263232 92404 263284 92410
rect 263232 92346 263284 92352
rect 263428 88126 263456 96902
rect 263416 88120 263468 88126
rect 263416 88062 263468 88068
rect 263140 85400 263192 85406
rect 263140 85342 263192 85348
rect 262956 17264 263008 17270
rect 262956 17206 263008 17212
rect 263520 12034 263548 96970
rect 263612 95674 263640 97446
rect 263796 96898 263824 100028
rect 263876 97640 263928 97646
rect 263876 97582 263928 97588
rect 263784 96892 263836 96898
rect 263784 96834 263836 96840
rect 263600 95668 263652 95674
rect 263600 95610 263652 95616
rect 263888 94246 263916 97582
rect 263980 96830 264008 100028
rect 263968 96824 264020 96830
rect 263968 96766 264020 96772
rect 264164 96694 264192 100028
rect 264440 96966 264468 100028
rect 264638 100014 264744 100042
rect 264428 96960 264480 96966
rect 264716 96948 264744 100014
rect 264808 97510 264836 100028
rect 264992 97646 265020 100028
rect 264980 97640 265032 97646
rect 264980 97582 265032 97588
rect 264796 97504 264848 97510
rect 264796 97446 264848 97452
rect 265072 97436 265124 97442
rect 265072 97378 265124 97384
rect 265084 97238 265112 97378
rect 265072 97232 265124 97238
rect 265072 97174 265124 97180
rect 264888 96960 264940 96966
rect 264716 96920 264836 96948
rect 264428 96902 264480 96908
rect 264612 96892 264664 96898
rect 264612 96834 264664 96840
rect 264152 96688 264204 96694
rect 264152 96630 264204 96636
rect 264244 94512 264296 94518
rect 264244 94454 264296 94460
rect 263876 94240 263928 94246
rect 263876 94182 263928 94188
rect 263508 12028 263560 12034
rect 263508 11970 263560 11976
rect 261760 5160 261812 5166
rect 261760 5102 261812 5108
rect 262864 5160 262916 5166
rect 262864 5102 262916 5108
rect 261484 4140 261536 4146
rect 261484 4082 261536 4088
rect 260748 3936 260800 3942
rect 260748 3878 260800 3884
rect 259460 3732 259512 3738
rect 259460 3674 259512 3680
rect 260104 3732 260156 3738
rect 260104 3674 260156 3680
rect 258092 2094 258304 2122
rect 258276 480 258304 2094
rect 259472 480 259500 3674
rect 260656 3324 260708 3330
rect 260656 3266 260708 3272
rect 260668 480 260696 3266
rect 261772 480 261800 5102
rect 264256 3806 264284 94454
rect 264624 92342 264652 96834
rect 264704 96824 264756 96830
rect 264704 96766 264756 96772
rect 264612 92336 264664 92342
rect 264612 92278 264664 92284
rect 264336 91792 264388 91798
rect 264336 91734 264388 91740
rect 262956 3800 263008 3806
rect 262956 3742 263008 3748
rect 264244 3800 264296 3806
rect 264244 3742 264296 3748
rect 262968 480 262996 3742
rect 264348 3330 264376 91734
rect 264716 86698 264744 96766
rect 264704 86692 264756 86698
rect 264704 86634 264756 86640
rect 264808 85270 264836 96920
rect 264888 96902 264940 96908
rect 264796 85264 264848 85270
rect 264796 85206 264848 85212
rect 264900 3874 264928 96902
rect 265176 96762 265204 100028
rect 265452 97442 265480 100028
rect 265440 97436 265492 97442
rect 265440 97378 265492 97384
rect 265636 97034 265664 100028
rect 265624 97028 265676 97034
rect 265624 96970 265676 96976
rect 265820 96966 265848 100028
rect 265808 96960 265860 96966
rect 265808 96902 265860 96908
rect 265900 96892 265952 96898
rect 265900 96834 265952 96840
rect 265164 96756 265216 96762
rect 265164 96698 265216 96704
rect 265912 8158 265940 96834
rect 266004 92206 266032 100028
rect 266084 96960 266136 96966
rect 266084 96902 266136 96908
rect 265992 92200 266044 92206
rect 265992 92142 266044 92148
rect 266096 11898 266124 96902
rect 266188 96898 266216 100028
rect 266464 97034 266492 100028
rect 266268 97028 266320 97034
rect 266268 96970 266320 96976
rect 266452 97028 266504 97034
rect 266452 96970 266504 96976
rect 266176 96892 266228 96898
rect 266176 96834 266228 96840
rect 266176 96756 266228 96762
rect 266176 96698 266228 96704
rect 266188 11966 266216 96698
rect 266280 93702 266308 96970
rect 266648 96830 266676 100028
rect 266832 96898 266860 100028
rect 267016 96966 267044 100028
rect 267200 97782 267228 100028
rect 267292 100014 267398 100042
rect 267188 97776 267240 97782
rect 267188 97718 267240 97724
rect 267004 96960 267056 96966
rect 267292 96948 267320 100014
rect 267464 97028 267516 97034
rect 267464 96970 267516 96976
rect 267004 96902 267056 96908
rect 267200 96920 267320 96948
rect 267372 96960 267424 96966
rect 266820 96892 266872 96898
rect 266820 96834 266872 96840
rect 266636 96824 266688 96830
rect 266636 96766 266688 96772
rect 267004 96688 267056 96694
rect 267004 96630 267056 96636
rect 266268 93696 266320 93702
rect 266268 93638 266320 93644
rect 267016 85338 267044 96630
rect 267004 85332 267056 85338
rect 267004 85274 267056 85280
rect 266176 11960 266228 11966
rect 266176 11902 266228 11908
rect 266084 11892 266136 11898
rect 266084 11834 266136 11840
rect 265900 8152 265952 8158
rect 265900 8094 265952 8100
rect 267200 8022 267228 96920
rect 267372 96902 267424 96908
rect 267280 96824 267332 96830
rect 267280 96766 267332 96772
rect 267292 89690 267320 96766
rect 267280 89684 267332 89690
rect 267280 89626 267332 89632
rect 267384 11762 267412 96902
rect 267476 11830 267504 96970
rect 267556 96892 267608 96898
rect 267556 96834 267608 96840
rect 267464 11824 267516 11830
rect 267464 11766 267516 11772
rect 267372 11756 267424 11762
rect 267372 11698 267424 11704
rect 267568 8090 267596 96834
rect 267660 92138 267688 100028
rect 267844 96898 267872 100028
rect 268028 96966 268056 100028
rect 268226 100014 268332 100042
rect 268200 97640 268252 97646
rect 268200 97582 268252 97588
rect 268016 96960 268068 96966
rect 268016 96902 268068 96908
rect 267832 96892 267884 96898
rect 267832 96834 267884 96840
rect 267832 96008 267884 96014
rect 267832 95950 267884 95956
rect 267648 92132 267700 92138
rect 267648 92074 267700 92080
rect 267740 22772 267792 22778
rect 267740 22714 267792 22720
rect 267556 8084 267608 8090
rect 267556 8026 267608 8032
rect 267188 8016 267240 8022
rect 267188 7958 267240 7964
rect 266544 7608 266596 7614
rect 266544 7550 266596 7556
rect 265348 5296 265400 5302
rect 265348 5238 265400 5244
rect 264888 3868 264940 3874
rect 264888 3810 264940 3816
rect 264336 3324 264388 3330
rect 264336 3266 264388 3272
rect 264152 3052 264204 3058
rect 264152 2994 264204 3000
rect 264164 480 264192 2994
rect 265360 480 265388 5238
rect 266556 480 266584 7550
rect 267752 480 267780 22714
rect 267844 3058 267872 95950
rect 268212 92274 268240 97582
rect 268304 96914 268332 100014
rect 268396 97238 268424 100028
rect 268384 97232 268436 97238
rect 268384 97174 268436 97180
rect 268672 97034 268700 100028
rect 268764 100014 268870 100042
rect 268660 97028 268712 97034
rect 268660 96970 268712 96976
rect 268304 96886 268700 96914
rect 268200 92268 268252 92274
rect 268200 92210 268252 92216
rect 268672 89622 268700 96886
rect 268660 89616 268712 89622
rect 268660 89558 268712 89564
rect 268764 86630 268792 100014
rect 269040 97986 269068 100028
rect 269028 97980 269080 97986
rect 269028 97922 269080 97928
rect 269224 97034 269252 100028
rect 269028 97028 269080 97034
rect 269028 96970 269080 96976
rect 269212 97028 269264 97034
rect 269212 96970 269264 96976
rect 268936 96960 268988 96966
rect 268936 96902 268988 96908
rect 268844 96892 268896 96898
rect 268844 96834 268896 96840
rect 268752 86624 268804 86630
rect 268752 86566 268804 86572
rect 268856 83842 268884 96834
rect 268844 83836 268896 83842
rect 268844 83778 268896 83784
rect 268948 7954 268976 96902
rect 268936 7948 268988 7954
rect 268936 7890 268988 7896
rect 269040 7886 269068 96970
rect 269408 96694 269436 100028
rect 269684 96966 269712 100028
rect 269672 96960 269724 96966
rect 269672 96902 269724 96908
rect 269868 96762 269896 100028
rect 269948 96892 270000 96898
rect 269948 96834 270000 96840
rect 269856 96756 269908 96762
rect 269856 96698 269908 96704
rect 269396 96688 269448 96694
rect 269396 96630 269448 96636
rect 269028 7880 269080 7886
rect 269028 7822 269080 7828
rect 269960 7682 269988 96834
rect 270052 88058 270080 100028
rect 270236 97646 270264 100028
rect 270224 97640 270276 97646
rect 270224 97582 270276 97588
rect 270316 97028 270368 97034
rect 270316 96970 270368 96976
rect 270132 96960 270184 96966
rect 270132 96902 270184 96908
rect 270040 88052 270092 88058
rect 270040 87994 270092 88000
rect 270144 82414 270172 96902
rect 270224 96756 270276 96762
rect 270224 96698 270276 96704
rect 270132 82408 270184 82414
rect 270132 82350 270184 82356
rect 270236 7750 270264 96698
rect 270328 7818 270356 96970
rect 270420 96898 270448 100028
rect 270408 96892 270460 96898
rect 270408 96834 270460 96840
rect 270696 96830 270724 100028
rect 270880 96966 270908 100028
rect 271064 99278 271092 100028
rect 271262 100014 271368 100042
rect 271052 99272 271104 99278
rect 271052 99214 271104 99220
rect 271052 97436 271104 97442
rect 271052 97378 271104 97384
rect 270868 96960 270920 96966
rect 270868 96902 270920 96908
rect 270684 96824 270736 96830
rect 270684 96766 270736 96772
rect 270408 96688 270460 96694
rect 270408 96630 270460 96636
rect 270420 93634 270448 96630
rect 271064 96490 271092 97378
rect 271144 97300 271196 97306
rect 271144 97242 271196 97248
rect 271052 96484 271104 96490
rect 271052 96426 271104 96432
rect 270408 93628 270460 93634
rect 270408 93570 270460 93576
rect 270316 7812 270368 7818
rect 270316 7754 270368 7760
rect 270224 7744 270276 7750
rect 270224 7686 270276 7692
rect 269948 7676 270000 7682
rect 269948 7618 270000 7624
rect 268844 5092 268896 5098
rect 268844 5034 268896 5040
rect 267832 3052 267884 3058
rect 267832 2994 267884 3000
rect 268856 480 268884 5034
rect 271156 3602 271184 97242
rect 271236 97164 271288 97170
rect 271236 97106 271288 97112
rect 271248 96614 271276 97106
rect 271340 96914 271368 100014
rect 271432 97238 271460 100028
rect 271616 99210 271644 100028
rect 271604 99204 271656 99210
rect 271604 99146 271656 99152
rect 271420 97232 271472 97238
rect 271420 97174 271472 97180
rect 271788 96960 271840 96966
rect 271340 96886 271736 96914
rect 271788 96902 271840 96908
rect 271604 96824 271656 96830
rect 271604 96766 271656 96772
rect 271248 96586 271368 96614
rect 271236 96484 271288 96490
rect 271236 96426 271288 96432
rect 271248 82482 271276 96426
rect 271340 82550 271368 96586
rect 271616 90982 271644 96766
rect 271604 90976 271656 90982
rect 271604 90918 271656 90924
rect 271708 86562 271736 96886
rect 271696 86556 271748 86562
rect 271696 86498 271748 86504
rect 271328 82544 271380 82550
rect 271328 82486 271380 82492
rect 271236 82476 271288 82482
rect 271236 82418 271288 82424
rect 271800 5098 271828 96902
rect 271892 96762 271920 100028
rect 272076 97034 272104 100028
rect 272260 99142 272288 100028
rect 272248 99136 272300 99142
rect 272248 99078 272300 99084
rect 272340 97912 272392 97918
rect 272340 97854 272392 97860
rect 272248 97844 272300 97850
rect 272248 97786 272300 97792
rect 272260 97510 272288 97786
rect 272352 97578 272380 97854
rect 272340 97572 272392 97578
rect 272340 97514 272392 97520
rect 272248 97504 272300 97510
rect 272248 97446 272300 97452
rect 272064 97028 272116 97034
rect 272064 96970 272116 96976
rect 272444 96966 272472 100028
rect 272432 96960 272484 96966
rect 272432 96902 272484 96908
rect 272628 96830 272656 100028
rect 272904 96898 272932 100028
rect 272984 96960 273036 96966
rect 272984 96902 273036 96908
rect 272892 96892 272944 96898
rect 272892 96834 272944 96840
rect 272616 96824 272668 96830
rect 272616 96766 272668 96772
rect 271880 96756 271932 96762
rect 271880 96698 271932 96704
rect 272892 96756 272944 96762
rect 272892 96698 272944 96704
rect 272904 87990 272932 96698
rect 272892 87984 272944 87990
rect 272892 87926 272944 87932
rect 272996 85202 273024 96902
rect 272984 85196 273036 85202
rect 272984 85138 273036 85144
rect 273088 13734 273116 100028
rect 273272 96966 273300 100028
rect 273456 99074 273484 100028
rect 273654 100014 273852 100042
rect 273930 100014 274036 100042
rect 273444 99068 273496 99074
rect 273444 99010 273496 99016
rect 273260 96960 273312 96966
rect 273260 96902 273312 96908
rect 273168 96892 273220 96898
rect 273168 96834 273220 96840
rect 273076 13728 273128 13734
rect 273076 13670 273128 13676
rect 273180 7614 273208 96834
rect 273824 89714 273852 100014
rect 273904 96960 273956 96966
rect 273904 96902 273956 96908
rect 273916 94466 273944 96902
rect 274008 94602 274036 100014
rect 274100 96694 274128 100028
rect 274298 100014 274404 100042
rect 274180 97096 274232 97102
rect 274178 97064 274180 97073
rect 274232 97064 274234 97073
rect 274178 96999 274234 97008
rect 274088 96688 274140 96694
rect 274088 96630 274140 96636
rect 274376 96370 274404 100014
rect 274468 98122 274496 100028
rect 274652 99006 274680 100028
rect 274640 99000 274692 99006
rect 274640 98942 274692 98948
rect 274456 98116 274508 98122
rect 274456 98058 274508 98064
rect 274928 96830 274956 100028
rect 274916 96824 274968 96830
rect 274916 96766 274968 96772
rect 275112 96694 275140 100028
rect 275296 98938 275324 100028
rect 275494 100014 275600 100042
rect 275284 98932 275336 98938
rect 275284 98874 275336 98880
rect 275572 97050 275600 100014
rect 275664 97374 275692 100028
rect 275652 97368 275704 97374
rect 275652 97310 275704 97316
rect 275572 97022 275876 97050
rect 275652 96960 275704 96966
rect 275652 96902 275704 96908
rect 274548 96688 274600 96694
rect 274548 96630 274600 96636
rect 275100 96688 275152 96694
rect 275100 96630 275152 96636
rect 274376 96342 274496 96370
rect 274008 94574 274404 94602
rect 273916 94438 274312 94466
rect 273824 89686 274220 89714
rect 274192 13666 274220 89686
rect 274284 80918 274312 94438
rect 274272 80912 274324 80918
rect 274272 80854 274324 80860
rect 274376 80850 274404 94574
rect 274364 80844 274416 80850
rect 274364 80786 274416 80792
rect 274180 13660 274232 13666
rect 274180 13602 274232 13608
rect 274468 13598 274496 96342
rect 274560 92002 274588 96630
rect 275664 92070 275692 96902
rect 275744 96688 275796 96694
rect 275744 96630 275796 96636
rect 275652 92064 275704 92070
rect 275652 92006 275704 92012
rect 274548 91996 274600 92002
rect 274548 91938 274600 91944
rect 275756 80782 275784 96630
rect 275744 80776 275796 80782
rect 275744 80718 275796 80724
rect 274456 13592 274508 13598
rect 274456 13534 274508 13540
rect 275848 13462 275876 97022
rect 275940 96966 275968 100028
rect 275928 96960 275980 96966
rect 275928 96902 275980 96908
rect 276124 96830 276152 100028
rect 276308 96966 276336 100028
rect 276492 98870 276520 100028
rect 276480 98864 276532 98870
rect 276480 98806 276532 98812
rect 276572 97300 276624 97306
rect 276572 97242 276624 97248
rect 276296 96960 276348 96966
rect 276296 96902 276348 96908
rect 275928 96824 275980 96830
rect 275928 96766 275980 96772
rect 276112 96824 276164 96830
rect 276112 96766 276164 96772
rect 275940 13530 275968 96766
rect 276584 89714 276612 97242
rect 276676 96898 276704 100028
rect 276874 100014 277072 100042
rect 277150 100014 277256 100042
rect 276848 97368 276900 97374
rect 276848 97310 276900 97316
rect 276664 96892 276716 96898
rect 276664 96834 276716 96840
rect 276860 91934 276888 97310
rect 276940 96688 276992 96694
rect 276940 96630 276992 96636
rect 276848 91928 276900 91934
rect 276848 91870 276900 91876
rect 276584 89686 276704 89714
rect 276676 82346 276704 89686
rect 276664 82340 276716 82346
rect 276664 82282 276716 82288
rect 275928 13524 275980 13530
rect 275928 13466 275980 13472
rect 275836 13456 275888 13462
rect 275836 13398 275888 13404
rect 276952 13258 276980 96630
rect 277044 86494 277072 100014
rect 277228 97374 277256 100014
rect 277216 97368 277268 97374
rect 277216 97310 277268 97316
rect 277216 96892 277268 96898
rect 277216 96834 277268 96840
rect 277124 96824 277176 96830
rect 277124 96766 277176 96772
rect 277032 86488 277084 86494
rect 277032 86430 277084 86436
rect 277136 13394 277164 96766
rect 277124 13388 277176 13394
rect 277124 13330 277176 13336
rect 277228 13326 277256 96834
rect 277320 96694 277348 100028
rect 277504 96694 277532 100028
rect 277702 100014 277808 100042
rect 277886 100014 278084 100042
rect 277308 96688 277360 96694
rect 277308 96630 277360 96636
rect 277492 96688 277544 96694
rect 277492 96630 277544 96636
rect 277780 93566 277808 100014
rect 277952 97640 278004 97646
rect 277952 97582 278004 97588
rect 277964 97374 277992 97582
rect 277952 97368 278004 97374
rect 277952 97310 278004 97316
rect 278056 94586 278084 100014
rect 278148 98054 278176 100028
rect 278332 99374 278360 100028
rect 278332 99346 278452 99374
rect 278228 98116 278280 98122
rect 278228 98058 278280 98064
rect 278136 98048 278188 98054
rect 278136 97990 278188 97996
rect 278136 97504 278188 97510
rect 278136 97446 278188 97452
rect 278148 97238 278176 97446
rect 278240 97238 278268 98058
rect 278320 97436 278372 97442
rect 278320 97378 278372 97384
rect 278136 97232 278188 97238
rect 278136 97174 278188 97180
rect 278228 97232 278280 97238
rect 278228 97174 278280 97180
rect 278332 97050 278360 97378
rect 278240 97034 278360 97050
rect 278228 97028 278360 97034
rect 278280 97022 278360 97028
rect 278228 96970 278280 96976
rect 278424 96694 278452 99346
rect 278320 96688 278372 96694
rect 278320 96630 278372 96636
rect 278412 96688 278464 96694
rect 278412 96630 278464 96636
rect 278044 94580 278096 94586
rect 278044 94522 278096 94528
rect 278228 94512 278280 94518
rect 278228 94454 278280 94460
rect 277768 93560 277820 93566
rect 277768 93502 277820 93508
rect 277216 13320 277268 13326
rect 277216 13262 277268 13268
rect 276940 13252 276992 13258
rect 276940 13194 276992 13200
rect 273168 7608 273220 7614
rect 273168 7550 273220 7556
rect 271788 5092 271840 5098
rect 271788 5034 271840 5040
rect 278240 4146 278268 94454
rect 278332 16574 278360 96630
rect 278412 94580 278464 94586
rect 278412 94522 278464 94528
rect 278424 86426 278452 94522
rect 278412 86420 278464 86426
rect 278412 86362 278464 86368
rect 278516 85134 278544 100028
rect 278608 100014 278714 100042
rect 278608 94518 278636 100014
rect 278884 99346 278912 100028
rect 278872 99340 278924 99346
rect 278872 99282 278924 99288
rect 278688 97164 278740 97170
rect 278688 97106 278740 97112
rect 278700 97073 278728 97106
rect 278686 97064 278742 97073
rect 279160 97034 279188 100028
rect 279344 97481 279372 100028
rect 279542 100014 279648 100042
rect 279726 100014 279832 100042
rect 279910 100014 280108 100042
rect 279330 97472 279386 97481
rect 279330 97407 279386 97416
rect 278686 96999 278742 97008
rect 279148 97028 279200 97034
rect 279148 96970 279200 96976
rect 278688 96688 278740 96694
rect 278688 96630 278740 96636
rect 278596 94512 278648 94518
rect 278596 94454 278648 94460
rect 278700 90914 278728 96630
rect 279620 91866 279648 100014
rect 279804 99374 279832 100014
rect 279804 99346 280016 99374
rect 279608 91860 279660 91866
rect 279608 91802 279660 91808
rect 278688 90908 278740 90914
rect 278688 90850 278740 90856
rect 278504 85128 278556 85134
rect 278504 85070 278556 85076
rect 278332 16546 278452 16574
rect 277124 4140 277176 4146
rect 277124 4082 277176 4088
rect 278228 4140 278280 4146
rect 278228 4082 278280 4088
rect 276020 3800 276072 3806
rect 276020 3742 276072 3748
rect 271236 3664 271288 3670
rect 271236 3606 271288 3612
rect 271052 3596 271104 3602
rect 271052 3538 271104 3544
rect 271144 3596 271196 3602
rect 271144 3538 271196 3544
rect 271064 3398 271092 3538
rect 270040 3392 270092 3398
rect 270040 3334 270092 3340
rect 271052 3392 271104 3398
rect 271052 3334 271104 3340
rect 270052 480 270080 3334
rect 271248 480 271276 3606
rect 274824 3596 274876 3602
rect 274824 3538 274876 3544
rect 272432 3392 272484 3398
rect 272432 3334 272484 3340
rect 272444 480 272472 3334
rect 273628 3324 273680 3330
rect 273628 3266 273680 3272
rect 273640 480 273668 3266
rect 274836 480 274864 3538
rect 276032 480 276060 3742
rect 277136 480 277164 4082
rect 278424 3806 278452 16546
rect 279988 13190 280016 99346
rect 279976 13184 280028 13190
rect 279976 13126 280028 13132
rect 279516 5024 279568 5030
rect 279516 4966 279568 4972
rect 278412 3800 278464 3806
rect 278412 3742 278464 3748
rect 278320 3732 278372 3738
rect 278320 3674 278372 3680
rect 278332 480 278360 3674
rect 279528 480 279556 4966
rect 280080 3738 280108 100014
rect 280172 96966 280200 100028
rect 280160 96960 280212 96966
rect 280160 96902 280212 96908
rect 280356 96830 280384 100028
rect 280540 97345 280568 100028
rect 280526 97336 280582 97345
rect 280526 97271 280582 97280
rect 280344 96824 280396 96830
rect 280344 96766 280396 96772
rect 280724 96694 280752 100028
rect 280908 96898 280936 100028
rect 281000 100014 281106 100042
rect 281276 100014 281382 100042
rect 280896 96892 280948 96898
rect 280896 96834 280948 96840
rect 280712 96688 280764 96694
rect 280712 96630 280764 96636
rect 280068 3732 280120 3738
rect 280068 3674 280120 3680
rect 281000 3670 281028 100014
rect 281172 97028 281224 97034
rect 281172 96970 281224 96976
rect 281184 96830 281212 96970
rect 281080 96824 281132 96830
rect 281080 96766 281132 96772
rect 281172 96824 281224 96830
rect 281172 96766 281224 96772
rect 281092 13122 281120 96766
rect 281172 96688 281224 96694
rect 281172 96630 281224 96636
rect 281080 13116 281132 13122
rect 281080 13058 281132 13064
rect 281184 9042 281212 96630
rect 281172 9036 281224 9042
rect 281172 8978 281224 8984
rect 281276 8974 281304 100014
rect 281356 96960 281408 96966
rect 281356 96902 281408 96908
rect 281368 9110 281396 96902
rect 281448 96892 281500 96898
rect 281448 96834 281500 96840
rect 281460 89486 281488 96834
rect 281552 96694 281580 100028
rect 281736 97102 281764 100028
rect 281724 97096 281776 97102
rect 281724 97038 281776 97044
rect 281540 96688 281592 96694
rect 281540 96630 281592 96636
rect 281920 96286 281948 100028
rect 281908 96280 281960 96286
rect 281908 96222 281960 96228
rect 282104 90778 282132 100028
rect 282394 100014 282500 100042
rect 282368 97980 282420 97986
rect 282368 97922 282420 97928
rect 282184 97232 282236 97238
rect 282184 97174 282236 97180
rect 282196 96898 282224 97174
rect 282380 97034 282408 97922
rect 282368 97028 282420 97034
rect 282368 96970 282420 96976
rect 282184 96892 282236 96898
rect 282184 96834 282236 96840
rect 282276 96824 282328 96830
rect 282276 96766 282328 96772
rect 282092 90772 282144 90778
rect 282092 90714 282144 90720
rect 282184 90364 282236 90370
rect 282184 90306 282236 90312
rect 281448 89480 281500 89486
rect 281448 89422 281500 89428
rect 281356 9104 281408 9110
rect 281356 9046 281408 9052
rect 281264 8968 281316 8974
rect 281264 8910 281316 8916
rect 280988 3664 281040 3670
rect 280988 3606 281040 3612
rect 281908 3596 281960 3602
rect 281908 3538 281960 3544
rect 280712 3528 280764 3534
rect 280712 3470 280764 3476
rect 280724 480 280752 3470
rect 281920 480 281948 3538
rect 282196 3534 282224 90306
rect 282288 85066 282316 96766
rect 282276 85060 282328 85066
rect 282276 85002 282328 85008
rect 282472 24138 282500 100014
rect 282564 96150 282592 100028
rect 282656 100014 282762 100042
rect 282656 99374 282684 100014
rect 282656 99346 282776 99374
rect 282644 97368 282696 97374
rect 282644 97310 282696 97316
rect 282656 97209 282684 97310
rect 282642 97200 282698 97209
rect 282642 97135 282698 97144
rect 282552 96144 282604 96150
rect 282552 96086 282604 96092
rect 282748 90846 282776 99346
rect 282932 96694 282960 100028
rect 283012 97300 283064 97306
rect 283012 97242 283064 97248
rect 283024 97209 283052 97242
rect 283010 97200 283066 97209
rect 283010 97135 283066 97144
rect 282828 96688 282880 96694
rect 282828 96630 282880 96636
rect 282920 96688 282972 96694
rect 282920 96630 282972 96636
rect 282736 90840 282788 90846
rect 282736 90782 282788 90788
rect 282840 84194 282868 96630
rect 283116 96218 283144 100028
rect 283392 98802 283420 100028
rect 283380 98796 283432 98802
rect 283380 98738 283432 98744
rect 283576 96830 283604 100028
rect 283656 97368 283708 97374
rect 283656 97310 283708 97316
rect 283668 96898 283696 97310
rect 283656 96892 283708 96898
rect 283656 96834 283708 96840
rect 283564 96824 283616 96830
rect 283564 96766 283616 96772
rect 283760 96354 283788 100028
rect 283840 96892 283892 96898
rect 283840 96834 283892 96840
rect 283748 96348 283800 96354
rect 283748 96290 283800 96296
rect 283104 96212 283156 96218
rect 283104 96154 283156 96160
rect 282748 84166 282868 84194
rect 282748 83774 282776 84166
rect 282736 83768 282788 83774
rect 282736 83710 282788 83716
rect 283852 83706 283880 96834
rect 283944 90710 283972 100028
rect 284128 96898 284156 100028
rect 284300 97096 284352 97102
rect 284300 97038 284352 97044
rect 284116 96892 284168 96898
rect 284116 96834 284168 96840
rect 284024 96824 284076 96830
rect 284024 96766 284076 96772
rect 283932 90704 283984 90710
rect 283932 90646 283984 90652
rect 284036 84930 284064 96766
rect 284312 96694 284340 97038
rect 284116 96688 284168 96694
rect 284116 96630 284168 96636
rect 284300 96688 284352 96694
rect 284300 96630 284352 96636
rect 284128 84998 284156 96630
rect 284404 96422 284432 100028
rect 284588 96830 284616 100028
rect 284786 100014 284892 100042
rect 284576 96824 284628 96830
rect 284576 96766 284628 96772
rect 284392 96416 284444 96422
rect 284392 96358 284444 96364
rect 284392 95940 284444 95946
rect 284392 95882 284444 95888
rect 284116 84992 284168 84998
rect 284116 84934 284168 84940
rect 284024 84924 284076 84930
rect 284024 84866 284076 84872
rect 283840 83700 283892 83706
rect 283840 83642 283892 83648
rect 282460 24132 282512 24138
rect 282460 24074 282512 24080
rect 284300 17264 284352 17270
rect 284300 17206 284352 17212
rect 284312 3534 284340 17206
rect 284404 3602 284432 95882
rect 284864 93854 284892 100014
rect 284956 96490 284984 100028
rect 285140 96898 285168 100028
rect 285232 100014 285430 100042
rect 285128 96892 285180 96898
rect 285128 96834 285180 96840
rect 284944 96484 284996 96490
rect 284944 96426 284996 96432
rect 284864 93826 285168 93854
rect 285140 83638 285168 93826
rect 285128 83632 285180 83638
rect 285128 83574 285180 83580
rect 285232 17270 285260 100014
rect 285404 96892 285456 96898
rect 285404 96834 285456 96840
rect 285312 96824 285364 96830
rect 285312 96766 285364 96772
rect 285324 90642 285352 96766
rect 285312 90636 285364 90642
rect 285312 90578 285364 90584
rect 285416 89418 285444 96834
rect 285600 96082 285628 100028
rect 285784 96898 285812 100028
rect 285772 96892 285824 96898
rect 285772 96834 285824 96840
rect 285968 96830 285996 100028
rect 285956 96824 286008 96830
rect 285956 96766 286008 96772
rect 285588 96076 285640 96082
rect 285588 96018 285640 96024
rect 286152 96014 286180 100028
rect 286336 97102 286364 100028
rect 286520 100014 286626 100042
rect 286324 97096 286376 97102
rect 286324 97038 286376 97044
rect 286416 96892 286468 96898
rect 286416 96834 286468 96840
rect 286140 96008 286192 96014
rect 286140 95950 286192 95956
rect 286428 90574 286456 96834
rect 286416 90568 286468 90574
rect 286416 90510 286468 90516
rect 285404 89412 285456 89418
rect 285404 89354 285456 89360
rect 286520 21418 286548 100014
rect 286796 98054 286824 100028
rect 286888 100014 286994 100042
rect 286784 98048 286836 98054
rect 286784 97990 286836 97996
rect 286692 97096 286744 97102
rect 286692 97038 286744 97044
rect 286784 97096 286836 97102
rect 286784 97038 286836 97044
rect 286600 96824 286652 96830
rect 286600 96766 286652 96772
rect 286508 21412 286560 21418
rect 286508 21354 286560 21360
rect 285220 17264 285272 17270
rect 285220 17206 285272 17212
rect 286612 16574 286640 96766
rect 286704 89282 286732 97038
rect 286796 96762 286824 97038
rect 286784 96756 286836 96762
rect 286784 96698 286836 96704
rect 286888 89350 286916 100014
rect 286968 98048 287020 98054
rect 286968 97990 287020 97996
rect 286980 94926 287008 97990
rect 287164 96898 287192 100028
rect 287152 96892 287204 96898
rect 287152 96834 287204 96840
rect 287348 95538 287376 100028
rect 287638 100014 287744 100042
rect 287822 100014 287928 100042
rect 287336 95532 287388 95538
rect 287336 95474 287388 95480
rect 286968 94920 287020 94926
rect 286968 94862 287020 94868
rect 287716 90506 287744 100014
rect 287900 96914 287928 100014
rect 287992 97170 288020 100028
rect 288084 100014 288190 100042
rect 287980 97164 288032 97170
rect 287980 97106 288032 97112
rect 287900 96886 288020 96914
rect 287888 96824 287940 96830
rect 287888 96766 287940 96772
rect 287704 90500 287756 90506
rect 287704 90442 287756 90448
rect 286876 89344 286928 89350
rect 286876 89286 286928 89292
rect 286692 89276 286744 89282
rect 286692 89218 286744 89224
rect 287900 18630 287928 96766
rect 287888 18624 287940 18630
rect 287888 18566 287940 18572
rect 286612 16546 286732 16574
rect 284484 6588 284536 6594
rect 284484 6530 284536 6536
rect 284392 3596 284444 3602
rect 284392 3538 284444 3544
rect 282184 3528 282236 3534
rect 282184 3470 282236 3476
rect 283104 3528 283156 3534
rect 283104 3470 283156 3476
rect 284300 3528 284352 3534
rect 284300 3470 284352 3476
rect 283116 480 283144 3470
rect 284496 762 284524 6530
rect 286704 5030 286732 16546
rect 287992 6254 288020 96886
rect 288084 89146 288112 100014
rect 288256 97164 288308 97170
rect 288256 97106 288308 97112
rect 288164 96892 288216 96898
rect 288164 96834 288216 96840
rect 288072 89140 288124 89146
rect 288072 89082 288124 89088
rect 288176 82278 288204 96834
rect 288268 94994 288296 97106
rect 288360 96830 288388 100028
rect 288636 96898 288664 100028
rect 288820 97170 288848 100028
rect 288808 97164 288860 97170
rect 288808 97106 288860 97112
rect 288624 96892 288676 96898
rect 288624 96834 288676 96840
rect 289004 96830 289032 100028
rect 288348 96824 288400 96830
rect 288348 96766 288400 96772
rect 288992 96824 289044 96830
rect 288992 96766 289044 96772
rect 289188 96762 289216 100028
rect 289268 96892 289320 96898
rect 289268 96834 289320 96840
rect 289176 96756 289228 96762
rect 289176 96698 289228 96704
rect 288256 94988 288308 94994
rect 288256 94930 288308 94936
rect 288164 82272 288216 82278
rect 288164 82214 288216 82220
rect 287796 6248 287848 6254
rect 287796 6190 287848 6196
rect 287980 6248 288032 6254
rect 287980 6190 288032 6196
rect 286692 5024 286744 5030
rect 286692 4966 286744 4972
rect 286600 4956 286652 4962
rect 286600 4898 286652 4904
rect 284668 4140 284720 4146
rect 284668 4082 284720 4088
rect 284680 3738 284708 4082
rect 284668 3732 284720 3738
rect 284668 3674 284720 3680
rect 285404 3528 285456 3534
rect 285404 3470 285456 3476
rect 284404 734 284524 762
rect 284404 626 284432 734
rect 284312 598 284432 626
rect 284312 480 284340 598
rect 285416 480 285444 3470
rect 286612 480 286640 4898
rect 287808 480 287836 6190
rect 289280 4962 289308 96834
rect 289372 89078 289400 100028
rect 289464 100014 289662 100042
rect 289360 89072 289412 89078
rect 289360 89014 289412 89020
rect 289464 14482 289492 100014
rect 289728 97164 289780 97170
rect 289728 97106 289780 97112
rect 289544 96824 289596 96830
rect 289544 96766 289596 96772
rect 289556 14550 289584 96766
rect 289636 96756 289688 96762
rect 289636 96698 289688 96704
rect 289544 14544 289596 14550
rect 289544 14486 289596 14492
rect 289452 14476 289504 14482
rect 289452 14418 289504 14424
rect 289268 4956 289320 4962
rect 289268 4898 289320 4904
rect 289648 4894 289676 96698
rect 289740 91798 289768 97106
rect 289832 95985 289860 100028
rect 290016 98734 290044 100028
rect 290004 98728 290056 98734
rect 290004 98670 290056 98676
rect 290200 96762 290228 100028
rect 290188 96756 290240 96762
rect 290188 96698 290240 96704
rect 289818 95976 289874 95985
rect 289818 95911 289874 95920
rect 290384 94790 290412 100028
rect 290568 96898 290596 100028
rect 290752 100014 290858 100042
rect 290556 96892 290608 96898
rect 290556 96834 290608 96840
rect 290372 94784 290424 94790
rect 290372 94726 290424 94732
rect 289728 91792 289780 91798
rect 289728 91734 289780 91740
rect 290752 84862 290780 100014
rect 290924 96892 290976 96898
rect 290924 96834 290976 96840
rect 290832 96756 290884 96762
rect 290832 96698 290884 96704
rect 290740 84856 290792 84862
rect 290740 84798 290792 84804
rect 290844 83570 290872 96698
rect 290936 90438 290964 96834
rect 291028 94722 291056 100028
rect 291212 96762 291240 100028
rect 291396 96898 291424 100028
rect 291384 96892 291436 96898
rect 291384 96834 291436 96840
rect 291200 96756 291252 96762
rect 291200 96698 291252 96704
rect 291016 94716 291068 94722
rect 291016 94658 291068 94664
rect 291580 94654 291608 100028
rect 291856 96830 291884 100028
rect 291936 96892 291988 96898
rect 291936 96834 291988 96840
rect 291844 96824 291896 96830
rect 291844 96766 291896 96772
rect 291568 94648 291620 94654
rect 291568 94590 291620 94596
rect 290924 90432 290976 90438
rect 290924 90374 290976 90380
rect 290832 83564 290884 83570
rect 290832 83506 290884 83512
rect 291948 6186 291976 96834
rect 292040 26926 292068 100028
rect 292224 97170 292252 100028
rect 292316 100014 292422 100042
rect 292212 97164 292264 97170
rect 292212 97106 292264 97112
rect 292316 96914 292344 100014
rect 292488 97164 292540 97170
rect 292488 97106 292540 97112
rect 292224 96886 292344 96914
rect 292120 96756 292172 96762
rect 292120 96698 292172 96704
rect 292132 89214 292160 96698
rect 292120 89208 292172 89214
rect 292120 89150 292172 89156
rect 292224 87786 292252 96886
rect 292304 96824 292356 96830
rect 292304 96766 292356 96772
rect 292316 87854 292344 96766
rect 292500 94858 292528 97106
rect 292592 96830 292620 100028
rect 292580 96824 292632 96830
rect 292580 96766 292632 96772
rect 292488 94852 292540 94858
rect 292488 94794 292540 94800
rect 292868 94586 292896 100028
rect 293052 96898 293080 100028
rect 293040 96892 293092 96898
rect 293040 96834 293092 96840
rect 292856 94580 292908 94586
rect 292856 94522 292908 94528
rect 292304 87848 292356 87854
rect 292304 87790 292356 87796
rect 292212 87780 292264 87786
rect 292212 87722 292264 87728
rect 293236 82210 293264 100028
rect 293328 100014 293434 100042
rect 293328 95062 293356 100014
rect 293408 96892 293460 96898
rect 293408 96834 293460 96840
rect 293500 96892 293552 96898
rect 293500 96834 293552 96840
rect 293316 95056 293368 95062
rect 293316 94998 293368 95004
rect 293420 93498 293448 96834
rect 293408 93492 293460 93498
rect 293408 93434 293460 93440
rect 293224 82204 293276 82210
rect 293224 82146 293276 82152
rect 292028 26920 292080 26926
rect 292028 26862 292080 26868
rect 293512 22778 293540 96834
rect 293604 89010 293632 100028
rect 293880 96898 293908 100028
rect 293868 96892 293920 96898
rect 293868 96834 293920 96840
rect 293684 96824 293736 96830
rect 293684 96766 293736 96772
rect 293592 89004 293644 89010
rect 293592 88946 293644 88952
rect 293696 83502 293724 96766
rect 294064 95849 294092 100028
rect 294262 100014 294368 100042
rect 294446 100014 294552 100042
rect 294340 95946 294368 100014
rect 294328 95940 294380 95946
rect 294328 95882 294380 95888
rect 294050 95840 294106 95849
rect 294050 95775 294106 95784
rect 294524 93854 294552 100014
rect 294616 96898 294644 100028
rect 294906 100014 295012 100042
rect 294604 96892 294656 96898
rect 294604 96834 294656 96840
rect 294880 96756 294932 96762
rect 294880 96698 294932 96704
rect 294524 93826 294828 93854
rect 293684 83496 293736 83502
rect 293684 83438 293736 83444
rect 294800 82142 294828 93826
rect 294788 82136 294840 82142
rect 294788 82078 294840 82084
rect 294892 28286 294920 96698
rect 294984 87922 295012 100014
rect 295076 96762 295104 100028
rect 295168 100014 295274 100042
rect 295064 96756 295116 96762
rect 295064 96698 295116 96704
rect 295064 95940 295116 95946
rect 295064 95882 295116 95888
rect 294972 87916 295024 87922
rect 294972 87858 295024 87864
rect 295076 87718 295104 95882
rect 295168 93362 295196 100014
rect 295444 96898 295472 100028
rect 295248 96892 295300 96898
rect 295248 96834 295300 96840
rect 295432 96892 295484 96898
rect 295432 96834 295484 96840
rect 295260 93430 295288 96834
rect 295628 96830 295656 100028
rect 295616 96824 295668 96830
rect 295616 96766 295668 96772
rect 295812 96762 295840 100028
rect 295984 98048 296036 98054
rect 295984 97990 296036 97996
rect 295800 96756 295852 96762
rect 295800 96698 295852 96704
rect 295340 95940 295392 95946
rect 295340 95882 295392 95888
rect 295352 95538 295380 95882
rect 295340 95532 295392 95538
rect 295340 95474 295392 95480
rect 295996 95130 296024 97990
rect 296088 97170 296116 100028
rect 296180 100014 296286 100042
rect 296364 100014 296470 100042
rect 296548 100014 296654 100042
rect 296076 97164 296128 97170
rect 296076 97106 296128 97112
rect 296076 96892 296128 96898
rect 296076 96834 296128 96840
rect 295984 95124 296036 95130
rect 295984 95066 296036 95072
rect 295248 93424 295300 93430
rect 295248 93366 295300 93372
rect 295156 93356 295208 93362
rect 295156 93298 295208 93304
rect 296088 90370 296116 96834
rect 296076 90364 296128 90370
rect 296076 90306 296128 90312
rect 295064 87712 295116 87718
rect 295064 87654 295116 87660
rect 294880 28280 294932 28286
rect 294880 28222 294932 28228
rect 296180 25566 296208 100014
rect 296364 98054 296392 100014
rect 296352 98048 296404 98054
rect 296352 97990 296404 97996
rect 296352 97164 296404 97170
rect 296352 97106 296404 97112
rect 296260 96824 296312 96830
rect 296260 96766 296312 96772
rect 296168 25560 296220 25566
rect 296168 25502 296220 25508
rect 293500 22772 293552 22778
rect 293500 22714 293552 22720
rect 291384 6180 291436 6186
rect 291384 6122 291436 6128
rect 291936 6180 291988 6186
rect 291936 6122 291988 6128
rect 290188 5228 290240 5234
rect 290188 5170 290240 5176
rect 288992 4888 289044 4894
rect 288992 4830 289044 4836
rect 289636 4888 289688 4894
rect 289636 4830 289688 4836
rect 289004 480 289032 4830
rect 290200 480 290228 5170
rect 291396 480 291424 6122
rect 296272 4826 296300 96766
rect 296364 87650 296392 97106
rect 296548 96914 296576 100014
rect 296628 97164 296680 97170
rect 296628 97106 296680 97112
rect 296456 96886 296576 96914
rect 296352 87644 296404 87650
rect 296352 87586 296404 87592
rect 296456 86290 296484 96886
rect 296536 96756 296588 96762
rect 296536 96698 296588 96704
rect 296548 93294 296576 96698
rect 296640 96694 296668 97106
rect 296824 96830 296852 100028
rect 297100 98666 297128 100028
rect 297088 98660 297140 98666
rect 297088 98602 297140 98608
rect 296812 96824 296864 96830
rect 296812 96766 296864 96772
rect 296628 96688 296680 96694
rect 296628 96630 296680 96636
rect 297284 94518 297312 100028
rect 297482 100014 297588 100042
rect 297560 96914 297588 100014
rect 297652 97034 297680 100028
rect 297640 97028 297692 97034
rect 297640 96970 297692 96976
rect 297560 96886 297772 96914
rect 297640 96824 297692 96830
rect 297640 96766 297692 96772
rect 297272 94512 297324 94518
rect 297272 94454 297324 94460
rect 296536 93288 296588 93294
rect 296536 93230 296588 93236
rect 297652 86358 297680 96766
rect 297640 86352 297692 86358
rect 297640 86294 297692 86300
rect 296444 86284 296496 86290
rect 296444 86226 296496 86232
rect 297744 80714 297772 96886
rect 297836 89554 297864 100028
rect 298112 97034 298140 100028
rect 298008 97028 298060 97034
rect 298008 96970 298060 96976
rect 298100 97028 298152 97034
rect 298100 96970 298152 96976
rect 298020 93226 298048 96970
rect 298296 96830 298324 100028
rect 298480 96898 298508 100028
rect 298664 96966 298692 100028
rect 298862 100014 298968 100042
rect 298652 96960 298704 96966
rect 298652 96902 298704 96908
rect 298468 96892 298520 96898
rect 298468 96834 298520 96840
rect 298284 96824 298336 96830
rect 298284 96766 298336 96772
rect 298008 93220 298060 93226
rect 298008 93162 298060 93168
rect 297824 89548 297876 89554
rect 297824 89490 297876 89496
rect 297732 80708 297784 80714
rect 297732 80650 297784 80656
rect 298100 10328 298152 10334
rect 298100 10270 298152 10276
rect 297272 6520 297324 6526
rect 297272 6462 297324 6468
rect 293684 4820 293736 4826
rect 293684 4762 293736 4768
rect 296260 4820 296312 4826
rect 296260 4762 296312 4768
rect 292580 4140 292632 4146
rect 292580 4082 292632 4088
rect 292592 480 292620 4082
rect 293696 480 293724 4762
rect 294880 3460 294932 3466
rect 294880 3402 294932 3408
rect 294892 480 294920 3402
rect 296076 3392 296128 3398
rect 296076 3334 296128 3340
rect 296088 480 296116 3334
rect 297284 480 297312 6462
rect 298112 490 298140 10270
rect 298940 3466 298968 100014
rect 299124 97209 299152 100028
rect 299110 97200 299166 97209
rect 299110 97135 299166 97144
rect 299112 97028 299164 97034
rect 299112 96970 299164 96976
rect 299020 96960 299072 96966
rect 299020 96902 299072 96908
rect 299032 15910 299060 96902
rect 299124 15978 299152 96970
rect 299204 96892 299256 96898
rect 299204 96834 299256 96840
rect 299112 15972 299164 15978
rect 299112 15914 299164 15920
rect 299020 15904 299072 15910
rect 299020 15846 299072 15852
rect 299216 10334 299244 96834
rect 299204 10328 299256 10334
rect 299204 10270 299256 10276
rect 298928 3460 298980 3466
rect 298928 3402 298980 3408
rect 299308 3262 299336 100028
rect 299492 99414 299520 100028
rect 299690 100014 299796 100042
rect 299768 99906 299796 100014
rect 299952 99906 299980 100150
rect 299768 99878 299980 99906
rect 299480 99408 299532 99414
rect 299480 99350 299532 99356
rect 304264 97232 304316 97238
rect 304264 97174 304316 97180
rect 299388 96824 299440 96830
rect 299388 96766 299440 96772
rect 299400 93158 299428 96766
rect 301504 96756 301556 96762
rect 301504 96698 301556 96704
rect 299664 95736 299716 95742
rect 299664 95678 299716 95684
rect 299480 95668 299532 95674
rect 299480 95610 299532 95616
rect 299388 93152 299440 93158
rect 299388 93094 299440 93100
rect 299492 3482 299520 95610
rect 299572 95600 299624 95606
rect 299572 95542 299624 95548
rect 299584 4146 299612 95542
rect 299676 16574 299704 95678
rect 301516 80986 301544 96698
rect 302884 96688 302936 96694
rect 302884 96630 302936 96636
rect 302332 95804 302384 95810
rect 302332 95746 302384 95752
rect 302240 94172 302292 94178
rect 302240 94114 302292 94120
rect 301504 80980 301556 80986
rect 301504 80922 301556 80928
rect 300860 19984 300912 19990
rect 300860 19926 300912 19932
rect 300872 16574 300900 19926
rect 299676 16546 299796 16574
rect 300872 16546 301544 16574
rect 299572 4140 299624 4146
rect 299572 4082 299624 4088
rect 299492 3454 299704 3482
rect 299296 3256 299348 3262
rect 299296 3198 299348 3204
rect 298296 598 298508 626
rect 298296 490 298324 598
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298112 462 298324 490
rect 298480 480 298508 598
rect 299676 480 299704 3454
rect 299768 3398 299796 16546
rect 300768 3528 300820 3534
rect 300768 3470 300820 3476
rect 299756 3392 299808 3398
rect 299756 3334 299808 3340
rect 300780 480 300808 3470
rect 301516 490 301544 16546
rect 302252 3346 302280 94114
rect 302344 3534 302372 95746
rect 302896 79354 302924 96630
rect 303620 90160 303672 90166
rect 303620 90102 303672 90108
rect 302884 79348 302936 79354
rect 302884 79290 302936 79296
rect 303632 16574 303660 90102
rect 303632 16546 303936 16574
rect 302332 3528 302384 3534
rect 302332 3470 302384 3476
rect 302252 3318 303200 3346
rect 301792 598 302004 626
rect 301792 490 301820 598
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301516 462 301820 490
rect 301976 480 302004 598
rect 303172 480 303200 3318
rect 303908 490 303936 16546
rect 304276 5302 304304 97174
rect 305656 33114 305684 300154
rect 306380 94308 306432 94314
rect 306380 94250 306432 94256
rect 305644 33108 305696 33114
rect 305644 33050 305696 33056
rect 304264 5296 304316 5302
rect 304264 5238 304316 5244
rect 305552 4072 305604 4078
rect 305552 4014 305604 4020
rect 304184 598 304396 626
rect 304184 490 304212 598
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 303908 462 304212 490
rect 304368 480 304396 598
rect 305564 480 305592 4014
rect 306392 490 306420 94250
rect 307036 86970 307064 300222
rect 309140 94376 309192 94382
rect 309140 94318 309192 94324
rect 307024 86964 307076 86970
rect 307024 86906 307076 86912
rect 307024 85468 307076 85474
rect 307024 85410 307076 85416
rect 307036 3398 307064 85410
rect 309152 16574 309180 94318
rect 309796 73166 309824 301378
rect 313924 300144 313976 300150
rect 313924 300086 313976 300092
rect 313936 113150 313964 300086
rect 316696 227050 316724 302942
rect 318064 298512 318116 298518
rect 318064 298454 318116 298460
rect 316684 227044 316736 227050
rect 316684 226986 316736 226992
rect 318076 194478 318104 298454
rect 322204 298308 322256 298314
rect 322204 298250 322256 298256
rect 320824 294024 320876 294030
rect 320824 293966 320876 293972
rect 318064 194472 318116 194478
rect 318064 194414 318116 194420
rect 320836 122806 320864 293966
rect 322216 195974 322244 298250
rect 324964 295928 325016 295934
rect 324964 295870 325016 295876
rect 324976 267714 325004 295870
rect 352564 295860 352616 295866
rect 352564 295802 352616 295808
rect 352576 270502 352604 295802
rect 359464 291236 359516 291242
rect 359464 291178 359516 291184
rect 353944 285728 353996 285734
rect 353944 285670 353996 285676
rect 352564 270496 352616 270502
rect 352564 270438 352616 270444
rect 324964 267708 325016 267714
rect 324964 267650 325016 267656
rect 353956 266257 353984 285670
rect 356704 281580 356756 281586
rect 356704 281522 356756 281528
rect 353942 266248 353998 266257
rect 353942 266183 353998 266192
rect 356716 266121 356744 281522
rect 358084 280152 358136 280158
rect 358084 280094 358136 280100
rect 358096 278798 358124 280094
rect 358084 278792 358136 278798
rect 358084 278734 358136 278740
rect 358096 271114 358124 278734
rect 358084 271108 358136 271114
rect 358084 271050 358136 271056
rect 356702 266112 356758 266121
rect 356702 266047 356758 266056
rect 358912 223916 358964 223922
rect 358912 223858 358964 223864
rect 358924 222154 358952 223858
rect 358912 222148 358964 222154
rect 358912 222090 358964 222096
rect 359372 198756 359424 198762
rect 359372 198698 359424 198704
rect 359384 197062 359412 198698
rect 359372 197056 359424 197062
rect 359372 196998 359424 197004
rect 322204 195968 322256 195974
rect 322204 195910 322256 195916
rect 359372 152040 359424 152046
rect 359372 151982 359424 151988
rect 359004 151904 359056 151910
rect 359004 151846 359056 151852
rect 359016 146266 359044 151846
rect 359384 150414 359412 151982
rect 359372 150408 359424 150414
rect 359372 150350 359424 150356
rect 359004 146260 359056 146266
rect 359004 146202 359056 146208
rect 320824 122800 320876 122806
rect 320824 122742 320876 122748
rect 359476 122738 359504 291178
rect 360212 280158 360240 340054
rect 362880 337793 362908 340068
rect 364904 337793 364932 340068
rect 362866 337784 362922 337793
rect 362866 337719 362922 337728
rect 364890 337784 364946 337793
rect 364890 337719 364946 337728
rect 366928 337414 366956 340068
rect 366916 337408 366968 337414
rect 366916 337350 366968 337356
rect 368952 335374 368980 340068
rect 368940 335368 368992 335374
rect 368940 335310 368992 335316
rect 360200 280152 360252 280158
rect 360200 280094 360252 280100
rect 369044 277250 369072 344986
rect 369124 335368 369176 335374
rect 369124 335310 369176 335316
rect 369136 282914 369164 335310
rect 369398 297392 369454 297401
rect 369398 297327 369454 297336
rect 369306 296848 369362 296857
rect 369412 296818 369440 297327
rect 369306 296783 369362 296792
rect 369400 296812 369452 296818
rect 369320 296750 369348 296783
rect 369400 296754 369452 296760
rect 369308 296744 369360 296750
rect 369308 296686 369360 296692
rect 369306 296304 369362 296313
rect 369306 296239 369362 296248
rect 369320 295866 369348 296239
rect 369308 295860 369360 295866
rect 369308 295802 369360 295808
rect 369136 282886 369256 282914
rect 369044 277234 369164 277250
rect 369044 277228 369176 277234
rect 369044 277222 369124 277228
rect 369124 277170 369176 277176
rect 369228 273254 369256 282886
rect 369308 277228 369360 277234
rect 369308 277170 369360 277176
rect 369320 277137 369348 277170
rect 369306 277128 369362 277137
rect 369306 277063 369362 277072
rect 369136 273226 369256 273254
rect 360660 271108 360712 271114
rect 360660 271050 360712 271056
rect 360672 268682 360700 271050
rect 369136 268682 369164 273226
rect 360672 268668 360962 268682
rect 368966 268668 369164 268682
rect 360672 268654 360976 268668
rect 360948 265742 360976 268654
rect 368952 268654 369164 268668
rect 362880 267889 362908 268124
rect 362866 267880 362922 267889
rect 362866 267815 362922 267824
rect 362880 266354 362908 267815
rect 362868 266348 362920 266354
rect 362868 266290 362920 266296
rect 364904 266286 364932 268124
rect 364892 266280 364944 266286
rect 364890 266248 364892 266257
rect 364944 266248 364946 266257
rect 364890 266183 364946 266192
rect 364904 266157 364932 266183
rect 366928 266150 366956 268124
rect 368952 266218 368980 268654
rect 369320 267734 369348 277063
rect 369964 273873 369992 345199
rect 370056 274961 370084 346831
rect 370226 295624 370282 295633
rect 370226 295559 370282 295568
rect 370240 295390 370268 295559
rect 370228 295384 370280 295390
rect 370228 295326 370280 295332
rect 370136 295248 370188 295254
rect 370136 295190 370188 295196
rect 370148 295089 370176 295190
rect 370134 295080 370190 295089
rect 370134 295015 370190 295024
rect 370042 274952 370098 274961
rect 370042 274887 370098 274896
rect 369950 273864 370006 273873
rect 369950 273799 370006 273808
rect 369044 267706 369348 267734
rect 368940 266212 368992 266218
rect 368940 266154 368992 266160
rect 366916 266144 366968 266150
rect 366916 266086 366968 266092
rect 360936 265736 360988 265742
rect 360936 265678 360988 265684
rect 360948 264994 360976 265678
rect 360200 264988 360252 264994
rect 360200 264930 360252 264936
rect 360936 264988 360988 264994
rect 360936 264930 360988 264936
rect 359556 224120 359608 224126
rect 359556 224062 359608 224068
rect 359568 213926 359596 224062
rect 359740 224052 359792 224058
rect 359740 223994 359792 224000
rect 359648 223984 359700 223990
rect 359648 223926 359700 223932
rect 359660 216646 359688 223926
rect 359752 219434 359780 223994
rect 359740 219428 359792 219434
rect 359740 219370 359792 219376
rect 359648 216640 359700 216646
rect 359648 216582 359700 216588
rect 360212 215294 360240 264930
rect 360212 215266 360608 215294
rect 359556 213920 359608 213926
rect 359556 213862 359608 213868
rect 359556 205692 359608 205698
rect 359556 205634 359608 205640
rect 359568 196994 359596 205634
rect 359648 202904 359700 202910
rect 359648 202846 359700 202852
rect 359660 197130 359688 202846
rect 359648 197124 359700 197130
rect 359648 197066 359700 197072
rect 359556 196988 359608 196994
rect 359556 196930 359608 196936
rect 360580 196058 360608 215266
rect 369044 205306 369072 267706
rect 369124 266212 369176 266218
rect 369124 266154 369176 266160
rect 369136 210610 369164 266154
rect 370148 260846 370176 295015
rect 370240 267034 370268 295326
rect 370332 277409 370360 349279
rect 370502 347712 370558 347721
rect 370502 347647 370558 347656
rect 370410 340232 370466 340241
rect 370410 340167 370466 340176
rect 370318 277400 370374 277409
rect 370318 277335 370374 277344
rect 370424 268297 370452 340167
rect 370516 275777 370544 347647
rect 370594 346080 370650 346089
rect 370594 346015 370650 346024
rect 370502 275768 370558 275777
rect 370502 275703 370558 275712
rect 370608 274145 370636 346015
rect 371240 298104 371292 298110
rect 371240 298046 371292 298052
rect 371252 297809 371280 298046
rect 371238 297800 371294 297809
rect 371238 297735 371294 297744
rect 371240 297424 371292 297430
rect 371240 297366 371292 297372
rect 371252 297265 371280 297366
rect 371238 297256 371294 297265
rect 371238 297191 371294 297200
rect 371238 296712 371294 296721
rect 371238 296647 371240 296656
rect 371292 296647 371294 296656
rect 371240 296618 371292 296624
rect 371238 296168 371294 296177
rect 371238 296103 371294 296112
rect 371252 295934 371280 296103
rect 371240 295928 371292 295934
rect 371240 295870 371292 295876
rect 371252 295594 371280 295870
rect 371240 295588 371292 295594
rect 371240 295530 371292 295536
rect 371240 294024 371292 294030
rect 371238 293992 371240 294001
rect 371292 293992 371294 294001
rect 371238 293927 371294 293936
rect 371238 293448 371294 293457
rect 371238 293383 371294 293392
rect 371252 293282 371280 293383
rect 371240 293276 371292 293282
rect 371240 293218 371292 293224
rect 371240 292936 371292 292942
rect 371238 292904 371240 292913
rect 371292 292904 371294 292913
rect 371238 292839 371294 292848
rect 371240 291916 371292 291922
rect 371240 291858 371292 291864
rect 371252 291825 371280 291858
rect 371238 291816 371294 291825
rect 371238 291751 371294 291760
rect 371238 291272 371294 291281
rect 371238 291207 371240 291216
rect 371292 291207 371294 291216
rect 371240 291178 371292 291184
rect 371240 290488 371292 290494
rect 371240 290430 371292 290436
rect 371252 290193 371280 290430
rect 371238 290184 371294 290193
rect 371238 290119 371294 290128
rect 371238 289096 371294 289105
rect 371238 289031 371240 289040
rect 371292 289031 371294 289040
rect 371240 289002 371292 289008
rect 371240 288380 371292 288386
rect 371240 288322 371292 288328
rect 371252 287609 371280 288322
rect 371238 287600 371294 287609
rect 371238 287535 371294 287544
rect 371344 286634 371372 351863
rect 371882 350296 371938 350305
rect 371882 350231 371938 350240
rect 371606 348256 371662 348265
rect 371606 348191 371608 348200
rect 371660 348191 371662 348200
rect 371608 348162 371660 348168
rect 371790 343904 371846 343913
rect 371790 343839 371846 343848
rect 371422 343360 371478 343369
rect 371422 343295 371478 343304
rect 371160 286606 371372 286634
rect 371160 286226 371188 286606
rect 371332 286476 371384 286482
rect 371332 286418 371384 286424
rect 371160 286198 371280 286226
rect 371252 279993 371280 286198
rect 371344 285977 371372 286418
rect 371330 285968 371386 285977
rect 371330 285903 371386 285912
rect 371238 279984 371294 279993
rect 371238 279919 371294 279928
rect 370686 275224 370742 275233
rect 370686 275159 370742 275168
rect 370594 274136 370650 274145
rect 370594 274071 370650 274080
rect 370410 268288 370466 268297
rect 370410 268223 370466 268232
rect 370424 267734 370452 268223
rect 370424 267706 370636 267734
rect 370228 267028 370280 267034
rect 370228 266970 370280 266976
rect 370136 260840 370188 260846
rect 370136 260782 370188 260788
rect 370504 247716 370556 247722
rect 370504 247658 370556 247664
rect 370516 241534 370544 247658
rect 370504 241528 370556 241534
rect 370504 241470 370556 241476
rect 370320 240780 370372 240786
rect 370320 240722 370372 240728
rect 369216 235272 369268 235278
rect 369216 235214 369268 235220
rect 369228 231742 369256 235214
rect 369216 231736 369268 231742
rect 369216 231678 369268 231684
rect 369228 229094 369256 231678
rect 369400 229764 369452 229770
rect 369400 229706 369452 229712
rect 369412 229158 369440 229706
rect 369400 229152 369452 229158
rect 369400 229094 369452 229100
rect 370332 229094 370360 240722
rect 369228 229066 369348 229094
rect 369320 220697 369348 229066
rect 369306 220688 369362 220697
rect 369306 220623 369362 220632
rect 369412 220561 369440 229094
rect 370332 229066 370452 229094
rect 370228 228404 370280 228410
rect 370228 228346 370280 228352
rect 369952 225684 370004 225690
rect 369952 225626 370004 225632
rect 369860 224392 369912 224398
rect 369860 224334 369912 224340
rect 369398 220552 369454 220561
rect 369398 220487 369454 220496
rect 369872 220153 369900 224334
rect 369858 220144 369914 220153
rect 369858 220079 369914 220088
rect 369872 219706 369900 220079
rect 369860 219700 369912 219706
rect 369860 219642 369912 219648
rect 369860 219564 369912 219570
rect 369860 219506 369912 219512
rect 369872 219434 369900 219506
rect 369860 219428 369912 219434
rect 369860 219370 369912 219376
rect 369872 219065 369900 219370
rect 369858 219056 369914 219065
rect 369858 218991 369914 219000
rect 369964 218929 369992 225626
rect 370136 225616 370188 225622
rect 370136 225558 370188 225564
rect 370044 224324 370096 224330
rect 370044 224266 370096 224272
rect 369950 218920 370006 218929
rect 369950 218855 369952 218864
rect 370004 218855 370006 218864
rect 369952 218826 370004 218832
rect 369964 218795 369992 218826
rect 370056 218754 370084 224266
rect 370044 218748 370096 218754
rect 370044 218690 370096 218696
rect 370056 218521 370084 218690
rect 370042 218512 370098 218521
rect 370042 218447 370098 218456
rect 370148 218006 370176 225558
rect 370240 219570 370268 228346
rect 370320 224256 370372 224262
rect 370320 224198 370372 224204
rect 370228 219564 370280 219570
rect 370228 219506 370280 219512
rect 370136 218000 370188 218006
rect 370136 217942 370188 217948
rect 370332 217025 370360 224198
rect 370424 221377 370452 229066
rect 370516 221921 370544 241470
rect 370502 221912 370558 221921
rect 370502 221847 370558 221856
rect 370410 221368 370466 221377
rect 370410 221303 370466 221312
rect 370424 220930 370452 221303
rect 370412 220924 370464 220930
rect 370412 220866 370464 220872
rect 370412 218000 370464 218006
rect 370412 217942 370464 217948
rect 370424 217569 370452 217942
rect 370410 217560 370466 217569
rect 370410 217495 370466 217504
rect 370318 217016 370374 217025
rect 370318 216951 370320 216960
rect 370372 216951 370374 216960
rect 370320 216922 370372 216928
rect 370226 212256 370282 212265
rect 370226 212191 370282 212200
rect 370240 211818 370268 212191
rect 370228 211812 370280 211818
rect 370228 211754 370280 211760
rect 369136 210582 369256 210610
rect 369044 205278 369164 205306
rect 369136 205222 369164 205278
rect 369124 205216 369176 205222
rect 369124 205158 369176 205164
rect 369228 202874 369256 210582
rect 370134 210080 370190 210089
rect 370134 210015 370190 210024
rect 369858 209264 369914 209273
rect 369858 209199 369914 209208
rect 369308 205216 369360 205222
rect 369306 205184 369308 205193
rect 369360 205184 369362 205193
rect 369306 205119 369362 205128
rect 369136 202846 369256 202874
rect 364522 196072 364578 196081
rect 360580 196030 360962 196058
rect 360580 180794 360608 196030
rect 362880 194585 362908 196044
rect 369136 196058 369164 202846
rect 369872 196722 369900 209199
rect 369950 203008 370006 203017
rect 369950 202943 370006 202952
rect 369860 196716 369912 196722
rect 369860 196658 369912 196664
rect 369872 196110 369900 196658
rect 364578 196044 364918 196058
rect 364578 196030 364932 196044
rect 364522 196007 364578 196016
rect 364904 194585 364932 196030
rect 362866 194576 362922 194585
rect 362866 194511 362922 194520
rect 364890 194576 364946 194585
rect 364890 194511 364946 194520
rect 366928 194478 366956 196044
rect 368966 196030 369164 196058
rect 369860 196104 369912 196110
rect 369860 196046 369912 196052
rect 366916 194472 366968 194478
rect 366916 194414 366968 194420
rect 360212 180766 360608 180794
rect 359556 151972 359608 151978
rect 359556 151914 359608 151920
rect 359568 143546 359596 151914
rect 359556 143540 359608 143546
rect 359556 143482 359608 143488
rect 360212 132494 360240 180766
rect 360212 132466 360608 132494
rect 360580 124794 360608 132466
rect 369044 124794 369072 196030
rect 369768 175160 369820 175166
rect 369768 175102 369820 175108
rect 369676 169720 369728 169726
rect 369676 169662 369728 169668
rect 369584 168360 369636 168366
rect 369584 168302 369636 168308
rect 369400 159996 369452 160002
rect 369400 159938 369452 159944
rect 369306 152960 369362 152969
rect 369228 152918 369306 152946
rect 369228 152522 369256 152918
rect 369306 152895 369362 152904
rect 369412 152810 369440 159938
rect 369492 156664 369544 156670
rect 369492 156606 369544 156612
rect 369320 152782 369440 152810
rect 369216 152516 369268 152522
rect 369216 152458 369268 152464
rect 369124 151972 369176 151978
rect 369124 151914 369176 151920
rect 369136 131458 369164 151914
rect 369228 135250 369256 152458
rect 369320 152046 369348 152782
rect 369308 152040 369360 152046
rect 369308 151982 369360 151988
rect 369216 135244 369268 135250
rect 369216 135186 369268 135192
rect 369320 132433 369348 151982
rect 369504 151910 369532 156606
rect 369596 153066 369624 168302
rect 369688 153134 369716 169662
rect 369780 153202 369808 175102
rect 369964 161474 369992 202943
rect 370148 202774 370176 210015
rect 370240 209774 370268 211754
rect 370240 209746 370360 209774
rect 370136 202768 370188 202774
rect 370136 202710 370188 202716
rect 370042 201920 370098 201929
rect 370042 201855 370098 201864
rect 370056 164218 370084 201855
rect 370148 184890 370176 202710
rect 370332 197198 370360 209746
rect 370502 208992 370558 209001
rect 370502 208927 370558 208936
rect 370320 197192 370372 197198
rect 370320 197134 370372 197140
rect 370516 195294 370544 208927
rect 370608 196217 370636 267706
rect 370700 203153 370728 275159
rect 370778 274136 370834 274145
rect 370778 274071 370834 274080
rect 370686 203144 370742 203153
rect 370686 203079 370742 203088
rect 370792 202065 370820 274071
rect 371054 273592 371110 273601
rect 371054 273527 371110 273536
rect 371068 273222 371096 273527
rect 371056 273216 371108 273222
rect 371056 273158 371108 273164
rect 371436 271697 371464 343295
rect 371514 341728 371570 341737
rect 371514 341663 371570 341672
rect 371422 271688 371478 271697
rect 371422 271623 371478 271632
rect 371528 271522 371556 341663
rect 371698 341184 371754 341193
rect 371698 341119 371754 341128
rect 371606 340640 371662 340649
rect 371606 340575 371662 340584
rect 371620 276418 371648 340575
rect 371608 276412 371660 276418
rect 371608 276354 371660 276360
rect 371606 276312 371662 276321
rect 371606 276247 371662 276256
rect 371620 276078 371648 276247
rect 371608 276072 371660 276078
rect 371608 276014 371660 276020
rect 371516 271516 371568 271522
rect 371516 271458 371568 271464
rect 371712 271402 371740 341119
rect 371804 271969 371832 343839
rect 371896 286618 371924 350231
rect 372158 349888 372214 349897
rect 372158 349823 372214 349832
rect 371974 344992 372030 345001
rect 371974 344927 372030 344936
rect 371884 286612 371936 286618
rect 371884 286554 371936 286560
rect 371882 286512 371938 286521
rect 371882 286447 371938 286456
rect 371896 286414 371924 286447
rect 371884 286408 371936 286414
rect 371884 286350 371936 286356
rect 371884 285660 371936 285666
rect 371884 285602 371936 285608
rect 371896 285433 371924 285602
rect 371882 285424 371938 285433
rect 371882 285359 371938 285368
rect 371884 285116 371936 285122
rect 371884 285058 371936 285064
rect 371896 284889 371924 285058
rect 371882 284880 371938 284889
rect 371882 284815 371938 284824
rect 371884 284368 371936 284374
rect 371882 284336 371884 284345
rect 371936 284336 371938 284345
rect 371882 284271 371938 284280
rect 371882 283792 371938 283801
rect 371882 283727 371938 283736
rect 371896 283626 371924 283727
rect 371884 283620 371936 283626
rect 371884 283562 371936 283568
rect 371882 283248 371938 283257
rect 371882 283183 371884 283192
rect 371936 283183 371938 283192
rect 371884 283154 371936 283160
rect 371884 282736 371936 282742
rect 371882 282704 371884 282713
rect 371936 282704 371938 282713
rect 371882 282639 371938 282648
rect 371884 282192 371936 282198
rect 371882 282160 371884 282169
rect 371936 282160 371938 282169
rect 371882 282095 371938 282104
rect 371988 273057 372016 344927
rect 372066 342816 372122 342825
rect 372066 342751 372122 342760
rect 371974 273048 372030 273057
rect 371974 272983 372030 272992
rect 371790 271960 371846 271969
rect 371790 271895 371846 271904
rect 371252 271374 371740 271402
rect 371252 269249 371280 271374
rect 371804 271266 371832 271895
rect 371882 271688 371938 271697
rect 371882 271623 371938 271632
rect 371344 271238 371832 271266
rect 371238 269240 371294 269249
rect 371238 269175 371294 269184
rect 370872 256760 370924 256766
rect 370872 256702 370924 256708
rect 370884 223582 370912 256702
rect 370872 223576 370924 223582
rect 370872 223518 370924 223524
rect 370962 211712 371018 211721
rect 370962 211647 371018 211656
rect 370870 208448 370926 208457
rect 370870 208383 370926 208392
rect 370778 202056 370834 202065
rect 370778 201991 370834 202000
rect 370594 196208 370650 196217
rect 370594 196143 370650 196152
rect 370778 196208 370834 196217
rect 370778 196143 370834 196152
rect 370504 195288 370556 195294
rect 370502 195256 370504 195265
rect 370556 195256 370558 195265
rect 370502 195191 370558 195200
rect 370516 195165 370544 195191
rect 370136 184884 370188 184890
rect 370136 184826 370188 184832
rect 370136 172508 370188 172514
rect 370136 172450 370188 172456
rect 370148 171154 370176 172450
rect 370136 171148 370188 171154
rect 370136 171090 370188 171096
rect 370044 164212 370096 164218
rect 370044 164154 370096 164160
rect 369872 161446 369992 161474
rect 369872 160070 369900 161446
rect 369860 160064 369912 160070
rect 369860 160006 369912 160012
rect 369768 153196 369820 153202
rect 369768 153138 369820 153144
rect 369676 153128 369728 153134
rect 369676 153070 369728 153076
rect 369584 153060 369636 153066
rect 369584 153002 369636 153008
rect 369596 152522 369624 153002
rect 369688 152794 369716 153070
rect 369676 152788 369728 152794
rect 369676 152730 369728 152736
rect 369584 152516 369636 152522
rect 369584 152458 369636 152464
rect 369492 151904 369544 151910
rect 369492 151846 369544 151852
rect 369400 135244 369452 135250
rect 369400 135186 369452 135192
rect 369412 135153 369440 135186
rect 369398 135144 369454 135153
rect 369398 135079 369454 135088
rect 369306 132424 369362 132433
rect 369306 132359 369362 132368
rect 369504 132025 369532 151846
rect 369780 151814 369808 153138
rect 369872 151978 369900 160006
rect 370044 154556 370096 154562
rect 370044 154498 370096 154504
rect 369952 152788 370004 152794
rect 369952 152730 370004 152736
rect 369860 151972 369912 151978
rect 369860 151914 369912 151920
rect 369780 151786 369900 151814
rect 369872 134609 369900 151786
rect 369858 134600 369914 134609
rect 369858 134535 369914 134544
rect 369964 133657 369992 152730
rect 370056 134065 370084 154498
rect 370148 153882 370176 171090
rect 370504 164212 370556 164218
rect 370504 164154 370556 164160
rect 370596 164212 370648 164218
rect 370596 164154 370648 164160
rect 370228 162716 370280 162722
rect 370228 162658 370280 162664
rect 370240 162178 370268 162658
rect 370228 162172 370280 162178
rect 370228 162114 370280 162120
rect 370136 153876 370188 153882
rect 370136 153818 370188 153824
rect 370148 135969 370176 153818
rect 370134 135960 370190 135969
rect 370134 135895 370190 135904
rect 370240 135425 370268 162114
rect 370320 152516 370372 152522
rect 370320 152458 370372 152464
rect 370226 135416 370282 135425
rect 370226 135351 370282 135360
rect 370042 134056 370098 134065
rect 370042 133991 370098 134000
rect 369950 133648 370006 133657
rect 369950 133583 370006 133592
rect 370332 132841 370360 152458
rect 370318 132832 370374 132841
rect 370318 132767 370374 132776
rect 369490 132016 369546 132025
rect 369490 131951 369546 131960
rect 369306 131472 369362 131481
rect 369136 131430 369306 131458
rect 369306 131407 369362 131416
rect 370240 130694 370268 130725
rect 370228 130688 370280 130694
rect 370226 130656 370228 130665
rect 370280 130656 370282 130665
rect 370226 130591 370282 130600
rect 369950 129840 370006 129849
rect 369950 129775 370006 129784
rect 369858 129160 369914 129169
rect 369858 129095 369860 129104
rect 369912 129095 369914 129104
rect 369860 129066 369912 129072
rect 369872 125186 369900 129066
rect 369860 125180 369912 125186
rect 369860 125122 369912 125128
rect 369964 125050 369992 129775
rect 370042 128616 370098 128625
rect 370042 128551 370098 128560
rect 369952 125044 370004 125050
rect 369952 124986 370004 124992
rect 370056 124982 370084 128551
rect 370134 127392 370190 127401
rect 370134 127327 370190 127336
rect 370044 124976 370096 124982
rect 370044 124918 370096 124924
rect 360580 124766 360962 124794
rect 368966 124766 369072 124794
rect 369950 124808 370006 124817
rect 369950 124743 370006 124752
rect 369858 124400 369914 124409
rect 369858 124335 369914 124344
rect 362788 124086 362894 124114
rect 364918 124086 365208 124114
rect 362788 124001 362816 124086
rect 365180 124001 365208 124086
rect 362774 123992 362830 124001
rect 362774 123927 362830 123936
rect 365166 123992 365222 124001
rect 365166 123927 365222 123936
rect 366928 122738 366956 124100
rect 359464 122732 359516 122738
rect 359464 122674 359516 122680
rect 366916 122732 366968 122738
rect 366916 122674 366968 122680
rect 313924 113144 313976 113150
rect 313924 113086 313976 113092
rect 369872 102134 369900 124335
rect 369964 123486 369992 124743
rect 369952 123480 370004 123486
rect 369952 123422 370004 123428
rect 370148 121446 370176 127327
rect 370240 125118 370268 130591
rect 370516 130121 370544 164154
rect 370608 154562 370636 164154
rect 370596 154556 370648 154562
rect 370596 154498 370648 154504
rect 370502 130112 370558 130121
rect 370502 130047 370558 130056
rect 370332 129062 370360 129093
rect 370320 129056 370372 129062
rect 370318 129024 370320 129033
rect 370372 129024 370374 129033
rect 370318 128959 370374 128968
rect 370332 125254 370360 128959
rect 370410 126304 370466 126313
rect 370410 126239 370466 126248
rect 370424 125934 370452 126239
rect 370412 125928 370464 125934
rect 370412 125870 370464 125876
rect 370320 125248 370372 125254
rect 370320 125190 370372 125196
rect 370228 125112 370280 125118
rect 370228 125054 370280 125060
rect 370424 123622 370452 125870
rect 370594 125760 370650 125769
rect 370594 125695 370650 125704
rect 370504 125520 370556 125526
rect 370504 125462 370556 125468
rect 370516 124817 370544 125462
rect 370502 124808 370558 124817
rect 370502 124743 370558 124752
rect 370412 123616 370464 123622
rect 370412 123558 370464 123564
rect 370136 121440 370188 121446
rect 370136 121382 370188 121388
rect 370608 111790 370636 125695
rect 370792 124914 370820 196143
rect 370884 190454 370912 208383
rect 370976 194546 371004 211647
rect 371252 197146 371280 269175
rect 371344 199889 371372 271238
rect 371516 271176 371568 271182
rect 371516 271118 371568 271124
rect 371792 271176 371844 271182
rect 371792 271118 371844 271124
rect 371528 269793 371556 271118
rect 371606 270328 371662 270337
rect 371606 270263 371662 270272
rect 371514 269784 371570 269793
rect 371514 269719 371570 269728
rect 371620 258074 371648 270263
rect 371528 258046 371648 258074
rect 371424 223576 371476 223582
rect 371424 223518 371476 223524
rect 371436 222465 371464 223518
rect 371422 222456 371478 222465
rect 371422 222391 371478 222400
rect 371422 213888 371478 213897
rect 371422 213823 371478 213832
rect 371436 213110 371464 213823
rect 371424 213104 371476 213110
rect 371424 213046 371476 213052
rect 371424 211880 371476 211886
rect 371424 211822 371476 211828
rect 371436 211721 371464 211822
rect 371422 211712 371478 211721
rect 371422 211647 371478 211656
rect 371422 205320 371478 205329
rect 371422 205255 371478 205264
rect 371436 204105 371464 205255
rect 371422 204096 371478 204105
rect 371422 204031 371478 204040
rect 371422 201376 371478 201385
rect 371422 201311 371478 201320
rect 371330 199880 371386 199889
rect 371330 199815 371386 199824
rect 371344 198937 371372 199815
rect 371330 198928 371386 198937
rect 371330 198863 371386 198872
rect 371330 197160 371386 197169
rect 371252 197118 371330 197146
rect 371330 197095 371386 197104
rect 371148 196104 371200 196110
rect 371146 196072 371148 196081
rect 371200 196072 371202 196081
rect 371146 196007 371202 196016
rect 370964 194540 371016 194546
rect 370964 194482 371016 194488
rect 370884 190426 371188 190454
rect 371160 185586 371188 190426
rect 371238 185600 371294 185609
rect 371160 185558 371238 185586
rect 371160 180794 371188 185558
rect 371238 185535 371294 185544
rect 370884 180766 371188 180794
rect 370884 175681 370912 180766
rect 370870 175672 370926 175681
rect 370870 175607 370926 175616
rect 370884 175234 370912 175607
rect 370872 175228 370924 175234
rect 370872 175170 370924 175176
rect 371146 162752 371202 162761
rect 371146 162687 371148 162696
rect 371200 162687 371202 162696
rect 371148 162658 371200 162664
rect 371240 147552 371292 147558
rect 371240 147494 371292 147500
rect 371252 147257 371280 147494
rect 371238 147248 371294 147257
rect 371238 147183 371294 147192
rect 371240 146736 371292 146742
rect 371238 146704 371240 146713
rect 371292 146704 371294 146713
rect 371238 146639 371294 146648
rect 371240 143540 371292 143546
rect 371240 143482 371292 143488
rect 371252 142497 371280 143482
rect 371238 142488 371294 142497
rect 371238 142423 371294 142432
rect 371240 142044 371292 142050
rect 371240 141986 371292 141992
rect 371252 140865 371280 141986
rect 371238 140856 371294 140865
rect 371238 140791 371294 140800
rect 371238 127936 371294 127945
rect 371238 127871 371294 127880
rect 370780 124908 370832 124914
rect 370780 124850 370832 124856
rect 370792 124273 370820 124850
rect 370778 124264 370834 124273
rect 370778 124199 370834 124208
rect 371252 124166 371280 127871
rect 371344 125322 371372 197095
rect 371436 129062 371464 201311
rect 371528 200114 371556 258046
rect 371606 225720 371662 225729
rect 371606 225655 371662 225664
rect 371620 225622 371648 225655
rect 371608 225616 371660 225622
rect 371608 225558 371660 225564
rect 371606 225176 371662 225185
rect 371606 225111 371662 225120
rect 371620 225010 371648 225111
rect 371608 225004 371660 225010
rect 371608 224946 371660 224952
rect 371606 224632 371662 224641
rect 371606 224567 371662 224576
rect 371620 223786 371648 224567
rect 371608 223780 371660 223786
rect 371608 223722 371660 223728
rect 371606 223544 371662 223553
rect 371606 223479 371608 223488
rect 371660 223479 371662 223488
rect 371608 223450 371660 223456
rect 371606 223000 371662 223009
rect 371606 222935 371662 222944
rect 371620 222698 371648 222935
rect 371608 222692 371660 222698
rect 371608 222634 371660 222640
rect 371608 216572 371660 216578
rect 371608 216514 371660 216520
rect 371620 216073 371648 216514
rect 371606 216064 371662 216073
rect 371606 215999 371662 216008
rect 371606 215520 371662 215529
rect 371606 215455 371662 215464
rect 371620 215354 371648 215455
rect 371608 215348 371660 215354
rect 371608 215290 371660 215296
rect 371698 214976 371754 214985
rect 371698 214911 371754 214920
rect 371608 214668 371660 214674
rect 371608 214610 371660 214616
rect 371620 214441 371648 214610
rect 371712 214606 371740 214911
rect 371700 214600 371752 214606
rect 371700 214542 371752 214548
rect 371606 214432 371662 214441
rect 371606 214367 371662 214376
rect 371606 213344 371662 213353
rect 371606 213279 371662 213288
rect 371700 213308 371752 213314
rect 371620 213246 371648 213279
rect 371700 213250 371752 213256
rect 371608 213240 371660 213246
rect 371608 213182 371660 213188
rect 371712 212809 371740 213250
rect 371698 212800 371754 212809
rect 371698 212735 371754 212744
rect 371698 207904 371754 207913
rect 371698 207839 371754 207848
rect 371608 206304 371660 206310
rect 371606 206272 371608 206281
rect 371660 206272 371662 206281
rect 371606 206207 371662 206216
rect 371712 206122 371740 207839
rect 371620 206094 371740 206122
rect 371620 203538 371648 206094
rect 371698 205864 371754 205873
rect 371698 205799 371700 205808
rect 371752 205799 371754 205808
rect 371700 205770 371752 205776
rect 371620 203510 371740 203538
rect 371608 201612 371660 201618
rect 371608 201554 371660 201560
rect 371620 201521 371648 201554
rect 371606 201512 371662 201521
rect 371606 201447 371662 201456
rect 371528 200086 371648 200114
rect 371620 198257 371648 200086
rect 371606 198248 371662 198257
rect 371606 198183 371662 198192
rect 371516 153196 371568 153202
rect 371516 153138 371568 153144
rect 371528 152697 371556 153138
rect 371514 152688 371570 152697
rect 371514 152623 371570 152632
rect 371516 151700 371568 151706
rect 371516 151642 371568 151648
rect 371528 150521 371556 151642
rect 371514 150512 371570 150521
rect 371514 150447 371570 150456
rect 371516 150340 371568 150346
rect 371516 150282 371568 150288
rect 371528 149433 371556 150282
rect 371514 149424 371570 149433
rect 371514 149359 371570 149368
rect 371516 146192 371568 146198
rect 371516 146134 371568 146140
rect 371528 145625 371556 146134
rect 371514 145616 371570 145625
rect 371514 145551 371570 145560
rect 371516 144900 371568 144906
rect 371516 144842 371568 144848
rect 371528 144129 371556 144842
rect 371514 144120 371570 144129
rect 371514 144055 371570 144064
rect 371516 142112 371568 142118
rect 371516 142054 371568 142060
rect 371528 141409 371556 142054
rect 371514 141400 371570 141409
rect 371514 141335 371570 141344
rect 371516 139392 371568 139398
rect 371516 139334 371568 139340
rect 371528 138145 371556 139334
rect 371514 138136 371570 138145
rect 371514 138071 371570 138080
rect 371424 129056 371476 129062
rect 371424 128998 371476 129004
rect 371620 125934 371648 198183
rect 371712 172514 371740 203510
rect 371804 201385 371832 271118
rect 371790 201376 371846 201385
rect 371790 201311 371846 201320
rect 371896 199345 371924 271623
rect 371988 271182 372016 272983
rect 371976 271176 372028 271182
rect 371976 271118 372028 271124
rect 372080 270881 372108 342751
rect 372172 278730 372200 349823
rect 372250 344448 372306 344457
rect 372250 344383 372306 344392
rect 372160 278724 372212 278730
rect 372160 278666 372212 278672
rect 372172 277953 372200 278666
rect 372158 277944 372214 277953
rect 372158 277879 372214 277888
rect 372160 276412 372212 276418
rect 372160 276354 372212 276360
rect 372066 270872 372122 270881
rect 372066 270807 372122 270816
rect 372080 258074 372108 270807
rect 372172 268705 372200 276354
rect 372264 272513 372292 344383
rect 372434 342272 372490 342281
rect 372434 342207 372490 342216
rect 372344 294636 372396 294642
rect 372344 294578 372396 294584
rect 372356 294545 372384 294578
rect 372342 294536 372398 294545
rect 372342 294471 372398 294480
rect 372342 292360 372398 292369
rect 372342 292295 372398 292304
rect 372356 291854 372384 292295
rect 372344 291848 372396 291854
rect 372344 291790 372396 291796
rect 372342 290728 372398 290737
rect 372342 290663 372398 290672
rect 372356 290562 372384 290663
rect 372344 290556 372396 290562
rect 372344 290498 372396 290504
rect 372342 289640 372398 289649
rect 372342 289575 372398 289584
rect 372356 288998 372384 289575
rect 372344 288992 372396 288998
rect 372344 288934 372396 288940
rect 372342 288144 372398 288153
rect 372342 288079 372398 288088
rect 372356 287094 372384 288079
rect 372344 287088 372396 287094
rect 372344 287030 372396 287036
rect 372344 286612 372396 286618
rect 372344 286554 372396 286560
rect 372356 278361 372384 286554
rect 372342 278352 372398 278361
rect 372342 278287 372398 278296
rect 372356 277506 372384 278287
rect 372344 277500 372396 277506
rect 372344 277442 372396 277448
rect 372250 272504 372306 272513
rect 372250 272439 372306 272448
rect 372158 268696 372214 268705
rect 372158 268631 372214 268640
rect 372172 268394 372200 268631
rect 372160 268388 372212 268394
rect 372160 268330 372212 268336
rect 372264 258074 372292 272439
rect 372448 270337 372476 342207
rect 372632 294642 372660 366438
rect 372802 362672 372858 362681
rect 372802 362607 372858 362616
rect 372710 346624 372766 346633
rect 372710 346559 372766 346568
rect 372620 294636 372672 294642
rect 372620 294578 372672 294584
rect 372526 287056 372582 287065
rect 372526 286991 372582 287000
rect 372540 286346 372568 286991
rect 372528 286340 372580 286346
rect 372528 286282 372580 286288
rect 372526 279984 372582 279993
rect 372526 279919 372582 279928
rect 372434 270328 372490 270337
rect 372434 270263 372490 270272
rect 372342 269784 372398 269793
rect 372342 269719 372398 269728
rect 371988 258046 372108 258074
rect 372172 258046 372292 258074
rect 371882 199336 371938 199345
rect 371882 199271 371938 199280
rect 371790 198792 371846 198801
rect 371790 198727 371846 198736
rect 371700 172508 371752 172514
rect 371700 172450 371752 172456
rect 371700 154556 371752 154562
rect 371700 154498 371752 154504
rect 371712 153785 371740 154498
rect 371698 153776 371754 153785
rect 371698 153711 371754 153720
rect 371700 153400 371752 153406
rect 371700 153342 371752 153348
rect 371712 153241 371740 153342
rect 371698 153232 371754 153241
rect 371698 153167 371754 153176
rect 371700 153128 371752 153134
rect 371700 153070 371752 153076
rect 371712 152153 371740 153070
rect 371698 152144 371754 152153
rect 371698 152079 371754 152088
rect 371700 151768 371752 151774
rect 371700 151710 371752 151716
rect 371712 151609 371740 151710
rect 371698 151600 371754 151609
rect 371698 151535 371754 151544
rect 371700 151088 371752 151094
rect 371698 151056 371700 151065
rect 371752 151056 371754 151065
rect 371698 150991 371754 151000
rect 371700 150408 371752 150414
rect 371700 150350 371752 150356
rect 371712 149977 371740 150350
rect 371698 149968 371754 149977
rect 371698 149903 371754 149912
rect 371700 149048 371752 149054
rect 371700 148990 371752 148996
rect 371712 148889 371740 148990
rect 371698 148880 371754 148889
rect 371698 148815 371754 148824
rect 371700 148436 371752 148442
rect 371700 148378 371752 148384
rect 371712 148345 371740 148378
rect 371698 148336 371754 148345
rect 371698 148271 371754 148280
rect 371700 148232 371752 148238
rect 371700 148174 371752 148180
rect 371712 147801 371740 148174
rect 371698 147792 371754 147801
rect 371698 147727 371754 147736
rect 371698 146160 371754 146169
rect 371698 146095 371700 146104
rect 371752 146095 371754 146104
rect 371700 146066 371752 146072
rect 371700 145104 371752 145110
rect 371698 145072 371700 145081
rect 371752 145072 371754 145081
rect 371698 145007 371754 145016
rect 371700 144560 371752 144566
rect 371698 144528 371700 144537
rect 371752 144528 371754 144537
rect 371698 144463 371754 144472
rect 371700 143472 371752 143478
rect 371700 143414 371752 143420
rect 371712 143041 371740 143414
rect 371698 143032 371754 143041
rect 371698 142967 371754 142976
rect 371700 141976 371752 141982
rect 371698 141944 371700 141953
rect 371752 141944 371754 141953
rect 371698 141879 371754 141888
rect 371700 140684 371752 140690
rect 371700 140626 371752 140632
rect 371712 140321 371740 140626
rect 371698 140312 371754 140321
rect 371698 140247 371754 140256
rect 371700 139256 371752 139262
rect 371698 139224 371700 139233
rect 371752 139224 371754 139233
rect 371698 139159 371754 139168
rect 371700 138916 371752 138922
rect 371700 138858 371752 138864
rect 371712 138689 371740 138858
rect 371698 138680 371754 138689
rect 371698 138615 371754 138624
rect 371804 126857 371832 198727
rect 371896 158030 371924 199271
rect 371988 198801 372016 258046
rect 372066 216472 372122 216481
rect 372066 216407 372068 216416
rect 372120 216407 372122 216416
rect 372068 216378 372120 216384
rect 372068 204264 372120 204270
rect 372066 204232 372068 204241
rect 372120 204232 372122 204241
rect 372066 204167 372122 204176
rect 372066 203688 372122 203697
rect 372066 203623 372122 203632
rect 372080 201521 372108 203623
rect 372066 201512 372122 201521
rect 372066 201447 372122 201456
rect 372172 200433 372200 258046
rect 372252 224256 372304 224262
rect 372252 224198 372304 224204
rect 372264 224097 372292 224198
rect 372250 224088 372306 224097
rect 372250 224023 372306 224032
rect 372356 209774 372384 269719
rect 372356 209746 372476 209774
rect 372158 200424 372214 200433
rect 372158 200359 372214 200368
rect 372172 200114 372200 200359
rect 372080 200086 372200 200114
rect 371974 198792 372030 198801
rect 371974 198727 372030 198736
rect 372080 162246 372108 200086
rect 372158 198928 372214 198937
rect 372158 198863 372214 198872
rect 372068 162240 372120 162246
rect 372068 162182 372120 162188
rect 372080 161474 372108 162182
rect 371988 161446 372108 161474
rect 371884 158024 371936 158030
rect 371884 157966 371936 157972
rect 371896 127401 371924 157966
rect 371988 128625 372016 161446
rect 372172 155242 372200 198863
rect 372448 197713 372476 209746
rect 372540 207913 372568 279919
rect 372724 277394 372752 346559
rect 372816 290562 372844 362607
rect 372896 355020 372948 355026
rect 372896 354962 372948 354968
rect 372804 290556 372856 290562
rect 372804 290498 372856 290504
rect 372816 288590 372844 288621
rect 372804 288584 372856 288590
rect 372802 288552 372804 288561
rect 372856 288552 372858 288561
rect 372802 288487 372858 288496
rect 372632 277366 372752 277394
rect 372632 274689 372660 277366
rect 372618 274680 372674 274689
rect 372618 274615 372674 274624
rect 372526 207904 372582 207913
rect 372526 207839 372582 207848
rect 372526 202600 372582 202609
rect 372632 202586 372660 274615
rect 372712 225072 372764 225078
rect 372710 225040 372712 225049
rect 372764 225040 372766 225049
rect 372710 224975 372766 224984
rect 372710 223952 372766 223961
rect 372710 223887 372712 223896
rect 372764 223887 372766 223896
rect 372712 223858 372764 223864
rect 372816 223854 372844 288487
rect 372908 283218 372936 354962
rect 374012 295594 374040 367474
rect 375380 365832 375432 365838
rect 375380 365774 375432 365780
rect 374460 364744 374512 364750
rect 374460 364686 374512 364692
rect 374276 360392 374328 360398
rect 374276 360334 374328 360340
rect 374184 354204 374236 354210
rect 374184 354146 374236 354152
rect 374092 353320 374144 353326
rect 374092 353262 374144 353268
rect 373356 295588 373408 295594
rect 373356 295530 373408 295536
rect 374000 295588 374052 295594
rect 374000 295530 374052 295536
rect 373264 291848 373316 291854
rect 373264 291790 373316 291796
rect 372896 283212 372948 283218
rect 372896 283154 372948 283160
rect 372988 278724 373040 278730
rect 372988 278666 373040 278672
rect 372896 268388 372948 268394
rect 372896 268330 372948 268336
rect 372804 223848 372856 223854
rect 372804 223790 372856 223796
rect 372816 216442 372844 223790
rect 372804 216436 372856 216442
rect 372804 216378 372856 216384
rect 372582 202570 372660 202586
rect 372582 202564 372672 202570
rect 372582 202558 372620 202564
rect 372526 202535 372582 202544
rect 372620 202506 372672 202512
rect 372908 200114 372936 268330
rect 373000 205834 373028 278666
rect 373276 229158 373304 291790
rect 373264 229152 373316 229158
rect 373264 229094 373316 229100
rect 373276 219502 373304 229094
rect 373368 224262 373396 295530
rect 374104 282198 374132 353262
rect 374196 282742 374224 354146
rect 374288 289066 374316 360334
rect 374368 348220 374420 348226
rect 374368 348162 374420 348168
rect 374276 289060 374328 289066
rect 374276 289002 374328 289008
rect 374184 282736 374236 282742
rect 374184 282678 374236 282684
rect 374092 282192 374144 282198
rect 374092 282134 374144 282140
rect 374276 282192 374328 282198
rect 374276 282134 374328 282140
rect 374184 277500 374236 277506
rect 374184 277442 374236 277448
rect 374000 276072 374052 276078
rect 374000 276014 374052 276020
rect 373356 224256 373408 224262
rect 373356 224198 373408 224204
rect 373264 219496 373316 219502
rect 373264 219438 373316 219444
rect 373356 218884 373408 218890
rect 373356 218826 373408 218832
rect 373172 212016 373224 212022
rect 373172 211958 373224 211964
rect 373184 211177 373212 211958
rect 373170 211168 373226 211177
rect 373170 211103 373226 211112
rect 373092 210662 373120 210693
rect 373080 210656 373132 210662
rect 373078 210624 373080 210633
rect 373132 210624 373134 210633
rect 373078 210559 373134 210568
rect 372988 205828 373040 205834
rect 372988 205770 373040 205776
rect 372632 200086 372936 200114
rect 372434 197704 372490 197713
rect 372434 197639 372490 197648
rect 372160 155236 372212 155242
rect 372160 155178 372212 155184
rect 372068 144832 372120 144838
rect 372068 144774 372120 144780
rect 372080 143585 372108 144774
rect 372066 143576 372122 143585
rect 372066 143511 372122 143520
rect 372172 142154 372200 155178
rect 372080 142126 372200 142154
rect 371974 128616 372030 128625
rect 371974 128551 372030 128560
rect 372080 127945 372108 142126
rect 372066 127936 372122 127945
rect 372066 127871 372122 127880
rect 371882 127392 371938 127401
rect 371882 127327 371938 127336
rect 371790 126848 371846 126857
rect 371790 126783 371846 126792
rect 371804 126002 371832 126783
rect 372448 126070 372476 197639
rect 372526 196616 372582 196625
rect 372632 196602 372660 200086
rect 372582 196574 372660 196602
rect 372526 196551 372582 196560
rect 372436 126064 372488 126070
rect 372436 126006 372488 126012
rect 371792 125996 371844 126002
rect 371792 125938 371844 125944
rect 371608 125928 371660 125934
rect 371608 125870 371660 125876
rect 371332 125316 371384 125322
rect 371332 125258 371384 125264
rect 371344 125225 371372 125258
rect 371330 125216 371386 125225
rect 371330 125151 371386 125160
rect 371240 124160 371292 124166
rect 371240 124102 371292 124108
rect 370596 111784 370648 111790
rect 370596 111726 370648 111732
rect 371344 109002 371372 125151
rect 371804 118658 371832 125938
rect 372448 125769 372476 126006
rect 372434 125760 372490 125769
rect 372434 125695 372490 125704
rect 372632 125526 372660 196574
rect 372712 194540 372764 194546
rect 372712 194482 372764 194488
rect 372724 139777 372752 194482
rect 373000 164218 373028 205770
rect 373092 193254 373120 210559
rect 373184 202706 373212 211103
rect 373172 202700 373224 202706
rect 373172 202642 373224 202648
rect 373264 202564 373316 202570
rect 373264 202506 373316 202512
rect 373080 193248 373132 193254
rect 373080 193190 373132 193196
rect 372988 164212 373040 164218
rect 372988 164154 373040 164160
rect 373276 162178 373304 202506
rect 373264 162172 373316 162178
rect 373264 162114 373316 162120
rect 372710 139768 372766 139777
rect 372710 139703 372766 139712
rect 373276 130694 373304 162114
rect 373368 146742 373396 218826
rect 373816 205624 373868 205630
rect 373816 205566 373868 205572
rect 373828 175166 373856 205566
rect 374012 204270 374040 276014
rect 374196 206310 374224 277442
rect 374184 206304 374236 206310
rect 374184 206246 374236 206252
rect 374196 205630 374224 206246
rect 374184 205624 374236 205630
rect 374184 205566 374236 205572
rect 374000 204264 374052 204270
rect 374000 204206 374052 204212
rect 374012 202874 374040 204206
rect 373920 202846 374040 202874
rect 373816 175160 373868 175166
rect 373816 175102 373868 175108
rect 373920 160002 373948 202846
rect 374288 202774 374316 282134
rect 374380 276078 374408 348162
rect 374472 292942 374500 364686
rect 375392 294030 375420 365774
rect 375748 363724 375800 363730
rect 375748 363666 375800 363672
rect 375564 360460 375616 360466
rect 375564 360402 375616 360408
rect 375472 360256 375524 360262
rect 375472 360198 375524 360204
rect 375380 294024 375432 294030
rect 375380 293966 375432 293972
rect 374460 292936 374512 292942
rect 374460 292878 374512 292884
rect 374920 292936 374972 292942
rect 374920 292878 374972 292884
rect 374736 288992 374788 288998
rect 374736 288934 374788 288940
rect 374644 285116 374696 285122
rect 374644 285058 374696 285064
rect 374552 282736 374604 282742
rect 374552 282678 374604 282684
rect 374368 276072 374420 276078
rect 374368 276014 374420 276020
rect 374368 273216 374420 273222
rect 374368 273158 374420 273164
rect 374276 202768 374328 202774
rect 374276 202710 374328 202716
rect 374380 201618 374408 273158
rect 374460 225004 374512 225010
rect 374460 224946 374512 224952
rect 374000 201612 374052 201618
rect 374000 201554 374052 201560
rect 374368 201612 374420 201618
rect 374368 201554 374420 201560
rect 373908 159996 373960 160002
rect 373908 159938 373960 159944
rect 373356 146736 373408 146742
rect 373356 146678 373408 146684
rect 373264 130688 373316 130694
rect 373264 130630 373316 130636
rect 374012 129130 374040 201554
rect 374092 193248 374144 193254
rect 374092 193190 374144 193196
rect 374104 187678 374132 193190
rect 374092 187672 374144 187678
rect 374092 187614 374144 187620
rect 374104 138922 374132 187614
rect 374276 184884 374328 184890
rect 374276 184826 374328 184832
rect 374288 139398 374316 184826
rect 374472 153406 374500 224946
rect 374564 210662 374592 282678
rect 374656 213314 374684 285058
rect 374748 218006 374776 288934
rect 374932 231742 374960 292878
rect 375392 241534 375420 293966
rect 375484 288998 375512 360198
rect 375472 288992 375524 288998
rect 375472 288934 375524 288940
rect 375576 288590 375604 360402
rect 375656 357740 375708 357746
rect 375656 357682 375708 357688
rect 375564 288584 375616 288590
rect 375564 288526 375616 288532
rect 375668 286482 375696 357682
rect 375760 291922 375788 363666
rect 376772 296682 376800 368562
rect 381084 368552 381136 368558
rect 381084 368494 381136 368500
rect 380992 367124 381044 367130
rect 380992 367066 381044 367072
rect 378232 365900 378284 365906
rect 378232 365842 378284 365848
rect 377036 363044 377088 363050
rect 377036 362986 377088 362992
rect 376852 361616 376904 361622
rect 376852 361558 376904 361564
rect 376760 296676 376812 296682
rect 376760 296618 376812 296624
rect 376772 295458 376800 296618
rect 376760 295452 376812 295458
rect 376760 295394 376812 295400
rect 375748 291916 375800 291922
rect 375748 291858 375800 291864
rect 376024 291236 376076 291242
rect 376024 291178 376076 291184
rect 375748 289060 375800 289066
rect 375748 289002 375800 289008
rect 375656 286476 375708 286482
rect 375656 286418 375708 286424
rect 375668 285734 375696 286418
rect 375656 285728 375708 285734
rect 375656 285670 375708 285676
rect 375472 283212 375524 283218
rect 375472 283154 375524 283160
rect 375380 241528 375432 241534
rect 375380 241470 375432 241476
rect 374920 231736 374972 231742
rect 374920 231678 374972 231684
rect 374932 220794 374960 231678
rect 375392 222154 375420 241470
rect 375380 222148 375432 222154
rect 375380 222090 375432 222096
rect 374920 220788 374972 220794
rect 374920 220730 374972 220736
rect 374828 219496 374880 219502
rect 374828 219438 374880 219444
rect 374736 218000 374788 218006
rect 374736 217942 374788 217948
rect 374644 213308 374696 213314
rect 374644 213250 374696 213256
rect 374552 210656 374604 210662
rect 374552 210598 374604 210604
rect 374642 204776 374698 204785
rect 374642 204711 374698 204720
rect 374550 201512 374606 201521
rect 374550 201447 374606 201456
rect 374564 156670 374592 201447
rect 374656 168366 374684 204711
rect 374734 204096 374790 204105
rect 374734 204031 374790 204040
rect 374748 169726 374776 204031
rect 374736 169720 374788 169726
rect 374736 169662 374788 169668
rect 374644 168360 374696 168366
rect 374644 168302 374696 168308
rect 374552 156664 374604 156670
rect 374552 156606 374604 156612
rect 374460 153400 374512 153406
rect 374460 153342 374512 153348
rect 374840 148442 374868 219438
rect 374920 216980 374972 216986
rect 374920 216922 374972 216928
rect 374828 148436 374880 148442
rect 374828 148378 374880 148384
rect 374932 145110 374960 216922
rect 375484 212022 375512 283154
rect 375564 222692 375616 222698
rect 375564 222634 375616 222640
rect 375472 212016 375524 212022
rect 375472 211958 375524 211964
rect 375380 202700 375432 202706
rect 375380 202642 375432 202648
rect 375392 196654 375420 202642
rect 375380 196648 375432 196654
rect 375380 196590 375432 196596
rect 374920 145104 374972 145110
rect 374920 145046 374972 145052
rect 374276 139392 374328 139398
rect 374276 139334 374328 139340
rect 375392 139262 375420 196590
rect 375576 151094 375604 222634
rect 375656 220720 375708 220726
rect 375656 220662 375708 220668
rect 375668 219706 375696 220662
rect 375656 219700 375708 219706
rect 375656 219642 375708 219648
rect 375564 151088 375616 151094
rect 375564 151030 375616 151036
rect 375668 148238 375696 219642
rect 375760 216986 375788 289002
rect 376036 219434 376064 291178
rect 376760 290556 376812 290562
rect 376760 290498 376812 290504
rect 376116 286408 376168 286414
rect 376116 286350 376168 286356
rect 376024 219428 376076 219434
rect 376024 219370 376076 219376
rect 376036 218074 376064 219370
rect 376024 218068 376076 218074
rect 376024 218010 376076 218016
rect 375748 216980 375800 216986
rect 375748 216922 375800 216928
rect 375840 216436 375892 216442
rect 375840 216378 375892 216384
rect 375748 213104 375800 213110
rect 375748 213046 375800 213052
rect 375760 196994 375788 213046
rect 375748 196988 375800 196994
rect 375748 196930 375800 196936
rect 375656 148232 375708 148238
rect 375656 148174 375708 148180
rect 375760 141982 375788 196930
rect 375852 144566 375880 216378
rect 376128 214674 376156 286350
rect 376772 218890 376800 290498
rect 376864 290494 376892 361558
rect 376944 354816 376996 354822
rect 376944 354758 376996 354764
rect 376852 290488 376904 290494
rect 376852 290430 376904 290436
rect 376760 218884 376812 218890
rect 376760 218826 376812 218832
rect 376864 218754 376892 290430
rect 376956 283626 376984 354758
rect 377048 291242 377076 362986
rect 378140 356244 378192 356250
rect 378140 356186 378192 356192
rect 377128 352640 377180 352646
rect 377128 352582 377180 352588
rect 377036 291236 377088 291242
rect 377036 291178 377088 291184
rect 377140 288386 377168 352582
rect 377404 295384 377456 295390
rect 377404 295326 377456 295332
rect 377128 288380 377180 288386
rect 377128 288322 377180 288328
rect 376944 283620 376996 283626
rect 376944 283562 376996 283568
rect 377220 283620 377272 283626
rect 377220 283562 377272 283568
rect 377128 224256 377180 224262
rect 377128 224198 377180 224204
rect 376944 224188 376996 224194
rect 376944 224130 376996 224136
rect 376852 218748 376904 218754
rect 376852 218690 376904 218696
rect 376864 218090 376892 218690
rect 376772 218062 376892 218090
rect 376116 214668 376168 214674
rect 376116 214610 376168 214616
rect 376772 146130 376800 218062
rect 376852 218000 376904 218006
rect 376852 217942 376904 217948
rect 376864 146198 376892 217942
rect 376956 214606 376984 224130
rect 377036 222080 377088 222086
rect 377036 222022 377088 222028
rect 377048 220930 377076 222022
rect 377036 220924 377088 220930
rect 377036 220866 377088 220872
rect 376944 214600 376996 214606
rect 376944 214542 376996 214548
rect 376852 146192 376904 146198
rect 376852 146134 376904 146140
rect 376760 146124 376812 146130
rect 376760 146066 376812 146072
rect 375840 144560 375892 144566
rect 375840 144502 375892 144508
rect 376956 143478 376984 214542
rect 377048 150346 377076 220866
rect 377140 153134 377168 224198
rect 377232 211886 377260 283562
rect 377416 223514 377444 295326
rect 378152 285122 378180 356186
rect 378244 295254 378272 365842
rect 378324 364404 378376 364410
rect 378324 364346 378376 364352
rect 378232 295248 378284 295254
rect 378232 295190 378284 295196
rect 378244 294778 378272 295190
rect 378232 294772 378284 294778
rect 378232 294714 378284 294720
rect 378232 294636 378284 294642
rect 378232 294578 378284 294584
rect 378140 285116 378192 285122
rect 378140 285058 378192 285064
rect 378140 284368 378192 284374
rect 378140 284310 378192 284316
rect 377404 223508 377456 223514
rect 377404 223450 377456 223456
rect 377220 211880 377272 211886
rect 377220 211822 377272 211828
rect 378152 211818 378180 284310
rect 378244 223582 378272 294578
rect 378336 293282 378364 364346
rect 378416 362976 378468 362982
rect 378416 362918 378468 362924
rect 378324 293276 378376 293282
rect 378324 293218 378376 293224
rect 378336 292602 378364 293218
rect 378324 292596 378376 292602
rect 378324 292538 378376 292544
rect 378324 291916 378376 291922
rect 378324 291858 378376 291864
rect 378232 223576 378284 223582
rect 378232 223518 378284 223524
rect 378336 220946 378364 291858
rect 378428 291854 378456 362918
rect 379520 359508 379572 359514
rect 379520 359450 379572 359456
rect 379532 297430 379560 359450
rect 379612 352572 379664 352578
rect 379612 352514 379664 352520
rect 379520 297424 379572 297430
rect 379520 297366 379572 297372
rect 378508 292596 378560 292602
rect 378508 292538 378560 292544
rect 378416 291848 378468 291854
rect 378416 291790 378468 291796
rect 378416 222148 378468 222154
rect 378416 222090 378468 222096
rect 378244 220918 378364 220946
rect 378244 220726 378272 220918
rect 378324 220788 378376 220794
rect 378324 220730 378376 220736
rect 378232 220720 378284 220726
rect 378232 220662 378284 220668
rect 378232 218068 378284 218074
rect 378232 218010 378284 218016
rect 378140 211812 378192 211818
rect 378140 211754 378192 211760
rect 377128 153128 377180 153134
rect 377128 153070 377180 153076
rect 377036 150340 377088 150346
rect 377036 150282 377088 150288
rect 376944 143472 376996 143478
rect 376944 143414 376996 143420
rect 375748 141976 375800 141982
rect 375748 141918 375800 141924
rect 378152 140690 378180 211754
rect 378244 147558 378272 218010
rect 378336 149054 378364 220730
rect 378428 150414 378456 222090
rect 378520 222086 378548 292538
rect 379532 225010 379560 297366
rect 379624 286346 379652 352514
rect 380900 295452 380952 295458
rect 380900 295394 380952 295400
rect 380912 287054 380940 295394
rect 381004 295390 381032 367066
rect 381096 298110 381124 368494
rect 383660 358828 383712 358834
rect 383660 358770 383712 358776
rect 382464 357468 382516 357474
rect 382464 357410 382516 357416
rect 381176 356176 381228 356182
rect 381176 356118 381228 356124
rect 381084 298104 381136 298110
rect 381084 298046 381136 298052
rect 381096 297498 381124 298046
rect 381084 297492 381136 297498
rect 381084 297434 381136 297440
rect 380992 295384 381044 295390
rect 380992 295326 381044 295332
rect 381084 294772 381136 294778
rect 381084 294714 381136 294720
rect 380912 287026 381032 287054
rect 379612 286340 379664 286346
rect 379612 286282 379664 286288
rect 379520 225004 379572 225010
rect 379520 224946 379572 224952
rect 379624 224262 379652 286282
rect 380900 285728 380952 285734
rect 380900 285670 380952 285676
rect 379612 224256 379664 224262
rect 379612 224198 379664 224204
rect 379520 224052 379572 224058
rect 379520 223994 379572 224000
rect 379532 223786 379560 223994
rect 379520 223780 379572 223786
rect 379520 223722 379572 223728
rect 378508 222080 378560 222086
rect 378508 222022 378560 222028
rect 379532 153202 379560 223722
rect 379612 214668 379664 214674
rect 379612 214610 379664 214616
rect 379624 197266 379652 214610
rect 380912 213466 380940 285670
rect 381004 224058 381032 287026
rect 380992 224052 381044 224058
rect 380992 223994 381044 224000
rect 380992 223576 381044 223582
rect 380992 223518 381044 223524
rect 380820 213438 380940 213466
rect 380820 213110 380848 213438
rect 380900 213308 380952 213314
rect 380900 213250 380952 213256
rect 380808 213104 380860 213110
rect 380808 213046 380860 213052
rect 379612 197260 379664 197266
rect 379612 197202 379664 197208
rect 379520 153196 379572 153202
rect 379520 153138 379572 153144
rect 378416 150408 378468 150414
rect 378416 150350 378468 150356
rect 378324 149048 378376 149054
rect 378324 148990 378376 148996
rect 378232 147552 378284 147558
rect 378232 147494 378284 147500
rect 379624 143546 379652 197202
rect 380912 197062 380940 213250
rect 380900 197056 380952 197062
rect 380900 196998 380952 197004
rect 379612 143540 379664 143546
rect 379612 143482 379664 143488
rect 380912 142050 380940 196998
rect 381004 151706 381032 223518
rect 381096 222698 381124 294714
rect 381188 285666 381216 356118
rect 382280 356108 382332 356114
rect 382280 356050 382332 356056
rect 381176 285660 381228 285666
rect 381176 285602 381228 285608
rect 381188 284442 381216 285602
rect 381176 284436 381228 284442
rect 381176 284378 381228 284384
rect 382292 284374 382320 356050
rect 382372 297492 382424 297498
rect 382372 297434 382424 297440
rect 382280 284368 382332 284374
rect 382280 284310 382332 284316
rect 382384 225622 382412 297434
rect 382476 286414 382504 357410
rect 383672 288538 383700 358770
rect 396736 327758 396764 699654
rect 396724 327752 396776 327758
rect 396724 327694 396776 327700
rect 429212 305794 429240 703582
rect 429672 703474 429700 703582
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494072 703582 494652 703610
rect 429856 703474 429884 703520
rect 429672 703446 429884 703474
rect 462332 699718 462360 703520
rect 478524 700534 478552 703520
rect 478512 700528 478564 700534
rect 478512 700470 478564 700476
rect 461584 699712 461636 699718
rect 461584 699654 461636 699660
rect 462320 699712 462372 699718
rect 462320 699654 462372 699660
rect 445206 369472 445262 369481
rect 445206 369407 445262 369416
rect 445220 368558 445248 369407
rect 445208 368552 445260 368558
rect 445208 368494 445260 368500
rect 452844 368552 452896 368558
rect 452844 368494 452896 368500
rect 445666 368384 445722 368393
rect 445666 368319 445722 368328
rect 445680 367266 445708 368319
rect 445668 367260 445720 367266
rect 445668 367202 445720 367208
rect 452660 367260 452712 367266
rect 452660 367202 452712 367208
rect 445666 367160 445722 367169
rect 445722 367118 445800 367146
rect 445666 367095 445722 367104
rect 444930 366072 444986 366081
rect 444930 366007 444986 366016
rect 444944 365770 444972 366007
rect 444932 365764 444984 365770
rect 444932 365706 444984 365712
rect 444930 364848 444986 364857
rect 444930 364783 444986 364792
rect 444944 364682 444972 364783
rect 444932 364676 444984 364682
rect 444932 364618 444984 364624
rect 444562 363760 444618 363769
rect 444562 363695 444618 363704
rect 444576 363186 444604 363695
rect 444564 363180 444616 363186
rect 444564 363122 444616 363128
rect 444930 362536 444986 362545
rect 444930 362471 444986 362480
rect 444944 361622 444972 362471
rect 444932 361616 444984 361622
rect 444932 361558 444984 361564
rect 445668 360256 445720 360262
rect 445666 360224 445668 360233
rect 445720 360224 445722 360233
rect 445666 360159 445722 360168
rect 444470 359136 444526 359145
rect 444470 359071 444526 359080
rect 444484 358834 444512 359071
rect 444472 358828 444524 358834
rect 444472 358770 444524 358776
rect 444930 357912 444986 357921
rect 444930 357847 444986 357856
rect 444944 357474 444972 357847
rect 444932 357468 444984 357474
rect 444932 357410 444984 357416
rect 444562 356824 444618 356833
rect 444562 356759 444564 356768
rect 444616 356759 444618 356768
rect 444564 356730 444616 356736
rect 444378 355600 444434 355609
rect 444378 355535 444434 355544
rect 444392 355162 444420 355535
rect 444380 355156 444432 355162
rect 444380 355098 444432 355104
rect 444470 354512 444526 354521
rect 444470 354447 444526 354456
rect 444484 353394 444512 354447
rect 444472 353388 444524 353394
rect 444472 353330 444524 353336
rect 444378 353288 444434 353297
rect 444378 353223 444434 353232
rect 444392 352034 444420 353223
rect 444380 352028 444432 352034
rect 444380 351970 444432 351976
rect 444562 350976 444618 350985
rect 444562 350911 444618 350920
rect 444378 349888 444434 349897
rect 444378 349823 444434 349832
rect 431972 340054 432952 340082
rect 434732 340054 434884 340082
rect 436112 340054 436908 340082
rect 438932 340054 438992 340082
rect 440956 340054 441292 340082
rect 429200 305788 429252 305794
rect 429200 305730 429252 305736
rect 383580 288510 383700 288538
rect 383580 287094 383608 288510
rect 383660 288380 383712 288386
rect 383660 288322 383712 288328
rect 382648 287088 382700 287094
rect 382648 287030 382700 287036
rect 383568 287088 383620 287094
rect 383568 287030 383620 287036
rect 382464 286408 382516 286414
rect 382464 286350 382516 286356
rect 382556 284436 382608 284442
rect 382556 284378 382608 284384
rect 382372 225616 382424 225622
rect 382372 225558 382424 225564
rect 381176 223508 381228 223514
rect 381176 223450 381228 223456
rect 381084 222692 381136 222698
rect 381084 222634 381136 222640
rect 381188 151774 381216 223450
rect 382280 215348 382332 215354
rect 382280 215290 382332 215296
rect 381176 151768 381228 151774
rect 381176 151710 381228 151716
rect 380992 151700 381044 151706
rect 380992 151642 381044 151648
rect 382292 144838 382320 215290
rect 382384 154562 382412 225558
rect 382464 224188 382516 224194
rect 382464 224130 382516 224136
rect 382476 216578 382504 224130
rect 382464 216572 382516 216578
rect 382464 216514 382516 216520
rect 382568 213246 382596 284378
rect 382660 224194 382688 287030
rect 382648 224188 382700 224194
rect 382648 224130 382700 224136
rect 383672 223990 383700 288322
rect 431972 287054 432000 340054
rect 434732 299130 434760 340054
rect 434720 299124 434772 299130
rect 434720 299066 434772 299072
rect 436112 297634 436140 340054
rect 438964 337482 438992 340054
rect 438952 337476 439004 337482
rect 438952 337418 439004 337424
rect 441264 336802 441292 340054
rect 441252 336796 441304 336802
rect 441252 336738 441304 336744
rect 441620 336796 441672 336802
rect 441620 336738 441672 336744
rect 436100 297628 436152 297634
rect 436100 297570 436152 297576
rect 431972 287026 432552 287054
rect 432524 268682 432552 287026
rect 432524 268654 432952 268682
rect 432616 265742 432644 268654
rect 441632 268138 441660 336738
rect 443644 299736 443696 299742
rect 443644 299678 443696 299684
rect 441712 299124 441764 299130
rect 441712 299066 441764 299072
rect 434884 268110 435220 268138
rect 436908 268110 437244 268138
rect 435192 266354 435220 268110
rect 437216 267734 437244 268110
rect 438918 268002 438946 268124
rect 440956 268110 441660 268138
rect 438872 267974 438946 268002
rect 437216 267706 437428 267734
rect 435180 266348 435232 266354
rect 435180 266290 435232 266296
rect 436008 266348 436060 266354
rect 436008 266290 436060 266296
rect 431960 265736 432012 265742
rect 431960 265678 432012 265684
rect 432604 265736 432656 265742
rect 432604 265678 432656 265684
rect 383660 223984 383712 223990
rect 383660 223926 383712 223932
rect 383672 216646 383700 223926
rect 382648 216640 382700 216646
rect 382648 216582 382700 216588
rect 383660 216640 383712 216646
rect 383660 216582 383712 216588
rect 382660 215354 382688 216582
rect 383752 216572 383804 216578
rect 383752 216514 383804 216520
rect 382648 215348 382700 215354
rect 382648 215290 382700 215296
rect 382556 213240 382608 213246
rect 382556 213182 382608 213188
rect 382568 200114 382596 213182
rect 382476 200086 382596 200114
rect 382476 197130 382504 200086
rect 382464 197124 382516 197130
rect 382464 197066 382516 197072
rect 382372 154556 382424 154562
rect 382372 154498 382424 154504
rect 382280 144832 382332 144838
rect 382280 144774 382332 144780
rect 382476 142118 382504 197066
rect 383764 144906 383792 216514
rect 431972 209774 432000 265678
rect 436020 227798 436048 266290
rect 437400 266286 437428 267706
rect 437388 266280 437440 266286
rect 437388 266222 437440 266228
rect 436008 227792 436060 227798
rect 436008 227734 436060 227740
rect 437400 226302 437428 266222
rect 438872 265674 438900 267974
rect 441356 266218 441384 268110
rect 441724 266354 441752 299066
rect 441804 297628 441856 297634
rect 441804 297570 441856 297576
rect 441712 266348 441764 266354
rect 441712 266290 441764 266296
rect 441816 266286 441844 297570
rect 441804 266280 441856 266286
rect 441540 266218 441660 266234
rect 441804 266222 441856 266228
rect 441344 266212 441396 266218
rect 441344 266154 441396 266160
rect 441528 266212 441660 266218
rect 441580 266206 441660 266212
rect 441528 266154 441580 266160
rect 438860 265668 438912 265674
rect 438860 265610 438912 265616
rect 437388 226296 437440 226302
rect 437388 226238 437440 226244
rect 431972 209746 432552 209774
rect 432524 196058 432552 209746
rect 441632 196874 441660 266206
rect 441896 227792 441948 227798
rect 441896 227734 441948 227740
rect 441712 226296 441764 226302
rect 441712 226238 441764 226244
rect 441724 223802 441752 226238
rect 441802 225040 441858 225049
rect 441802 224975 441804 224984
rect 441856 224975 441858 224984
rect 441804 224946 441856 224952
rect 441802 223952 441858 223961
rect 441802 223887 441804 223896
rect 441856 223887 441858 223896
rect 441804 223858 441856 223864
rect 441724 223774 441844 223802
rect 441712 223644 441764 223650
rect 441712 223586 441764 223592
rect 441540 196846 441660 196874
rect 441540 196058 441568 196846
rect 432524 196030 432952 196058
rect 434884 196030 435220 196058
rect 436908 196030 437428 196058
rect 432524 180794 432552 196030
rect 435192 193662 435220 196030
rect 437400 194546 437428 196030
rect 438780 196030 438932 196058
rect 440956 196030 441568 196058
rect 438780 195974 438808 196030
rect 438768 195968 438820 195974
rect 438768 195910 438820 195916
rect 437388 194540 437440 194546
rect 437388 194482 437440 194488
rect 436008 194472 436060 194478
rect 436008 194414 436060 194420
rect 436020 193662 436048 194414
rect 435180 193656 435232 193662
rect 435180 193598 435232 193604
rect 436008 193656 436060 193662
rect 436008 193598 436060 193604
rect 431972 180766 432552 180794
rect 383752 144900 383804 144906
rect 383752 144842 383804 144848
rect 382464 142112 382516 142118
rect 382464 142054 382516 142060
rect 380900 142044 380952 142050
rect 380900 141986 380952 141992
rect 378140 140684 378192 140690
rect 378140 140626 378192 140632
rect 375380 139256 375432 139262
rect 375380 139198 375432 139204
rect 374092 138916 374144 138922
rect 374092 138858 374144 138864
rect 431972 132494 432000 180766
rect 436020 155922 436048 193598
rect 436008 155916 436060 155922
rect 436008 155858 436060 155864
rect 437400 153610 437428 194482
rect 441356 193214 441384 196030
rect 441724 194478 441752 223586
rect 441816 194546 441844 223774
rect 441908 223650 441936 227734
rect 441896 223644 441948 223650
rect 441896 223586 441948 223592
rect 441804 194540 441856 194546
rect 441804 194482 441856 194488
rect 441712 194472 441764 194478
rect 441712 194414 441764 194420
rect 441356 193186 441660 193214
rect 437388 153604 437440 153610
rect 437388 153546 437440 153552
rect 431972 132466 432552 132494
rect 374000 129124 374052 129130
rect 374000 129066 374052 129072
rect 427820 129124 427872 129130
rect 427820 129066 427872 129072
rect 372620 125520 372672 125526
rect 372620 125462 372672 125468
rect 427832 125458 427860 129066
rect 430580 129056 430632 129062
rect 430580 128998 430632 129004
rect 427820 125452 427872 125458
rect 427820 125394 427872 125400
rect 430592 125390 430620 128998
rect 430580 125384 430632 125390
rect 430580 125326 430632 125332
rect 432524 124794 432552 132466
rect 441632 125594 441660 193186
rect 441712 155916 441764 155922
rect 441712 155858 441764 155864
rect 441356 125566 441660 125594
rect 441356 124794 441384 125566
rect 441620 125520 441672 125526
rect 441618 125488 441620 125497
rect 441672 125488 441674 125497
rect 441618 125423 441674 125432
rect 432524 124766 432952 124794
rect 440956 124766 441384 124794
rect 434884 124086 435220 124114
rect 436908 124086 437244 124114
rect 435192 122670 435220 124086
rect 437216 122738 437244 124086
rect 438918 123842 438946 124100
rect 438872 123814 438946 123842
rect 438872 122806 438900 123814
rect 438860 122800 438912 122806
rect 438860 122742 438912 122748
rect 437204 122732 437256 122738
rect 437204 122674 437256 122680
rect 441724 122670 441752 155858
rect 441896 153604 441948 153610
rect 441896 153546 441948 153552
rect 441908 142154 441936 153546
rect 443656 153202 443684 299678
rect 444392 278730 444420 349823
rect 444470 347576 444526 347585
rect 444470 347511 444526 347520
rect 444380 278724 444432 278730
rect 444380 278666 444432 278672
rect 444484 275641 444512 347511
rect 444576 280090 444604 350911
rect 444654 348664 444710 348673
rect 444654 348599 444710 348608
rect 444564 280084 444616 280090
rect 444564 280026 444616 280032
rect 444668 277394 444696 348599
rect 445206 346352 445262 346361
rect 445206 346287 445262 346296
rect 445220 345642 445248 346287
rect 445208 345636 445260 345642
rect 445208 345578 445260 345584
rect 445666 345264 445722 345273
rect 445666 345199 445722 345208
rect 445680 345166 445708 345199
rect 445668 345160 445720 345166
rect 445668 345102 445720 345108
rect 445666 344040 445722 344049
rect 445666 343975 445722 343984
rect 445680 343670 445708 343975
rect 445668 343664 445720 343670
rect 445668 343606 445720 343612
rect 445666 342952 445722 342961
rect 445666 342887 445722 342896
rect 445680 342310 445708 342887
rect 445668 342304 445720 342310
rect 445668 342246 445720 342252
rect 445114 341728 445170 341737
rect 445114 341663 445170 341672
rect 445128 341018 445156 341663
rect 445116 341012 445168 341018
rect 445116 340954 445168 340960
rect 444746 340640 444802 340649
rect 444746 340575 444802 340584
rect 444760 340270 444788 340575
rect 444748 340264 444800 340270
rect 444748 340206 444800 340212
rect 445666 297528 445722 297537
rect 445666 297463 445722 297472
rect 445680 297022 445708 297463
rect 445668 297016 445720 297022
rect 445668 296958 445720 296964
rect 445666 296440 445722 296449
rect 445666 296375 445722 296384
rect 445680 296002 445708 296375
rect 445668 295996 445720 296002
rect 445668 295938 445720 295944
rect 445668 295248 445720 295254
rect 445772 295225 445800 367118
rect 448612 365764 448664 365770
rect 448612 365706 448664 365712
rect 447416 363180 447468 363186
rect 447416 363122 447468 363128
rect 445850 361448 445906 361457
rect 445850 361383 445906 361392
rect 445668 295190 445720 295196
rect 445758 295216 445814 295225
rect 445680 294137 445708 295190
rect 445758 295151 445814 295160
rect 445666 294128 445722 294137
rect 445666 294063 445722 294072
rect 445772 294030 445800 295151
rect 445760 294024 445812 294030
rect 445760 293966 445812 293972
rect 445668 292936 445720 292942
rect 445666 292904 445668 292913
rect 445720 292904 445722 292913
rect 445666 292839 445722 292848
rect 445666 291816 445722 291825
rect 445666 291751 445722 291760
rect 445680 291242 445708 291751
rect 445668 291236 445720 291242
rect 445668 291178 445720 291184
rect 445668 290624 445720 290630
rect 445666 290592 445668 290601
rect 445720 290592 445722 290601
rect 445666 290527 445722 290536
rect 445666 289504 445722 289513
rect 445864 289474 445892 361383
rect 447232 358828 447284 358834
rect 447232 358770 447284 358776
rect 446036 355156 446088 355162
rect 446036 355098 446088 355104
rect 445942 352200 445998 352209
rect 445942 352135 445998 352144
rect 445666 289439 445668 289448
rect 445720 289439 445722 289448
rect 445852 289468 445904 289474
rect 445668 289410 445720 289416
rect 445852 289410 445904 289416
rect 445668 288380 445720 288386
rect 445668 288322 445720 288328
rect 445680 288289 445708 288322
rect 445666 288280 445722 288289
rect 445666 288215 445722 288224
rect 445116 288108 445168 288114
rect 445116 288050 445168 288056
rect 445128 287201 445156 288050
rect 445114 287192 445170 287201
rect 445114 287127 445170 287136
rect 445666 285968 445722 285977
rect 445666 285903 445722 285912
rect 445680 285734 445708 285903
rect 445668 285728 445720 285734
rect 445668 285670 445720 285676
rect 445668 284912 445720 284918
rect 445666 284880 445668 284889
rect 445720 284880 445722 284889
rect 445666 284815 445722 284824
rect 445484 283688 445536 283694
rect 445482 283656 445484 283665
rect 445536 283656 445538 283665
rect 445482 283591 445538 283600
rect 445390 282568 445446 282577
rect 445390 282503 445392 282512
rect 445444 282503 445446 282512
rect 445392 282474 445444 282480
rect 445116 281512 445168 281518
rect 445116 281454 445168 281460
rect 445128 281353 445156 281454
rect 445114 281344 445170 281353
rect 445114 281279 445170 281288
rect 445956 280634 445984 352135
rect 446048 283694 446076 355098
rect 447140 352028 447192 352034
rect 447140 351970 447192 351976
rect 446128 340264 446180 340270
rect 446128 340206 446180 340212
rect 446036 283688 446088 283694
rect 446036 283630 446088 283636
rect 446048 282946 446076 283630
rect 446036 282940 446088 282946
rect 446036 282882 446088 282888
rect 444748 280628 444800 280634
rect 444748 280570 444800 280576
rect 445944 280628 445996 280634
rect 445944 280570 445996 280576
rect 444760 280265 444788 280570
rect 444746 280256 444802 280265
rect 444746 280191 444802 280200
rect 444840 280084 444892 280090
rect 444840 280026 444892 280032
rect 444852 279041 444880 280026
rect 444838 279032 444894 279041
rect 444838 278967 444894 278976
rect 444576 277366 444696 277394
rect 444576 276729 444604 277366
rect 444562 276720 444618 276729
rect 444562 276655 444618 276664
rect 444470 275632 444526 275641
rect 444470 275567 444526 275576
rect 444378 206952 444434 206961
rect 444378 206887 444434 206896
rect 443644 153196 443696 153202
rect 443644 153138 443696 153144
rect 441816 142126 441936 142154
rect 441816 122738 441844 142126
rect 444392 142118 444420 206887
rect 444484 203561 444512 275567
rect 444576 204649 444604 276655
rect 444746 208176 444802 208185
rect 444746 208111 444802 208120
rect 444760 207942 444788 208111
rect 444748 207936 444800 207942
rect 444748 207878 444800 207884
rect 444852 206961 444880 278967
rect 445116 278724 445168 278730
rect 445116 278666 445168 278672
rect 445128 277953 445156 278666
rect 445114 277944 445170 277953
rect 445114 277879 445170 277888
rect 444838 206952 444894 206961
rect 444838 206887 444894 206896
rect 445128 205873 445156 277879
rect 445576 274644 445628 274650
rect 445576 274586 445628 274592
rect 445588 273329 445616 274586
rect 445666 274408 445722 274417
rect 445666 274343 445722 274352
rect 445574 273320 445630 273329
rect 445680 273290 445708 274343
rect 445574 273255 445630 273264
rect 445668 273284 445720 273290
rect 445668 273226 445720 273232
rect 445668 272536 445720 272542
rect 445668 272478 445720 272484
rect 445680 272105 445708 272478
rect 445666 272096 445722 272105
rect 445666 272031 445722 272040
rect 445666 271008 445722 271017
rect 445666 270943 445722 270952
rect 445680 270638 445708 270943
rect 445668 270632 445720 270638
rect 445668 270574 445720 270580
rect 445666 269784 445722 269793
rect 445666 269719 445722 269728
rect 445680 269142 445708 269719
rect 445668 269136 445720 269142
rect 445668 269078 445720 269084
rect 445666 268696 445722 268705
rect 445722 268654 445800 268682
rect 445666 268631 445722 268640
rect 445772 267734 445800 268654
rect 446140 267734 446168 340206
rect 446404 302728 446456 302734
rect 446404 302670 446456 302676
rect 445772 267706 446168 267734
rect 445576 225616 445628 225622
rect 445576 225558 445628 225564
rect 445588 225457 445616 225558
rect 445574 225448 445630 225457
rect 445574 225383 445630 225392
rect 445668 223168 445720 223174
rect 445666 223136 445668 223145
rect 445720 223136 445722 223145
rect 445666 223071 445722 223080
rect 445666 222048 445722 222057
rect 445666 221983 445722 221992
rect 445680 221270 445708 221983
rect 445668 221264 445720 221270
rect 445668 221206 445720 221212
rect 445666 220824 445722 220833
rect 445666 220759 445668 220768
rect 445720 220759 445722 220768
rect 445668 220730 445720 220736
rect 445666 219736 445722 219745
rect 445666 219671 445722 219680
rect 445680 219638 445708 219671
rect 445668 219632 445720 219638
rect 445668 219574 445720 219580
rect 445482 218512 445538 218521
rect 445482 218447 445484 218456
rect 445536 218447 445538 218456
rect 445484 218418 445536 218424
rect 445666 217424 445722 217433
rect 445666 217359 445668 217368
rect 445720 217359 445722 217368
rect 445668 217330 445720 217336
rect 445666 216200 445722 216209
rect 445666 216135 445668 216144
rect 445720 216135 445722 216144
rect 445668 216106 445720 216112
rect 445482 215112 445538 215121
rect 445482 215047 445538 215056
rect 445496 214810 445524 215047
rect 445484 214804 445536 214810
rect 445484 214746 445536 214752
rect 445668 213920 445720 213926
rect 445666 213888 445668 213897
rect 445720 213888 445722 213897
rect 445666 213823 445722 213832
rect 445666 212800 445722 212809
rect 445666 212735 445668 212744
rect 445720 212735 445722 212744
rect 445668 212706 445720 212712
rect 445484 211608 445536 211614
rect 445482 211576 445484 211585
rect 445536 211576 445538 211585
rect 445482 211511 445538 211520
rect 445392 210520 445444 210526
rect 445390 210488 445392 210497
rect 445444 210488 445446 210497
rect 445390 210423 445446 210432
rect 445206 209264 445262 209273
rect 445206 209199 445208 209208
rect 445260 209199 445262 209208
rect 445208 209170 445260 209176
rect 444654 205864 444710 205873
rect 444654 205799 444710 205808
rect 445114 205864 445170 205873
rect 445114 205799 445170 205808
rect 444562 204640 444618 204649
rect 444562 204575 444618 204584
rect 444470 203552 444526 203561
rect 444470 203487 444526 203496
rect 444484 158030 444512 203487
rect 444472 158024 444524 158030
rect 444472 157966 444524 157972
rect 444380 142112 444432 142118
rect 444380 142054 444432 142060
rect 444380 141976 444432 141982
rect 444378 141944 444380 141953
rect 444432 141944 444434 141953
rect 444378 141879 444434 141888
rect 444380 140480 444432 140486
rect 444380 140422 444432 140428
rect 444392 139641 444420 140422
rect 444378 139632 444434 139641
rect 444378 139567 444434 139576
rect 444380 138644 444432 138650
rect 444380 138586 444432 138592
rect 444392 138553 444420 138586
rect 444378 138544 444434 138553
rect 444378 138479 444434 138488
rect 444380 137352 444432 137358
rect 444378 137320 444380 137329
rect 444432 137320 444434 137329
rect 444378 137255 444434 137264
rect 444484 131617 444512 157966
rect 444576 155242 444604 204575
rect 444668 162246 444696 205799
rect 445666 202328 445722 202337
rect 445666 202263 445722 202272
rect 445680 201550 445708 202263
rect 445668 201544 445720 201550
rect 445668 201486 445720 201492
rect 445666 201240 445722 201249
rect 445666 201175 445722 201184
rect 445680 200190 445708 201175
rect 445668 200184 445720 200190
rect 445668 200126 445720 200132
rect 445666 200016 445722 200025
rect 445666 199951 445722 199960
rect 445680 199510 445708 199951
rect 445668 199504 445720 199510
rect 445668 199446 445720 199452
rect 445666 198928 445722 198937
rect 445666 198863 445722 198872
rect 445680 198830 445708 198863
rect 445668 198824 445720 198830
rect 445720 198784 445800 198812
rect 445668 198766 445720 198772
rect 445668 197804 445720 197810
rect 445668 197746 445720 197752
rect 445680 197713 445708 197746
rect 445666 197704 445722 197713
rect 445666 197639 445722 197648
rect 444656 162240 444708 162246
rect 444656 162182 444708 162188
rect 444564 155236 444616 155242
rect 444564 155178 444616 155184
rect 444576 132705 444604 155178
rect 444668 133929 444696 162182
rect 444748 156664 444800 156670
rect 444748 156606 444800 156612
rect 444760 140865 444788 156606
rect 445668 154556 445720 154562
rect 445668 154498 445720 154504
rect 444932 153876 444984 153882
rect 444932 153818 444984 153824
rect 444838 152416 444894 152425
rect 444838 152351 444894 152360
rect 444852 151910 444880 152351
rect 444840 151904 444892 151910
rect 444840 151846 444892 151852
rect 444840 151360 444892 151366
rect 444840 151302 444892 151308
rect 444852 151201 444880 151302
rect 444838 151192 444894 151201
rect 444838 151127 444894 151136
rect 444944 150113 444972 153818
rect 445680 153513 445708 154498
rect 445666 153504 445722 153513
rect 445666 153439 445722 153448
rect 444930 150104 444986 150113
rect 444930 150039 444986 150048
rect 445300 148912 445352 148918
rect 445298 148880 445300 148889
rect 445352 148880 445354 148889
rect 445298 148815 445354 148824
rect 445576 148164 445628 148170
rect 445576 148106 445628 148112
rect 445588 147801 445616 148106
rect 445574 147792 445630 147801
rect 445574 147727 445630 147736
rect 444840 146600 444892 146606
rect 444838 146568 444840 146577
rect 444892 146568 444894 146577
rect 444838 146503 444894 146512
rect 445484 146056 445536 146062
rect 445484 145998 445536 146004
rect 445496 145489 445524 145998
rect 445482 145480 445538 145489
rect 445482 145415 445538 145424
rect 445116 144764 445168 144770
rect 445116 144706 445168 144712
rect 445128 144265 445156 144706
rect 445114 144256 445170 144265
rect 445114 144191 445170 144200
rect 445116 143200 445168 143206
rect 445114 143168 445116 143177
rect 445168 143168 445170 143177
rect 445114 143103 445170 143112
rect 444840 142112 444892 142118
rect 444840 142054 444892 142060
rect 444746 140856 444802 140865
rect 444746 140791 444802 140800
rect 444746 136232 444802 136241
rect 444746 136167 444802 136176
rect 444654 133920 444710 133929
rect 444654 133855 444710 133864
rect 444562 132696 444618 132705
rect 444562 132631 444618 132640
rect 444470 131608 444526 131617
rect 444470 131543 444526 131552
rect 443920 130416 443972 130422
rect 442998 130384 443054 130393
rect 442998 130319 443054 130328
rect 443918 130384 443920 130393
rect 443972 130384 443974 130393
rect 443918 130319 443974 130328
rect 441894 126440 441950 126449
rect 441894 126375 441950 126384
rect 441908 125322 441936 126375
rect 443012 126002 443040 130319
rect 443642 129296 443698 129305
rect 443642 129231 443698 129240
rect 443656 128382 443684 129231
rect 443644 128376 443696 128382
rect 443644 128318 443696 128324
rect 443090 128072 443146 128081
rect 443090 128007 443146 128016
rect 443104 126070 443132 128007
rect 443092 126064 443144 126070
rect 443092 126006 443144 126012
rect 443000 125996 443052 126002
rect 443000 125938 443052 125944
rect 443656 125934 443684 128318
rect 444380 128104 444432 128110
rect 444378 128072 444380 128081
rect 444432 128072 444434 128081
rect 444378 128007 444434 128016
rect 444380 126676 444432 126682
rect 444380 126618 444432 126624
rect 443644 125928 443696 125934
rect 443644 125870 443696 125876
rect 444392 125769 444420 126618
rect 444378 125760 444434 125769
rect 444378 125695 444434 125704
rect 444760 125458 444788 136167
rect 444852 135017 444880 142054
rect 444838 135008 444894 135017
rect 444838 134943 444894 134952
rect 444748 125452 444800 125458
rect 444748 125394 444800 125400
rect 444852 125390 444880 134943
rect 445666 126984 445722 126993
rect 445772 126970 445800 198784
rect 445864 196625 445892 267706
rect 446128 218952 446180 218958
rect 446128 218894 446180 218900
rect 446140 218482 446168 218894
rect 446128 218476 446180 218482
rect 446128 218418 446180 218424
rect 446036 212492 446088 212498
rect 446036 212434 446088 212440
rect 446048 211614 446076 212434
rect 446036 211608 446088 211614
rect 446036 211550 446088 211556
rect 445944 207936 445996 207942
rect 445944 207878 445996 207884
rect 445850 196616 445906 196625
rect 445850 196551 445906 196560
rect 445722 126942 445800 126970
rect 445666 126919 445722 126928
rect 444840 125384 444892 125390
rect 444840 125326 444892 125332
rect 441896 125316 441948 125322
rect 441896 125258 441948 125264
rect 441894 124944 441950 124953
rect 445864 124914 445892 196551
rect 445956 136241 445984 207878
rect 446048 160138 446076 211550
rect 446140 175234 446168 218418
rect 446416 193186 446444 302670
rect 446496 292936 446548 292942
rect 446496 292878 446548 292884
rect 446508 220794 446536 292878
rect 446680 284912 446732 284918
rect 446680 284854 446732 284860
rect 446588 281512 446640 281518
rect 446588 281454 446640 281460
rect 446496 220788 446548 220794
rect 446496 220730 446548 220736
rect 446600 209234 446628 281454
rect 446692 212770 446720 284854
rect 447152 281518 447180 351970
rect 447244 288114 447272 358770
rect 447324 353388 447376 353394
rect 447324 353330 447376 353336
rect 447232 288108 447284 288114
rect 447232 288050 447284 288056
rect 447336 287054 447364 353330
rect 447428 291242 447456 363122
rect 447968 302796 448020 302802
rect 447968 302738 448020 302744
rect 447784 297016 447836 297022
rect 447784 296958 447836 296964
rect 447796 296886 447824 296958
rect 447784 296880 447836 296886
rect 447784 296822 447836 296828
rect 447416 291236 447468 291242
rect 447416 291178 447468 291184
rect 447244 287026 447364 287054
rect 447244 282538 447272 287026
rect 447232 282532 447284 282538
rect 447232 282474 447284 282480
rect 447140 281512 447192 281518
rect 447140 281454 447192 281460
rect 447140 280628 447192 280634
rect 447140 280570 447192 280576
rect 446680 212764 446732 212770
rect 446680 212706 446732 212712
rect 446588 209228 446640 209234
rect 446588 209170 446640 209176
rect 446600 208418 446628 209170
rect 446588 208412 446640 208418
rect 446588 208354 446640 208360
rect 447152 207942 447180 280570
rect 447244 210526 447272 282474
rect 447796 225622 447824 296822
rect 447876 288380 447928 288386
rect 447876 288322 447928 288328
rect 447784 225616 447836 225622
rect 447784 225558 447836 225564
rect 447508 223576 447560 223582
rect 447508 223518 447560 223524
rect 447520 223174 447548 223518
rect 447508 223168 447560 223174
rect 447508 223110 447560 223116
rect 447324 213920 447376 213926
rect 447324 213862 447376 213868
rect 447232 210520 447284 210526
rect 447232 210462 447284 210468
rect 447140 207936 447192 207942
rect 447140 207878 447192 207884
rect 447140 197804 447192 197810
rect 447140 197746 447192 197752
rect 446404 193180 446456 193186
rect 446404 193122 446456 193128
rect 446128 175228 446180 175234
rect 446128 175170 446180 175176
rect 446036 160132 446088 160138
rect 446036 160074 446088 160080
rect 446048 140486 446076 160074
rect 446140 146606 446168 175170
rect 446128 146600 446180 146606
rect 446128 146542 446180 146548
rect 446036 140480 446088 140486
rect 446036 140422 446088 140428
rect 445942 136232 445998 136241
rect 445942 136167 445998 136176
rect 447152 126682 447180 197746
rect 447244 162178 447272 210462
rect 447232 162172 447284 162178
rect 447232 162114 447284 162120
rect 447244 138650 447272 162114
rect 447336 160070 447364 213862
rect 447416 208412 447468 208418
rect 447416 208354 447468 208360
rect 447428 164286 447456 208354
rect 447520 185609 447548 223110
rect 447888 216170 447916 288322
rect 447980 233238 448008 302738
rect 448624 295254 448652 365706
rect 449992 364676 450044 364682
rect 449992 364618 450044 364624
rect 449900 360256 449952 360262
rect 449900 360198 449952 360204
rect 448888 357468 448940 357474
rect 448888 357410 448940 357416
rect 448704 356788 448756 356794
rect 448704 356730 448756 356736
rect 448612 295248 448664 295254
rect 448612 295190 448664 295196
rect 448624 294098 448652 295190
rect 448612 294092 448664 294098
rect 448612 294034 448664 294040
rect 448612 291168 448664 291174
rect 448612 291110 448664 291116
rect 448624 290630 448652 291110
rect 448612 290624 448664 290630
rect 448612 290566 448664 290572
rect 448520 288108 448572 288114
rect 448520 288050 448572 288056
rect 447968 233232 448020 233238
rect 447968 233174 448020 233180
rect 447876 216164 447928 216170
rect 447876 216106 447928 216112
rect 447888 215354 447916 216106
rect 447876 215348 447928 215354
rect 447876 215290 447928 215296
rect 448532 214810 448560 288050
rect 448624 218958 448652 290566
rect 448716 284918 448744 356730
rect 448796 341012 448848 341018
rect 448796 340954 448848 340960
rect 448704 284912 448756 284918
rect 448704 284854 448756 284860
rect 448704 282940 448756 282946
rect 448704 282882 448756 282888
rect 448612 218952 448664 218958
rect 448612 218894 448664 218900
rect 448520 214804 448572 214810
rect 448520 214746 448572 214752
rect 448612 212764 448664 212770
rect 448612 212706 448664 212712
rect 448520 201544 448572 201550
rect 448520 201486 448572 201492
rect 447506 185600 447562 185609
rect 447506 185535 447562 185544
rect 447416 164280 447468 164286
rect 447416 164222 447468 164228
rect 447324 160064 447376 160070
rect 447324 160006 447376 160012
rect 447336 141982 447364 160006
rect 447324 141976 447376 141982
rect 447324 141918 447376 141924
rect 447232 138644 447284 138650
rect 447232 138586 447284 138592
rect 447428 137358 447456 164222
rect 447520 151366 447548 185535
rect 447508 151360 447560 151366
rect 447508 151302 447560 151308
rect 447416 137352 447468 137358
rect 447416 137294 447468 137300
rect 448532 130422 448560 201486
rect 448624 156670 448652 212706
rect 448716 212498 448744 282882
rect 448808 269142 448836 340954
rect 448900 285734 448928 357410
rect 449164 299600 449216 299606
rect 449164 299542 449216 299548
rect 448888 285728 448940 285734
rect 448888 285670 448940 285676
rect 448796 269136 448848 269142
rect 448796 269078 448848 269084
rect 448888 220788 448940 220794
rect 448888 220730 448940 220736
rect 448796 215348 448848 215354
rect 448796 215290 448848 215296
rect 448704 212492 448756 212498
rect 448704 212434 448756 212440
rect 448808 171134 448836 215290
rect 448900 173233 448928 220730
rect 448886 173224 448942 173233
rect 448886 173159 448942 173168
rect 448716 171106 448836 171134
rect 448716 169726 448744 171106
rect 448704 169720 448756 169726
rect 448704 169662 448756 169668
rect 448612 156664 448664 156670
rect 448612 156606 448664 156612
rect 448716 144770 448744 169662
rect 448900 148918 448928 173159
rect 448888 148912 448940 148918
rect 448888 148854 448940 148860
rect 448704 144764 448756 144770
rect 448704 144706 448756 144712
rect 448520 130416 448572 130422
rect 448520 130358 448572 130364
rect 449176 126954 449204 299542
rect 449912 288386 449940 360198
rect 450004 292942 450032 364618
rect 450084 361616 450136 361622
rect 450084 361558 450136 361564
rect 449992 292936 450044 292942
rect 449992 292878 450044 292884
rect 450096 291174 450124 361558
rect 450176 345636 450228 345642
rect 450176 345578 450228 345584
rect 450084 291168 450136 291174
rect 450084 291110 450136 291116
rect 450084 289468 450136 289474
rect 450084 289410 450136 289416
rect 449900 288380 449952 288386
rect 449900 288322 449952 288328
rect 449900 285728 449952 285734
rect 449900 285670 449952 285676
rect 449256 274644 449308 274650
rect 449256 274586 449308 274592
rect 449268 200190 449296 274586
rect 449912 213926 449940 285670
rect 450096 219434 450124 289410
rect 450188 273290 450216 345578
rect 451372 342304 451424 342310
rect 451372 342246 451424 342252
rect 450544 299668 450596 299674
rect 450544 299610 450596 299616
rect 450268 294024 450320 294030
rect 450268 293966 450320 293972
rect 450176 273284 450228 273290
rect 450176 273226 450228 273232
rect 450280 223582 450308 293966
rect 450268 223576 450320 223582
rect 450268 223518 450320 223524
rect 450176 220040 450228 220046
rect 450176 219982 450228 219988
rect 450188 219638 450216 219982
rect 450176 219632 450228 219638
rect 450176 219574 450228 219580
rect 450004 219406 450124 219434
rect 450004 217394 450032 219406
rect 449992 217388 450044 217394
rect 449992 217330 450044 217336
rect 449900 213920 449952 213926
rect 449900 213862 449952 213868
rect 449256 200184 449308 200190
rect 449256 200126 449308 200132
rect 449900 199504 449952 199510
rect 449900 199446 449952 199452
rect 449912 128110 449940 199446
rect 450004 164218 450032 217330
rect 450084 214804 450136 214810
rect 450084 214746 450136 214752
rect 450096 168366 450124 214746
rect 450188 171737 450216 219574
rect 450556 206990 450584 299610
rect 451280 291236 451332 291242
rect 451280 291178 451332 291184
rect 451292 220046 451320 291178
rect 451384 270638 451412 342246
rect 452672 296002 452700 367202
rect 452752 345160 452804 345166
rect 452752 345102 452804 345108
rect 452660 295996 452712 296002
rect 452660 295938 452712 295944
rect 452672 295390 452700 295938
rect 452660 295384 452712 295390
rect 452660 295326 452712 295332
rect 452660 294092 452712 294098
rect 452660 294034 452712 294040
rect 451372 270632 451424 270638
rect 451372 270574 451424 270580
rect 451280 220040 451332 220046
rect 451280 219982 451332 219988
rect 450544 206984 450596 206990
rect 450544 206926 450596 206932
rect 451384 198830 451412 270574
rect 452672 221270 452700 294034
rect 452764 274650 452792 345102
rect 452856 296886 452884 368494
rect 454040 343664 454092 343670
rect 454040 343606 454092 343612
rect 453304 302388 453356 302394
rect 453304 302330 453356 302336
rect 452844 296880 452896 296886
rect 452844 296822 452896 296828
rect 452752 274644 452804 274650
rect 452752 274586 452804 274592
rect 452936 273284 452988 273290
rect 452936 273226 452988 273232
rect 452844 269136 452896 269142
rect 452844 269078 452896 269084
rect 452752 223916 452804 223922
rect 452752 223858 452804 223864
rect 451464 221264 451516 221270
rect 451464 221206 451516 221212
rect 452660 221264 452712 221270
rect 452660 221206 452712 221212
rect 451372 198824 451424 198830
rect 451372 198766 451424 198772
rect 450174 171728 450230 171737
rect 450174 171663 450230 171672
rect 450084 168360 450136 168366
rect 450084 168302 450136 168308
rect 449992 164212 450044 164218
rect 449992 164154 450044 164160
rect 450004 146062 450032 164154
rect 449992 146056 450044 146062
rect 449992 145998 450044 146004
rect 450096 143206 450124 168302
rect 450188 148170 450216 171663
rect 451476 153882 451504 221206
rect 452660 200184 452712 200190
rect 452660 200126 452712 200132
rect 451464 153876 451516 153882
rect 451464 153818 451516 153824
rect 450176 148164 450228 148170
rect 450176 148106 450228 148112
rect 450084 143200 450136 143206
rect 450084 143142 450136 143148
rect 452672 128382 452700 200126
rect 452764 151910 452792 223858
rect 452856 197810 452884 269078
rect 452948 201550 452976 273226
rect 452936 201544 452988 201550
rect 452936 201486 452988 201492
rect 452844 197804 452896 197810
rect 452844 197746 452896 197752
rect 452752 151904 452804 151910
rect 452752 151846 452804 151852
rect 452660 128376 452712 128382
rect 452660 128318 452712 128324
rect 449900 128104 449952 128110
rect 449900 128046 449952 128052
rect 449164 126948 449216 126954
rect 449164 126890 449216 126896
rect 447140 126676 447192 126682
rect 447140 126618 447192 126624
rect 441894 124879 441896 124888
rect 441948 124879 441950 124888
rect 445852 124908 445904 124914
rect 441896 124850 441948 124856
rect 445852 124850 445904 124856
rect 441804 122732 441856 122738
rect 441804 122674 441856 122680
rect 435180 122664 435232 122670
rect 435180 122606 435232 122612
rect 441712 122664 441764 122670
rect 441712 122606 441764 122612
rect 371792 118652 371844 118658
rect 371792 118594 371844 118600
rect 371332 108996 371384 109002
rect 371332 108938 371384 108944
rect 369860 102128 369912 102134
rect 369860 102070 369912 102076
rect 414664 99340 414716 99346
rect 414664 99282 414716 99288
rect 413284 99272 413336 99278
rect 413284 99214 413336 99220
rect 348424 98592 348476 98598
rect 348424 98534 348476 98540
rect 345664 98524 345716 98530
rect 345664 98466 345716 98472
rect 342904 98456 342956 98462
rect 342904 98398 342956 98404
rect 323676 97980 323728 97986
rect 323676 97922 323728 97928
rect 309876 97912 309928 97918
rect 309876 97854 309928 97860
rect 309784 73160 309836 73166
rect 309784 73102 309836 73108
rect 309152 16546 309824 16574
rect 307944 4004 307996 4010
rect 307944 3946 307996 3952
rect 307024 3392 307076 3398
rect 307024 3334 307076 3340
rect 306576 598 306788 626
rect 306576 490 306604 598
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306392 462 306604 490
rect 306760 480 306788 598
rect 307956 480 307984 3946
rect 309048 3392 309100 3398
rect 309048 3334 309100 3340
rect 309060 480 309088 3334
rect 309796 490 309824 16546
rect 309888 5234 309916 97854
rect 322204 97164 322256 97170
rect 322204 97106 322256 97112
rect 312544 97096 312596 97102
rect 312544 97038 312596 97044
rect 310520 90228 310572 90234
rect 310520 90170 310572 90176
rect 310532 16574 310560 90170
rect 312556 35222 312584 97038
rect 320180 96620 320232 96626
rect 320180 96562 320232 96568
rect 313280 95872 313332 95878
rect 313280 95814 313332 95820
rect 312544 35216 312596 35222
rect 312544 35158 312596 35164
rect 311900 29640 311952 29646
rect 311900 29582 311952 29588
rect 311912 16574 311940 29582
rect 313292 16574 313320 95814
rect 316040 94240 316092 94246
rect 316040 94182 316092 94188
rect 313924 87576 313976 87582
rect 313924 87518 313976 87524
rect 310532 16546 311480 16574
rect 311912 16546 312216 16574
rect 313292 16546 313872 16574
rect 309876 5228 309928 5234
rect 309876 5170 309928 5176
rect 310072 598 310284 626
rect 310072 490 310100 598
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 309796 462 310100 490
rect 310256 480 310284 598
rect 311452 480 311480 16546
rect 312188 490 312216 16546
rect 312464 598 312676 626
rect 312464 490 312492 598
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312188 462 312492 490
rect 312648 480 312676 598
rect 313844 480 313872 16546
rect 313936 3398 313964 87518
rect 316052 3398 316080 94182
rect 317420 91656 317472 91662
rect 317420 91598 317472 91604
rect 316132 86216 316184 86222
rect 316132 86158 316184 86164
rect 316144 16574 316172 86158
rect 316144 16546 316264 16574
rect 313924 3392 313976 3398
rect 313924 3334 313976 3340
rect 315028 3392 315080 3398
rect 315028 3334 315080 3340
rect 316040 3392 316092 3398
rect 316040 3334 316092 3340
rect 315040 480 315068 3334
rect 316236 480 316264 16546
rect 317432 6914 317460 91598
rect 318064 84040 318116 84046
rect 318064 83982 318116 83988
rect 318076 16574 318104 83982
rect 320192 16574 320220 96562
rect 321560 90296 321612 90302
rect 321560 90238 321612 90244
rect 321572 16574 321600 90238
rect 322216 37942 322244 97106
rect 323584 88868 323636 88874
rect 323584 88810 323636 88816
rect 322204 37936 322256 37942
rect 322204 37878 322256 37884
rect 322940 33788 322992 33794
rect 322940 33730 322992 33736
rect 318076 16546 318196 16574
rect 320192 16546 320496 16574
rect 321572 16546 322152 16574
rect 317432 6886 318104 6914
rect 317328 3392 317380 3398
rect 317328 3334 317380 3340
rect 317340 480 317368 3334
rect 318076 490 318104 6886
rect 318168 3398 318196 16546
rect 318156 3392 318208 3398
rect 318156 3334 318208 3340
rect 319720 3392 319772 3398
rect 319720 3334 319772 3340
rect 318352 598 318564 626
rect 318352 490 318380 598
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318076 462 318380 490
rect 318536 480 318564 598
rect 319732 480 319760 3334
rect 320468 490 320496 16546
rect 320744 598 320956 626
rect 320744 490 320772 598
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320468 462 320772 490
rect 320928 480 320956 598
rect 322124 480 322152 16546
rect 322952 490 322980 33730
rect 323596 3398 323624 88810
rect 323688 33794 323716 97922
rect 341524 97844 341576 97850
rect 341524 97786 341576 97792
rect 336004 96552 336056 96558
rect 336004 96494 336056 96500
rect 324412 94444 324464 94450
rect 324412 94386 324464 94392
rect 323676 33788 323728 33794
rect 323676 33730 323728 33736
rect 323584 3392 323636 3398
rect 323584 3334 323636 3340
rect 323136 598 323348 626
rect 323136 490 323164 598
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 322952 462 323164 490
rect 323320 480 323348 598
rect 324424 480 324452 94386
rect 333980 93084 334032 93090
rect 333980 93026 334032 93032
rect 331220 93016 331272 93022
rect 331220 92958 331272 92964
rect 327080 92948 327132 92954
rect 327080 92890 327132 92896
rect 324964 83972 325016 83978
rect 324964 83914 325016 83920
rect 324976 3126 325004 83914
rect 327092 16574 327120 92890
rect 328460 88324 328512 88330
rect 328460 88266 328512 88272
rect 328472 16574 328500 88266
rect 329840 31068 329892 31074
rect 329840 31010 329892 31016
rect 329852 16574 329880 31010
rect 327092 16546 328040 16574
rect 328472 16546 328776 16574
rect 329852 16546 330432 16574
rect 325608 3392 325660 3398
rect 325608 3334 325660 3340
rect 324964 3120 325016 3126
rect 324964 3062 325016 3068
rect 325620 480 325648 3334
rect 326804 3120 326856 3126
rect 326804 3062 326856 3068
rect 326816 480 326844 3062
rect 328012 480 328040 16546
rect 328748 490 328776 16546
rect 329024 598 329236 626
rect 329024 490 329052 598
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 328748 462 329052 490
rect 329208 480 329236 598
rect 330404 480 330432 16546
rect 331232 490 331260 92958
rect 331864 88936 331916 88942
rect 331864 88878 331916 88884
rect 331876 3398 331904 88878
rect 332692 85400 332744 85406
rect 332692 85342 332744 85348
rect 332704 11694 332732 85342
rect 333992 16574 334020 93026
rect 335360 88256 335412 88262
rect 335360 88198 335412 88204
rect 335372 16574 335400 88198
rect 333992 16546 334664 16574
rect 335372 16546 335952 16574
rect 332692 11688 332744 11694
rect 332692 11630 332744 11636
rect 333888 11688 333940 11694
rect 333888 11630 333940 11636
rect 331864 3392 331916 3398
rect 331864 3334 331916 3340
rect 332692 3392 332744 3398
rect 332692 3334 332744 3340
rect 331416 598 331628 626
rect 331416 490 331444 598
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331232 462 331444 490
rect 331600 480 331628 598
rect 332704 480 332732 3334
rect 333900 480 333928 11630
rect 334636 490 334664 16546
rect 335924 3210 335952 16546
rect 336016 3398 336044 96494
rect 338120 93832 338172 93838
rect 338120 93774 338172 93780
rect 338132 16574 338160 93774
rect 339500 86896 339552 86902
rect 339500 86838 339552 86844
rect 338132 16546 338712 16574
rect 336004 3392 336056 3398
rect 336004 3334 336056 3340
rect 337476 3392 337528 3398
rect 337476 3334 337528 3340
rect 335924 3182 336320 3210
rect 334912 598 335124 626
rect 334912 490 334940 598
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 334636 462 334940 490
rect 335096 480 335124 598
rect 336292 480 336320 3182
rect 337488 480 337516 3334
rect 338684 480 338712 16546
rect 339512 490 339540 86838
rect 340972 16040 341024 16046
rect 340972 15982 341024 15988
rect 339696 598 339908 626
rect 339696 490 339724 598
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339512 462 339724 490
rect 339880 480 339908 598
rect 340984 480 341012 15982
rect 341536 6458 341564 97786
rect 342916 16574 342944 98398
rect 342916 16546 343036 16574
rect 342904 12164 342956 12170
rect 342904 12106 342956 12112
rect 342168 6588 342220 6594
rect 342168 6530 342220 6536
rect 341524 6452 341576 6458
rect 341524 6394 341576 6400
rect 342180 480 342208 6530
rect 342916 490 342944 12106
rect 343008 3398 343036 16546
rect 345676 3398 345704 98466
rect 347044 97708 347096 97714
rect 347044 97650 347096 97656
rect 346952 12096 347004 12102
rect 346952 12038 347004 12044
rect 345756 6520 345808 6526
rect 345756 6462 345808 6468
rect 342996 3392 343048 3398
rect 342996 3334 343048 3340
rect 344560 3392 344612 3398
rect 344560 3334 344612 3340
rect 345664 3392 345716 3398
rect 345664 3334 345716 3340
rect 343192 598 343404 626
rect 343192 490 343220 598
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 342916 462 343220 490
rect 343376 480 343404 598
rect 344572 480 344600 3334
rect 345768 480 345796 6462
rect 346964 480 346992 12038
rect 347056 3330 347084 97650
rect 348436 3398 348464 98534
rect 352564 97776 352616 97782
rect 352564 97718 352616 97724
rect 352576 6322 352604 97718
rect 369124 97640 369176 97646
rect 369124 97582 369176 97588
rect 358820 95192 358872 95198
rect 358820 95134 358872 95140
rect 356060 91724 356112 91730
rect 356060 91666 356112 91672
rect 353300 91044 353352 91050
rect 353300 90986 353352 90992
rect 353312 16574 353340 90986
rect 356072 16574 356100 91666
rect 357440 88188 357492 88194
rect 357440 88130 357492 88136
rect 357452 16574 357480 88130
rect 358832 16574 358860 95134
rect 362960 93764 363012 93770
rect 362960 93706 363012 93712
rect 360200 86828 360252 86834
rect 360200 86770 360252 86776
rect 360212 16574 360240 86770
rect 360844 83904 360896 83910
rect 360844 83846 360896 83852
rect 353312 16546 353616 16574
rect 356072 16546 356376 16574
rect 357452 16546 357572 16574
rect 358832 16546 359504 16574
rect 360212 16546 360792 16574
rect 352840 6384 352892 6390
rect 352840 6326 352892 6332
rect 352564 6316 352616 6322
rect 352564 6258 352616 6264
rect 349252 3936 349304 3942
rect 349252 3878 349304 3884
rect 348056 3392 348108 3398
rect 348056 3334 348108 3340
rect 348424 3392 348476 3398
rect 348424 3334 348476 3340
rect 347044 3324 347096 3330
rect 347044 3266 347096 3272
rect 348068 480 348096 3334
rect 349264 480 349292 3878
rect 351644 3392 351696 3398
rect 351644 3334 351696 3340
rect 350448 3324 350500 3330
rect 350448 3266 350500 3272
rect 350460 480 350488 3266
rect 351656 480 351684 3334
rect 352852 480 352880 6326
rect 353588 490 353616 16546
rect 355232 5160 355284 5166
rect 355232 5102 355284 5108
rect 353864 598 354076 626
rect 353864 490 353892 598
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 353588 462 353892 490
rect 354048 480 354076 598
rect 355244 480 355272 5102
rect 356348 480 356376 16546
rect 357544 480 357572 16546
rect 358728 5296 358780 5302
rect 358728 5238 358780 5244
rect 358740 480 358768 5238
rect 359476 490 359504 16546
rect 360764 2938 360792 16546
rect 360856 3126 360884 83846
rect 362972 16574 363000 93706
rect 364984 92472 365036 92478
rect 364984 92414 365036 92420
rect 363604 86760 363656 86766
rect 363604 86702 363656 86708
rect 362972 16546 363552 16574
rect 360844 3120 360896 3126
rect 360844 3062 360896 3068
rect 362316 3120 362368 3126
rect 362316 3062 362368 3068
rect 360764 2910 361160 2938
rect 359752 598 359964 626
rect 359752 490 359780 598
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359476 462 359780 490
rect 359936 480 359964 598
rect 361132 480 361160 2910
rect 362328 480 362356 3062
rect 363524 480 363552 16546
rect 363616 4146 363644 86702
rect 363604 4140 363656 4146
rect 363604 4082 363656 4088
rect 364616 4140 364668 4146
rect 364616 4082 364668 4088
rect 364628 480 364656 4082
rect 364996 3398 365024 92414
rect 367744 88120 367796 88126
rect 367744 88062 367796 88068
rect 365812 82544 365864 82550
rect 365812 82486 365864 82492
rect 364984 3392 365036 3398
rect 364984 3334 365036 3340
rect 365824 480 365852 82486
rect 367756 16574 367784 88062
rect 367756 16546 367876 16574
rect 367744 12028 367796 12034
rect 367744 11970 367796 11976
rect 367008 3392 367060 3398
rect 367008 3334 367060 3340
rect 367020 480 367048 3334
rect 367756 490 367784 11970
rect 367848 3398 367876 16546
rect 367836 3392 367888 3398
rect 367836 3334 367888 3340
rect 369136 2922 369164 97582
rect 377404 97572 377456 97578
rect 377404 97514 377456 97520
rect 369860 92404 369912 92410
rect 369860 92346 369912 92352
rect 369872 16574 369900 92346
rect 374000 92336 374052 92342
rect 374000 92278 374052 92284
rect 369872 16546 370176 16574
rect 369400 3392 369452 3398
rect 369400 3334 369452 3340
rect 369124 2916 369176 2922
rect 369124 2858 369176 2864
rect 368032 598 368244 626
rect 368032 490 368060 598
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 367756 462 368060 490
rect 368216 480 368244 598
rect 369412 480 369440 3334
rect 370148 490 370176 16546
rect 374012 6914 374040 92278
rect 374092 86692 374144 86698
rect 374092 86634 374144 86640
rect 374104 11694 374132 86634
rect 375380 85332 375432 85338
rect 375380 85274 375432 85280
rect 375392 16574 375420 85274
rect 375392 16546 376064 16574
rect 374092 11688 374144 11694
rect 374092 11630 374144 11636
rect 375288 11688 375340 11694
rect 375288 11630 375340 11636
rect 374012 6886 374132 6914
rect 372896 5228 372948 5234
rect 372896 5170 372948 5176
rect 371700 2916 371752 2922
rect 371700 2858 371752 2864
rect 370424 598 370636 626
rect 370424 490 370452 598
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370148 462 370452 490
rect 370608 480 370636 598
rect 371712 480 371740 2858
rect 372908 480 372936 5170
rect 374104 480 374132 6886
rect 375300 480 375328 11630
rect 376036 490 376064 16546
rect 377416 5166 377444 97514
rect 388444 97504 388496 97510
rect 388444 97446 388496 97452
rect 382924 93696 382976 93702
rect 382924 93638 382976 93644
rect 380900 92268 380952 92274
rect 380900 92210 380952 92216
rect 378140 85264 378192 85270
rect 378140 85206 378192 85212
rect 378152 16574 378180 85206
rect 380912 16574 380940 92210
rect 382280 82476 382332 82482
rect 382280 82418 382332 82424
rect 378152 16546 378456 16574
rect 380912 16546 381216 16574
rect 377404 5160 377456 5166
rect 377404 5102 377456 5108
rect 377680 3868 377732 3874
rect 377680 3810 377732 3816
rect 376312 598 376524 626
rect 376312 490 376340 598
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376036 462 376340 490
rect 376496 480 376524 598
rect 377692 480 377720 3810
rect 378428 490 378456 16546
rect 379980 6452 380032 6458
rect 379980 6394 380032 6400
rect 378704 598 378916 626
rect 378704 490 378732 598
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378428 462 378732 490
rect 378888 480 378916 598
rect 379992 480 380020 6394
rect 381188 480 381216 16546
rect 382292 3398 382320 82418
rect 382372 11960 382424 11966
rect 382372 11902 382424 11908
rect 382280 3392 382332 3398
rect 382280 3334 382332 3340
rect 382384 480 382412 11902
rect 382936 3262 382964 93638
rect 385684 92200 385736 92206
rect 385684 92142 385736 92148
rect 385592 11892 385644 11898
rect 385592 11834 385644 11840
rect 383568 3392 383620 3398
rect 383568 3334 383620 3340
rect 382924 3256 382976 3262
rect 382924 3198 382976 3204
rect 383580 480 383608 3334
rect 384764 3256 384816 3262
rect 384764 3198 384816 3204
rect 384776 480 384804 3198
rect 385604 3074 385632 11834
rect 385696 3194 385724 92142
rect 388260 8152 388312 8158
rect 388260 8094 388312 8100
rect 385684 3188 385736 3194
rect 385684 3130 385736 3136
rect 387156 3188 387208 3194
rect 387156 3130 387208 3136
rect 385604 3046 386000 3074
rect 385972 480 386000 3046
rect 387168 480 387196 3130
rect 388272 480 388300 8094
rect 388456 6390 388484 97446
rect 393964 97436 394016 97442
rect 393964 97378 394016 97384
rect 389824 89684 389876 89690
rect 389824 89626 389876 89632
rect 389456 11824 389508 11830
rect 389456 11766 389508 11772
rect 388444 6384 388496 6390
rect 388444 6326 388496 6332
rect 389468 480 389496 11766
rect 389836 3398 389864 89626
rect 392584 82408 392636 82414
rect 392584 82350 392636 82356
rect 392596 16574 392624 82350
rect 392596 16546 392716 16574
rect 392584 11756 392636 11762
rect 392584 11698 392636 11704
rect 391848 8084 391900 8090
rect 391848 8026 391900 8032
rect 389824 3392 389876 3398
rect 389824 3334 389876 3340
rect 390652 3392 390704 3398
rect 390652 3334 390704 3340
rect 390664 480 390692 3334
rect 391860 480 391888 8026
rect 392596 490 392624 11698
rect 392688 3874 392716 16546
rect 393976 6322 394004 97378
rect 411904 97368 411956 97374
rect 411904 97310 411956 97316
rect 407212 93628 407264 93634
rect 407212 93570 407264 93576
rect 396080 92132 396132 92138
rect 396080 92074 396132 92080
rect 395344 83836 395396 83842
rect 395344 83778 395396 83784
rect 395252 8016 395304 8022
rect 395252 7958 395304 7964
rect 394240 6452 394292 6458
rect 394240 6394 394292 6400
rect 393964 6316 394016 6322
rect 393964 6258 394016 6264
rect 392676 3868 392728 3874
rect 392676 3810 392728 3816
rect 392872 598 393084 626
rect 392872 490 392900 598
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 392596 462 392900 490
rect 393056 480 393084 598
rect 394252 480 394280 6394
rect 395264 3482 395292 7958
rect 395356 3942 395384 83778
rect 395344 3936 395396 3942
rect 395344 3878 395396 3884
rect 395264 3454 395384 3482
rect 395356 480 395384 3454
rect 396092 490 396120 92074
rect 406384 90976 406436 90982
rect 406384 90918 406436 90924
rect 398840 89616 398892 89622
rect 398840 89558 398892 89564
rect 397736 3936 397788 3942
rect 397736 3878 397788 3884
rect 396368 598 396580 626
rect 396368 490 396396 598
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396092 462 396396 490
rect 396552 480 396580 598
rect 397748 480 397776 3878
rect 398852 3398 398880 89558
rect 402980 86624 403032 86630
rect 402980 86566 403032 86572
rect 400220 82340 400272 82346
rect 400220 82282 400272 82288
rect 400232 16574 400260 82282
rect 402992 16574 403020 86566
rect 404360 80980 404412 80986
rect 404360 80922 404412 80928
rect 400232 16546 400904 16574
rect 402992 16546 403664 16574
rect 398932 7948 398984 7954
rect 398932 7890 398984 7896
rect 398840 3392 398892 3398
rect 398840 3334 398892 3340
rect 398944 480 398972 7890
rect 400128 3392 400180 3398
rect 400128 3334 400180 3340
rect 400140 480 400168 3334
rect 400876 490 400904 16546
rect 402520 7880 402572 7886
rect 402520 7822 402572 7828
rect 401152 598 401364 626
rect 401152 490 401180 598
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 400876 462 401180 490
rect 401336 480 401364 598
rect 402532 480 402560 7822
rect 403636 480 403664 16546
rect 404372 490 404400 80922
rect 406016 7812 406068 7818
rect 406016 7754 406068 7760
rect 404648 598 404860 626
rect 404648 490 404676 598
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404372 462 404676 490
rect 404832 480 404860 598
rect 406028 480 406056 7754
rect 406396 4146 406424 90918
rect 406384 4140 406436 4146
rect 406384 4082 406436 4088
rect 407224 480 407252 93570
rect 409880 88052 409932 88058
rect 409880 87994 409932 88000
rect 409892 16574 409920 87994
rect 409892 16546 410840 16574
rect 409604 7744 409656 7750
rect 409604 7686 409656 7692
rect 408408 3868 408460 3874
rect 408408 3810 408460 3816
rect 408420 480 408448 3810
rect 409616 480 409644 7686
rect 410812 480 410840 16546
rect 411916 5166 411944 97310
rect 413100 7676 413152 7682
rect 413100 7618 413152 7624
rect 411812 5160 411864 5166
rect 411812 5102 411864 5108
rect 411904 5160 411956 5166
rect 411904 5102 411956 5108
rect 411824 2666 411852 5102
rect 411824 2638 411944 2666
rect 411916 480 411944 2638
rect 413112 480 413140 7618
rect 413296 3194 413324 99214
rect 414296 4140 414348 4146
rect 414296 4082 414348 4088
rect 413284 3188 413336 3194
rect 413284 3130 413336 3136
rect 414308 480 414336 4082
rect 414676 3874 414704 99282
rect 417424 99204 417476 99210
rect 417424 99146 417476 99152
rect 416780 86556 416832 86562
rect 416780 86498 416832 86504
rect 416792 6914 416820 86498
rect 417436 16574 417464 99146
rect 421564 99136 421616 99142
rect 421564 99078 421616 99084
rect 418804 97300 418856 97306
rect 418804 97242 418856 97248
rect 417436 16546 417556 16574
rect 416792 6886 417464 6914
rect 415492 5092 415544 5098
rect 415492 5034 415544 5040
rect 414664 3868 414716 3874
rect 414664 3810 414716 3816
rect 415504 480 415532 5034
rect 416688 3188 416740 3194
rect 416688 3130 416740 3136
rect 416700 480 416728 3130
rect 417436 490 417464 6886
rect 417528 2922 417556 16546
rect 418816 6390 418844 97242
rect 420920 87984 420972 87990
rect 420920 87926 420972 87932
rect 418988 6520 419040 6526
rect 418988 6462 419040 6468
rect 418804 6384 418856 6390
rect 418804 6326 418856 6332
rect 417516 2916 417568 2922
rect 417516 2858 417568 2864
rect 417712 598 417924 626
rect 417712 490 417740 598
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417436 462 417740 490
rect 417896 480 417924 598
rect 419000 480 419028 6462
rect 420184 2916 420236 2922
rect 420184 2858 420236 2864
rect 420196 480 420224 2858
rect 420932 490 420960 87926
rect 421576 3330 421604 99078
rect 430580 99068 430632 99074
rect 430580 99010 430632 99016
rect 428464 92064 428516 92070
rect 428464 92006 428516 92012
rect 425704 86488 425756 86494
rect 425704 86430 425756 86436
rect 423772 85196 423824 85202
rect 423772 85138 423824 85144
rect 423784 11762 423812 85138
rect 425060 35216 425112 35222
rect 425060 35158 425112 35164
rect 423772 11756 423824 11762
rect 423772 11698 423824 11704
rect 424968 11756 425020 11762
rect 424968 11698 425020 11704
rect 422576 6452 422628 6458
rect 422576 6394 422628 6400
rect 421564 3324 421616 3330
rect 421564 3266 421616 3272
rect 421208 598 421420 626
rect 421208 490 421236 598
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 420932 462 421236 490
rect 421392 480 421420 598
rect 422588 480 422616 6394
rect 423772 3324 423824 3330
rect 423772 3266 423824 3272
rect 423784 480 423812 3266
rect 424980 480 425008 11698
rect 425072 6914 425100 35158
rect 425716 16574 425744 86430
rect 425716 16546 425836 16574
rect 425072 6886 425744 6914
rect 425716 490 425744 6886
rect 425808 3942 425836 16546
rect 428372 13728 428424 13734
rect 428372 13670 428424 13676
rect 427268 7608 427320 7614
rect 427268 7550 427320 7556
rect 425796 3936 425848 3942
rect 425796 3878 425848 3884
rect 425992 598 426204 626
rect 425992 490 426020 598
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 425716 462 426020 490
rect 426176 480 426204 598
rect 427280 480 427308 7550
rect 428384 3482 428412 13670
rect 428476 4010 428504 92006
rect 429200 80912 429252 80918
rect 429200 80854 429252 80860
rect 428464 4004 428516 4010
rect 428464 3946 428516 3952
rect 428384 3454 428504 3482
rect 428476 480 428504 3454
rect 429212 490 429240 80854
rect 430592 16574 430620 99010
rect 435364 99000 435416 99006
rect 435364 98942 435416 98948
rect 432604 91996 432656 92002
rect 432604 91938 432656 91944
rect 431224 80844 431276 80850
rect 431224 80786 431276 80792
rect 430592 16546 430896 16574
rect 429488 598 429700 626
rect 429488 490 429516 598
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429212 462 429516 490
rect 429672 480 429700 598
rect 430868 480 430896 16546
rect 431236 3330 431264 80786
rect 432052 13660 432104 13666
rect 432052 13602 432104 13608
rect 431224 3324 431276 3330
rect 431224 3266 431276 3272
rect 432064 480 432092 13602
rect 432616 3398 432644 91938
rect 435088 13592 435140 13598
rect 435088 13534 435140 13540
rect 432604 3392 432656 3398
rect 432604 3334 432656 3340
rect 434444 3392 434496 3398
rect 434444 3334 434496 3340
rect 433248 3324 433300 3330
rect 433248 3266 433300 3272
rect 433260 480 433288 3266
rect 434456 480 434484 3334
rect 435100 490 435128 13534
rect 435376 3398 435404 98942
rect 439504 98932 439556 98938
rect 439504 98874 439556 98880
rect 436742 97472 436798 97481
rect 436742 97407 436798 97416
rect 436652 5160 436704 5166
rect 436652 5102 436704 5108
rect 435364 3392 435416 3398
rect 435364 3334 435416 3340
rect 436664 2666 436692 5102
rect 436756 5098 436784 97407
rect 439136 13524 439188 13530
rect 439136 13466 439188 13472
rect 436744 5092 436796 5098
rect 436744 5034 436796 5040
rect 437940 3392 437992 3398
rect 437940 3334 437992 3340
rect 436664 2638 436784 2666
rect 435376 598 435588 626
rect 435376 490 435404 598
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435100 462 435404 490
rect 435560 480 435588 598
rect 436756 480 436784 2638
rect 437952 480 437980 3334
rect 439148 480 439176 13466
rect 439516 3398 439544 98874
rect 448520 98864 448572 98870
rect 448520 98806 448572 98812
rect 443642 97336 443698 97345
rect 443642 97271 443698 97280
rect 440332 80776 440384 80782
rect 440332 80718 440384 80724
rect 439504 3392 439556 3398
rect 439504 3334 439556 3340
rect 440344 480 440372 80718
rect 442632 13456 442684 13462
rect 442632 13398 442684 13404
rect 441528 3392 441580 3398
rect 441528 3334 441580 3340
rect 441540 480 441568 3334
rect 442644 480 442672 13398
rect 443656 5166 443684 97271
rect 446404 91928 446456 91934
rect 446404 91870 446456 91876
rect 445760 13388 445812 13394
rect 445760 13330 445812 13336
rect 443828 6384 443880 6390
rect 443828 6326 443880 6332
rect 443644 5160 443696 5166
rect 443644 5102 443696 5108
rect 443840 480 443868 6326
rect 445024 4004 445076 4010
rect 445024 3946 445076 3952
rect 445036 480 445064 3946
rect 445772 490 445800 13330
rect 446416 2990 446444 91870
rect 447140 79348 447192 79354
rect 447140 79290 447192 79296
rect 447152 16574 447180 79290
rect 448532 16574 448560 98806
rect 453316 20670 453344 302330
rect 454052 272542 454080 343606
rect 461596 323610 461624 699654
rect 461584 323604 461636 323610
rect 461584 323546 461636 323552
rect 494072 304502 494100 703582
rect 494624 703474 494652 703582
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 494808 703474 494836 703520
rect 494624 703446 494836 703474
rect 527192 699718 527220 703520
rect 543476 700330 543504 703520
rect 559668 702434 559696 703520
rect 558932 702406 559696 702434
rect 543464 700324 543516 700330
rect 543464 700266 543516 700272
rect 526444 699712 526496 699718
rect 526444 699654 526496 699660
rect 527180 699712 527232 699718
rect 527180 699654 527232 699660
rect 526456 305658 526484 699654
rect 526444 305652 526496 305658
rect 526444 305594 526496 305600
rect 494060 304496 494112 304502
rect 494060 304438 494112 304444
rect 558932 304434 558960 702406
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 580184 696998 580212 697167
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 580170 683904 580226 683913
rect 580170 683839 580226 683848
rect 580184 683194 580212 683839
rect 580172 683188 580224 683194
rect 580172 683130 580224 683136
rect 580172 670744 580224 670750
rect 580170 670712 580172 670721
rect 580224 670712 580226 670721
rect 580170 670647 580226 670656
rect 580170 644056 580226 644065
rect 580170 643991 580226 644000
rect 580184 643142 580212 643991
rect 580172 643136 580224 643142
rect 580172 643078 580224 643084
rect 580170 630864 580226 630873
rect 580170 630799 580226 630808
rect 580184 630698 580212 630799
rect 580172 630692 580224 630698
rect 580172 630634 580224 630640
rect 580170 617536 580226 617545
rect 580170 617471 580226 617480
rect 580184 616894 580212 617471
rect 580172 616888 580224 616894
rect 580172 616830 580224 616836
rect 579802 591016 579858 591025
rect 579802 590951 579858 590960
rect 579816 590714 579844 590951
rect 579804 590708 579856 590714
rect 579804 590650 579856 590656
rect 580170 577688 580226 577697
rect 580170 577623 580226 577632
rect 580184 576910 580212 577623
rect 580172 576904 580224 576910
rect 580172 576846 580224 576852
rect 579802 564360 579858 564369
rect 579802 564295 579858 564304
rect 579816 563106 579844 564295
rect 579804 563100 579856 563106
rect 579804 563042 579856 563048
rect 580170 537840 580226 537849
rect 580170 537775 580226 537784
rect 580184 536858 580212 537775
rect 580172 536852 580224 536858
rect 580172 536794 580224 536800
rect 580170 524512 580226 524521
rect 580170 524447 580172 524456
rect 580224 524447 580226 524456
rect 580172 524418 580224 524424
rect 580170 511320 580226 511329
rect 580170 511255 580226 511264
rect 580184 510678 580212 511255
rect 580172 510672 580224 510678
rect 580172 510614 580224 510620
rect 580170 484664 580226 484673
rect 580170 484599 580226 484608
rect 580184 484430 580212 484599
rect 580172 484424 580224 484430
rect 580172 484366 580224 484372
rect 579986 471472 580042 471481
rect 579986 471407 580042 471416
rect 580000 470626 580028 471407
rect 579988 470620 580040 470626
rect 579988 470562 580040 470568
rect 580170 458144 580226 458153
rect 580170 458079 580226 458088
rect 580184 456822 580212 458079
rect 580172 456816 580224 456822
rect 580172 456758 580224 456764
rect 580170 431624 580226 431633
rect 580170 431559 580226 431568
rect 580184 430642 580212 431559
rect 580172 430636 580224 430642
rect 580172 430578 580224 430584
rect 580170 418296 580226 418305
rect 580170 418231 580226 418240
rect 580184 418198 580212 418231
rect 580172 418192 580224 418198
rect 580172 418134 580224 418140
rect 580170 404968 580226 404977
rect 580170 404903 580226 404912
rect 580184 404394 580212 404903
rect 580172 404388 580224 404394
rect 580172 404330 580224 404336
rect 580170 378448 580226 378457
rect 580170 378383 580226 378392
rect 580184 378214 580212 378383
rect 580172 378208 580224 378214
rect 580172 378150 580224 378156
rect 580262 365120 580318 365129
rect 580262 365055 580318 365064
rect 580170 325272 580226 325281
rect 580170 325207 580226 325216
rect 580184 324358 580212 325207
rect 580172 324352 580224 324358
rect 580172 324294 580224 324300
rect 580170 312080 580226 312089
rect 580170 312015 580226 312024
rect 580184 311914 580212 312015
rect 580172 311908 580224 311914
rect 580172 311850 580224 311856
rect 558920 304428 558972 304434
rect 558920 304370 558972 304376
rect 580276 304366 580304 365055
rect 580354 351928 580410 351937
rect 580354 351863 580410 351872
rect 580264 304360 580316 304366
rect 580264 304302 580316 304308
rect 580368 304298 580396 351863
rect 580356 304292 580408 304298
rect 580356 304234 580408 304240
rect 464344 302660 464396 302666
rect 464344 302602 464396 302608
rect 461584 302592 461636 302598
rect 461584 302534 461636 302540
rect 457444 302524 457496 302530
rect 457444 302466 457496 302472
rect 454684 302456 454736 302462
rect 454684 302398 454736 302404
rect 454132 295384 454184 295390
rect 454132 295326 454184 295332
rect 454040 272536 454092 272542
rect 454040 272478 454092 272484
rect 454052 199510 454080 272478
rect 454144 223922 454172 295326
rect 454224 225616 454276 225622
rect 454224 225558 454276 225564
rect 454132 223916 454184 223922
rect 454132 223858 454184 223864
rect 454040 199504 454092 199510
rect 454040 199446 454092 199452
rect 454236 154562 454264 225558
rect 454224 154556 454276 154562
rect 454224 154498 454276 154504
rect 453396 86420 453448 86426
rect 453396 86362 453448 86368
rect 453304 20664 453356 20670
rect 453304 20606 453356 20612
rect 447152 16546 447456 16574
rect 448532 16546 448652 16574
rect 446404 2984 446456 2990
rect 446404 2926 446456 2932
rect 446048 598 446260 626
rect 446048 490 446076 598
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 445772 462 446076 490
rect 446232 480 446260 598
rect 447428 480 447456 16546
rect 448624 480 448652 16546
rect 449808 13320 449860 13326
rect 449808 13262 449860 13268
rect 449820 480 449848 13262
rect 453304 13252 453356 13258
rect 453304 13194 453356 13200
rect 450912 3936 450964 3942
rect 450912 3878 450964 3884
rect 450924 480 450952 3878
rect 452108 2984 452160 2990
rect 452108 2926 452160 2932
rect 452120 480 452148 2926
rect 453316 480 453344 13194
rect 453408 3330 453436 86362
rect 454696 60722 454724 302398
rect 457456 100706 457484 302466
rect 461596 179382 461624 302534
rect 464356 259418 464384 302602
rect 465724 301164 465776 301170
rect 465724 301106 465776 301112
rect 464344 259412 464396 259418
rect 464344 259354 464396 259360
rect 461584 179376 461636 179382
rect 461584 179318 461636 179324
rect 465736 139398 465764 301106
rect 582472 300960 582524 300966
rect 582472 300902 582524 300908
rect 582380 300892 582432 300898
rect 582380 300834 582432 300840
rect 580170 298752 580226 298761
rect 580170 298687 580226 298696
rect 580184 298246 580212 298687
rect 580172 298240 580224 298246
rect 580172 298182 580224 298188
rect 580264 298172 580316 298178
rect 580264 298114 580316 298120
rect 580276 272241 580304 298114
rect 580262 272232 580318 272241
rect 580262 272167 580318 272176
rect 580172 259412 580224 259418
rect 580172 259354 580224 259360
rect 580184 258913 580212 259354
rect 580170 258904 580226 258913
rect 580170 258839 580226 258848
rect 580172 245608 580224 245614
rect 580170 245576 580172 245585
rect 580224 245576 580226 245585
rect 580170 245511 580226 245520
rect 579988 233232 580040 233238
rect 579988 233174 580040 233180
rect 580000 232393 580028 233174
rect 579986 232384 580042 232393
rect 579986 232319 580042 232328
rect 580264 227044 580316 227050
rect 580264 226986 580316 226992
rect 580276 219065 580304 226986
rect 580262 219056 580318 219065
rect 580262 218991 580318 219000
rect 579804 206984 579856 206990
rect 579804 206926 579856 206932
rect 579816 205737 579844 206926
rect 579802 205728 579858 205737
rect 579802 205663 579858 205672
rect 580172 193180 580224 193186
rect 580172 193122 580224 193128
rect 580184 192545 580212 193122
rect 580170 192536 580226 192545
rect 580170 192471 580226 192480
rect 580172 179376 580224 179382
rect 580172 179318 580224 179324
rect 580184 179217 580212 179318
rect 580170 179208 580226 179217
rect 580170 179143 580226 179152
rect 580172 167000 580224 167006
rect 580172 166942 580224 166948
rect 580184 165889 580212 166942
rect 580170 165880 580226 165889
rect 580170 165815 580226 165824
rect 580172 153196 580224 153202
rect 580172 153138 580224 153144
rect 580184 152697 580212 153138
rect 580170 152688 580226 152697
rect 580170 152623 580226 152632
rect 465724 139392 465776 139398
rect 580172 139392 580224 139398
rect 465724 139334 465776 139340
rect 580170 139360 580172 139369
rect 580224 139360 580226 139369
rect 580170 139295 580226 139304
rect 580172 126948 580224 126954
rect 580172 126890 580224 126896
rect 580184 126041 580212 126890
rect 580170 126032 580226 126041
rect 580170 125967 580226 125976
rect 579804 113144 579856 113150
rect 579804 113086 579856 113092
rect 579816 112849 579844 113086
rect 579802 112840 579858 112849
rect 579802 112775 579858 112784
rect 457444 100700 457496 100706
rect 457444 100642 457496 100648
rect 580172 100700 580224 100706
rect 580172 100642 580224 100648
rect 580184 99521 580212 100642
rect 580170 99512 580226 99521
rect 580170 99447 580226 99456
rect 486424 98796 486476 98802
rect 486424 98738 486476 98744
rect 461584 96484 461636 96490
rect 461584 96426 461636 96432
rect 454776 93560 454828 93566
rect 454776 93502 454828 93508
rect 454684 60716 454736 60722
rect 454684 60658 454736 60664
rect 454500 3800 454552 3806
rect 454500 3742 454552 3748
rect 453396 3324 453448 3330
rect 453396 3266 453448 3272
rect 454512 480 454540 3742
rect 454788 3398 454816 93502
rect 457444 90908 457496 90914
rect 457444 90850 457496 90856
rect 456892 33788 456944 33794
rect 456892 33730 456944 33736
rect 456904 16574 456932 33730
rect 456904 16546 457392 16574
rect 454776 3392 454828 3398
rect 454776 3334 454828 3340
rect 455696 3392 455748 3398
rect 455696 3334 455748 3340
rect 455708 480 455736 3334
rect 456892 3324 456944 3330
rect 456892 3266 456944 3272
rect 456904 480 456932 3266
rect 457364 3210 457392 16546
rect 457456 3398 457484 90850
rect 459560 85128 459612 85134
rect 459560 85070 459612 85076
rect 459572 16574 459600 85070
rect 459572 16546 459968 16574
rect 457444 3392 457496 3398
rect 457444 3334 457496 3340
rect 459192 3392 459244 3398
rect 459192 3334 459244 3340
rect 457364 3182 458128 3210
rect 458100 480 458128 3182
rect 459204 480 459232 3334
rect 459940 490 459968 16546
rect 461596 3942 461624 96426
rect 468484 96416 468536 96422
rect 468484 96358 468536 96364
rect 465724 95124 465776 95130
rect 465724 95066 465776 95072
rect 464344 91860 464396 91866
rect 464344 91802 464396 91808
rect 463700 85060 463752 85066
rect 463700 85002 463752 85008
rect 463712 16574 463740 85002
rect 463712 16546 464016 16574
rect 461584 3936 461636 3942
rect 461584 3878 461636 3884
rect 462780 3868 462832 3874
rect 462780 3810 462832 3816
rect 461584 3732 461636 3738
rect 461584 3674 461636 3680
rect 460216 598 460428 626
rect 460216 490 460244 598
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 459940 462 460244 490
rect 460400 480 460428 598
rect 461596 480 461624 3674
rect 462792 480 462820 3810
rect 463988 480 464016 16546
rect 464356 2990 464384 91802
rect 465172 5092 465224 5098
rect 465172 5034 465224 5040
rect 464344 2984 464396 2990
rect 464344 2926 464396 2932
rect 465184 480 465212 5034
rect 465736 3806 465764 95066
rect 467104 89548 467156 89554
rect 467104 89490 467156 89496
rect 467116 16574 467144 89490
rect 467116 16546 467236 16574
rect 467104 13184 467156 13190
rect 467104 13126 467156 13132
rect 465724 3800 465776 3806
rect 465724 3742 465776 3748
rect 467116 3482 467144 13126
rect 467208 3738 467236 16546
rect 468496 3874 468524 96358
rect 472624 96348 472676 96354
rect 472624 96290 472676 96296
rect 471244 90840 471296 90846
rect 471244 90782 471296 90788
rect 470600 13116 470652 13122
rect 470600 13058 470652 13064
rect 469864 9104 469916 9110
rect 469864 9046 469916 9052
rect 468484 3868 468536 3874
rect 468484 3810 468536 3816
rect 467196 3732 467248 3738
rect 467196 3674 467248 3680
rect 468668 3664 468720 3670
rect 468668 3606 468720 3612
rect 467116 3454 467512 3482
rect 466276 2984 466328 2990
rect 466276 2926 466328 2932
rect 466288 480 466316 2926
rect 467484 480 467512 3454
rect 468680 480 468708 3606
rect 469876 480 469904 9046
rect 470612 490 470640 13058
rect 471256 4146 471284 90782
rect 472256 5160 472308 5166
rect 472256 5102 472308 5108
rect 471244 4140 471296 4146
rect 471244 4082 471296 4088
rect 470888 598 471100 626
rect 470888 490 470916 598
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 470612 462 470916 490
rect 471072 480 471100 598
rect 472268 480 472296 5102
rect 472636 4010 472664 96290
rect 479524 96280 479576 96286
rect 479524 96222 479576 96228
rect 475384 96212 475436 96218
rect 475384 96154 475436 96160
rect 472716 89480 472768 89486
rect 472716 89422 472768 89428
rect 472624 4004 472676 4010
rect 472624 3946 472676 3952
rect 472728 3602 472756 89422
rect 473452 9036 473504 9042
rect 473452 8978 473504 8984
rect 472716 3596 472768 3602
rect 472716 3538 472768 3544
rect 473464 480 473492 8978
rect 475396 4078 475424 96154
rect 477500 83768 477552 83774
rect 477500 83710 477552 83716
rect 477512 16574 477540 83710
rect 478880 37936 478932 37942
rect 478880 37878 478932 37884
rect 477512 16546 478184 16574
rect 476948 8968 477000 8974
rect 476948 8910 477000 8916
rect 475844 4140 475896 4146
rect 475844 4082 475896 4088
rect 475384 4072 475436 4078
rect 475384 4014 475436 4020
rect 475856 3670 475884 4082
rect 475752 3664 475804 3670
rect 475752 3606 475804 3612
rect 475844 3664 475896 3670
rect 475844 3606 475896 3612
rect 474556 3596 474608 3602
rect 474556 3538 474608 3544
rect 474568 480 474596 3538
rect 475764 480 475792 3606
rect 476960 480 476988 8910
rect 478156 480 478184 16546
rect 478892 490 478920 37878
rect 479536 4146 479564 96222
rect 483020 96144 483072 96150
rect 483020 96086 483072 96092
rect 481640 90772 481692 90778
rect 481640 90714 481692 90720
rect 481652 6914 481680 90714
rect 481732 24132 481784 24138
rect 481732 24074 481784 24080
rect 481744 16574 481772 24074
rect 483032 16574 483060 96086
rect 485044 95056 485096 95062
rect 485044 94998 485096 95004
rect 481744 16546 482416 16574
rect 483032 16546 484072 16574
rect 481652 6886 481772 6914
rect 479524 4140 479576 4146
rect 479524 4082 479576 4088
rect 480536 4140 480588 4146
rect 480536 4082 480588 4088
rect 479168 598 479380 626
rect 479168 490 479196 598
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 478892 462 479196 490
rect 479352 480 479380 598
rect 480548 480 480576 4082
rect 481744 480 481772 6886
rect 482388 490 482416 16546
rect 482664 598 482876 626
rect 482664 490 482692 598
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482388 462 482692 490
rect 482848 480 482876 598
rect 484044 480 484072 16546
rect 485056 3602 485084 94998
rect 485780 84992 485832 84998
rect 485780 84934 485832 84940
rect 485792 16574 485820 84934
rect 485792 16546 486372 16574
rect 485228 3664 485280 3670
rect 485228 3606 485280 3612
rect 485044 3596 485096 3602
rect 485044 3538 485096 3544
rect 485240 480 485268 3606
rect 486344 3482 486372 16546
rect 486436 3602 486464 98738
rect 525064 98728 525116 98734
rect 525064 98670 525116 98676
rect 500960 96076 501012 96082
rect 500960 96018 501012 96024
rect 489184 94988 489236 94994
rect 489184 94930 489236 94936
rect 487620 4072 487672 4078
rect 487620 4014 487672 4020
rect 486424 3596 486476 3602
rect 486424 3538 486476 3544
rect 486344 3454 486464 3482
rect 486436 480 486464 3454
rect 487632 480 487660 4014
rect 489196 3670 489224 94930
rect 490564 90704 490616 90710
rect 490564 90646 490616 90652
rect 490012 84924 490064 84930
rect 490012 84866 490064 84872
rect 490024 6914 490052 84866
rect 489932 6886 490052 6914
rect 489184 3664 489236 3670
rect 489184 3606 489236 3612
rect 488816 3596 488868 3602
rect 488816 3538 488868 3544
rect 488828 480 488856 3538
rect 489932 480 489960 6886
rect 490576 3398 490604 90646
rect 493324 90636 493376 90642
rect 493324 90578 493376 90584
rect 492680 83700 492732 83706
rect 492680 83642 492732 83648
rect 492692 16574 492720 83642
rect 492692 16546 493088 16574
rect 491116 4004 491168 4010
rect 491116 3946 491168 3952
rect 490564 3392 490616 3398
rect 490564 3334 490616 3340
rect 491128 480 491156 3946
rect 492312 3392 492364 3398
rect 492312 3334 492364 3340
rect 492324 480 492352 3334
rect 493060 490 493088 16546
rect 493336 2990 493364 90578
rect 500224 90568 500276 90574
rect 500224 90510 500276 90516
rect 497464 89412 497516 89418
rect 497464 89354 497516 89360
rect 496820 83632 496872 83638
rect 496820 83574 496872 83580
rect 496832 16574 496860 83574
rect 496832 16546 497136 16574
rect 494704 3868 494756 3874
rect 494704 3810 494756 3816
rect 493324 2984 493376 2990
rect 493324 2926 493376 2932
rect 493336 598 493548 626
rect 493336 490 493364 598
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493060 462 493364 490
rect 493520 480 493548 598
rect 494716 480 494744 3810
rect 495900 2984 495952 2990
rect 495900 2926 495952 2932
rect 495912 480 495940 2926
rect 497108 480 497136 16546
rect 497476 3398 497504 89354
rect 499580 17264 499632 17270
rect 499580 17206 499632 17212
rect 499592 6914 499620 17206
rect 500236 16574 500264 90510
rect 500972 16574 501000 96018
rect 502984 96008 503036 96014
rect 502984 95950 503036 95956
rect 500236 16546 500356 16574
rect 500972 16546 501368 16574
rect 499592 6886 500264 6914
rect 498200 3936 498252 3942
rect 498200 3878 498252 3884
rect 497464 3392 497516 3398
rect 497464 3334 497516 3340
rect 498212 480 498240 3878
rect 499396 3392 499448 3398
rect 499396 3334 499448 3340
rect 499408 480 499436 3334
rect 500236 3074 500264 6886
rect 500328 3262 500356 16546
rect 500316 3256 500368 3262
rect 500316 3198 500368 3204
rect 500236 3046 500632 3074
rect 500604 480 500632 3046
rect 501340 490 501368 16546
rect 502996 3398 503024 95950
rect 512000 95940 512052 95946
rect 512000 95882 512052 95888
rect 507860 94920 507912 94926
rect 507860 94862 507912 94868
rect 504364 89344 504416 89350
rect 504364 89286 504416 89292
rect 504180 5024 504232 5030
rect 504180 4966 504232 4972
rect 502984 3392 503036 3398
rect 502984 3334 503036 3340
rect 502984 3256 503036 3262
rect 502984 3198 503036 3204
rect 501616 598 501828 626
rect 501616 490 501644 598
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501340 462 501644 490
rect 501800 480 501828 598
rect 502996 480 503024 3198
rect 504192 480 504220 4966
rect 504376 2990 504404 89286
rect 506480 89276 506532 89282
rect 506480 89218 506532 89224
rect 505376 3392 505428 3398
rect 505376 3334 505428 3340
rect 504364 2984 504416 2990
rect 504364 2926 504416 2932
rect 505388 480 505416 3334
rect 506492 480 506520 89218
rect 506572 21412 506624 21418
rect 506572 21354 506624 21360
rect 506584 16574 506612 21354
rect 507872 16574 507900 94862
rect 511264 90500 511316 90506
rect 511264 90442 511316 90448
rect 510620 82272 510672 82278
rect 510620 82214 510672 82220
rect 510632 16574 510660 82214
rect 506584 16546 507256 16574
rect 507872 16546 508912 16574
rect 510632 16546 511212 16574
rect 507228 490 507256 16546
rect 507504 598 507716 626
rect 507504 490 507532 598
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507228 462 507532 490
rect 507688 480 507716 598
rect 508884 480 508912 16546
rect 510068 2984 510120 2990
rect 510068 2926 510120 2932
rect 511184 2938 511212 16546
rect 511276 3058 511304 90442
rect 511264 3052 511316 3058
rect 511264 2994 511316 3000
rect 510080 480 510108 2926
rect 511184 2910 511304 2938
rect 511276 480 511304 2910
rect 512012 490 512040 95882
rect 519544 94852 519596 94858
rect 519544 94794 519596 94800
rect 518164 89208 518216 89214
rect 518164 89150 518216 89156
rect 515404 89140 515456 89146
rect 515404 89082 515456 89088
rect 514760 6248 514812 6254
rect 514760 6190 514812 6196
rect 513564 3052 513616 3058
rect 513564 2994 513616 3000
rect 512288 598 512500 626
rect 512288 490 512316 598
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512012 462 512316 490
rect 512472 480 512500 598
rect 513576 480 513604 2994
rect 514772 480 514800 6190
rect 515416 3398 515444 89082
rect 517520 18624 517572 18630
rect 517520 18566 517572 18572
rect 517532 16574 517560 18566
rect 517532 16546 517928 16574
rect 515956 3664 516008 3670
rect 515956 3606 516008 3612
rect 515404 3392 515456 3398
rect 515404 3334 515456 3340
rect 515968 480 515996 3606
rect 517152 3392 517204 3398
rect 517152 3334 517204 3340
rect 517164 480 517192 3334
rect 517900 490 517928 16546
rect 518176 3670 518204 89150
rect 519556 16574 519584 94794
rect 520280 91792 520332 91798
rect 520280 91734 520332 91740
rect 519556 16546 519676 16574
rect 519544 4956 519596 4962
rect 519544 4898 519596 4904
rect 518164 3664 518216 3670
rect 518164 3606 518216 3612
rect 518176 598 518388 626
rect 518176 490 518204 598
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 517900 462 518204 490
rect 518360 480 518388 598
rect 519556 480 519584 4898
rect 519648 3874 519676 16546
rect 519636 3868 519688 3874
rect 519636 3810 519688 3816
rect 520292 490 520320 91734
rect 522304 89072 522356 89078
rect 522304 89014 522356 89020
rect 521844 14544 521896 14550
rect 521844 14486 521896 14492
rect 520568 598 520780 626
rect 520568 490 520596 598
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520292 462 520596 490
rect 520752 480 520780 598
rect 521856 480 521884 14486
rect 522316 3398 522344 89014
rect 525076 16574 525104 98670
rect 568580 98660 568632 98666
rect 568580 98602 568632 98608
rect 525798 95976 525854 95985
rect 525798 95911 525854 95920
rect 525812 16574 525840 95911
rect 550638 95840 550694 95849
rect 550638 95775 550694 95784
rect 529940 94784 529992 94790
rect 529940 94726 529992 94732
rect 529204 90432 529256 90438
rect 529204 90374 529256 90380
rect 528560 83564 528612 83570
rect 528560 83506 528612 83512
rect 525076 16546 525196 16574
rect 525812 16546 526208 16574
rect 525064 14476 525116 14482
rect 525064 14418 525116 14424
rect 523040 4888 523092 4894
rect 523040 4830 523092 4836
rect 522304 3392 522356 3398
rect 522304 3334 522356 3340
rect 523052 480 523080 4830
rect 524236 3392 524288 3398
rect 524236 3334 524288 3340
rect 524248 480 524276 3334
rect 525076 2802 525104 14418
rect 525168 2922 525196 16546
rect 525156 2916 525208 2922
rect 525156 2858 525208 2864
rect 525076 2774 525472 2802
rect 525444 480 525472 2774
rect 526180 490 526208 16546
rect 527824 2916 527876 2922
rect 527824 2858 527876 2864
rect 526456 598 526668 626
rect 526456 490 526484 598
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526180 462 526484 490
rect 526640 480 526668 598
rect 527836 480 527864 2858
rect 528572 490 528600 83506
rect 529216 3670 529244 90374
rect 529952 16574 529980 94726
rect 532700 94716 532752 94722
rect 532700 94658 532752 94664
rect 530584 84856 530636 84862
rect 530584 84798 530636 84804
rect 529952 16546 530164 16574
rect 529112 3664 529164 3670
rect 529112 3606 529164 3612
rect 529204 3664 529256 3670
rect 529204 3606 529256 3612
rect 529124 3330 529152 3606
rect 529112 3324 529164 3330
rect 529112 3266 529164 3272
rect 528848 598 529060 626
rect 528848 490 528876 598
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528572 462 528876 490
rect 529032 480 529060 598
rect 530136 480 530164 16546
rect 530596 3398 530624 84798
rect 532712 16574 532740 94658
rect 536840 94648 536892 94654
rect 536840 94590 536892 94596
rect 536104 87916 536156 87922
rect 536104 87858 536156 87864
rect 532712 16546 533752 16574
rect 531320 3664 531372 3670
rect 531320 3606 531372 3612
rect 530584 3392 530636 3398
rect 530584 3334 530636 3340
rect 531332 480 531360 3606
rect 532516 3392 532568 3398
rect 532516 3334 532568 3340
rect 532528 480 532556 3334
rect 533724 480 533752 16546
rect 536012 6180 536064 6186
rect 536012 6122 536064 6128
rect 534908 3324 534960 3330
rect 534908 3266 534960 3272
rect 534920 480 534948 3266
rect 536024 3074 536052 6122
rect 536116 3670 536144 87858
rect 536852 16574 536880 94590
rect 543740 94580 543792 94586
rect 543740 94522 543792 94528
rect 543004 93492 543056 93498
rect 543004 93434 543056 93440
rect 538220 87848 538272 87854
rect 538220 87790 538272 87796
rect 538232 16574 538260 87790
rect 540244 87780 540296 87786
rect 540244 87722 540296 87728
rect 539692 26920 539744 26926
rect 539692 26862 539744 26868
rect 536852 16546 537248 16574
rect 538232 16546 538444 16574
rect 536104 3664 536156 3670
rect 536104 3606 536156 3612
rect 536024 3046 536144 3074
rect 536116 480 536144 3046
rect 537220 480 537248 16546
rect 538416 480 538444 16546
rect 539704 6914 539732 26862
rect 539612 6886 539732 6914
rect 539612 480 539640 6886
rect 540256 3398 540284 87722
rect 542360 83496 542412 83502
rect 542360 83438 542412 83444
rect 542372 16574 542400 83438
rect 542372 16546 542768 16574
rect 540796 3868 540848 3874
rect 540796 3810 540848 3816
rect 540244 3392 540296 3398
rect 540244 3334 540296 3340
rect 540808 480 540836 3810
rect 541992 3392 542044 3398
rect 541992 3334 542044 3340
rect 542004 480 542032 3334
rect 542740 490 542768 16546
rect 543016 2990 543044 93434
rect 543752 16574 543780 94522
rect 547972 89004 548024 89010
rect 547972 88946 548024 88952
rect 547144 87712 547196 87718
rect 547144 87654 547196 87660
rect 546500 82204 546552 82210
rect 546500 82146 546552 82152
rect 546512 16574 546540 82146
rect 543752 16546 544424 16574
rect 546512 16546 546724 16574
rect 543004 2984 543056 2990
rect 543004 2926 543056 2932
rect 543016 598 543228 626
rect 543016 490 543044 598
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 542740 462 543044 490
rect 543200 480 543228 598
rect 544396 480 544424 16546
rect 545488 2984 545540 2990
rect 545488 2926 545540 2932
rect 545500 480 545528 2926
rect 546696 480 546724 16546
rect 547156 3874 547184 87654
rect 547984 16574 548012 88946
rect 548524 22772 548576 22778
rect 548524 22714 548576 22720
rect 547984 16546 548472 16574
rect 547144 3868 547196 3874
rect 547144 3810 547196 3816
rect 547880 3596 547932 3602
rect 547880 3538 547932 3544
rect 547892 480 547920 3538
rect 548444 626 548472 16546
rect 548536 3330 548564 22714
rect 550652 16574 550680 95775
rect 565084 94512 565136 94518
rect 565084 94454 565136 94460
rect 554780 93424 554832 93430
rect 554780 93366 554832 93372
rect 553400 82136 553452 82142
rect 553400 82078 553452 82084
rect 553412 16574 553440 82078
rect 554792 16574 554820 93366
rect 557540 93356 557592 93362
rect 557540 93298 557592 93304
rect 556804 90364 556856 90370
rect 556804 90306 556856 90312
rect 556252 28280 556304 28286
rect 556252 28222 556304 28228
rect 556264 16574 556292 28222
rect 550652 16546 551048 16574
rect 553412 16546 553808 16574
rect 554792 16546 555004 16574
rect 556264 16546 556752 16574
rect 548524 3324 548576 3330
rect 548524 3266 548576 3272
rect 550272 3324 550324 3330
rect 550272 3266 550324 3272
rect 548444 598 548656 626
rect 548628 490 548656 598
rect 548904 598 549116 626
rect 548904 490 548932 598
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 548628 462 548932 490
rect 549088 480 549116 598
rect 550284 480 550312 3266
rect 551020 490 551048 16546
rect 552664 3868 552716 3874
rect 552664 3810 552716 3816
rect 551296 598 551508 626
rect 551296 490 551324 598
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551020 462 551324 490
rect 551480 480 551508 598
rect 552676 480 552704 3810
rect 553780 480 553808 16546
rect 554976 480 555004 16546
rect 556160 3664 556212 3670
rect 556160 3606 556212 3612
rect 556172 480 556200 3606
rect 556724 626 556752 16546
rect 556816 3262 556844 90306
rect 557552 16574 557580 93298
rect 561680 93288 561732 93294
rect 561680 93230 561732 93236
rect 560944 87644 560996 87650
rect 560944 87586 560996 87592
rect 557552 16546 558592 16574
rect 556804 3256 556856 3262
rect 556804 3198 556856 3204
rect 556724 598 556936 626
rect 556908 490 556936 598
rect 557184 598 557396 626
rect 557184 490 557212 598
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 556908 462 557212 490
rect 557368 480 557396 598
rect 558564 480 558592 16546
rect 560852 4820 560904 4826
rect 560852 4762 560904 4768
rect 559748 3256 559800 3262
rect 559748 3198 559800 3204
rect 559760 480 559788 3198
rect 560864 480 560892 4762
rect 560956 3602 560984 87586
rect 561692 16574 561720 93230
rect 564532 25560 564584 25566
rect 564532 25502 564584 25508
rect 561692 16546 562088 16574
rect 560944 3596 560996 3602
rect 560944 3538 560996 3544
rect 562060 480 562088 16546
rect 564544 6914 564572 25502
rect 564452 6886 564572 6914
rect 563244 3596 563296 3602
rect 563244 3538 563296 3544
rect 563256 480 563284 3538
rect 564452 480 564480 6886
rect 565096 3602 565124 94454
rect 566464 86352 566516 86358
rect 566464 86294 566516 86300
rect 565820 86284 565872 86290
rect 565820 86226 565872 86232
rect 565832 6914 565860 86226
rect 566476 16574 566504 86294
rect 568592 16574 568620 98602
rect 580262 97200 580318 97209
rect 580262 97135 580318 97144
rect 572812 93220 572864 93226
rect 572812 93162 572864 93168
rect 571340 80708 571392 80714
rect 571340 80650 571392 80656
rect 571352 16574 571380 80650
rect 566476 16546 566596 16574
rect 568592 16546 568712 16574
rect 571352 16546 571564 16574
rect 565832 6886 566504 6914
rect 565636 3800 565688 3806
rect 565636 3742 565688 3748
rect 565084 3596 565136 3602
rect 565084 3538 565136 3544
rect 565648 480 565676 3742
rect 566476 3482 566504 6886
rect 566568 4146 566596 16546
rect 566556 4140 566608 4146
rect 566556 4082 566608 4088
rect 568028 4140 568080 4146
rect 568028 4082 568080 4088
rect 566476 3454 566872 3482
rect 566844 480 566872 3454
rect 568040 480 568068 4082
rect 568684 490 568712 16546
rect 570328 3596 570380 3602
rect 570328 3538 570380 3544
rect 568960 598 569172 626
rect 568960 490 568988 598
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 568684 462 568988 490
rect 569144 480 569172 598
rect 570340 480 570368 3538
rect 571536 480 571564 16546
rect 572824 6914 572852 93162
rect 575480 93152 575532 93158
rect 575480 93094 575532 93100
rect 575492 16574 575520 93094
rect 580172 86964 580224 86970
rect 580172 86906 580224 86912
rect 580184 86193 580212 86906
rect 580170 86184 580226 86193
rect 580170 86119 580226 86128
rect 579988 73160 580040 73166
rect 579988 73102 580040 73108
rect 580000 73001 580028 73102
rect 579986 72992 580042 73001
rect 579986 72927 580042 72936
rect 580172 60716 580224 60722
rect 580172 60658 580224 60664
rect 580184 59673 580212 60658
rect 580170 59664 580226 59673
rect 580170 59599 580226 59608
rect 580170 33144 580226 33153
rect 580170 33079 580172 33088
rect 580224 33079 580226 33088
rect 580172 33050 580224 33056
rect 580172 20664 580224 20670
rect 580172 20606 580224 20612
rect 580184 19825 580212 20606
rect 580170 19816 580226 19825
rect 580170 19751 580226 19760
rect 575492 16546 575888 16574
rect 575112 15972 575164 15978
rect 575112 15914 575164 15920
rect 572732 6886 572852 6914
rect 572732 480 572760 6886
rect 573916 3732 573968 3738
rect 573916 3674 573968 3680
rect 573928 480 573956 3674
rect 575124 480 575152 15914
rect 575860 490 575888 16546
rect 578608 15904 578660 15910
rect 578608 15846 578660 15852
rect 576952 10328 577004 10334
rect 576952 10270 577004 10276
rect 576136 598 576348 626
rect 576136 490 576164 598
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 575860 462 576164 490
rect 576320 480 576348 598
rect 576964 490 576992 10270
rect 577240 598 577452 626
rect 577240 490 577268 598
rect 576278 -960 576390 480
rect 576964 462 577268 490
rect 577424 480 577452 598
rect 578620 480 578648 15846
rect 580276 3534 580304 97135
rect 582392 6633 582420 300834
rect 582484 46345 582512 300902
rect 582470 46336 582526 46345
rect 582470 46271 582526 46280
rect 582378 6624 582434 6633
rect 582378 6559 582434 6568
rect 580264 3528 580316 3534
rect 580264 3470 580316 3476
rect 582196 3528 582248 3534
rect 582196 3470 582248 3476
rect 581000 3460 581052 3466
rect 581000 3402 581052 3408
rect 581012 480 581040 3402
rect 582208 480 582236 3470
rect 583392 3392 583444 3398
rect 583392 3334 583444 3340
rect 583404 480 583432 3334
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 3422 671200 3478 671256
rect 3422 658144 3478 658200
rect 3422 632068 3424 632088
rect 3424 632068 3476 632088
rect 3476 632068 3478 632088
rect 3422 632032 3478 632068
rect 3146 619112 3202 619168
rect 3238 606056 3294 606112
rect 3330 579944 3386 580000
rect 3422 566888 3478 566944
rect 3422 553832 3478 553888
rect 3422 527856 3478 527912
rect 3422 514820 3478 514856
rect 3422 514800 3424 514820
rect 3424 514800 3476 514820
rect 3476 514800 3478 514820
rect 3054 501744 3110 501800
rect 3422 475632 3478 475688
rect 3238 462576 3294 462632
rect 3146 449520 3202 449576
rect 3422 423544 3478 423600
rect 3146 410488 3202 410544
rect 3422 397468 3424 397488
rect 3424 397468 3476 397488
rect 3476 397468 3478 397488
rect 3422 397432 3478 397468
rect 3422 371320 3478 371376
rect 3146 358400 3202 358456
rect 3330 345344 3386 345400
rect 3422 319232 3478 319288
rect 3238 306176 3294 306232
rect 2870 293120 2926 293176
rect 3238 267144 3294 267200
rect 3330 214920 3386 214976
rect 3054 201864 3110 201920
rect 3606 254088 3662 254144
rect 3514 241032 3570 241088
rect 3422 188808 3478 188864
rect 3238 162832 3294 162888
rect 3422 149776 3478 149832
rect 3238 136720 3294 136776
rect 3422 110608 3478 110664
rect 3422 97552 3478 97608
rect 3146 84632 3202 84688
rect 2778 71612 2780 71632
rect 2780 71612 2832 71632
rect 2832 71612 2834 71632
rect 2778 71576 2834 71612
rect 3054 58520 3110 58576
rect 3422 45500 3424 45520
rect 3424 45500 3476 45520
rect 3476 45500 3478 45520
rect 3422 45464 3478 45500
rect 3146 32408 3202 32464
rect 3422 19352 3478 19408
rect 3422 6432 3478 6488
rect 32402 97144 32458 97200
rect 39302 97416 39358 97472
rect 38566 97280 38622 97336
rect 50342 97552 50398 97608
rect 171690 174800 171746 174856
rect 171506 173576 171562 173632
rect 171782 170448 171838 170504
rect 171874 168136 171930 168192
rect 171966 164464 172022 164520
rect 172426 189896 172482 189952
rect 172426 188672 172482 188728
rect 172426 187312 172482 187368
rect 172426 186088 172482 186144
rect 172426 184764 172428 184784
rect 172428 184764 172480 184784
rect 172480 184764 172482 184784
rect 172426 184728 172482 184764
rect 172334 184320 172390 184376
rect 172426 182960 172482 183016
rect 172426 181736 172482 181792
rect 172058 163512 172114 163568
rect 171782 162288 171838 162344
rect 171598 153720 171654 153776
rect 171230 153176 171286 153232
rect 171506 149912 171562 149968
rect 171690 149404 171692 149424
rect 171692 149404 171744 149424
rect 171744 149404 171746 149424
rect 171690 149368 171746 149404
rect 171690 148280 171746 148336
rect 171690 147736 171746 147792
rect 171874 150492 171876 150512
rect 171876 150492 171928 150512
rect 171928 150492 171930 150512
rect 171874 150456 171930 150492
rect 171874 148860 171876 148880
rect 171876 148860 171928 148880
rect 171928 148860 171930 148880
rect 171874 148824 171930 148860
rect 171874 146648 171930 146704
rect 172426 180548 172428 180568
rect 172428 180548 172480 180568
rect 172480 180548 172482 180568
rect 172426 180512 172482 180548
rect 172426 179188 172428 179208
rect 172428 179188 172480 179208
rect 172480 179188 172482 179208
rect 172426 179152 172482 179188
rect 172334 177948 172390 177984
rect 172334 177928 172336 177948
rect 172336 177928 172388 177948
rect 172388 177928 172390 177948
rect 172426 177384 172482 177440
rect 172426 176024 172482 176080
rect 172426 172352 172482 172408
rect 172426 171028 172428 171048
rect 172428 171028 172480 171048
rect 172480 171028 172482 171048
rect 172426 170992 172482 171028
rect 172426 169088 172482 169144
rect 172426 166640 172482 166696
rect 172426 164056 172482 164112
rect 172242 160928 172298 160984
rect 172426 152632 172482 152688
rect 172334 152088 172390 152144
rect 172426 151580 172428 151600
rect 172428 151580 172480 151600
rect 172480 151580 172482 151600
rect 172426 151544 172482 151580
rect 172334 151000 172390 151056
rect 172426 147192 172482 147248
rect 172242 146124 172298 146160
rect 172242 146104 172244 146124
rect 172244 146104 172296 146124
rect 172296 146104 172298 146124
rect 172426 145560 172482 145616
rect 172334 145016 172390 145072
rect 172426 144472 172482 144528
rect 172150 144064 172206 144120
rect 171782 143520 171838 143576
rect 171874 142976 171930 143032
rect 171690 142432 171746 142488
rect 171506 141888 171562 141944
rect 171782 141344 171838 141400
rect 172426 140800 172482 140856
rect 171690 140256 171746 140312
rect 171690 139748 171692 139768
rect 171692 139748 171744 139768
rect 171744 139748 171746 139768
rect 171690 139712 171746 139748
rect 171598 138624 171654 138680
rect 171506 138080 171562 138136
rect 172058 137536 172114 137592
rect 172426 139168 172482 139224
rect 172334 136992 172390 137048
rect 172426 136448 172482 136504
rect 172242 135904 172298 135960
rect 171690 135360 171746 135416
rect 172242 134272 172298 134328
rect 171230 133864 171286 133920
rect 172426 134816 172482 134872
rect 172426 133320 172482 133376
rect 172334 132776 172390 132832
rect 171138 132232 171194 132288
rect 172426 131724 172428 131744
rect 172428 131724 172480 131744
rect 172480 131724 172482 131744
rect 172426 131688 172482 131724
rect 171506 131144 171562 131200
rect 172334 130600 172390 130656
rect 171874 130076 171930 130112
rect 171874 130056 171876 130076
rect 171876 130056 171928 130076
rect 171928 130056 171930 130076
rect 172058 128968 172114 129024
rect 171874 128424 171930 128480
rect 171782 127336 171838 127392
rect 171690 124616 171746 124672
rect 171966 127880 172022 127936
rect 172426 129512 172482 129568
rect 172242 126792 172298 126848
rect 172334 126248 172390 126304
rect 172426 125740 172428 125760
rect 172428 125740 172480 125760
rect 172480 125740 172482 125760
rect 172426 125704 172482 125740
rect 172426 125160 172482 125216
rect 172150 124228 172206 124264
rect 172150 124208 172152 124228
rect 172152 124208 172204 124228
rect 172204 124208 172206 124228
rect 198554 298832 198610 298888
rect 197910 294480 197966 294536
rect 198094 292304 198150 292360
rect 197358 290128 197414 290184
rect 197634 287952 197690 288008
rect 197358 285776 197414 285832
rect 197358 283600 197414 283656
rect 197358 281424 197414 281480
rect 197358 279248 197414 279304
rect 197542 277072 197598 277128
rect 198370 274916 198426 274952
rect 198370 274896 198372 274916
rect 198372 274896 198424 274916
rect 198424 274896 198426 274916
rect 197358 272720 197414 272776
rect 197358 270564 197414 270600
rect 197358 270544 197360 270564
rect 197360 270544 197412 270564
rect 197412 270544 197414 270564
rect 197726 268368 197782 268424
rect 197358 266192 197414 266248
rect 197910 264016 197966 264072
rect 198646 261860 198702 261896
rect 198646 261840 198648 261860
rect 198648 261840 198700 261860
rect 198700 261840 198702 261860
rect 197726 259664 197782 259720
rect 198094 257488 198150 257544
rect 197358 255332 197414 255368
rect 197358 255312 197360 255332
rect 197360 255312 197412 255332
rect 197412 255312 197414 255332
rect 197358 253136 197414 253192
rect 198002 250960 198058 251016
rect 197358 244432 197414 244488
rect 197726 242256 197782 242312
rect 197358 240080 197414 240136
rect 197358 237904 197414 237960
rect 197542 235728 197598 235784
rect 197634 231376 197690 231432
rect 197358 229200 197414 229256
rect 197358 222672 197414 222728
rect 197542 220496 197598 220552
rect 197910 216144 197966 216200
rect 197358 213988 197414 214024
rect 197358 213968 197360 213988
rect 197360 213968 197412 213988
rect 197412 213968 197414 213988
rect 197726 211792 197782 211848
rect 197358 209616 197414 209672
rect 197358 207440 197414 207496
rect 197542 205264 197598 205320
rect 197358 203088 197414 203144
rect 197358 200912 197414 200968
rect 197358 198756 197414 198792
rect 197358 198736 197360 198756
rect 197360 198736 197412 198756
rect 197412 198736 197414 198756
rect 197358 196560 197414 196616
rect 197358 192208 197414 192264
rect 197542 190032 197598 190088
rect 197358 187856 197414 187912
rect 197358 185680 197414 185736
rect 197358 181328 197414 181384
rect 197542 179152 197598 179208
rect 197358 176976 197414 177032
rect 197634 174800 197690 174856
rect 197358 172624 197414 172680
rect 198186 248784 198242 248840
rect 198094 246608 198150 246664
rect 197358 170448 197414 170504
rect 198186 233552 198242 233608
rect 198738 227024 198794 227080
rect 198278 224848 198334 224904
rect 198462 218320 198518 218376
rect 198646 194404 198702 194440
rect 198646 194384 198648 194404
rect 198648 194384 198700 194404
rect 198700 194384 198702 194404
rect 198186 183504 198242 183560
rect 197910 168272 197966 168328
rect 198002 163920 198058 163976
rect 197358 161744 197414 161800
rect 197358 159568 197414 159624
rect 197358 157412 197414 157448
rect 197358 157392 197360 157412
rect 197360 157392 197412 157412
rect 197412 157392 197414 157412
rect 198462 166116 198518 166152
rect 198462 166096 198464 166116
rect 198464 166096 198516 166116
rect 198516 166096 198518 166116
rect 198278 155216 198334 155272
rect 198094 153040 198150 153096
rect 197726 146532 197782 146568
rect 197726 146512 197728 146532
rect 197728 146512 197780 146532
rect 197780 146512 197782 146532
rect 197358 144336 197414 144392
rect 197358 142180 197414 142216
rect 197358 142160 197360 142180
rect 197360 142160 197412 142180
rect 197412 142160 197414 142180
rect 198370 150864 198426 150920
rect 198278 148688 198334 148744
rect 198278 139984 198334 140040
rect 197542 137808 197598 137864
rect 198094 135632 198150 135688
rect 197542 133456 197598 133512
rect 197910 131280 197966 131336
rect 197358 129104 197414 129160
rect 197358 126948 197414 126984
rect 197358 126928 197360 126948
rect 197360 126928 197412 126948
rect 197412 126928 197414 126948
rect 198554 124752 198610 124808
rect 217046 299512 217102 299568
rect 218058 299512 218114 299568
rect 218058 299376 218114 299432
rect 218794 299376 218850 299432
rect 217138 299276 217140 299296
rect 217140 299276 217192 299296
rect 217192 299276 217194 299296
rect 217138 299240 217194 299276
rect 219898 299276 219900 299296
rect 219900 299276 219952 299296
rect 219952 299276 219954 299296
rect 219898 299240 219954 299276
rect 199842 296656 199898 296712
rect 198002 122576 198058 122632
rect 197542 120400 197598 120456
rect 197542 116048 197598 116104
rect 197358 113872 197414 113928
rect 197358 111732 197360 111752
rect 197360 111732 197412 111752
rect 197412 111732 197414 111752
rect 197358 111696 197414 111732
rect 198094 118224 198150 118280
rect 198002 109520 198058 109576
rect 198554 107344 198610 107400
rect 197542 105168 197598 105224
rect 197910 102992 197966 103048
rect 197542 100952 197598 101008
rect 371698 369688 371754 369744
rect 371606 368620 371662 368656
rect 371606 368600 371608 368620
rect 371608 368600 371660 368620
rect 371660 368600 371662 368620
rect 371882 369144 371938 369200
rect 371606 368056 371662 368112
rect 371514 367512 371570 367568
rect 371606 366968 371662 367024
rect 371238 365880 371294 365936
rect 371606 365336 371662 365392
rect 371238 364792 371294 364848
rect 371698 364248 371754 364304
rect 371606 363724 371662 363760
rect 371606 363704 371608 363724
rect 371608 363704 371660 363724
rect 371660 363704 371662 363724
rect 371422 363160 371478 363216
rect 371422 362072 371478 362128
rect 371514 361528 371570 361584
rect 371698 360984 371754 361040
rect 371606 360460 371662 360496
rect 371606 360440 371608 360460
rect 371608 360440 371660 360460
rect 371660 360440 371662 360460
rect 371330 360032 371386 360088
rect 372526 366424 372582 366480
rect 372066 359488 372122 359544
rect 371514 358400 371570 358456
rect 371422 357856 371478 357912
rect 371238 357312 371294 357368
rect 371330 356768 371386 356824
rect 371422 356224 371478 356280
rect 371698 355680 371754 355736
rect 371238 355136 371294 355192
rect 371514 354592 371570 354648
rect 371698 354048 371754 354104
rect 372250 358944 372306 359000
rect 371330 351872 371386 351928
rect 370318 349288 370374 349344
rect 369306 348472 369362 348528
rect 370042 346840 370098 346896
rect 369950 345208 370006 345264
rect 302790 298308 302846 298344
rect 302790 298288 302792 298308
rect 302792 298288 302844 298308
rect 302844 298288 302846 298308
rect 302422 295160 302478 295216
rect 302330 291896 302386 291952
rect 302790 285676 302792 285696
rect 302792 285676 302844 285696
rect 302844 285676 302846 285696
rect 302790 285640 302846 285676
rect 302422 282376 302478 282432
rect 302606 279248 302662 279304
rect 302974 288768 303030 288824
rect 302882 272856 302938 272912
rect 302330 269728 302386 269784
rect 302422 266600 302478 266656
rect 303066 276120 303122 276176
rect 302514 263336 302570 263392
rect 302790 260208 302846 260264
rect 302790 257080 302846 257136
rect 302882 253816 302938 253872
rect 303158 250688 303214 250744
rect 303066 247560 303122 247616
rect 302974 244296 303030 244352
rect 302790 241168 302846 241224
rect 302882 231648 302938 231704
rect 302790 228384 302846 228440
rect 302790 225256 302846 225312
rect 303158 238040 303214 238096
rect 303250 234776 303306 234832
rect 302790 222148 302846 222184
rect 302790 222128 302792 222148
rect 302792 222128 302844 222148
rect 302844 222128 302846 222148
rect 302790 218864 302846 218920
rect 302790 215736 302846 215792
rect 302790 212608 302846 212664
rect 302882 209344 302938 209400
rect 302330 206216 302386 206272
rect 302790 203088 302846 203144
rect 302514 199824 302570 199880
rect 302698 196696 302754 196752
rect 302422 193568 302478 193624
rect 302698 187176 302754 187232
rect 302790 184048 302846 184104
rect 303066 190304 303122 190360
rect 302974 180784 303030 180840
rect 302882 177656 302938 177712
rect 302238 174528 302294 174584
rect 302790 171264 302846 171320
rect 302698 168136 302754 168192
rect 302606 164872 302662 164928
rect 302974 161744 303030 161800
rect 302790 158616 302846 158672
rect 302882 155352 302938 155408
rect 302790 152224 302846 152280
rect 302790 149096 302846 149152
rect 302790 145832 302846 145888
rect 302790 142704 302846 142760
rect 302882 139576 302938 139632
rect 302790 130056 302846 130112
rect 302606 126792 302662 126848
rect 302974 136312 303030 136368
rect 303066 133184 303122 133240
rect 302698 123664 302754 123720
rect 302790 120536 302846 120592
rect 302790 117272 302846 117328
rect 302330 111016 302386 111072
rect 302790 107752 302846 107808
rect 302974 114144 303030 114200
rect 302882 104624 302938 104680
rect 302790 101496 302846 101552
rect 203522 97416 203578 97472
rect 204902 97144 204958 97200
rect 206098 97552 206154 97608
rect 206558 97280 206614 97336
rect 274178 97044 274180 97064
rect 274180 97044 274232 97064
rect 274232 97044 274234 97064
rect 274178 97008 274234 97044
rect 278686 97008 278742 97064
rect 279330 97416 279386 97472
rect 280526 97280 280582 97336
rect 282642 97144 282698 97200
rect 283010 97144 283066 97200
rect 289818 95920 289874 95976
rect 294050 95784 294106 95840
rect 299110 97144 299166 97200
rect 353942 266192 353998 266248
rect 356702 266056 356758 266112
rect 362866 337728 362922 337784
rect 364890 337728 364946 337784
rect 369398 297336 369454 297392
rect 369306 296792 369362 296848
rect 369306 296248 369362 296304
rect 369306 277072 369362 277128
rect 362866 267824 362922 267880
rect 364890 266228 364892 266248
rect 364892 266228 364944 266248
rect 364944 266228 364946 266248
rect 364890 266192 364946 266228
rect 370226 295568 370282 295624
rect 370134 295024 370190 295080
rect 370042 274896 370098 274952
rect 369950 273808 370006 273864
rect 370502 347656 370558 347712
rect 370410 340176 370466 340232
rect 370318 277344 370374 277400
rect 370594 346024 370650 346080
rect 370502 275712 370558 275768
rect 371238 297744 371294 297800
rect 371238 297200 371294 297256
rect 371238 296676 371294 296712
rect 371238 296656 371240 296676
rect 371240 296656 371292 296676
rect 371292 296656 371294 296676
rect 371238 296112 371294 296168
rect 371238 293972 371240 293992
rect 371240 293972 371292 293992
rect 371292 293972 371294 293992
rect 371238 293936 371294 293972
rect 371238 293392 371294 293448
rect 371238 292884 371240 292904
rect 371240 292884 371292 292904
rect 371292 292884 371294 292904
rect 371238 292848 371294 292884
rect 371238 291760 371294 291816
rect 371238 291236 371294 291272
rect 371238 291216 371240 291236
rect 371240 291216 371292 291236
rect 371292 291216 371294 291236
rect 371238 290128 371294 290184
rect 371238 289060 371294 289096
rect 371238 289040 371240 289060
rect 371240 289040 371292 289060
rect 371292 289040 371294 289060
rect 371238 287544 371294 287600
rect 371882 350240 371938 350296
rect 371606 348220 371662 348256
rect 371606 348200 371608 348220
rect 371608 348200 371660 348220
rect 371660 348200 371662 348220
rect 371790 343848 371846 343904
rect 371422 343304 371478 343360
rect 371330 285912 371386 285968
rect 371238 279928 371294 279984
rect 370686 275168 370742 275224
rect 370594 274080 370650 274136
rect 370410 268232 370466 268288
rect 369306 220632 369362 220688
rect 369398 220496 369454 220552
rect 369858 220088 369914 220144
rect 369858 219000 369914 219056
rect 369950 218884 370006 218920
rect 369950 218864 369952 218884
rect 369952 218864 370004 218884
rect 370004 218864 370006 218884
rect 370042 218456 370098 218512
rect 370502 221856 370558 221912
rect 370410 221312 370466 221368
rect 370410 217504 370466 217560
rect 370318 216980 370374 217016
rect 370318 216960 370320 216980
rect 370320 216960 370372 216980
rect 370372 216960 370374 216980
rect 370226 212200 370282 212256
rect 370134 210024 370190 210080
rect 369858 209208 369914 209264
rect 369306 205164 369308 205184
rect 369308 205164 369360 205184
rect 369360 205164 369362 205184
rect 369306 205128 369362 205164
rect 364522 196016 364578 196072
rect 369950 202952 370006 203008
rect 362866 194520 362922 194576
rect 364890 194520 364946 194576
rect 369306 152904 369362 152960
rect 370042 201864 370098 201920
rect 370502 208936 370558 208992
rect 370778 274080 370834 274136
rect 370686 203088 370742 203144
rect 371054 273536 371110 273592
rect 371514 341672 371570 341728
rect 371422 271632 371478 271688
rect 371698 341128 371754 341184
rect 371606 340584 371662 340640
rect 371606 276256 371662 276312
rect 372158 349832 372214 349888
rect 371974 344936 372030 344992
rect 371882 286456 371938 286512
rect 371882 285368 371938 285424
rect 371882 284824 371938 284880
rect 371882 284316 371884 284336
rect 371884 284316 371936 284336
rect 371936 284316 371938 284336
rect 371882 284280 371938 284316
rect 371882 283736 371938 283792
rect 371882 283212 371938 283248
rect 371882 283192 371884 283212
rect 371884 283192 371936 283212
rect 371936 283192 371938 283212
rect 371882 282684 371884 282704
rect 371884 282684 371936 282704
rect 371936 282684 371938 282704
rect 371882 282648 371938 282684
rect 371882 282140 371884 282160
rect 371884 282140 371936 282160
rect 371936 282140 371938 282160
rect 371882 282104 371938 282140
rect 372066 342760 372122 342816
rect 371974 272992 372030 273048
rect 371790 271904 371846 271960
rect 371882 271632 371938 271688
rect 371238 269184 371294 269240
rect 370962 211656 371018 211712
rect 370870 208392 370926 208448
rect 370778 202000 370834 202056
rect 370594 196152 370650 196208
rect 370778 196152 370834 196208
rect 370502 195236 370504 195256
rect 370504 195236 370556 195256
rect 370556 195236 370558 195256
rect 370502 195200 370558 195236
rect 369398 135088 369454 135144
rect 369306 132368 369362 132424
rect 369858 134544 369914 134600
rect 370134 135904 370190 135960
rect 370226 135360 370282 135416
rect 370042 134000 370098 134056
rect 369950 133592 370006 133648
rect 370318 132776 370374 132832
rect 369490 131960 369546 132016
rect 369306 131416 369362 131472
rect 370226 130636 370228 130656
rect 370228 130636 370280 130656
rect 370280 130636 370282 130656
rect 370226 130600 370282 130636
rect 369950 129784 370006 129840
rect 369858 129124 369914 129160
rect 369858 129104 369860 129124
rect 369860 129104 369912 129124
rect 369912 129104 369914 129124
rect 370042 128560 370098 128616
rect 370134 127336 370190 127392
rect 369950 124752 370006 124808
rect 369858 124344 369914 124400
rect 362774 123936 362830 123992
rect 365166 123936 365222 123992
rect 370502 130056 370558 130112
rect 370318 129004 370320 129024
rect 370320 129004 370372 129024
rect 370372 129004 370374 129024
rect 370318 128968 370374 129004
rect 370410 126248 370466 126304
rect 370594 125704 370650 125760
rect 370502 124752 370558 124808
rect 371606 270272 371662 270328
rect 371514 269728 371570 269784
rect 371422 222400 371478 222456
rect 371422 213832 371478 213888
rect 371422 211656 371478 211712
rect 371422 205264 371478 205320
rect 371422 204040 371478 204096
rect 371422 201320 371478 201376
rect 371330 199824 371386 199880
rect 371330 198872 371386 198928
rect 371330 197104 371386 197160
rect 371146 196052 371148 196072
rect 371148 196052 371200 196072
rect 371200 196052 371202 196072
rect 371146 196016 371202 196052
rect 371238 185544 371294 185600
rect 370870 175616 370926 175672
rect 371146 162716 371202 162752
rect 371146 162696 371148 162716
rect 371148 162696 371200 162716
rect 371200 162696 371202 162716
rect 371238 147192 371294 147248
rect 371238 146684 371240 146704
rect 371240 146684 371292 146704
rect 371292 146684 371294 146704
rect 371238 146648 371294 146684
rect 371238 142432 371294 142488
rect 371238 140800 371294 140856
rect 371238 127880 371294 127936
rect 370778 124208 370834 124264
rect 371606 225664 371662 225720
rect 371606 225120 371662 225176
rect 371606 224576 371662 224632
rect 371606 223508 371662 223544
rect 371606 223488 371608 223508
rect 371608 223488 371660 223508
rect 371660 223488 371662 223508
rect 371606 222944 371662 223000
rect 371606 216008 371662 216064
rect 371606 215464 371662 215520
rect 371698 214920 371754 214976
rect 371606 214376 371662 214432
rect 371606 213288 371662 213344
rect 371698 212744 371754 212800
rect 371698 207848 371754 207904
rect 371606 206252 371608 206272
rect 371608 206252 371660 206272
rect 371660 206252 371662 206272
rect 371606 206216 371662 206252
rect 371698 205828 371754 205864
rect 371698 205808 371700 205828
rect 371700 205808 371752 205828
rect 371752 205808 371754 205828
rect 371606 201456 371662 201512
rect 371606 198192 371662 198248
rect 371514 152632 371570 152688
rect 371514 150456 371570 150512
rect 371514 149368 371570 149424
rect 371514 145560 371570 145616
rect 371514 144064 371570 144120
rect 371514 141344 371570 141400
rect 371514 138080 371570 138136
rect 371790 201320 371846 201376
rect 372250 344392 372306 344448
rect 372158 277888 372214 277944
rect 372066 270816 372122 270872
rect 372434 342216 372490 342272
rect 372342 294480 372398 294536
rect 372342 292304 372398 292360
rect 372342 290672 372398 290728
rect 372342 289584 372398 289640
rect 372342 288088 372398 288144
rect 372342 278296 372398 278352
rect 372250 272448 372306 272504
rect 372158 268640 372214 268696
rect 372802 362616 372858 362672
rect 372710 346568 372766 346624
rect 372526 287000 372582 287056
rect 372526 279928 372582 279984
rect 372434 270272 372490 270328
rect 372342 269728 372398 269784
rect 371882 199280 371938 199336
rect 371790 198736 371846 198792
rect 371698 153720 371754 153776
rect 371698 153176 371754 153232
rect 371698 152088 371754 152144
rect 371698 151544 371754 151600
rect 371698 151036 371700 151056
rect 371700 151036 371752 151056
rect 371752 151036 371754 151056
rect 371698 151000 371754 151036
rect 371698 149912 371754 149968
rect 371698 148824 371754 148880
rect 371698 148280 371754 148336
rect 371698 147736 371754 147792
rect 371698 146124 371754 146160
rect 371698 146104 371700 146124
rect 371700 146104 371752 146124
rect 371752 146104 371754 146124
rect 371698 145052 371700 145072
rect 371700 145052 371752 145072
rect 371752 145052 371754 145072
rect 371698 145016 371754 145052
rect 371698 144508 371700 144528
rect 371700 144508 371752 144528
rect 371752 144508 371754 144528
rect 371698 144472 371754 144508
rect 371698 142976 371754 143032
rect 371698 141924 371700 141944
rect 371700 141924 371752 141944
rect 371752 141924 371754 141944
rect 371698 141888 371754 141924
rect 371698 140256 371754 140312
rect 371698 139204 371700 139224
rect 371700 139204 371752 139224
rect 371752 139204 371754 139224
rect 371698 139168 371754 139204
rect 371698 138624 371754 138680
rect 372066 216436 372122 216472
rect 372066 216416 372068 216436
rect 372068 216416 372120 216436
rect 372120 216416 372122 216436
rect 372066 204212 372068 204232
rect 372068 204212 372120 204232
rect 372120 204212 372122 204232
rect 372066 204176 372122 204212
rect 372066 203632 372122 203688
rect 372066 201456 372122 201512
rect 372250 224032 372306 224088
rect 372158 200368 372214 200424
rect 371974 198736 372030 198792
rect 372158 198872 372214 198928
rect 372802 288532 372804 288552
rect 372804 288532 372856 288552
rect 372856 288532 372858 288552
rect 372802 288496 372858 288532
rect 372618 274624 372674 274680
rect 372526 207848 372582 207904
rect 372526 202544 372582 202600
rect 372710 225020 372712 225040
rect 372712 225020 372764 225040
rect 372764 225020 372766 225040
rect 372710 224984 372766 225020
rect 372710 223916 372766 223952
rect 372710 223896 372712 223916
rect 372712 223896 372764 223916
rect 372764 223896 372766 223916
rect 373170 211112 373226 211168
rect 373078 210604 373080 210624
rect 373080 210604 373132 210624
rect 373132 210604 373134 210624
rect 373078 210568 373134 210604
rect 372434 197648 372490 197704
rect 372066 143520 372122 143576
rect 371974 128560 372030 128616
rect 372066 127880 372122 127936
rect 371882 127336 371938 127392
rect 371790 126792 371846 126848
rect 372526 196560 372582 196616
rect 371330 125160 371386 125216
rect 372434 125704 372490 125760
rect 372710 139712 372766 139768
rect 374642 204720 374698 204776
rect 374550 201456 374606 201512
rect 374734 204040 374790 204096
rect 445206 369416 445262 369472
rect 445666 368328 445722 368384
rect 445666 367104 445722 367160
rect 444930 366016 444986 366072
rect 444930 364792 444986 364848
rect 444562 363704 444618 363760
rect 444930 362480 444986 362536
rect 445666 360204 445668 360224
rect 445668 360204 445720 360224
rect 445720 360204 445722 360224
rect 445666 360168 445722 360204
rect 444470 359080 444526 359136
rect 444930 357856 444986 357912
rect 444562 356788 444618 356824
rect 444562 356768 444564 356788
rect 444564 356768 444616 356788
rect 444616 356768 444618 356788
rect 444378 355544 444434 355600
rect 444470 354456 444526 354512
rect 444378 353232 444434 353288
rect 444562 350920 444618 350976
rect 444378 349832 444434 349888
rect 441802 225004 441858 225040
rect 441802 224984 441804 225004
rect 441804 224984 441856 225004
rect 441856 224984 441858 225004
rect 441802 223916 441858 223952
rect 441802 223896 441804 223916
rect 441804 223896 441856 223916
rect 441856 223896 441858 223916
rect 441618 125468 441620 125488
rect 441620 125468 441672 125488
rect 441672 125468 441674 125488
rect 441618 125432 441674 125468
rect 444470 347520 444526 347576
rect 444654 348608 444710 348664
rect 445206 346296 445262 346352
rect 445666 345208 445722 345264
rect 445666 343984 445722 344040
rect 445666 342896 445722 342952
rect 445114 341672 445170 341728
rect 444746 340584 444802 340640
rect 445666 297472 445722 297528
rect 445666 296384 445722 296440
rect 445850 361392 445906 361448
rect 445758 295160 445814 295216
rect 445666 294072 445722 294128
rect 445666 292884 445668 292904
rect 445668 292884 445720 292904
rect 445720 292884 445722 292904
rect 445666 292848 445722 292884
rect 445666 291760 445722 291816
rect 445666 290572 445668 290592
rect 445668 290572 445720 290592
rect 445720 290572 445722 290592
rect 445666 290536 445722 290572
rect 445666 289468 445722 289504
rect 445942 352144 445998 352200
rect 445666 289448 445668 289468
rect 445668 289448 445720 289468
rect 445720 289448 445722 289468
rect 445666 288224 445722 288280
rect 445114 287136 445170 287192
rect 445666 285912 445722 285968
rect 445666 284860 445668 284880
rect 445668 284860 445720 284880
rect 445720 284860 445722 284880
rect 445666 284824 445722 284860
rect 445482 283636 445484 283656
rect 445484 283636 445536 283656
rect 445536 283636 445538 283656
rect 445482 283600 445538 283636
rect 445390 282532 445446 282568
rect 445390 282512 445392 282532
rect 445392 282512 445444 282532
rect 445444 282512 445446 282532
rect 445114 281288 445170 281344
rect 444746 280200 444802 280256
rect 444838 278976 444894 279032
rect 444562 276664 444618 276720
rect 444470 275576 444526 275632
rect 444378 206896 444434 206952
rect 444746 208120 444802 208176
rect 445114 277888 445170 277944
rect 444838 206896 444894 206952
rect 445666 274352 445722 274408
rect 445574 273264 445630 273320
rect 445666 272040 445722 272096
rect 445666 270952 445722 271008
rect 445666 269728 445722 269784
rect 445666 268640 445722 268696
rect 445574 225392 445630 225448
rect 445666 223116 445668 223136
rect 445668 223116 445720 223136
rect 445720 223116 445722 223136
rect 445666 223080 445722 223116
rect 445666 221992 445722 222048
rect 445666 220788 445722 220824
rect 445666 220768 445668 220788
rect 445668 220768 445720 220788
rect 445720 220768 445722 220788
rect 445666 219680 445722 219736
rect 445482 218476 445538 218512
rect 445482 218456 445484 218476
rect 445484 218456 445536 218476
rect 445536 218456 445538 218476
rect 445666 217388 445722 217424
rect 445666 217368 445668 217388
rect 445668 217368 445720 217388
rect 445720 217368 445722 217388
rect 445666 216164 445722 216200
rect 445666 216144 445668 216164
rect 445668 216144 445720 216164
rect 445720 216144 445722 216164
rect 445482 215056 445538 215112
rect 445666 213868 445668 213888
rect 445668 213868 445720 213888
rect 445720 213868 445722 213888
rect 445666 213832 445722 213868
rect 445666 212764 445722 212800
rect 445666 212744 445668 212764
rect 445668 212744 445720 212764
rect 445720 212744 445722 212764
rect 445482 211556 445484 211576
rect 445484 211556 445536 211576
rect 445536 211556 445538 211576
rect 445482 211520 445538 211556
rect 445390 210468 445392 210488
rect 445392 210468 445444 210488
rect 445444 210468 445446 210488
rect 445390 210432 445446 210468
rect 445206 209228 445262 209264
rect 445206 209208 445208 209228
rect 445208 209208 445260 209228
rect 445260 209208 445262 209228
rect 444654 205808 444710 205864
rect 445114 205808 445170 205864
rect 444562 204584 444618 204640
rect 444470 203496 444526 203552
rect 444378 141924 444380 141944
rect 444380 141924 444432 141944
rect 444432 141924 444434 141944
rect 444378 141888 444434 141924
rect 444378 139576 444434 139632
rect 444378 138488 444434 138544
rect 444378 137300 444380 137320
rect 444380 137300 444432 137320
rect 444432 137300 444434 137320
rect 444378 137264 444434 137300
rect 445666 202272 445722 202328
rect 445666 201184 445722 201240
rect 445666 199960 445722 200016
rect 445666 198872 445722 198928
rect 445666 197648 445722 197704
rect 444838 152360 444894 152416
rect 444838 151136 444894 151192
rect 445666 153448 445722 153504
rect 444930 150048 444986 150104
rect 445298 148860 445300 148880
rect 445300 148860 445352 148880
rect 445352 148860 445354 148880
rect 445298 148824 445354 148860
rect 445574 147736 445630 147792
rect 444838 146548 444840 146568
rect 444840 146548 444892 146568
rect 444892 146548 444894 146568
rect 444838 146512 444894 146548
rect 445482 145424 445538 145480
rect 445114 144200 445170 144256
rect 445114 143148 445116 143168
rect 445116 143148 445168 143168
rect 445168 143148 445170 143168
rect 445114 143112 445170 143148
rect 444746 140800 444802 140856
rect 444746 136176 444802 136232
rect 444654 133864 444710 133920
rect 444562 132640 444618 132696
rect 444470 131552 444526 131608
rect 442998 130328 443054 130384
rect 443918 130364 443920 130384
rect 443920 130364 443972 130384
rect 443972 130364 443974 130384
rect 443918 130328 443974 130364
rect 441894 126384 441950 126440
rect 443642 129240 443698 129296
rect 443090 128016 443146 128072
rect 444378 128052 444380 128072
rect 444380 128052 444432 128072
rect 444432 128052 444434 128072
rect 444378 128016 444434 128052
rect 444378 125704 444434 125760
rect 444838 134952 444894 135008
rect 445666 126928 445722 126984
rect 445850 196560 445906 196616
rect 441894 124908 441950 124944
rect 445942 136176 445998 136232
rect 447506 185544 447562 185600
rect 448886 173168 448942 173224
rect 450174 171672 450230 171728
rect 441894 124888 441896 124908
rect 441896 124888 441948 124908
rect 441948 124888 441950 124908
rect 436742 97416 436798 97472
rect 443642 97280 443698 97336
rect 580170 697176 580226 697232
rect 580170 683848 580226 683904
rect 580170 670692 580172 670712
rect 580172 670692 580224 670712
rect 580224 670692 580226 670712
rect 580170 670656 580226 670692
rect 580170 644000 580226 644056
rect 580170 630808 580226 630864
rect 580170 617480 580226 617536
rect 579802 590960 579858 591016
rect 580170 577632 580226 577688
rect 579802 564304 579858 564360
rect 580170 537784 580226 537840
rect 580170 524476 580226 524512
rect 580170 524456 580172 524476
rect 580172 524456 580224 524476
rect 580224 524456 580226 524476
rect 580170 511264 580226 511320
rect 580170 484608 580226 484664
rect 579986 471416 580042 471472
rect 580170 458088 580226 458144
rect 580170 431568 580226 431624
rect 580170 418240 580226 418296
rect 580170 404912 580226 404968
rect 580170 378392 580226 378448
rect 580262 365064 580318 365120
rect 580170 325216 580226 325272
rect 580170 312024 580226 312080
rect 580354 351872 580410 351928
rect 580170 298696 580226 298752
rect 580262 272176 580318 272232
rect 580170 258848 580226 258904
rect 580170 245556 580172 245576
rect 580172 245556 580224 245576
rect 580224 245556 580226 245576
rect 580170 245520 580226 245556
rect 579986 232328 580042 232384
rect 580262 219000 580318 219056
rect 579802 205672 579858 205728
rect 580170 192480 580226 192536
rect 580170 179152 580226 179208
rect 580170 165824 580226 165880
rect 580170 152632 580226 152688
rect 580170 139340 580172 139360
rect 580172 139340 580224 139360
rect 580224 139340 580226 139360
rect 580170 139304 580226 139340
rect 580170 125976 580226 126032
rect 579802 112784 579858 112840
rect 580170 99456 580226 99512
rect 525798 95920 525854 95976
rect 550638 95784 550694 95840
rect 580262 97144 580318 97200
rect 580170 86128 580226 86184
rect 579986 72936 580042 72992
rect 580170 59608 580226 59664
rect 580170 33108 580226 33144
rect 580170 33088 580172 33108
rect 580172 33088 580224 33108
rect 580224 33088 580226 33108
rect 580170 19760 580226 19816
rect 582470 46280 582526 46336
rect 582378 6568 582434 6624
<< metal3 >>
rect -960 697220 480 697460
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 580165 683906 580231 683909
rect 583520 683906 584960 683996
rect 580165 683904 584960 683906
rect 580165 683848 580170 683904
rect 580226 683848 584960 683904
rect 580165 683846 584960 683848
rect 580165 683843 580231 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3417 671258 3483 671261
rect -960 671256 3483 671258
rect -960 671200 3422 671256
rect 3478 671200 3483 671256
rect -960 671198 3483 671200
rect -960 671108 480 671198
rect 3417 671195 3483 671198
rect 580165 670714 580231 670717
rect 583520 670714 584960 670804
rect 580165 670712 584960 670714
rect 580165 670656 580170 670712
rect 580226 670656 584960 670712
rect 580165 670654 584960 670656
rect 580165 670651 580231 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3417 658202 3483 658205
rect -960 658200 3483 658202
rect -960 658144 3422 658200
rect 3478 658144 3483 658200
rect -960 658142 3483 658144
rect -960 658052 480 658142
rect 3417 658139 3483 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 580165 644058 580231 644061
rect 583520 644058 584960 644148
rect 580165 644056 584960 644058
rect 580165 644000 580170 644056
rect 580226 644000 584960 644056
rect 580165 643998 584960 644000
rect 580165 643995 580231 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 3417 632090 3483 632093
rect -960 632088 3483 632090
rect -960 632032 3422 632088
rect 3478 632032 3483 632088
rect -960 632030 3483 632032
rect -960 631940 480 632030
rect 3417 632027 3483 632030
rect 580165 630866 580231 630869
rect 583520 630866 584960 630956
rect 580165 630864 584960 630866
rect 580165 630808 580170 630864
rect 580226 630808 584960 630864
rect 580165 630806 584960 630808
rect 580165 630803 580231 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3141 619170 3207 619173
rect -960 619168 3207 619170
rect -960 619112 3146 619168
rect 3202 619112 3207 619168
rect -960 619110 3207 619112
rect -960 619020 480 619110
rect 3141 619107 3207 619110
rect 580165 617538 580231 617541
rect 583520 617538 584960 617628
rect 580165 617536 584960 617538
rect 580165 617480 580170 617536
rect 580226 617480 584960 617536
rect 580165 617478 584960 617480
rect 580165 617475 580231 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3233 606114 3299 606117
rect -960 606112 3299 606114
rect -960 606056 3238 606112
rect 3294 606056 3299 606112
rect -960 606054 3299 606056
rect -960 605964 480 606054
rect 3233 606051 3299 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 579797 591018 579863 591021
rect 583520 591018 584960 591108
rect 579797 591016 584960 591018
rect 579797 590960 579802 591016
rect 579858 590960 584960 591016
rect 579797 590958 584960 590960
rect 579797 590955 579863 590958
rect 583520 590868 584960 590958
rect -960 580002 480 580092
rect 3325 580002 3391 580005
rect -960 580000 3391 580002
rect -960 579944 3330 580000
rect 3386 579944 3391 580000
rect -960 579942 3391 579944
rect -960 579852 480 579942
rect 3325 579939 3391 579942
rect 580165 577690 580231 577693
rect 583520 577690 584960 577780
rect 580165 577688 584960 577690
rect 580165 577632 580170 577688
rect 580226 577632 584960 577688
rect 580165 577630 584960 577632
rect 580165 577627 580231 577630
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 3417 566946 3483 566949
rect -960 566944 3483 566946
rect -960 566888 3422 566944
rect 3478 566888 3483 566944
rect -960 566886 3483 566888
rect -960 566796 480 566886
rect 3417 566883 3483 566886
rect 579797 564362 579863 564365
rect 583520 564362 584960 564452
rect 579797 564360 584960 564362
rect 579797 564304 579802 564360
rect 579858 564304 584960 564360
rect 579797 564302 584960 564304
rect 579797 564299 579863 564302
rect 583520 564212 584960 564302
rect -960 553890 480 553980
rect 3417 553890 3483 553893
rect -960 553888 3483 553890
rect -960 553832 3422 553888
rect 3478 553832 3483 553888
rect -960 553830 3483 553832
rect -960 553740 480 553830
rect 3417 553827 3483 553830
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 580165 537842 580231 537845
rect 583520 537842 584960 537932
rect 580165 537840 584960 537842
rect 580165 537784 580170 537840
rect 580226 537784 584960 537840
rect 580165 537782 584960 537784
rect 580165 537779 580231 537782
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect 3417 527914 3483 527917
rect -960 527912 3483 527914
rect -960 527856 3422 527912
rect 3478 527856 3483 527912
rect -960 527854 3483 527856
rect -960 527764 480 527854
rect 3417 527851 3483 527854
rect 580165 524514 580231 524517
rect 583520 524514 584960 524604
rect 580165 524512 584960 524514
rect 580165 524456 580170 524512
rect 580226 524456 584960 524512
rect 580165 524454 584960 524456
rect 580165 524451 580231 524454
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 3417 514858 3483 514861
rect -960 514856 3483 514858
rect -960 514800 3422 514856
rect 3478 514800 3483 514856
rect -960 514798 3483 514800
rect -960 514708 480 514798
rect 3417 514795 3483 514798
rect 580165 511322 580231 511325
rect 583520 511322 584960 511412
rect 580165 511320 584960 511322
rect 580165 511264 580170 511320
rect 580226 511264 584960 511320
rect 580165 511262 584960 511264
rect 580165 511259 580231 511262
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect 3049 501802 3115 501805
rect -960 501800 3115 501802
rect -960 501744 3054 501800
rect 3110 501744 3115 501800
rect -960 501742 3115 501744
rect -960 501652 480 501742
rect 3049 501739 3115 501742
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 580165 484666 580231 484669
rect 583520 484666 584960 484756
rect 580165 484664 584960 484666
rect 580165 484608 580170 484664
rect 580226 484608 584960 484664
rect 580165 484606 584960 484608
rect 580165 484603 580231 484606
rect 583520 484516 584960 484606
rect -960 475690 480 475780
rect 3417 475690 3483 475693
rect -960 475688 3483 475690
rect -960 475632 3422 475688
rect 3478 475632 3483 475688
rect -960 475630 3483 475632
rect -960 475540 480 475630
rect 3417 475627 3483 475630
rect 579981 471474 580047 471477
rect 583520 471474 584960 471564
rect 579981 471472 584960 471474
rect 579981 471416 579986 471472
rect 580042 471416 584960 471472
rect 579981 471414 584960 471416
rect 579981 471411 580047 471414
rect 583520 471324 584960 471414
rect -960 462634 480 462724
rect 3233 462634 3299 462637
rect -960 462632 3299 462634
rect -960 462576 3238 462632
rect 3294 462576 3299 462632
rect -960 462574 3299 462576
rect -960 462484 480 462574
rect 3233 462571 3299 462574
rect 580165 458146 580231 458149
rect 583520 458146 584960 458236
rect 580165 458144 584960 458146
rect 580165 458088 580170 458144
rect 580226 458088 584960 458144
rect 580165 458086 584960 458088
rect 580165 458083 580231 458086
rect 583520 457996 584960 458086
rect -960 449578 480 449668
rect 3141 449578 3207 449581
rect -960 449576 3207 449578
rect -960 449520 3146 449576
rect 3202 449520 3207 449576
rect -960 449518 3207 449520
rect -960 449428 480 449518
rect 3141 449515 3207 449518
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 580165 431626 580231 431629
rect 583520 431626 584960 431716
rect 580165 431624 584960 431626
rect 580165 431568 580170 431624
rect 580226 431568 584960 431624
rect 580165 431566 584960 431568
rect 580165 431563 580231 431566
rect 583520 431476 584960 431566
rect -960 423602 480 423692
rect 3417 423602 3483 423605
rect -960 423600 3483 423602
rect -960 423544 3422 423600
rect 3478 423544 3483 423600
rect -960 423542 3483 423544
rect -960 423452 480 423542
rect 3417 423539 3483 423542
rect 580165 418298 580231 418301
rect 583520 418298 584960 418388
rect 580165 418296 584960 418298
rect 580165 418240 580170 418296
rect 580226 418240 584960 418296
rect 580165 418238 584960 418240
rect 580165 418235 580231 418238
rect 583520 418148 584960 418238
rect -960 410546 480 410636
rect 3141 410546 3207 410549
rect -960 410544 3207 410546
rect -960 410488 3146 410544
rect 3202 410488 3207 410544
rect -960 410486 3207 410488
rect -960 410396 480 410486
rect 3141 410483 3207 410486
rect 580165 404970 580231 404973
rect 583520 404970 584960 405060
rect 580165 404968 584960 404970
rect 580165 404912 580170 404968
rect 580226 404912 584960 404968
rect 580165 404910 584960 404912
rect 580165 404907 580231 404910
rect 583520 404820 584960 404910
rect -960 397490 480 397580
rect 3417 397490 3483 397493
rect -960 397488 3483 397490
rect -960 397432 3422 397488
rect 3478 397432 3483 397488
rect -960 397430 3483 397432
rect -960 397340 480 397430
rect 3417 397427 3483 397430
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 580165 378450 580231 378453
rect 583520 378450 584960 378540
rect 580165 378448 584960 378450
rect 580165 378392 580170 378448
rect 580226 378392 584960 378448
rect 580165 378390 584960 378392
rect 580165 378387 580231 378390
rect 583520 378300 584960 378390
rect -960 371378 480 371468
rect 3417 371378 3483 371381
rect -960 371376 3483 371378
rect -960 371320 3422 371376
rect 3478 371320 3483 371376
rect -960 371318 3483 371320
rect -960 371228 480 371318
rect 3417 371315 3483 371318
rect 371693 369746 371759 369749
rect 369932 369744 371759 369746
rect 369932 369688 371698 369744
rect 371754 369688 371759 369744
rect 369932 369686 371759 369688
rect 371693 369683 371759 369686
rect 445201 369474 445267 369477
rect 441876 369472 445267 369474
rect 441876 369416 445206 369472
rect 445262 369416 445267 369472
rect 441876 369414 445267 369416
rect 445201 369411 445267 369414
rect 371877 369202 371943 369205
rect 369932 369200 371943 369202
rect 369932 369144 371882 369200
rect 371938 369144 371943 369200
rect 369932 369142 371943 369144
rect 371877 369139 371943 369142
rect 371601 368658 371667 368661
rect 369932 368656 371667 368658
rect 369932 368600 371606 368656
rect 371662 368600 371667 368656
rect 369932 368598 371667 368600
rect 371601 368595 371667 368598
rect 445661 368386 445727 368389
rect 441876 368384 445727 368386
rect 441876 368328 445666 368384
rect 445722 368328 445727 368384
rect 441876 368326 445727 368328
rect 445661 368323 445727 368326
rect 371601 368114 371667 368117
rect 369932 368112 371667 368114
rect 369932 368056 371606 368112
rect 371662 368056 371667 368112
rect 369932 368054 371667 368056
rect 371601 368051 371667 368054
rect 371509 367570 371575 367573
rect 369932 367568 371575 367570
rect 369932 367512 371514 367568
rect 371570 367512 371575 367568
rect 369932 367510 371575 367512
rect 371509 367507 371575 367510
rect 445661 367162 445727 367165
rect 441876 367160 445727 367162
rect 441876 367104 445666 367160
rect 445722 367104 445727 367160
rect 441876 367102 445727 367104
rect 445661 367099 445727 367102
rect 371601 367026 371667 367029
rect 369932 367024 371667 367026
rect 369932 366968 371606 367024
rect 371662 366968 371667 367024
rect 369932 366966 371667 366968
rect 371601 366963 371667 366966
rect 372521 366482 372587 366485
rect 369932 366480 372587 366482
rect 369932 366424 372526 366480
rect 372582 366424 372587 366480
rect 369932 366422 372587 366424
rect 372521 366419 372587 366422
rect 444925 366074 444991 366077
rect 441876 366072 444991 366074
rect 441876 366016 444930 366072
rect 444986 366016 444991 366072
rect 441876 366014 444991 366016
rect 444925 366011 444991 366014
rect 371233 365938 371299 365941
rect 369932 365936 371299 365938
rect 369932 365880 371238 365936
rect 371294 365880 371299 365936
rect 369932 365878 371299 365880
rect 371233 365875 371299 365878
rect 371601 365394 371667 365397
rect 369932 365392 371667 365394
rect 369932 365336 371606 365392
rect 371662 365336 371667 365392
rect 369932 365334 371667 365336
rect 371601 365331 371667 365334
rect 580257 365122 580323 365125
rect 583520 365122 584960 365212
rect 580257 365120 584960 365122
rect 580257 365064 580262 365120
rect 580318 365064 584960 365120
rect 580257 365062 584960 365064
rect 580257 365059 580323 365062
rect 583520 364972 584960 365062
rect 371233 364850 371299 364853
rect 444925 364850 444991 364853
rect 369932 364848 371299 364850
rect 369932 364792 371238 364848
rect 371294 364792 371299 364848
rect 369932 364790 371299 364792
rect 441876 364848 444991 364850
rect 441876 364792 444930 364848
rect 444986 364792 444991 364848
rect 441876 364790 444991 364792
rect 371233 364787 371299 364790
rect 444925 364787 444991 364790
rect 371693 364306 371759 364309
rect 369932 364304 371759 364306
rect 369932 364248 371698 364304
rect 371754 364248 371759 364304
rect 369932 364246 371759 364248
rect 371693 364243 371759 364246
rect 371601 363762 371667 363765
rect 444557 363762 444623 363765
rect 369932 363760 371667 363762
rect 369932 363704 371606 363760
rect 371662 363704 371667 363760
rect 369932 363702 371667 363704
rect 441876 363760 444623 363762
rect 441876 363704 444562 363760
rect 444618 363704 444623 363760
rect 441876 363702 444623 363704
rect 371601 363699 371667 363702
rect 444557 363699 444623 363702
rect 371417 363218 371483 363221
rect 369932 363216 371483 363218
rect 369932 363160 371422 363216
rect 371478 363160 371483 363216
rect 369932 363158 371483 363160
rect 371417 363155 371483 363158
rect 372797 362674 372863 362677
rect 369932 362672 372863 362674
rect 369932 362616 372802 362672
rect 372858 362616 372863 362672
rect 369932 362614 372863 362616
rect 372797 362611 372863 362614
rect 444925 362538 444991 362541
rect 441876 362536 444991 362538
rect 441876 362480 444930 362536
rect 444986 362480 444991 362536
rect 441876 362478 444991 362480
rect 444925 362475 444991 362478
rect 371417 362130 371483 362133
rect 369932 362128 371483 362130
rect 369932 362072 371422 362128
rect 371478 362072 371483 362128
rect 369932 362070 371483 362072
rect 371417 362067 371483 362070
rect 371509 361586 371575 361589
rect 369932 361584 371575 361586
rect 369932 361528 371514 361584
rect 371570 361528 371575 361584
rect 369932 361526 371575 361528
rect 371509 361523 371575 361526
rect 445845 361450 445911 361453
rect 441876 361448 445911 361450
rect 441876 361392 445850 361448
rect 445906 361392 445911 361448
rect 441876 361390 445911 361392
rect 445845 361387 445911 361390
rect 371693 361042 371759 361045
rect 369932 361040 371759 361042
rect 369932 360984 371698 361040
rect 371754 360984 371759 361040
rect 369932 360982 371759 360984
rect 371693 360979 371759 360982
rect 371601 360498 371667 360501
rect 369932 360496 371667 360498
rect 369932 360440 371606 360496
rect 371662 360440 371667 360496
rect 369932 360438 371667 360440
rect 371601 360435 371667 360438
rect 445661 360226 445727 360229
rect 441876 360224 445727 360226
rect 441876 360168 445666 360224
rect 445722 360168 445727 360224
rect 441876 360166 445727 360168
rect 445661 360163 445727 360166
rect 371325 360090 371391 360093
rect 369932 360088 371391 360090
rect 369932 360032 371330 360088
rect 371386 360032 371391 360088
rect 369932 360030 371391 360032
rect 371325 360027 371391 360030
rect 372061 359546 372127 359549
rect 369932 359544 372127 359546
rect 369932 359488 372066 359544
rect 372122 359488 372127 359544
rect 369932 359486 372127 359488
rect 372061 359483 372127 359486
rect 444465 359138 444531 359141
rect 441876 359136 444531 359138
rect 441876 359080 444470 359136
rect 444526 359080 444531 359136
rect 441876 359078 444531 359080
rect 444465 359075 444531 359078
rect 372245 359002 372311 359005
rect 369932 359000 372311 359002
rect 369932 358944 372250 359000
rect 372306 358944 372311 359000
rect 369932 358942 372311 358944
rect 372245 358939 372311 358942
rect -960 358458 480 358548
rect 3141 358458 3207 358461
rect 371509 358458 371575 358461
rect -960 358456 3207 358458
rect -960 358400 3146 358456
rect 3202 358400 3207 358456
rect -960 358398 3207 358400
rect 369932 358456 371575 358458
rect 369932 358400 371514 358456
rect 371570 358400 371575 358456
rect 369932 358398 371575 358400
rect -960 358308 480 358398
rect 3141 358395 3207 358398
rect 371509 358395 371575 358398
rect 371417 357914 371483 357917
rect 444925 357914 444991 357917
rect 369932 357912 371483 357914
rect 369932 357856 371422 357912
rect 371478 357856 371483 357912
rect 369932 357854 371483 357856
rect 441876 357912 444991 357914
rect 441876 357856 444930 357912
rect 444986 357856 444991 357912
rect 441876 357854 444991 357856
rect 371417 357851 371483 357854
rect 444925 357851 444991 357854
rect 371233 357370 371299 357373
rect 369932 357368 371299 357370
rect 369932 357312 371238 357368
rect 371294 357312 371299 357368
rect 369932 357310 371299 357312
rect 371233 357307 371299 357310
rect 371325 356826 371391 356829
rect 444557 356826 444623 356829
rect 369932 356824 371391 356826
rect 369932 356768 371330 356824
rect 371386 356768 371391 356824
rect 369932 356766 371391 356768
rect 441876 356824 444623 356826
rect 441876 356768 444562 356824
rect 444618 356768 444623 356824
rect 441876 356766 444623 356768
rect 371325 356763 371391 356766
rect 444557 356763 444623 356766
rect 371417 356282 371483 356285
rect 369932 356280 371483 356282
rect 369932 356224 371422 356280
rect 371478 356224 371483 356280
rect 369932 356222 371483 356224
rect 371417 356219 371483 356222
rect 371693 355738 371759 355741
rect 369932 355736 371759 355738
rect 369932 355680 371698 355736
rect 371754 355680 371759 355736
rect 369932 355678 371759 355680
rect 371693 355675 371759 355678
rect 444373 355602 444439 355605
rect 441876 355600 444439 355602
rect 441876 355544 444378 355600
rect 444434 355544 444439 355600
rect 441876 355542 444439 355544
rect 444373 355539 444439 355542
rect 371233 355194 371299 355197
rect 369932 355192 371299 355194
rect 369932 355136 371238 355192
rect 371294 355136 371299 355192
rect 369932 355134 371299 355136
rect 371233 355131 371299 355134
rect 371509 354650 371575 354653
rect 369932 354648 371575 354650
rect 369932 354592 371514 354648
rect 371570 354592 371575 354648
rect 369932 354590 371575 354592
rect 371509 354587 371575 354590
rect 444465 354514 444531 354517
rect 441876 354512 444531 354514
rect 441876 354456 444470 354512
rect 444526 354456 444531 354512
rect 441876 354454 444531 354456
rect 444465 354451 444531 354454
rect 371693 354106 371759 354109
rect 369932 354104 371759 354106
rect 369932 354048 371698 354104
rect 371754 354048 371759 354104
rect 369932 354046 371759 354048
rect 371693 354043 371759 354046
rect 371918 353562 371924 353564
rect 369932 353502 371924 353562
rect 371918 353500 371924 353502
rect 371988 353500 371994 353564
rect 444373 353290 444439 353293
rect 441876 353288 444439 353290
rect 441876 353232 444378 353288
rect 444434 353232 444439 353288
rect 441876 353230 444439 353232
rect 444373 353227 444439 353230
rect 371734 353018 371740 353020
rect 369932 352958 371740 353018
rect 371734 352956 371740 352958
rect 371804 352956 371810 353020
rect 372102 352474 372108 352476
rect 369932 352414 372108 352474
rect 372102 352412 372108 352414
rect 372172 352412 372178 352476
rect 445937 352202 446003 352205
rect 441876 352200 446003 352202
rect 441876 352144 445942 352200
rect 445998 352144 446003 352200
rect 441876 352142 446003 352144
rect 445937 352139 446003 352142
rect 371325 351930 371391 351933
rect 369932 351928 371391 351930
rect 369932 351872 371330 351928
rect 371386 351872 371391 351928
rect 369932 351870 371391 351872
rect 371325 351867 371391 351870
rect 580349 351930 580415 351933
rect 583520 351930 584960 352020
rect 580349 351928 584960 351930
rect 580349 351872 580354 351928
rect 580410 351872 584960 351928
rect 580349 351870 584960 351872
rect 580349 351867 580415 351870
rect 583520 351780 584960 351870
rect 371550 351386 371556 351388
rect 369932 351326 371556 351386
rect 371550 351324 371556 351326
rect 371620 351324 371626 351388
rect 444557 350978 444623 350981
rect 441876 350976 444623 350978
rect 441876 350920 444562 350976
rect 444618 350920 444623 350976
rect 441876 350918 444623 350920
rect 444557 350915 444623 350918
rect 371182 350842 371188 350844
rect 369932 350782 371188 350842
rect 371182 350780 371188 350782
rect 371252 350780 371258 350844
rect 371877 350298 371943 350301
rect 369932 350296 371943 350298
rect 369932 350240 371882 350296
rect 371938 350240 371943 350296
rect 369932 350238 371943 350240
rect 371877 350235 371943 350238
rect 372153 349890 372219 349893
rect 444373 349890 444439 349893
rect 369932 349888 372219 349890
rect 369932 349832 372158 349888
rect 372214 349832 372219 349888
rect 369932 349830 372219 349832
rect 441876 349888 444439 349890
rect 441876 349832 444378 349888
rect 444434 349832 444439 349888
rect 441876 349830 444439 349832
rect 372153 349827 372219 349830
rect 444373 349827 444439 349830
rect 370313 349346 370379 349349
rect 369932 349344 370379 349346
rect 369932 349288 370318 349344
rect 370374 349288 370379 349344
rect 369932 349286 370379 349288
rect 370313 349283 370379 349286
rect 369350 348533 369410 348772
rect 444649 348666 444715 348669
rect 441876 348664 444715 348666
rect 441876 348608 444654 348664
rect 444710 348608 444715 348664
rect 441876 348606 444715 348608
rect 444649 348603 444715 348606
rect 369301 348528 369410 348533
rect 369301 348472 369306 348528
rect 369362 348472 369410 348528
rect 369301 348470 369410 348472
rect 369301 348467 369367 348470
rect 371601 348258 371667 348261
rect 369932 348256 371667 348258
rect 369932 348200 371606 348256
rect 371662 348200 371667 348256
rect 369932 348198 371667 348200
rect 371601 348195 371667 348198
rect 370497 347714 370563 347717
rect 369932 347712 370563 347714
rect 369932 347656 370502 347712
rect 370558 347656 370563 347712
rect 369932 347654 370563 347656
rect 370497 347651 370563 347654
rect 444465 347578 444531 347581
rect 441876 347576 444531 347578
rect 441876 347520 444470 347576
rect 444526 347520 444531 347576
rect 441876 347518 444531 347520
rect 444465 347515 444531 347518
rect 369902 346898 369962 347140
rect 370037 346898 370103 346901
rect 369902 346896 370103 346898
rect 369902 346840 370042 346896
rect 370098 346840 370103 346896
rect 369902 346838 370103 346840
rect 370037 346835 370103 346838
rect 372705 346626 372771 346629
rect 369932 346624 372771 346626
rect 369932 346568 372710 346624
rect 372766 346568 372771 346624
rect 369932 346566 372771 346568
rect 372705 346563 372771 346566
rect 445201 346354 445267 346357
rect 441876 346352 445267 346354
rect 441876 346296 445206 346352
rect 445262 346296 445267 346352
rect 441876 346294 445267 346296
rect 445201 346291 445267 346294
rect 370589 346082 370655 346085
rect 369932 346080 370655 346082
rect 369932 346024 370594 346080
rect 370650 346024 370655 346080
rect 369932 346022 370655 346024
rect 370589 346019 370655 346022
rect -960 345402 480 345492
rect 3325 345402 3391 345405
rect -960 345400 3391 345402
rect -960 345344 3330 345400
rect 3386 345344 3391 345400
rect -960 345342 3391 345344
rect -960 345252 480 345342
rect 3325 345339 3391 345342
rect 369902 345269 369962 345508
rect 369902 345264 370011 345269
rect 445661 345266 445727 345269
rect 369902 345208 369950 345264
rect 370006 345208 370011 345264
rect 369902 345206 370011 345208
rect 441876 345264 445727 345266
rect 441876 345208 445666 345264
rect 445722 345208 445727 345264
rect 441876 345206 445727 345208
rect 369945 345203 370011 345206
rect 445661 345203 445727 345206
rect 371969 344994 372035 344997
rect 369932 344992 372035 344994
rect 369932 344936 371974 344992
rect 372030 344936 372035 344992
rect 369932 344934 372035 344936
rect 371969 344931 372035 344934
rect 372245 344450 372311 344453
rect 369932 344448 372311 344450
rect 369932 344392 372250 344448
rect 372306 344392 372311 344448
rect 369932 344390 372311 344392
rect 372245 344387 372311 344390
rect 445661 344042 445727 344045
rect 441876 344040 445727 344042
rect 441876 343984 445666 344040
rect 445722 343984 445727 344040
rect 441876 343982 445727 343984
rect 445661 343979 445727 343982
rect 371785 343906 371851 343909
rect 369932 343904 371851 343906
rect 369932 343848 371790 343904
rect 371846 343848 371851 343904
rect 369932 343846 371851 343848
rect 371785 343843 371851 343846
rect 371417 343362 371483 343365
rect 369932 343360 371483 343362
rect 369932 343304 371422 343360
rect 371478 343304 371483 343360
rect 369932 343302 371483 343304
rect 371417 343299 371483 343302
rect 445661 342954 445727 342957
rect 441876 342952 445727 342954
rect 441876 342896 445666 342952
rect 445722 342896 445727 342952
rect 441876 342894 445727 342896
rect 445661 342891 445727 342894
rect 372061 342818 372127 342821
rect 369932 342816 372127 342818
rect 369932 342760 372066 342816
rect 372122 342760 372127 342816
rect 369932 342758 372127 342760
rect 372061 342755 372127 342758
rect 372429 342274 372495 342277
rect 369932 342272 372495 342274
rect 369932 342216 372434 342272
rect 372490 342216 372495 342272
rect 369932 342214 372495 342216
rect 372429 342211 372495 342214
rect 371509 341730 371575 341733
rect 445109 341730 445175 341733
rect 369932 341728 371575 341730
rect 369932 341672 371514 341728
rect 371570 341672 371575 341728
rect 369932 341670 371575 341672
rect 441876 341728 445175 341730
rect 441876 341672 445114 341728
rect 445170 341672 445175 341728
rect 441876 341670 445175 341672
rect 371509 341667 371575 341670
rect 445109 341667 445175 341670
rect 371693 341186 371759 341189
rect 369932 341184 371759 341186
rect 369932 341128 371698 341184
rect 371754 341128 371759 341184
rect 369932 341126 371759 341128
rect 371693 341123 371759 341126
rect 371601 340642 371667 340645
rect 444741 340642 444807 340645
rect 369932 340640 371667 340642
rect 369932 340584 371606 340640
rect 371662 340584 371667 340640
rect 369932 340582 371667 340584
rect 441876 340640 444807 340642
rect 441876 340584 444746 340640
rect 444802 340584 444807 340640
rect 441876 340582 444807 340584
rect 371601 340579 371667 340582
rect 444741 340579 444807 340582
rect 370405 340234 370471 340237
rect 369932 340232 370471 340234
rect 369932 340176 370410 340232
rect 370466 340176 370471 340232
rect 369932 340174 370471 340176
rect 370405 340171 370471 340174
rect 583520 338452 584960 338692
rect 361614 337724 361620 337788
rect 361684 337786 361690 337788
rect 362861 337786 362927 337789
rect 361684 337784 362927 337786
rect 361684 337728 362866 337784
rect 362922 337728 362927 337784
rect 361684 337726 362927 337728
rect 361684 337724 361690 337726
rect 362861 337723 362927 337726
rect 364374 337724 364380 337788
rect 364444 337786 364450 337788
rect 364885 337786 364951 337789
rect 364444 337784 364951 337786
rect 364444 337728 364890 337784
rect 364946 337728 364951 337784
rect 364444 337726 364951 337728
rect 364444 337724 364450 337726
rect 364885 337723 364951 337726
rect -960 332196 480 332436
rect 580165 325274 580231 325277
rect 583520 325274 584960 325364
rect 580165 325272 584960 325274
rect 580165 325216 580170 325272
rect 580226 325216 584960 325272
rect 580165 325214 584960 325216
rect 580165 325211 580231 325214
rect 583520 325124 584960 325214
rect -960 319290 480 319380
rect 3417 319290 3483 319293
rect -960 319288 3483 319290
rect -960 319232 3422 319288
rect 3478 319232 3483 319288
rect -960 319230 3483 319232
rect -960 319140 480 319230
rect 3417 319227 3483 319230
rect 580165 312082 580231 312085
rect 583520 312082 584960 312172
rect 580165 312080 584960 312082
rect 580165 312024 580170 312080
rect 580226 312024 584960 312080
rect 580165 312022 584960 312024
rect 580165 312019 580231 312022
rect 583520 311932 584960 312022
rect -960 306234 480 306324
rect 3233 306234 3299 306237
rect -960 306232 3299 306234
rect -960 306176 3238 306232
rect 3294 306176 3299 306232
rect -960 306174 3299 306176
rect -960 306084 480 306174
rect 3233 306171 3299 306174
rect 217041 299570 217107 299573
rect 218053 299570 218119 299573
rect 217041 299568 218119 299570
rect 217041 299512 217046 299568
rect 217102 299512 218058 299568
rect 218114 299512 218119 299568
rect 217041 299510 218119 299512
rect 217041 299507 217107 299510
rect 218053 299507 218119 299510
rect 218053 299434 218119 299437
rect 218789 299434 218855 299437
rect 218053 299432 218855 299434
rect 218053 299376 218058 299432
rect 218114 299376 218794 299432
rect 218850 299376 218855 299432
rect 218053 299374 218855 299376
rect 218053 299371 218119 299374
rect 218789 299371 218855 299374
rect 217133 299298 217199 299301
rect 219893 299298 219959 299301
rect 217133 299296 219959 299298
rect 217133 299240 217138 299296
rect 217194 299240 219898 299296
rect 219954 299240 219959 299296
rect 217133 299238 219959 299240
rect 217133 299235 217199 299238
rect 219893 299235 219959 299238
rect 198549 298890 198615 298893
rect 198549 298888 200100 298890
rect 198549 298832 198554 298888
rect 198610 298832 200100 298888
rect 198549 298830 200100 298832
rect 198549 298827 198615 298830
rect 580165 298754 580231 298757
rect 583520 298754 584960 298844
rect 580165 298752 584960 298754
rect 580165 298696 580170 298752
rect 580226 298696 584960 298752
rect 580165 298694 584960 298696
rect 580165 298691 580231 298694
rect 583520 298604 584960 298694
rect 302785 298346 302851 298349
rect 299828 298344 302851 298346
rect 299828 298288 302790 298344
rect 302846 298288 302851 298344
rect 299828 298286 302851 298288
rect 302785 298283 302851 298286
rect 371233 297802 371299 297805
rect 369380 297800 371299 297802
rect 369380 297772 371238 297800
rect 369350 297744 371238 297772
rect 371294 297744 371299 297800
rect 369350 297742 371299 297744
rect 369350 297397 369410 297742
rect 371233 297739 371299 297742
rect 445661 297530 445727 297533
rect 441876 297528 445727 297530
rect 441876 297472 445666 297528
rect 445722 297472 445727 297528
rect 441876 297470 445727 297472
rect 445661 297467 445727 297470
rect 369350 297392 369459 297397
rect 369350 297336 369398 297392
rect 369454 297336 369459 297392
rect 369350 297334 369459 297336
rect 369393 297331 369459 297334
rect 371233 297258 371299 297261
rect 369380 297256 371299 297258
rect 369380 297228 371238 297256
rect 369350 297200 371238 297228
rect 371294 297200 371299 297256
rect 369350 297198 371299 297200
rect 369350 296853 369410 297198
rect 371233 297195 371299 297198
rect 369301 296848 369410 296853
rect 369301 296792 369306 296848
rect 369362 296792 369410 296848
rect 369301 296790 369410 296792
rect 369301 296787 369367 296790
rect 199837 296714 199903 296717
rect 371233 296714 371299 296717
rect 199837 296712 200100 296714
rect 199837 296656 199842 296712
rect 199898 296656 200100 296712
rect 369380 296712 371299 296714
rect 369380 296684 371238 296712
rect 199837 296654 200100 296656
rect 369350 296656 371238 296684
rect 371294 296656 371299 296712
rect 369350 296654 371299 296656
rect 199837 296651 199903 296654
rect 369350 296309 369410 296654
rect 371233 296651 371299 296654
rect 445661 296442 445727 296445
rect 441876 296440 445727 296442
rect 441876 296384 445666 296440
rect 445722 296384 445727 296440
rect 441876 296382 445727 296384
rect 445661 296379 445727 296382
rect 369301 296304 369410 296309
rect 369301 296248 369306 296304
rect 369362 296248 369410 296304
rect 369301 296246 369410 296248
rect 369301 296243 369367 296246
rect 371233 296170 371299 296173
rect 369932 296168 371299 296170
rect 369932 296112 371238 296168
rect 371294 296112 371299 296168
rect 369932 296110 371299 296112
rect 371233 296107 371299 296110
rect 370221 295626 370287 295629
rect 369932 295624 370287 295626
rect 369932 295568 370226 295624
rect 370282 295568 370287 295624
rect 369932 295566 370287 295568
rect 370221 295563 370287 295566
rect 302417 295218 302483 295221
rect 445753 295218 445819 295221
rect 299828 295216 302483 295218
rect 299828 295160 302422 295216
rect 302478 295160 302483 295216
rect 299828 295158 302483 295160
rect 441876 295216 445819 295218
rect 441876 295160 445758 295216
rect 445814 295160 445819 295216
rect 441876 295158 445819 295160
rect 302417 295155 302483 295158
rect 445753 295155 445819 295158
rect 370129 295082 370195 295085
rect 369932 295080 370195 295082
rect 369932 295024 370134 295080
rect 370190 295024 370195 295080
rect 369932 295022 370195 295024
rect 370129 295019 370195 295022
rect 197905 294538 197971 294541
rect 372337 294538 372403 294541
rect 197905 294536 200100 294538
rect 197905 294480 197910 294536
rect 197966 294480 200100 294536
rect 197905 294478 200100 294480
rect 369932 294536 372403 294538
rect 369932 294480 372342 294536
rect 372398 294480 372403 294536
rect 369932 294478 372403 294480
rect 197905 294475 197971 294478
rect 372337 294475 372403 294478
rect 445661 294130 445727 294133
rect 441876 294128 445727 294130
rect 441876 294072 445666 294128
rect 445722 294072 445727 294128
rect 441876 294070 445727 294072
rect 445661 294067 445727 294070
rect 371233 293994 371299 293997
rect 369932 293992 371299 293994
rect 369932 293936 371238 293992
rect 371294 293936 371299 293992
rect 369932 293934 371299 293936
rect 371233 293931 371299 293934
rect 371233 293450 371299 293453
rect 369932 293448 371299 293450
rect 369932 293392 371238 293448
rect 371294 293392 371299 293448
rect 369932 293390 371299 293392
rect 371233 293387 371299 293390
rect -960 293178 480 293268
rect 2865 293178 2931 293181
rect -960 293176 2931 293178
rect -960 293120 2870 293176
rect 2926 293120 2931 293176
rect -960 293118 2931 293120
rect -960 293028 480 293118
rect 2865 293115 2931 293118
rect 371233 292906 371299 292909
rect 445661 292906 445727 292909
rect 369932 292904 371299 292906
rect 369932 292848 371238 292904
rect 371294 292848 371299 292904
rect 369932 292846 371299 292848
rect 441876 292904 445727 292906
rect 441876 292848 445666 292904
rect 445722 292848 445727 292904
rect 441876 292846 445727 292848
rect 371233 292843 371299 292846
rect 445661 292843 445727 292846
rect 198089 292362 198155 292365
rect 372337 292362 372403 292365
rect 198089 292360 200100 292362
rect 198089 292304 198094 292360
rect 198150 292304 200100 292360
rect 198089 292302 200100 292304
rect 369932 292360 372403 292362
rect 369932 292304 372342 292360
rect 372398 292304 372403 292360
rect 369932 292302 372403 292304
rect 198089 292299 198155 292302
rect 372337 292299 372403 292302
rect 302325 291954 302391 291957
rect 299828 291952 302391 291954
rect 299828 291896 302330 291952
rect 302386 291896 302391 291952
rect 299828 291894 302391 291896
rect 302325 291891 302391 291894
rect 371233 291818 371299 291821
rect 445661 291818 445727 291821
rect 369932 291816 371299 291818
rect 369932 291760 371238 291816
rect 371294 291760 371299 291816
rect 369932 291758 371299 291760
rect 441876 291816 445727 291818
rect 441876 291760 445666 291816
rect 445722 291760 445727 291816
rect 441876 291758 445727 291760
rect 371233 291755 371299 291758
rect 445661 291755 445727 291758
rect 371233 291274 371299 291277
rect 369932 291272 371299 291274
rect 369932 291216 371238 291272
rect 371294 291216 371299 291272
rect 369932 291214 371299 291216
rect 371233 291211 371299 291214
rect 372337 290730 372403 290733
rect 369932 290728 372403 290730
rect 369932 290672 372342 290728
rect 372398 290672 372403 290728
rect 369932 290670 372403 290672
rect 372337 290667 372403 290670
rect 445661 290594 445727 290597
rect 441876 290592 445727 290594
rect 441876 290536 445666 290592
rect 445722 290536 445727 290592
rect 441876 290534 445727 290536
rect 445661 290531 445727 290534
rect 197353 290186 197419 290189
rect 371233 290186 371299 290189
rect 197353 290184 200100 290186
rect 197353 290128 197358 290184
rect 197414 290128 200100 290184
rect 197353 290126 200100 290128
rect 369932 290184 371299 290186
rect 369932 290128 371238 290184
rect 371294 290128 371299 290184
rect 369932 290126 371299 290128
rect 197353 290123 197419 290126
rect 371233 290123 371299 290126
rect 372337 289642 372403 289645
rect 369932 289640 372403 289642
rect 369932 289584 372342 289640
rect 372398 289584 372403 289640
rect 369932 289582 372403 289584
rect 372337 289579 372403 289582
rect 445661 289506 445727 289509
rect 441876 289504 445727 289506
rect 441876 289448 445666 289504
rect 445722 289448 445727 289504
rect 441876 289446 445727 289448
rect 445661 289443 445727 289446
rect 371233 289098 371299 289101
rect 369932 289096 371299 289098
rect 369932 289040 371238 289096
rect 371294 289040 371299 289096
rect 369932 289038 371299 289040
rect 371233 289035 371299 289038
rect 302969 288826 303035 288829
rect 299828 288824 303035 288826
rect 299828 288768 302974 288824
rect 303030 288768 303035 288824
rect 299828 288766 303035 288768
rect 302969 288763 303035 288766
rect 372797 288554 372863 288557
rect 369932 288552 372863 288554
rect 369932 288496 372802 288552
rect 372858 288496 372863 288552
rect 369932 288494 372863 288496
rect 372797 288491 372863 288494
rect 445661 288282 445727 288285
rect 441876 288280 445727 288282
rect 441876 288224 445666 288280
rect 445722 288224 445727 288280
rect 441876 288222 445727 288224
rect 445661 288219 445727 288222
rect 372337 288146 372403 288149
rect 369932 288144 372403 288146
rect 369932 288088 372342 288144
rect 372398 288088 372403 288144
rect 369932 288086 372403 288088
rect 372337 288083 372403 288086
rect 197629 288010 197695 288013
rect 197629 288008 200100 288010
rect 197629 287952 197634 288008
rect 197690 287952 200100 288008
rect 197629 287950 200100 287952
rect 197629 287947 197695 287950
rect 371233 287602 371299 287605
rect 369932 287600 371299 287602
rect 369932 287544 371238 287600
rect 371294 287544 371299 287600
rect 369932 287542 371299 287544
rect 371233 287539 371299 287542
rect 445109 287194 445175 287197
rect 441876 287192 445175 287194
rect 441876 287136 445114 287192
rect 445170 287136 445175 287192
rect 441876 287134 445175 287136
rect 445109 287131 445175 287134
rect 372521 287058 372587 287061
rect 369932 287056 372587 287058
rect 369932 287000 372526 287056
rect 372582 287000 372587 287056
rect 369932 286998 372587 287000
rect 372521 286995 372587 286998
rect 371877 286514 371943 286517
rect 369932 286512 371943 286514
rect 369932 286456 371882 286512
rect 371938 286456 371943 286512
rect 369932 286454 371943 286456
rect 371877 286451 371943 286454
rect 371325 285970 371391 285973
rect 445661 285970 445727 285973
rect 369932 285968 371391 285970
rect 369932 285912 371330 285968
rect 371386 285912 371391 285968
rect 369932 285910 371391 285912
rect 441876 285968 445727 285970
rect 441876 285912 445666 285968
rect 445722 285912 445727 285968
rect 441876 285910 445727 285912
rect 371325 285907 371391 285910
rect 445661 285907 445727 285910
rect 197353 285834 197419 285837
rect 197353 285832 200100 285834
rect 197353 285776 197358 285832
rect 197414 285776 200100 285832
rect 197353 285774 200100 285776
rect 197353 285771 197419 285774
rect 302785 285698 302851 285701
rect 299828 285696 302851 285698
rect 299828 285640 302790 285696
rect 302846 285640 302851 285696
rect 299828 285638 302851 285640
rect 302785 285635 302851 285638
rect 371877 285426 371943 285429
rect 369932 285424 371943 285426
rect 369932 285368 371882 285424
rect 371938 285368 371943 285424
rect 369932 285366 371943 285368
rect 371877 285363 371943 285366
rect 583520 285276 584960 285516
rect 371877 284882 371943 284885
rect 445661 284882 445727 284885
rect 369932 284880 371943 284882
rect 369932 284824 371882 284880
rect 371938 284824 371943 284880
rect 369932 284822 371943 284824
rect 441876 284880 445727 284882
rect 441876 284824 445666 284880
rect 445722 284824 445727 284880
rect 441876 284822 445727 284824
rect 371877 284819 371943 284822
rect 445661 284819 445727 284822
rect 371877 284338 371943 284341
rect 369932 284336 371943 284338
rect 369932 284280 371882 284336
rect 371938 284280 371943 284336
rect 369932 284278 371943 284280
rect 371877 284275 371943 284278
rect 371877 283794 371943 283797
rect 369932 283792 371943 283794
rect 369932 283736 371882 283792
rect 371938 283736 371943 283792
rect 369932 283734 371943 283736
rect 371877 283731 371943 283734
rect 197353 283658 197419 283661
rect 445477 283658 445543 283661
rect 197353 283656 200100 283658
rect 197353 283600 197358 283656
rect 197414 283600 200100 283656
rect 197353 283598 200100 283600
rect 441876 283656 445543 283658
rect 441876 283600 445482 283656
rect 445538 283600 445543 283656
rect 441876 283598 445543 283600
rect 197353 283595 197419 283598
rect 445477 283595 445543 283598
rect 371877 283250 371943 283253
rect 369932 283248 371943 283250
rect 369932 283192 371882 283248
rect 371938 283192 371943 283248
rect 369932 283190 371943 283192
rect 371877 283187 371943 283190
rect 371877 282706 371943 282709
rect 369932 282704 371943 282706
rect 369932 282648 371882 282704
rect 371938 282648 371943 282704
rect 369932 282646 371943 282648
rect 371877 282643 371943 282646
rect 445385 282570 445451 282573
rect 441876 282568 445451 282570
rect 441876 282512 445390 282568
rect 445446 282512 445451 282568
rect 441876 282510 445451 282512
rect 445385 282507 445451 282510
rect 302417 282434 302483 282437
rect 299828 282432 302483 282434
rect 299828 282376 302422 282432
rect 302478 282376 302483 282432
rect 299828 282374 302483 282376
rect 302417 282371 302483 282374
rect 371877 282162 371943 282165
rect 369932 282160 371943 282162
rect 369932 282104 371882 282160
rect 371938 282104 371943 282160
rect 369932 282102 371943 282104
rect 371877 282099 371943 282102
rect 371366 281618 371372 281620
rect 369932 281558 371372 281618
rect 371366 281556 371372 281558
rect 371436 281618 371442 281620
rect 371918 281618 371924 281620
rect 371436 281558 371924 281618
rect 371436 281556 371442 281558
rect 371918 281556 371924 281558
rect 371988 281556 371994 281620
rect 197353 281482 197419 281485
rect 197353 281480 200100 281482
rect 197353 281424 197358 281480
rect 197414 281424 200100 281480
rect 197353 281422 200100 281424
rect 197353 281419 197419 281422
rect 445109 281346 445175 281349
rect 441876 281344 445175 281346
rect 441876 281288 445114 281344
rect 445170 281288 445175 281344
rect 441876 281286 445175 281288
rect 445109 281283 445175 281286
rect 371734 281074 371740 281076
rect 369932 281014 371740 281074
rect 371734 281012 371740 281014
rect 371804 281012 371810 281076
rect 372102 280530 372108 280532
rect 369932 280470 372108 280530
rect 372102 280468 372108 280470
rect 372172 280468 372178 280532
rect 444741 280258 444807 280261
rect 441876 280256 444807 280258
rect -960 279972 480 280212
rect 441876 280200 444746 280256
rect 444802 280200 444807 280256
rect 441876 280198 444807 280200
rect 444741 280195 444807 280198
rect 371233 279986 371299 279989
rect 372521 279986 372587 279989
rect 369932 279984 372587 279986
rect 369932 279928 371238 279984
rect 371294 279928 372526 279984
rect 372582 279928 372587 279984
rect 369932 279926 372587 279928
rect 371233 279923 371299 279926
rect 372521 279923 372587 279926
rect 371550 279442 371556 279444
rect 369932 279382 371556 279442
rect 371550 279380 371556 279382
rect 371620 279380 371626 279444
rect 197353 279306 197419 279309
rect 302601 279306 302667 279309
rect 197353 279304 200100 279306
rect 197353 279248 197358 279304
rect 197414 279248 200100 279304
rect 197353 279246 200100 279248
rect 299828 279304 302667 279306
rect 299828 279248 302606 279304
rect 302662 279248 302667 279304
rect 299828 279246 302667 279248
rect 197353 279243 197419 279246
rect 302601 279243 302667 279246
rect 444833 279034 444899 279037
rect 441876 279032 444899 279034
rect 441876 278976 444838 279032
rect 444894 278976 444899 279032
rect 441876 278974 444899 278976
rect 444833 278971 444899 278974
rect 371182 278898 371188 278900
rect 369932 278838 371188 278898
rect 371182 278836 371188 278838
rect 371252 278836 371258 278900
rect 372337 278354 372403 278357
rect 369932 278352 372403 278354
rect 369932 278296 372342 278352
rect 372398 278296 372403 278352
rect 369932 278294 372403 278296
rect 372337 278291 372403 278294
rect 372153 277946 372219 277949
rect 445109 277946 445175 277949
rect 369932 277944 372219 277946
rect 369932 277888 372158 277944
rect 372214 277888 372219 277944
rect 369932 277886 372219 277888
rect 441876 277944 445175 277946
rect 441876 277888 445114 277944
rect 445170 277888 445175 277944
rect 441876 277886 445175 277888
rect 372153 277883 372219 277886
rect 445109 277883 445175 277886
rect 370313 277402 370379 277405
rect 369932 277400 370379 277402
rect 369932 277372 370318 277400
rect 369902 277344 370318 277372
rect 370374 277344 370379 277400
rect 369902 277342 370379 277344
rect 197537 277130 197603 277133
rect 369301 277130 369367 277133
rect 197537 277128 200100 277130
rect 197537 277072 197542 277128
rect 197598 277072 200100 277128
rect 197537 277070 200100 277072
rect 369301 277128 369410 277130
rect 369301 277072 369306 277128
rect 369362 277072 369410 277128
rect 197537 277067 197603 277070
rect 369301 277067 369410 277072
rect 369350 276828 369410 277067
rect 369902 276994 369962 277342
rect 370313 277339 370379 277342
rect 370078 276994 370084 276996
rect 369902 276934 370084 276994
rect 370078 276932 370084 276934
rect 370148 276932 370154 276996
rect 444557 276722 444623 276725
rect 441876 276720 444623 276722
rect 441876 276664 444562 276720
rect 444618 276664 444623 276720
rect 441876 276662 444623 276664
rect 444557 276659 444623 276662
rect 371601 276314 371667 276317
rect 369932 276312 371667 276314
rect 369932 276256 371606 276312
rect 371662 276256 371667 276312
rect 369932 276254 371667 276256
rect 371601 276251 371667 276254
rect 303061 276178 303127 276181
rect 299828 276176 303127 276178
rect 299828 276120 303066 276176
rect 303122 276120 303127 276176
rect 299828 276118 303127 276120
rect 303061 276115 303127 276118
rect 370497 275770 370563 275773
rect 369932 275768 370563 275770
rect 369932 275740 370502 275768
rect 369902 275712 370502 275740
rect 370558 275712 370563 275768
rect 369902 275710 370563 275712
rect 369902 275362 369962 275710
rect 370497 275707 370563 275710
rect 444465 275634 444531 275637
rect 441876 275632 444531 275634
rect 441876 275576 444470 275632
rect 444526 275576 444531 275632
rect 441876 275574 444531 275576
rect 444465 275571 444531 275574
rect 370262 275362 370268 275364
rect 369902 275302 370268 275362
rect 370262 275300 370268 275302
rect 370332 275300 370338 275364
rect 370681 275226 370747 275229
rect 369932 275224 370747 275226
rect 369932 275196 370686 275224
rect 369902 275168 370686 275196
rect 370742 275168 370747 275224
rect 369902 275166 370747 275168
rect 198365 274954 198431 274957
rect 369902 274954 369962 275166
rect 370681 275163 370747 275166
rect 370037 274954 370103 274957
rect 198365 274952 200100 274954
rect 198365 274896 198370 274952
rect 198426 274896 200100 274952
rect 198365 274894 200100 274896
rect 369902 274952 370103 274954
rect 369902 274896 370042 274952
rect 370098 274896 370103 274952
rect 369902 274894 370103 274896
rect 198365 274891 198431 274894
rect 370037 274891 370103 274894
rect 372613 274682 372679 274685
rect 369932 274680 372679 274682
rect 369932 274624 372618 274680
rect 372674 274624 372679 274680
rect 369932 274622 372679 274624
rect 372613 274619 372679 274622
rect 445661 274410 445727 274413
rect 441876 274408 445727 274410
rect 441876 274352 445666 274408
rect 445722 274352 445727 274408
rect 441876 274350 445727 274352
rect 445661 274347 445727 274350
rect 370589 274138 370655 274141
rect 370773 274138 370839 274141
rect 369932 274136 370839 274138
rect 369932 274080 370594 274136
rect 370650 274080 370778 274136
rect 370834 274080 370839 274136
rect 369932 274078 370839 274080
rect 370589 274075 370655 274078
rect 370773 274075 370839 274078
rect 369945 273866 370011 273869
rect 369902 273864 370011 273866
rect 369902 273808 369950 273864
rect 370006 273808 370011 273864
rect 369902 273803 370011 273808
rect 369902 273594 369962 273803
rect 371049 273594 371115 273597
rect 369902 273592 371115 273594
rect 369902 273564 371054 273592
rect 369932 273536 371054 273564
rect 371110 273536 371115 273592
rect 369932 273534 371115 273536
rect 371049 273531 371115 273534
rect 445569 273322 445635 273325
rect 441876 273320 445635 273322
rect 441876 273264 445574 273320
rect 445630 273264 445635 273320
rect 441876 273262 445635 273264
rect 445569 273259 445635 273262
rect 371969 273050 372035 273053
rect 369932 273048 372035 273050
rect 369932 272992 371974 273048
rect 372030 272992 372035 273048
rect 369932 272990 372035 272992
rect 371969 272987 372035 272990
rect 302877 272914 302943 272917
rect 299828 272912 302943 272914
rect 299828 272856 302882 272912
rect 302938 272856 302943 272912
rect 299828 272854 302943 272856
rect 302877 272851 302943 272854
rect 197353 272778 197419 272781
rect 197353 272776 200100 272778
rect 197353 272720 197358 272776
rect 197414 272720 200100 272776
rect 197353 272718 200100 272720
rect 197353 272715 197419 272718
rect 372245 272506 372311 272509
rect 369932 272504 372311 272506
rect 369932 272448 372250 272504
rect 372306 272448 372311 272504
rect 369932 272446 372311 272448
rect 372245 272443 372311 272446
rect 580257 272234 580323 272237
rect 583520 272234 584960 272324
rect 580257 272232 584960 272234
rect 580257 272176 580262 272232
rect 580318 272176 584960 272232
rect 580257 272174 584960 272176
rect 580257 272171 580323 272174
rect 445661 272098 445727 272101
rect 441876 272096 445727 272098
rect 441876 272040 445666 272096
rect 445722 272040 445727 272096
rect 583520 272084 584960 272174
rect 441876 272038 445727 272040
rect 445661 272035 445727 272038
rect 371785 271962 371851 271965
rect 369932 271960 371851 271962
rect 369932 271904 371790 271960
rect 371846 271904 371851 271960
rect 369932 271902 371851 271904
rect 371785 271899 371851 271902
rect 371417 271690 371483 271693
rect 371877 271690 371943 271693
rect 369902 271688 371943 271690
rect 369902 271632 371422 271688
rect 371478 271632 371882 271688
rect 371938 271632 371943 271688
rect 369902 271630 371943 271632
rect 369902 271388 369962 271630
rect 371417 271627 371483 271630
rect 371877 271627 371943 271630
rect 445661 271010 445727 271013
rect 441876 271008 445727 271010
rect 441876 270952 445666 271008
rect 445722 270952 445727 271008
rect 441876 270950 445727 270952
rect 445661 270947 445727 270950
rect 372061 270874 372127 270877
rect 369932 270872 372127 270874
rect 369932 270816 372066 270872
rect 372122 270816 372127 270872
rect 369932 270814 372127 270816
rect 372061 270811 372127 270814
rect 197353 270602 197419 270605
rect 197353 270600 200100 270602
rect 197353 270544 197358 270600
rect 197414 270544 200100 270600
rect 197353 270542 200100 270544
rect 197353 270539 197419 270542
rect 371601 270330 371667 270333
rect 372429 270330 372495 270333
rect 369932 270328 372495 270330
rect 369932 270272 371606 270328
rect 371662 270272 372434 270328
rect 372490 270272 372495 270328
rect 369932 270270 372495 270272
rect 371601 270267 371667 270270
rect 372429 270267 372495 270270
rect 302325 269786 302391 269789
rect 371509 269786 371575 269789
rect 372337 269786 372403 269789
rect 445661 269786 445727 269789
rect 299828 269784 302391 269786
rect 299828 269728 302330 269784
rect 302386 269728 302391 269784
rect 299828 269726 302391 269728
rect 369932 269784 372403 269786
rect 369932 269728 371514 269784
rect 371570 269728 372342 269784
rect 372398 269728 372403 269784
rect 369932 269726 372403 269728
rect 441876 269784 445727 269786
rect 441876 269728 445666 269784
rect 445722 269728 445727 269784
rect 441876 269726 445727 269728
rect 302325 269723 302391 269726
rect 371509 269723 371575 269726
rect 372337 269723 372403 269726
rect 445661 269723 445727 269726
rect 371233 269242 371299 269245
rect 369932 269240 371299 269242
rect 369932 269184 371238 269240
rect 371294 269184 371299 269240
rect 369932 269182 371299 269184
rect 371233 269179 371299 269182
rect 372153 268698 372219 268701
rect 445661 268698 445727 268701
rect 369932 268696 372219 268698
rect 369932 268640 372158 268696
rect 372214 268640 372219 268696
rect 369932 268638 372219 268640
rect 441876 268696 445727 268698
rect 441876 268640 445666 268696
rect 445722 268640 445727 268696
rect 441876 268638 445727 268640
rect 372153 268635 372219 268638
rect 445661 268635 445727 268638
rect 197721 268426 197787 268429
rect 197721 268424 200100 268426
rect 197721 268368 197726 268424
rect 197782 268368 200100 268424
rect 197721 268366 200100 268368
rect 197721 268363 197787 268366
rect 370405 268290 370471 268293
rect 369932 268288 370471 268290
rect 369932 268232 370410 268288
rect 370466 268232 370471 268288
rect 369932 268230 370471 268232
rect 370405 268227 370471 268230
rect 361614 267820 361620 267884
rect 361684 267882 361690 267884
rect 362861 267882 362927 267885
rect 361684 267880 362927 267882
rect 361684 267824 362866 267880
rect 362922 267824 362927 267880
rect 361684 267822 362927 267824
rect 361684 267820 361690 267822
rect 362861 267819 362927 267822
rect -960 267202 480 267292
rect 3233 267202 3299 267205
rect -960 267200 3299 267202
rect -960 267144 3238 267200
rect 3294 267144 3299 267200
rect -960 267142 3299 267144
rect -960 267052 480 267142
rect 3233 267139 3299 267142
rect 302417 266658 302483 266661
rect 299828 266656 302483 266658
rect 299828 266600 302422 266656
rect 302478 266600 302483 266656
rect 299828 266598 302483 266600
rect 302417 266595 302483 266598
rect 197353 266250 197419 266253
rect 353937 266250 354003 266253
rect 364374 266250 364380 266252
rect 197353 266248 200100 266250
rect 197353 266192 197358 266248
rect 197414 266192 200100 266248
rect 197353 266190 200100 266192
rect 353937 266248 364380 266250
rect 353937 266192 353942 266248
rect 353998 266192 364380 266248
rect 353937 266190 364380 266192
rect 197353 266187 197419 266190
rect 353937 266187 354003 266190
rect 364374 266188 364380 266190
rect 364444 266250 364450 266252
rect 364885 266250 364951 266253
rect 364444 266248 364951 266250
rect 364444 266192 364890 266248
rect 364946 266192 364951 266248
rect 364444 266190 364951 266192
rect 364444 266188 364450 266190
rect 364885 266187 364951 266190
rect 356697 266114 356763 266117
rect 361614 266114 361620 266116
rect 356697 266112 361620 266114
rect 356697 266056 356702 266112
rect 356758 266056 361620 266112
rect 356697 266054 361620 266056
rect 356697 266051 356763 266054
rect 361614 266052 361620 266054
rect 361684 266052 361690 266116
rect 197905 264074 197971 264077
rect 197905 264072 200100 264074
rect 197905 264016 197910 264072
rect 197966 264016 200100 264072
rect 197905 264014 200100 264016
rect 197905 264011 197971 264014
rect 302509 263394 302575 263397
rect 299828 263392 302575 263394
rect 299828 263336 302514 263392
rect 302570 263336 302575 263392
rect 299828 263334 302575 263336
rect 302509 263331 302575 263334
rect 198641 261898 198707 261901
rect 198641 261896 200100 261898
rect 198641 261840 198646 261896
rect 198702 261840 200100 261896
rect 198641 261838 200100 261840
rect 198641 261835 198707 261838
rect 302785 260266 302851 260269
rect 299828 260264 302851 260266
rect 299828 260208 302790 260264
rect 302846 260208 302851 260264
rect 299828 260206 302851 260208
rect 302785 260203 302851 260206
rect 197721 259722 197787 259725
rect 197721 259720 200100 259722
rect 197721 259664 197726 259720
rect 197782 259664 200100 259720
rect 197721 259662 200100 259664
rect 197721 259659 197787 259662
rect 580165 258906 580231 258909
rect 583520 258906 584960 258996
rect 580165 258904 584960 258906
rect 580165 258848 580170 258904
rect 580226 258848 584960 258904
rect 580165 258846 584960 258848
rect 580165 258843 580231 258846
rect 583520 258756 584960 258846
rect 198089 257546 198155 257549
rect 198089 257544 200100 257546
rect 198089 257488 198094 257544
rect 198150 257488 200100 257544
rect 198089 257486 200100 257488
rect 198089 257483 198155 257486
rect 302785 257138 302851 257141
rect 299828 257136 302851 257138
rect 299828 257080 302790 257136
rect 302846 257080 302851 257136
rect 299828 257078 302851 257080
rect 302785 257075 302851 257078
rect 197353 255370 197419 255373
rect 197353 255368 200100 255370
rect 197353 255312 197358 255368
rect 197414 255312 200100 255368
rect 197353 255310 200100 255312
rect 197353 255307 197419 255310
rect -960 254146 480 254236
rect 3601 254146 3667 254149
rect -960 254144 3667 254146
rect -960 254088 3606 254144
rect 3662 254088 3667 254144
rect -960 254086 3667 254088
rect -960 253996 480 254086
rect 3601 254083 3667 254086
rect 302877 253874 302943 253877
rect 299828 253872 302943 253874
rect 299828 253816 302882 253872
rect 302938 253816 302943 253872
rect 299828 253814 302943 253816
rect 302877 253811 302943 253814
rect 197353 253194 197419 253197
rect 197353 253192 200100 253194
rect 197353 253136 197358 253192
rect 197414 253136 200100 253192
rect 197353 253134 200100 253136
rect 197353 253131 197419 253134
rect 197997 251018 198063 251021
rect 197997 251016 200100 251018
rect 197997 250960 198002 251016
rect 198058 250960 200100 251016
rect 197997 250958 200100 250960
rect 197997 250955 198063 250958
rect 303153 250746 303219 250749
rect 299828 250744 303219 250746
rect 299828 250688 303158 250744
rect 303214 250688 303219 250744
rect 299828 250686 303219 250688
rect 303153 250683 303219 250686
rect 198181 248842 198247 248845
rect 198181 248840 200100 248842
rect 198181 248784 198186 248840
rect 198242 248784 200100 248840
rect 198181 248782 200100 248784
rect 198181 248779 198247 248782
rect 303061 247618 303127 247621
rect 299828 247616 303127 247618
rect 299828 247560 303066 247616
rect 303122 247560 303127 247616
rect 299828 247558 303127 247560
rect 303061 247555 303127 247558
rect 198089 246666 198155 246669
rect 198089 246664 200100 246666
rect 198089 246608 198094 246664
rect 198150 246608 200100 246664
rect 198089 246606 200100 246608
rect 198089 246603 198155 246606
rect 580165 245578 580231 245581
rect 583520 245578 584960 245668
rect 580165 245576 584960 245578
rect 580165 245520 580170 245576
rect 580226 245520 584960 245576
rect 580165 245518 584960 245520
rect 580165 245515 580231 245518
rect 583520 245428 584960 245518
rect 197353 244490 197419 244493
rect 197353 244488 200100 244490
rect 197353 244432 197358 244488
rect 197414 244432 200100 244488
rect 197353 244430 200100 244432
rect 197353 244427 197419 244430
rect 302969 244354 303035 244357
rect 299828 244352 303035 244354
rect 299828 244296 302974 244352
rect 303030 244296 303035 244352
rect 299828 244294 303035 244296
rect 302969 244291 303035 244294
rect 197721 242314 197787 242317
rect 197721 242312 200100 242314
rect 197721 242256 197726 242312
rect 197782 242256 200100 242312
rect 197721 242254 200100 242256
rect 197721 242251 197787 242254
rect 302785 241226 302851 241229
rect 299828 241224 302851 241226
rect -960 241090 480 241180
rect 299828 241168 302790 241224
rect 302846 241168 302851 241224
rect 299828 241166 302851 241168
rect 302785 241163 302851 241166
rect 3509 241090 3575 241093
rect -960 241088 3575 241090
rect -960 241032 3514 241088
rect 3570 241032 3575 241088
rect -960 241030 3575 241032
rect -960 240940 480 241030
rect 3509 241027 3575 241030
rect 197353 240138 197419 240141
rect 197353 240136 200100 240138
rect 197353 240080 197358 240136
rect 197414 240080 200100 240136
rect 197353 240078 200100 240080
rect 197353 240075 197419 240078
rect 303153 238098 303219 238101
rect 299828 238096 303219 238098
rect 299828 238040 303158 238096
rect 303214 238040 303219 238096
rect 299828 238038 303219 238040
rect 303153 238035 303219 238038
rect 197353 237962 197419 237965
rect 197353 237960 200100 237962
rect 197353 237904 197358 237960
rect 197414 237904 200100 237960
rect 197353 237902 200100 237904
rect 197353 237899 197419 237902
rect 197537 235786 197603 235789
rect 197537 235784 200100 235786
rect 197537 235728 197542 235784
rect 197598 235728 200100 235784
rect 197537 235726 200100 235728
rect 197537 235723 197603 235726
rect 303245 234834 303311 234837
rect 299828 234832 303311 234834
rect 299828 234776 303250 234832
rect 303306 234776 303311 234832
rect 299828 234774 303311 234776
rect 303245 234771 303311 234774
rect 198181 233610 198247 233613
rect 198181 233608 200100 233610
rect 198181 233552 198186 233608
rect 198242 233552 200100 233608
rect 198181 233550 200100 233552
rect 198181 233547 198247 233550
rect 579981 232386 580047 232389
rect 583520 232386 584960 232476
rect 579981 232384 584960 232386
rect 579981 232328 579986 232384
rect 580042 232328 584960 232384
rect 579981 232326 584960 232328
rect 579981 232323 580047 232326
rect 583520 232236 584960 232326
rect 302877 231706 302943 231709
rect 299828 231704 302943 231706
rect 299828 231648 302882 231704
rect 302938 231648 302943 231704
rect 299828 231646 302943 231648
rect 302877 231643 302943 231646
rect 197629 231434 197695 231437
rect 197629 231432 200100 231434
rect 197629 231376 197634 231432
rect 197690 231376 200100 231432
rect 197629 231374 200100 231376
rect 197629 231371 197695 231374
rect 197353 229258 197419 229261
rect 197353 229256 200100 229258
rect 197353 229200 197358 229256
rect 197414 229200 200100 229256
rect 197353 229198 200100 229200
rect 197353 229195 197419 229198
rect 302785 228442 302851 228445
rect 299828 228440 302851 228442
rect 299828 228384 302790 228440
rect 302846 228384 302851 228440
rect 299828 228382 302851 228384
rect 302785 228379 302851 228382
rect -960 227884 480 228124
rect 198733 227082 198799 227085
rect 198733 227080 200100 227082
rect 198733 227024 198738 227080
rect 198794 227024 200100 227080
rect 198733 227022 200100 227024
rect 198733 227019 198799 227022
rect 371601 225722 371667 225725
rect 369932 225720 371667 225722
rect 369932 225664 371606 225720
rect 371662 225664 371667 225720
rect 369932 225662 371667 225664
rect 371601 225659 371667 225662
rect 445569 225450 445635 225453
rect 441876 225448 445635 225450
rect 441876 225420 445574 225448
rect 441846 225392 445574 225420
rect 445630 225392 445635 225448
rect 441846 225390 445635 225392
rect 302785 225314 302851 225317
rect 299828 225312 302851 225314
rect 299828 225256 302790 225312
rect 302846 225256 302851 225312
rect 299828 225254 302851 225256
rect 302785 225251 302851 225254
rect 371601 225178 371667 225181
rect 369932 225176 371667 225178
rect 369932 225120 371606 225176
rect 371662 225120 371667 225176
rect 369932 225118 371667 225120
rect 371601 225115 371667 225118
rect 441846 225045 441906 225390
rect 445569 225387 445635 225390
rect 371366 224980 371372 225044
rect 371436 225042 371442 225044
rect 372705 225042 372771 225045
rect 371436 225040 372771 225042
rect 371436 224984 372710 225040
rect 372766 224984 372771 225040
rect 371436 224982 372771 224984
rect 371436 224980 371442 224982
rect 372705 224979 372771 224982
rect 441797 225040 441906 225045
rect 441797 224984 441802 225040
rect 441858 224984 441906 225040
rect 441797 224982 441906 224984
rect 441797 224979 441863 224982
rect 198273 224906 198339 224909
rect 198273 224904 200100 224906
rect 198273 224848 198278 224904
rect 198334 224848 200100 224904
rect 198273 224846 200100 224848
rect 198273 224843 198339 224846
rect 371601 224634 371667 224637
rect 369932 224632 371667 224634
rect 369932 224576 371606 224632
rect 371662 224576 371667 224632
rect 369932 224574 371667 224576
rect 371601 224571 371667 224574
rect 372245 224090 372311 224093
rect 369932 224088 372311 224090
rect 369932 224032 372250 224088
rect 372306 224032 372311 224088
rect 369932 224030 372311 224032
rect 372245 224027 372311 224030
rect 441846 223957 441906 224332
rect 371734 223892 371740 223956
rect 371804 223954 371810 223956
rect 372705 223954 372771 223957
rect 371804 223952 372771 223954
rect 371804 223896 372710 223952
rect 372766 223896 372771 223952
rect 371804 223894 372771 223896
rect 371804 223892 371810 223894
rect 372705 223891 372771 223894
rect 441797 223952 441906 223957
rect 441797 223896 441802 223952
rect 441858 223896 441906 223952
rect 441797 223894 441906 223896
rect 441797 223891 441863 223894
rect 371601 223546 371667 223549
rect 369932 223544 371667 223546
rect 369932 223488 371606 223544
rect 371662 223488 371667 223544
rect 369932 223486 371667 223488
rect 371601 223483 371667 223486
rect 445661 223138 445727 223141
rect 441876 223136 445727 223138
rect 441876 223080 445666 223136
rect 445722 223080 445727 223136
rect 441876 223078 445727 223080
rect 445661 223075 445727 223078
rect 371601 223002 371667 223005
rect 369932 223000 371667 223002
rect 369932 222944 371606 223000
rect 371662 222944 371667 223000
rect 369932 222942 371667 222944
rect 371601 222939 371667 222942
rect 197353 222730 197419 222733
rect 197353 222728 200100 222730
rect 197353 222672 197358 222728
rect 197414 222672 200100 222728
rect 197353 222670 200100 222672
rect 197353 222667 197419 222670
rect 371417 222458 371483 222461
rect 369932 222456 371483 222458
rect 369932 222400 371422 222456
rect 371478 222400 371483 222456
rect 369932 222398 371483 222400
rect 371417 222395 371483 222398
rect 302785 222186 302851 222189
rect 299828 222184 302851 222186
rect 299828 222128 302790 222184
rect 302846 222128 302851 222184
rect 299828 222126 302851 222128
rect 302785 222123 302851 222126
rect 445661 222050 445727 222053
rect 441876 222048 445727 222050
rect 441876 221992 445666 222048
rect 445722 221992 445727 222048
rect 441876 221990 445727 221992
rect 445661 221987 445727 221990
rect 370497 221914 370563 221917
rect 369932 221912 370563 221914
rect 369932 221856 370502 221912
rect 370558 221856 370563 221912
rect 369932 221854 370563 221856
rect 370497 221851 370563 221854
rect 370405 221370 370471 221373
rect 369932 221368 370471 221370
rect 369932 221312 370410 221368
rect 370466 221312 370471 221368
rect 369932 221310 370471 221312
rect 370405 221307 370471 221310
rect 445661 220826 445727 220829
rect 441876 220824 445727 220826
rect 369350 220693 369410 220796
rect 441876 220768 445666 220824
rect 445722 220768 445727 220824
rect 441876 220766 445727 220768
rect 445661 220763 445727 220766
rect 369301 220688 369410 220693
rect 369301 220632 369306 220688
rect 369362 220632 369410 220688
rect 369301 220630 369410 220632
rect 369301 220627 369367 220630
rect 197537 220554 197603 220557
rect 369393 220554 369459 220557
rect 197537 220552 200100 220554
rect 197537 220496 197542 220552
rect 197598 220496 200100 220552
rect 197537 220494 200100 220496
rect 369350 220552 369459 220554
rect 369350 220496 369398 220552
rect 369454 220496 369459 220552
rect 197537 220491 197603 220494
rect 369350 220491 369459 220496
rect 369350 220252 369410 220491
rect 369853 220146 369919 220149
rect 369853 220144 369962 220146
rect 369853 220088 369858 220144
rect 369914 220088 369962 220144
rect 369853 220083 369962 220088
rect 369902 219708 369962 220083
rect 445661 219738 445727 219741
rect 441876 219736 445727 219738
rect 441876 219680 445666 219736
rect 445722 219680 445727 219736
rect 441876 219678 445727 219680
rect 445661 219675 445727 219678
rect 369902 219061 369962 219164
rect 369853 219056 369962 219061
rect 369853 219000 369858 219056
rect 369914 219000 369962 219056
rect 369853 218998 369962 219000
rect 580257 219058 580323 219061
rect 583520 219058 584960 219148
rect 580257 219056 584960 219058
rect 580257 219000 580262 219056
rect 580318 219000 584960 219056
rect 580257 218998 584960 219000
rect 369853 218995 369919 218998
rect 580257 218995 580323 218998
rect 302785 218922 302851 218925
rect 369945 218922 370011 218925
rect 299828 218920 302851 218922
rect 299828 218864 302790 218920
rect 302846 218864 302851 218920
rect 299828 218862 302851 218864
rect 302785 218859 302851 218862
rect 369902 218920 370011 218922
rect 369902 218864 369950 218920
rect 370006 218864 370011 218920
rect 583520 218908 584960 218998
rect 369902 218859 370011 218864
rect 369902 218620 369962 218859
rect 370037 218514 370103 218517
rect 445477 218514 445543 218517
rect 369902 218512 370103 218514
rect 369902 218456 370042 218512
rect 370098 218456 370103 218512
rect 369902 218454 370103 218456
rect 441876 218512 445543 218514
rect 441876 218456 445482 218512
rect 445538 218456 445543 218512
rect 441876 218454 445543 218456
rect 198457 218378 198523 218381
rect 198457 218376 200100 218378
rect 198457 218320 198462 218376
rect 198518 218320 200100 218376
rect 198457 218318 200100 218320
rect 198457 218315 198523 218318
rect 369902 218076 369962 218454
rect 370037 218451 370103 218454
rect 445477 218451 445543 218454
rect 370405 217562 370471 217565
rect 369932 217560 370471 217562
rect 369932 217504 370410 217560
rect 370466 217504 370471 217560
rect 369932 217502 370471 217504
rect 370405 217499 370471 217502
rect 445661 217426 445727 217429
rect 441876 217424 445727 217426
rect 441876 217368 445666 217424
rect 445722 217368 445727 217424
rect 441876 217366 445727 217368
rect 445661 217363 445727 217366
rect 370313 217018 370379 217021
rect 369932 217016 370379 217018
rect 369932 216960 370318 217016
rect 370374 216960 370379 217016
rect 369932 216958 370379 216960
rect 370313 216955 370379 216958
rect 372061 216474 372127 216477
rect 369932 216472 372127 216474
rect 369932 216416 372066 216472
rect 372122 216416 372127 216472
rect 369932 216414 372127 216416
rect 372061 216411 372127 216414
rect 197905 216202 197971 216205
rect 445661 216202 445727 216205
rect 197905 216200 200100 216202
rect 197905 216144 197910 216200
rect 197966 216144 200100 216200
rect 197905 216142 200100 216144
rect 441876 216200 445727 216202
rect 441876 216144 445666 216200
rect 445722 216144 445727 216200
rect 441876 216142 445727 216144
rect 197905 216139 197971 216142
rect 445661 216139 445727 216142
rect 371601 216066 371667 216069
rect 369932 216064 371667 216066
rect 369932 216008 371606 216064
rect 371662 216008 371667 216064
rect 369932 216006 371667 216008
rect 371601 216003 371667 216006
rect 302785 215794 302851 215797
rect 299828 215792 302851 215794
rect 299828 215736 302790 215792
rect 302846 215736 302851 215792
rect 299828 215734 302851 215736
rect 302785 215731 302851 215734
rect 371601 215522 371667 215525
rect 369932 215520 371667 215522
rect 369932 215464 371606 215520
rect 371662 215464 371667 215520
rect 369932 215462 371667 215464
rect 371601 215459 371667 215462
rect 445477 215114 445543 215117
rect 441876 215112 445543 215114
rect -960 214978 480 215068
rect 441876 215056 445482 215112
rect 445538 215056 445543 215112
rect 441876 215054 445543 215056
rect 445477 215051 445543 215054
rect 3325 214978 3391 214981
rect 371693 214978 371759 214981
rect -960 214976 3391 214978
rect -960 214920 3330 214976
rect 3386 214920 3391 214976
rect -960 214918 3391 214920
rect 369932 214976 371759 214978
rect 369932 214920 371698 214976
rect 371754 214920 371759 214976
rect 369932 214918 371759 214920
rect -960 214828 480 214918
rect 3325 214915 3391 214918
rect 371693 214915 371759 214918
rect 371601 214434 371667 214437
rect 369932 214432 371667 214434
rect 369932 214376 371606 214432
rect 371662 214376 371667 214432
rect 369932 214374 371667 214376
rect 371601 214371 371667 214374
rect 197353 214026 197419 214029
rect 197353 214024 200100 214026
rect 197353 213968 197358 214024
rect 197414 213968 200100 214024
rect 197353 213966 200100 213968
rect 197353 213963 197419 213966
rect 371417 213890 371483 213893
rect 445661 213890 445727 213893
rect 369932 213888 371483 213890
rect 369932 213832 371422 213888
rect 371478 213832 371483 213888
rect 369932 213830 371483 213832
rect 441876 213888 445727 213890
rect 441876 213832 445666 213888
rect 445722 213832 445727 213888
rect 441876 213830 445727 213832
rect 371417 213827 371483 213830
rect 445661 213827 445727 213830
rect 371601 213346 371667 213349
rect 369932 213344 371667 213346
rect 369932 213288 371606 213344
rect 371662 213288 371667 213344
rect 369932 213286 371667 213288
rect 371601 213283 371667 213286
rect 371693 212802 371759 212805
rect 445661 212802 445727 212805
rect 369932 212800 371759 212802
rect 369932 212744 371698 212800
rect 371754 212744 371759 212800
rect 369932 212742 371759 212744
rect 441876 212800 445727 212802
rect 441876 212744 445666 212800
rect 445722 212744 445727 212800
rect 441876 212742 445727 212744
rect 371693 212739 371759 212742
rect 445661 212739 445727 212742
rect 302785 212666 302851 212669
rect 299828 212664 302851 212666
rect 299828 212608 302790 212664
rect 302846 212608 302851 212664
rect 299828 212606 302851 212608
rect 302785 212603 302851 212606
rect 370221 212258 370287 212261
rect 369932 212256 370287 212258
rect 369932 212200 370226 212256
rect 370282 212200 370287 212256
rect 369932 212198 370287 212200
rect 370221 212195 370287 212198
rect 197721 211850 197787 211853
rect 197721 211848 200100 211850
rect 197721 211792 197726 211848
rect 197782 211792 200100 211848
rect 197721 211790 200100 211792
rect 197721 211787 197787 211790
rect 370957 211714 371023 211717
rect 371417 211714 371483 211717
rect 369932 211712 371483 211714
rect 369932 211656 370962 211712
rect 371018 211656 371422 211712
rect 371478 211656 371483 211712
rect 369932 211654 371483 211656
rect 370957 211651 371023 211654
rect 371417 211651 371483 211654
rect 445477 211578 445543 211581
rect 441876 211576 445543 211578
rect 441876 211520 445482 211576
rect 445538 211520 445543 211576
rect 441876 211518 445543 211520
rect 445477 211515 445543 211518
rect 373165 211170 373231 211173
rect 369932 211168 373231 211170
rect 369932 211112 373170 211168
rect 373226 211112 373231 211168
rect 369932 211110 373231 211112
rect 373165 211107 373231 211110
rect 373073 210626 373139 210629
rect 369932 210624 373139 210626
rect 369932 210568 373078 210624
rect 373134 210568 373139 210624
rect 369932 210566 373139 210568
rect 373073 210563 373139 210566
rect 445385 210490 445451 210493
rect 441876 210488 445451 210490
rect 441876 210432 445390 210488
rect 445446 210432 445451 210488
rect 441876 210430 445451 210432
rect 445385 210427 445451 210430
rect 370129 210082 370195 210085
rect 369932 210080 370195 210082
rect 369932 210024 370134 210080
rect 370190 210024 370195 210080
rect 369932 210022 370195 210024
rect 370129 210019 370195 210022
rect 197353 209674 197419 209677
rect 197353 209672 200100 209674
rect 197353 209616 197358 209672
rect 197414 209616 200100 209672
rect 197353 209614 200100 209616
rect 197353 209611 197419 209614
rect 371366 209538 371372 209540
rect 369932 209508 371372 209538
rect 369902 209478 371372 209508
rect 302877 209402 302943 209405
rect 299828 209400 302943 209402
rect 299828 209344 302882 209400
rect 302938 209344 302943 209400
rect 299828 209342 302943 209344
rect 302877 209339 302943 209342
rect 369902 209269 369962 209478
rect 371366 209476 371372 209478
rect 371436 209476 371442 209540
rect 369853 209264 369962 209269
rect 445201 209266 445267 209269
rect 369853 209208 369858 209264
rect 369914 209208 369962 209264
rect 369853 209206 369962 209208
rect 441876 209264 445267 209266
rect 441876 209208 445206 209264
rect 445262 209208 445267 209264
rect 441876 209206 445267 209208
rect 369853 209203 369919 209206
rect 445201 209203 445267 209206
rect 370497 208994 370563 208997
rect 371734 208994 371740 208996
rect 369932 208992 371740 208994
rect 369932 208936 370502 208992
rect 370558 208936 371740 208992
rect 369932 208934 371740 208936
rect 370497 208931 370563 208934
rect 371734 208932 371740 208934
rect 371804 208932 371810 208996
rect 370865 208450 370931 208453
rect 371918 208450 371924 208452
rect 369932 208448 371924 208450
rect 369932 208392 370870 208448
rect 370926 208392 371924 208448
rect 369932 208390 371924 208392
rect 370865 208387 370931 208390
rect 371918 208388 371924 208390
rect 371988 208388 371994 208452
rect 444741 208178 444807 208181
rect 441876 208176 444807 208178
rect 441876 208120 444746 208176
rect 444802 208120 444807 208176
rect 441876 208118 444807 208120
rect 444741 208115 444807 208118
rect 371693 207906 371759 207909
rect 372521 207906 372587 207909
rect 369932 207904 372587 207906
rect 369932 207848 371698 207904
rect 371754 207848 372526 207904
rect 372582 207848 372587 207904
rect 369932 207846 372587 207848
rect 371693 207843 371759 207846
rect 372521 207843 372587 207846
rect 197353 207498 197419 207501
rect 197353 207496 200100 207498
rect 197353 207440 197358 207496
rect 197414 207440 200100 207496
rect 197353 207438 200100 207440
rect 197353 207435 197419 207438
rect 371550 207362 371556 207364
rect 369932 207302 371556 207362
rect 371550 207300 371556 207302
rect 371620 207362 371626 207364
rect 371918 207362 371924 207364
rect 371620 207302 371924 207362
rect 371620 207300 371626 207302
rect 371918 207300 371924 207302
rect 371988 207300 371994 207364
rect 444373 206954 444439 206957
rect 444833 206954 444899 206957
rect 441876 206952 444899 206954
rect 441876 206896 444378 206952
rect 444434 206896 444838 206952
rect 444894 206896 444899 206952
rect 441876 206894 444899 206896
rect 444373 206891 444439 206894
rect 444833 206891 444899 206894
rect 371182 206818 371188 206820
rect 369932 206758 371188 206818
rect 371182 206756 371188 206758
rect 371252 206818 371258 206820
rect 372286 206818 372292 206820
rect 371252 206758 372292 206818
rect 371252 206756 371258 206758
rect 372286 206756 372292 206758
rect 372356 206756 372362 206820
rect 302325 206274 302391 206277
rect 371601 206274 371667 206277
rect 299828 206272 302391 206274
rect 299828 206216 302330 206272
rect 302386 206216 302391 206272
rect 299828 206214 302391 206216
rect 369932 206272 371667 206274
rect 369932 206216 371606 206272
rect 371662 206216 371667 206272
rect 369932 206214 371667 206216
rect 302325 206211 302391 206214
rect 371601 206211 371667 206214
rect 371693 205866 371759 205869
rect 444649 205866 444715 205869
rect 445109 205866 445175 205869
rect 369932 205864 371759 205866
rect 369932 205808 371698 205864
rect 371754 205808 371759 205864
rect 369932 205806 371759 205808
rect 441876 205864 445175 205866
rect 441876 205808 444654 205864
rect 444710 205808 445114 205864
rect 445170 205808 445175 205864
rect 441876 205806 445175 205808
rect 371693 205803 371759 205806
rect 444649 205803 444715 205806
rect 445109 205803 445175 205806
rect 579797 205730 579863 205733
rect 583520 205730 584960 205820
rect 579797 205728 584960 205730
rect 579797 205672 579802 205728
rect 579858 205672 584960 205728
rect 579797 205670 584960 205672
rect 579797 205667 579863 205670
rect 583520 205580 584960 205670
rect 197537 205322 197603 205325
rect 370078 205322 370084 205324
rect 197537 205320 200100 205322
rect 197537 205264 197542 205320
rect 197598 205264 200100 205320
rect 197537 205262 200100 205264
rect 369932 205262 370084 205322
rect 197537 205259 197603 205262
rect 370078 205260 370084 205262
rect 370148 205322 370154 205324
rect 371417 205322 371483 205325
rect 370148 205320 371483 205322
rect 370148 205264 371422 205320
rect 371478 205264 371483 205320
rect 370148 205262 371483 205264
rect 370148 205260 370154 205262
rect 371417 205259 371483 205262
rect 369301 205186 369367 205189
rect 369301 205184 369410 205186
rect 369301 205128 369306 205184
rect 369362 205128 369410 205184
rect 369301 205123 369410 205128
rect 369350 204778 369410 205123
rect 374637 204778 374703 204781
rect 369350 204776 374703 204778
rect 369350 204748 374642 204776
rect 369380 204720 374642 204748
rect 374698 204720 374703 204776
rect 369380 204718 374703 204720
rect 374637 204715 374703 204718
rect 444557 204642 444623 204645
rect 441876 204640 444623 204642
rect 441876 204584 444562 204640
rect 444618 204584 444623 204640
rect 441876 204582 444623 204584
rect 444557 204579 444623 204582
rect 372061 204234 372127 204237
rect 369932 204232 372127 204234
rect 369932 204176 372066 204232
rect 372122 204176 372127 204232
rect 369932 204174 372127 204176
rect 372061 204171 372127 204174
rect 371417 204098 371483 204101
rect 374729 204098 374795 204101
rect 371417 204096 374795 204098
rect 371417 204040 371422 204096
rect 371478 204040 374734 204096
rect 374790 204040 374795 204096
rect 371417 204038 374795 204040
rect 371417 204035 371483 204038
rect 374729 204035 374795 204038
rect 370262 203690 370268 203692
rect 369932 203630 370268 203690
rect 370262 203628 370268 203630
rect 370332 203690 370338 203692
rect 372061 203690 372127 203693
rect 370332 203688 372127 203690
rect 370332 203632 372066 203688
rect 372122 203632 372127 203688
rect 370332 203630 372127 203632
rect 370332 203628 370338 203630
rect 372061 203627 372127 203630
rect 444465 203554 444531 203557
rect 441876 203552 444531 203554
rect 441876 203496 444470 203552
rect 444526 203496 444531 203552
rect 441876 203494 444531 203496
rect 444465 203491 444531 203494
rect 197353 203146 197419 203149
rect 302785 203146 302851 203149
rect 370681 203146 370747 203149
rect 197353 203144 200100 203146
rect 197353 203088 197358 203144
rect 197414 203088 200100 203144
rect 197353 203086 200100 203088
rect 299828 203144 302851 203146
rect 299828 203088 302790 203144
rect 302846 203088 302851 203144
rect 369932 203144 370747 203146
rect 369932 203116 370686 203144
rect 299828 203086 302851 203088
rect 197353 203083 197419 203086
rect 302785 203083 302851 203086
rect 369902 203088 370686 203116
rect 370742 203088 370747 203144
rect 369902 203086 370747 203088
rect 369902 203013 369962 203086
rect 370681 203083 370747 203086
rect 369902 203008 370011 203013
rect 369902 202952 369950 203008
rect 370006 202952 370011 203008
rect 369902 202950 370011 202952
rect 369945 202947 370011 202950
rect 372521 202602 372587 202605
rect 369932 202600 372587 202602
rect 369932 202544 372526 202600
rect 372582 202544 372587 202600
rect 369932 202542 372587 202544
rect 372521 202539 372587 202542
rect 445661 202330 445727 202333
rect 441876 202328 445727 202330
rect 441876 202272 445666 202328
rect 445722 202272 445727 202328
rect 441876 202270 445727 202272
rect 445661 202267 445727 202270
rect 370773 202058 370839 202061
rect 369932 202056 370839 202058
rect 369932 202028 370778 202056
rect -960 201922 480 202012
rect 369902 202000 370778 202028
rect 370834 202000 370839 202056
rect 369902 201998 370839 202000
rect 3049 201922 3115 201925
rect -960 201920 3115 201922
rect -960 201864 3054 201920
rect 3110 201864 3115 201920
rect -960 201862 3115 201864
rect 369902 201922 369962 201998
rect 370773 201995 370839 201998
rect 370037 201922 370103 201925
rect 369902 201920 370103 201922
rect 369902 201864 370042 201920
rect 370098 201864 370103 201920
rect 369902 201862 370103 201864
rect -960 201772 480 201862
rect 3049 201859 3115 201862
rect 370037 201859 370103 201862
rect 371601 201514 371667 201517
rect 369932 201512 371667 201514
rect 369932 201456 371606 201512
rect 371662 201456 371667 201512
rect 369932 201454 371667 201456
rect 371601 201451 371667 201454
rect 372061 201514 372127 201517
rect 374545 201514 374611 201517
rect 372061 201512 374611 201514
rect 372061 201456 372066 201512
rect 372122 201456 374550 201512
rect 374606 201456 374611 201512
rect 372061 201454 374611 201456
rect 372061 201451 372127 201454
rect 374545 201451 374611 201454
rect 371417 201378 371483 201381
rect 371785 201378 371851 201381
rect 369902 201376 371851 201378
rect 369902 201320 371422 201376
rect 371478 201320 371790 201376
rect 371846 201320 371851 201376
rect 369902 201318 371851 201320
rect 197353 200970 197419 200973
rect 197353 200968 200100 200970
rect 197353 200912 197358 200968
rect 197414 200912 200100 200968
rect 369902 200940 369962 201318
rect 371417 201315 371483 201318
rect 371785 201315 371851 201318
rect 445661 201242 445727 201245
rect 441876 201240 445727 201242
rect 441876 201184 445666 201240
rect 445722 201184 445727 201240
rect 441876 201182 445727 201184
rect 445661 201179 445727 201182
rect 197353 200910 200100 200912
rect 197353 200907 197419 200910
rect 372153 200426 372219 200429
rect 369932 200424 372219 200426
rect 369932 200368 372158 200424
rect 372214 200368 372219 200424
rect 369932 200366 372219 200368
rect 372153 200363 372219 200366
rect 445661 200018 445727 200021
rect 441876 200016 445727 200018
rect 441876 199960 445666 200016
rect 445722 199960 445727 200016
rect 441876 199958 445727 199960
rect 445661 199955 445727 199958
rect 302509 199882 302575 199885
rect 371325 199882 371391 199885
rect 299828 199880 302575 199882
rect 299828 199824 302514 199880
rect 302570 199824 302575 199880
rect 299828 199822 302575 199824
rect 369932 199880 371391 199882
rect 369932 199824 371330 199880
rect 371386 199824 371391 199880
rect 369932 199822 371391 199824
rect 302509 199819 302575 199822
rect 371325 199819 371391 199822
rect 371877 199338 371943 199341
rect 369932 199336 371943 199338
rect 369932 199280 371882 199336
rect 371938 199280 371943 199336
rect 369932 199278 371943 199280
rect 371877 199275 371943 199278
rect 371325 198930 371391 198933
rect 372153 198930 372219 198933
rect 445661 198930 445727 198933
rect 371325 198928 372219 198930
rect 371325 198872 371330 198928
rect 371386 198872 372158 198928
rect 372214 198872 372219 198928
rect 371325 198870 372219 198872
rect 441876 198928 445727 198930
rect 441876 198872 445666 198928
rect 445722 198872 445727 198928
rect 441876 198870 445727 198872
rect 371325 198867 371391 198870
rect 372153 198867 372219 198870
rect 445661 198867 445727 198870
rect 197353 198794 197419 198797
rect 371785 198794 371851 198797
rect 371969 198794 372035 198797
rect 197353 198792 200100 198794
rect 197353 198736 197358 198792
rect 197414 198736 200100 198792
rect 197353 198734 200100 198736
rect 369932 198792 372035 198794
rect 369932 198736 371790 198792
rect 371846 198736 371974 198792
rect 372030 198736 372035 198792
rect 369932 198734 372035 198736
rect 197353 198731 197419 198734
rect 371785 198731 371851 198734
rect 371969 198731 372035 198734
rect 371601 198250 371667 198253
rect 369932 198248 371667 198250
rect 369932 198192 371606 198248
rect 371662 198192 371667 198248
rect 369932 198190 371667 198192
rect 371601 198187 371667 198190
rect 372429 197706 372495 197709
rect 445661 197706 445727 197709
rect 369932 197704 372495 197706
rect 369932 197648 372434 197704
rect 372490 197648 372495 197704
rect 369932 197646 372495 197648
rect 441876 197704 445727 197706
rect 441876 197648 445666 197704
rect 445722 197648 445727 197704
rect 441876 197646 445727 197648
rect 372429 197643 372495 197646
rect 445661 197643 445727 197646
rect 371325 197162 371391 197165
rect 369932 197160 371391 197162
rect 369932 197104 371330 197160
rect 371386 197104 371391 197160
rect 369932 197102 371391 197104
rect 371325 197099 371391 197102
rect 302693 196754 302759 196757
rect 299828 196752 302759 196754
rect 299828 196696 302698 196752
rect 302754 196696 302759 196752
rect 299828 196694 302759 196696
rect 302693 196691 302759 196694
rect 197353 196618 197419 196621
rect 372521 196618 372587 196621
rect 445845 196618 445911 196621
rect 197353 196616 200100 196618
rect 197353 196560 197358 196616
rect 197414 196560 200100 196616
rect 197353 196558 200100 196560
rect 369932 196616 372587 196618
rect 369932 196560 372526 196616
rect 372582 196560 372587 196616
rect 369932 196558 372587 196560
rect 441876 196616 445911 196618
rect 441876 196560 445850 196616
rect 445906 196560 445911 196616
rect 441876 196558 445911 196560
rect 197353 196555 197419 196558
rect 372521 196555 372587 196558
rect 445845 196555 445911 196558
rect 370589 196210 370655 196213
rect 370773 196210 370839 196213
rect 369932 196208 370839 196210
rect 369932 196152 370594 196208
rect 370650 196152 370778 196208
rect 370834 196152 370839 196208
rect 369932 196150 370839 196152
rect 370589 196147 370655 196150
rect 370773 196147 370839 196150
rect 364374 196012 364380 196076
rect 364444 196074 364450 196076
rect 364517 196074 364583 196077
rect 364444 196072 364583 196074
rect 364444 196016 364522 196072
rect 364578 196016 364583 196072
rect 364444 196014 364583 196016
rect 364444 196012 364450 196014
rect 364517 196011 364583 196014
rect 371141 196074 371207 196077
rect 371366 196074 371372 196076
rect 371141 196072 371372 196074
rect 371141 196016 371146 196072
rect 371202 196016 371372 196072
rect 371141 196014 371372 196016
rect 371141 196011 371207 196014
rect 371366 196012 371372 196014
rect 371436 196012 371442 196076
rect 370497 195258 370563 195261
rect 372470 195258 372476 195260
rect 370497 195256 372476 195258
rect 370497 195200 370502 195256
rect 370558 195200 372476 195256
rect 370497 195198 372476 195200
rect 370497 195195 370563 195198
rect 372470 195196 372476 195198
rect 372540 195196 372546 195260
rect 361614 194516 361620 194580
rect 361684 194578 361690 194580
rect 362718 194578 362724 194580
rect 361684 194518 362724 194578
rect 361684 194516 361690 194518
rect 362718 194516 362724 194518
rect 362788 194578 362794 194580
rect 362861 194578 362927 194581
rect 362788 194576 362927 194578
rect 362788 194520 362866 194576
rect 362922 194520 362927 194576
rect 362788 194518 362927 194520
rect 362788 194516 362794 194518
rect 362861 194515 362927 194518
rect 364885 194578 364951 194581
rect 365294 194578 365300 194580
rect 364885 194576 365300 194578
rect 364885 194520 364890 194576
rect 364946 194520 365300 194576
rect 364885 194518 365300 194520
rect 364885 194515 364951 194518
rect 365294 194516 365300 194518
rect 365364 194516 365370 194580
rect 198641 194442 198707 194445
rect 198641 194440 200100 194442
rect 198641 194384 198646 194440
rect 198702 194384 200100 194440
rect 198641 194382 200100 194384
rect 198641 194379 198707 194382
rect 302417 193626 302483 193629
rect 299828 193624 302483 193626
rect 299828 193568 302422 193624
rect 302478 193568 302483 193624
rect 299828 193566 302483 193568
rect 302417 193563 302483 193566
rect 580165 192538 580231 192541
rect 583520 192538 584960 192628
rect 580165 192536 584960 192538
rect 580165 192480 580170 192536
rect 580226 192480 584960 192536
rect 580165 192478 584960 192480
rect 580165 192475 580231 192478
rect 583520 192388 584960 192478
rect 197353 192266 197419 192269
rect 197353 192264 200100 192266
rect 197353 192208 197358 192264
rect 197414 192208 200100 192264
rect 197353 192206 200100 192208
rect 197353 192203 197419 192206
rect 303061 190362 303127 190365
rect 299828 190360 303127 190362
rect 299828 190304 303066 190360
rect 303122 190304 303127 190360
rect 299828 190302 303127 190304
rect 303061 190299 303127 190302
rect 197537 190090 197603 190093
rect 197537 190088 200100 190090
rect 197537 190032 197542 190088
rect 197598 190032 200100 190088
rect 197537 190030 200100 190032
rect 197537 190027 197603 190030
rect 172421 189954 172487 189957
rect 169894 189952 172487 189954
rect 169894 189896 172426 189952
rect 172482 189896 172487 189952
rect 169894 189894 172487 189896
rect 169894 189448 169954 189894
rect 172421 189891 172487 189894
rect -960 188866 480 188956
rect 3417 188866 3483 188869
rect -960 188864 3483 188866
rect -960 188808 3422 188864
rect 3478 188808 3483 188864
rect -960 188806 3483 188808
rect -960 188716 480 188806
rect 3417 188803 3483 188806
rect 172421 188730 172487 188733
rect 169894 188728 172487 188730
rect 169894 188672 172426 188728
rect 172482 188672 172487 188728
rect 169894 188670 172487 188672
rect 169894 188360 169954 188670
rect 172421 188667 172487 188670
rect 197353 187914 197419 187917
rect 197353 187912 200100 187914
rect 197353 187856 197358 187912
rect 197414 187856 200100 187912
rect 197353 187854 200100 187856
rect 197353 187851 197419 187854
rect 172421 187370 172487 187373
rect 169894 187368 172487 187370
rect 169894 187312 172426 187368
rect 172482 187312 172487 187368
rect 169894 187310 172487 187312
rect 169894 187136 169954 187310
rect 172421 187307 172487 187310
rect 302693 187234 302759 187237
rect 299828 187232 302759 187234
rect 299828 187176 302698 187232
rect 302754 187176 302759 187232
rect 299828 187174 302759 187176
rect 302693 187171 302759 187174
rect 172421 186146 172487 186149
rect 169894 186144 172487 186146
rect 169894 186088 172426 186144
rect 172482 186088 172487 186144
rect 169894 186086 172487 186088
rect 169894 186048 169954 186086
rect 172421 186083 172487 186086
rect 197353 185738 197419 185741
rect 197353 185736 200100 185738
rect 197353 185680 197358 185736
rect 197414 185680 200100 185736
rect 197353 185678 200100 185680
rect 197353 185675 197419 185678
rect 371233 185602 371299 185605
rect 447501 185602 447567 185605
rect 371233 185600 447567 185602
rect 371233 185544 371238 185600
rect 371294 185544 447506 185600
rect 447562 185544 447567 185600
rect 371233 185542 447567 185544
rect 371233 185539 371299 185542
rect 447501 185539 447567 185542
rect 169894 184786 169954 184824
rect 172421 184786 172487 184789
rect 169894 184784 172487 184786
rect 169894 184728 172426 184784
rect 172482 184728 172487 184784
rect 169894 184726 172487 184728
rect 172421 184723 172487 184726
rect 172329 184378 172395 184381
rect 169894 184376 172395 184378
rect 169894 184320 172334 184376
rect 172390 184320 172395 184376
rect 169894 184318 172395 184320
rect 169894 183736 169954 184318
rect 172329 184315 172395 184318
rect 302785 184106 302851 184109
rect 299828 184104 302851 184106
rect 299828 184048 302790 184104
rect 302846 184048 302851 184104
rect 299828 184046 302851 184048
rect 302785 184043 302851 184046
rect 198181 183562 198247 183565
rect 198181 183560 200100 183562
rect 198181 183504 198186 183560
rect 198242 183504 200100 183560
rect 198181 183502 200100 183504
rect 198181 183499 198247 183502
rect 172421 183018 172487 183021
rect 169894 183016 172487 183018
rect 169894 182960 172426 183016
rect 172482 182960 172487 183016
rect 169894 182958 172487 182960
rect 169894 182512 169954 182958
rect 172421 182955 172487 182958
rect 172421 181794 172487 181797
rect 169894 181792 172487 181794
rect 169894 181736 172426 181792
rect 172482 181736 172487 181792
rect 169894 181734 172487 181736
rect 169894 181424 169954 181734
rect 172421 181731 172487 181734
rect 197353 181386 197419 181389
rect 197353 181384 200100 181386
rect 197353 181328 197358 181384
rect 197414 181328 200100 181384
rect 197353 181326 200100 181328
rect 197353 181323 197419 181326
rect 302969 180842 303035 180845
rect 299828 180840 303035 180842
rect 299828 180784 302974 180840
rect 303030 180784 303035 180840
rect 299828 180782 303035 180784
rect 302969 180779 303035 180782
rect 172421 180570 172487 180573
rect 169894 180568 172487 180570
rect 169894 180512 172426 180568
rect 172482 180512 172487 180568
rect 169894 180510 172487 180512
rect 169894 180200 169954 180510
rect 172421 180507 172487 180510
rect 172421 179210 172487 179213
rect 169894 179208 172487 179210
rect 169894 179152 172426 179208
rect 172482 179152 172487 179208
rect 169894 179150 172487 179152
rect 169894 179112 169954 179150
rect 172421 179147 172487 179150
rect 197537 179210 197603 179213
rect 580165 179210 580231 179213
rect 583520 179210 584960 179300
rect 197537 179208 200100 179210
rect 197537 179152 197542 179208
rect 197598 179152 200100 179208
rect 197537 179150 200100 179152
rect 580165 179208 584960 179210
rect 580165 179152 580170 179208
rect 580226 179152 584960 179208
rect 580165 179150 584960 179152
rect 197537 179147 197603 179150
rect 580165 179147 580231 179150
rect 583520 179060 584960 179150
rect 172329 177986 172395 177989
rect 169894 177984 172395 177986
rect 169894 177928 172334 177984
rect 172390 177928 172395 177984
rect 169894 177926 172395 177928
rect 169894 177888 169954 177926
rect 172329 177923 172395 177926
rect 302877 177714 302943 177717
rect 299828 177712 302943 177714
rect 299828 177656 302882 177712
rect 302938 177656 302943 177712
rect 299828 177654 302943 177656
rect 302877 177651 302943 177654
rect 172421 177442 172487 177445
rect 169894 177440 172487 177442
rect 169894 177384 172426 177440
rect 172482 177384 172487 177440
rect 169894 177382 172487 177384
rect 169894 176800 169954 177382
rect 172421 177379 172487 177382
rect 197353 177034 197419 177037
rect 197353 177032 200100 177034
rect 197353 176976 197358 177032
rect 197414 176976 200100 177032
rect 197353 176974 200100 176976
rect 197353 176971 197419 176974
rect 172421 176082 172487 176085
rect 169894 176080 172487 176082
rect -960 175796 480 176036
rect 169894 176024 172426 176080
rect 172482 176024 172487 176080
rect 169894 176022 172487 176024
rect 169894 175576 169954 176022
rect 172421 176019 172487 176022
rect 370865 175674 370931 175677
rect 371734 175674 371740 175676
rect 370865 175672 371740 175674
rect 370865 175616 370870 175672
rect 370926 175616 371740 175672
rect 370865 175614 371740 175616
rect 370865 175611 370931 175614
rect 371734 175612 371740 175614
rect 371804 175612 371810 175676
rect 372286 175266 372292 175268
rect 371926 175206 372292 175266
rect 371926 174996 371986 175206
rect 372286 175204 372292 175206
rect 372356 175204 372362 175268
rect 371918 174932 371924 174996
rect 371988 174932 371994 174996
rect 171685 174858 171751 174861
rect 169894 174856 171751 174858
rect 169894 174800 171690 174856
rect 171746 174800 171751 174856
rect 169894 174798 171751 174800
rect 169894 174488 169954 174798
rect 171685 174795 171751 174798
rect 197629 174858 197695 174861
rect 197629 174856 200100 174858
rect 197629 174800 197634 174856
rect 197690 174800 200100 174856
rect 197629 174798 200100 174800
rect 197629 174795 197695 174798
rect 302233 174586 302299 174589
rect 299828 174584 302299 174586
rect 299828 174528 302238 174584
rect 302294 174528 302299 174584
rect 299828 174526 302299 174528
rect 302233 174523 302299 174526
rect 171501 173634 171567 173637
rect 169894 173632 171567 173634
rect 169894 173576 171506 173632
rect 171562 173576 171567 173632
rect 169894 173574 171567 173576
rect 169894 173264 169954 173574
rect 171501 173571 171567 173574
rect 372286 173164 372292 173228
rect 372356 173226 372362 173228
rect 448881 173226 448947 173229
rect 372356 173224 448947 173226
rect 372356 173168 448886 173224
rect 448942 173168 448947 173224
rect 372356 173166 448947 173168
rect 372356 173164 372362 173166
rect 448881 173163 448947 173166
rect 197353 172682 197419 172685
rect 197353 172680 200100 172682
rect 197353 172624 197358 172680
rect 197414 172624 200100 172680
rect 197353 172622 200100 172624
rect 197353 172619 197419 172622
rect 172421 172410 172487 172413
rect 169894 172408 172487 172410
rect 169894 172352 172426 172408
rect 172482 172352 172487 172408
rect 169894 172350 172487 172352
rect 169894 172176 169954 172350
rect 172421 172347 172487 172350
rect 371918 171668 371924 171732
rect 371988 171730 371994 171732
rect 450169 171730 450235 171733
rect 371988 171728 450235 171730
rect 371988 171672 450174 171728
rect 450230 171672 450235 171728
rect 371988 171670 450235 171672
rect 371988 171668 371994 171670
rect 450169 171667 450235 171670
rect 302785 171322 302851 171325
rect 299828 171320 302851 171322
rect 299828 171264 302790 171320
rect 302846 171264 302851 171320
rect 299828 171262 302851 171264
rect 302785 171259 302851 171262
rect 172421 171050 172487 171053
rect 169894 171048 172487 171050
rect 169894 170992 172426 171048
rect 172482 170992 172487 171048
rect 169894 170990 172487 170992
rect 169894 170952 169954 170990
rect 172421 170987 172487 170990
rect 171777 170506 171843 170509
rect 169894 170504 171843 170506
rect 169894 170448 171782 170504
rect 171838 170448 171843 170504
rect 169894 170446 171843 170448
rect 169894 169864 169954 170446
rect 171777 170443 171843 170446
rect 197353 170506 197419 170509
rect 197353 170504 200100 170506
rect 197353 170448 197358 170504
rect 197414 170448 200100 170504
rect 197353 170446 200100 170448
rect 197353 170443 197419 170446
rect 172421 169146 172487 169149
rect 169894 169144 172487 169146
rect 169894 169088 172426 169144
rect 172482 169088 172487 169144
rect 169894 169086 172487 169088
rect 169894 168640 169954 169086
rect 172421 169083 172487 169086
rect 197905 168330 197971 168333
rect 197905 168328 200100 168330
rect 197905 168272 197910 168328
rect 197966 168272 200100 168328
rect 197905 168270 200100 168272
rect 197905 168267 197971 168270
rect 171869 168194 171935 168197
rect 302693 168194 302759 168197
rect 169894 168192 171935 168194
rect 169894 168136 171874 168192
rect 171930 168136 171935 168192
rect 169894 168134 171935 168136
rect 299828 168192 302759 168194
rect 299828 168136 302698 168192
rect 302754 168136 302759 168192
rect 299828 168134 302759 168136
rect 169894 167552 169954 168134
rect 171869 168131 171935 168134
rect 302693 168131 302759 168134
rect 172421 166698 172487 166701
rect 169894 166696 172487 166698
rect 169894 166640 172426 166696
rect 172482 166640 172487 166696
rect 169894 166638 172487 166640
rect 169894 166328 169954 166638
rect 172421 166635 172487 166638
rect 198457 166154 198523 166157
rect 198457 166152 200100 166154
rect 198457 166096 198462 166152
rect 198518 166096 200100 166152
rect 198457 166094 200100 166096
rect 198457 166091 198523 166094
rect 580165 165882 580231 165885
rect 583520 165882 584960 165972
rect 580165 165880 584960 165882
rect 580165 165824 580170 165880
rect 580226 165824 584960 165880
rect 580165 165822 584960 165824
rect 580165 165819 580231 165822
rect 583520 165732 584960 165822
rect 169894 164522 169954 165240
rect 302601 164930 302667 164933
rect 299828 164928 302667 164930
rect 299828 164872 302606 164928
rect 302662 164872 302667 164928
rect 299828 164870 302667 164872
rect 302601 164867 302667 164870
rect 171961 164522 172027 164525
rect 169894 164520 172027 164522
rect 169894 164464 171966 164520
rect 172022 164464 172027 164520
rect 169894 164462 172027 164464
rect 171961 164459 172027 164462
rect 172421 164114 172487 164117
rect 169894 164112 172487 164114
rect 169894 164056 172426 164112
rect 172482 164056 172487 164112
rect 169894 164054 172487 164056
rect 169894 164016 169954 164054
rect 172421 164051 172487 164054
rect 197997 163978 198063 163981
rect 197997 163976 200100 163978
rect 197997 163920 198002 163976
rect 198058 163920 200100 163976
rect 197997 163918 200100 163920
rect 197997 163915 198063 163918
rect 172053 163570 172119 163573
rect 169894 163568 172119 163570
rect 169894 163512 172058 163568
rect 172114 163512 172119 163568
rect 169894 163510 172119 163512
rect -960 162890 480 162980
rect 169894 162928 169954 163510
rect 172053 163507 172119 163510
rect 3233 162890 3299 162893
rect -960 162888 3299 162890
rect -960 162832 3238 162888
rect 3294 162832 3299 162888
rect -960 162830 3299 162832
rect -960 162740 480 162830
rect 3233 162827 3299 162830
rect 371141 162754 371207 162757
rect 372286 162754 372292 162756
rect 371141 162752 372292 162754
rect 371141 162696 371146 162752
rect 371202 162696 372292 162752
rect 371141 162694 372292 162696
rect 371141 162691 371207 162694
rect 372286 162692 372292 162694
rect 372356 162692 372362 162756
rect 171777 162346 171843 162349
rect 169894 162344 171843 162346
rect 169894 162288 171782 162344
rect 171838 162288 171843 162344
rect 169894 162286 171843 162288
rect 169894 161704 169954 162286
rect 171777 162283 171843 162286
rect 197353 161802 197419 161805
rect 302969 161802 303035 161805
rect 197353 161800 200100 161802
rect 197353 161744 197358 161800
rect 197414 161744 200100 161800
rect 197353 161742 200100 161744
rect 299828 161800 303035 161802
rect 299828 161744 302974 161800
rect 303030 161744 303035 161800
rect 299828 161742 303035 161744
rect 197353 161739 197419 161742
rect 302969 161739 303035 161742
rect 172237 160986 172303 160989
rect 169894 160984 172303 160986
rect 169894 160928 172242 160984
rect 172298 160928 172303 160984
rect 169894 160926 172303 160928
rect 169894 160616 169954 160926
rect 172237 160923 172303 160926
rect 197353 159626 197419 159629
rect 197353 159624 200100 159626
rect 197353 159568 197358 159624
rect 197414 159568 200100 159624
rect 197353 159566 200100 159568
rect 197353 159563 197419 159566
rect 302785 158674 302851 158677
rect 299828 158672 302851 158674
rect 299828 158616 302790 158672
rect 302846 158616 302851 158672
rect 299828 158614 302851 158616
rect 302785 158611 302851 158614
rect 197353 157450 197419 157453
rect 197353 157448 200100 157450
rect 197353 157392 197358 157448
rect 197414 157392 200100 157448
rect 197353 157390 200100 157392
rect 197353 157387 197419 157390
rect 302877 155410 302943 155413
rect 299828 155408 302943 155410
rect 299828 155352 302882 155408
rect 302938 155352 302943 155408
rect 299828 155350 302943 155352
rect 302877 155347 302943 155350
rect 198273 155274 198339 155277
rect 198273 155272 200100 155274
rect 198273 155216 198278 155272
rect 198334 155216 200100 155272
rect 198273 155214 200100 155216
rect 198273 155211 198339 155214
rect 171593 153778 171659 153781
rect 371693 153778 371759 153781
rect 169924 153776 171659 153778
rect 169924 153720 171598 153776
rect 171654 153720 171659 153776
rect 169924 153718 171659 153720
rect 369932 153776 371759 153778
rect 369932 153720 371698 153776
rect 371754 153720 371759 153776
rect 369932 153718 371759 153720
rect 171593 153715 171659 153718
rect 371693 153715 371759 153718
rect 445661 153506 445727 153509
rect 441876 153504 445727 153506
rect 441876 153448 445666 153504
rect 445722 153448 445727 153504
rect 441876 153446 445727 153448
rect 445661 153443 445727 153446
rect 171225 153234 171291 153237
rect 371693 153234 371759 153237
rect 169924 153232 171291 153234
rect 169924 153176 171230 153232
rect 171286 153176 171291 153232
rect 169924 153174 171291 153176
rect 369932 153232 371759 153234
rect 369932 153176 371698 153232
rect 371754 153176 371759 153232
rect 369932 153174 371759 153176
rect 171225 153171 171291 153174
rect 371693 153171 371759 153174
rect 198089 153098 198155 153101
rect 198089 153096 200100 153098
rect 198089 153040 198094 153096
rect 198150 153040 200100 153096
rect 198089 153038 200100 153040
rect 198089 153035 198155 153038
rect 369301 152962 369367 152965
rect 371918 152962 371924 152964
rect 369301 152960 371924 152962
rect 369301 152904 369306 152960
rect 369362 152904 371924 152960
rect 369301 152902 371924 152904
rect 369301 152899 369367 152902
rect 371918 152900 371924 152902
rect 371988 152900 371994 152964
rect 172421 152690 172487 152693
rect 371509 152690 371575 152693
rect 169924 152688 172487 152690
rect 169924 152632 172426 152688
rect 172482 152632 172487 152688
rect 169924 152630 172487 152632
rect 369932 152688 371575 152690
rect 369932 152632 371514 152688
rect 371570 152632 371575 152688
rect 369932 152630 371575 152632
rect 172421 152627 172487 152630
rect 371509 152627 371575 152630
rect 580165 152690 580231 152693
rect 583520 152690 584960 152780
rect 580165 152688 584960 152690
rect 580165 152632 580170 152688
rect 580226 152632 584960 152688
rect 580165 152630 584960 152632
rect 580165 152627 580231 152630
rect 583520 152540 584960 152630
rect 444833 152418 444899 152421
rect 441876 152416 444899 152418
rect 441876 152360 444838 152416
rect 444894 152360 444899 152416
rect 441876 152358 444899 152360
rect 444833 152355 444899 152358
rect 302785 152282 302851 152285
rect 299828 152280 302851 152282
rect 299828 152224 302790 152280
rect 302846 152224 302851 152280
rect 299828 152222 302851 152224
rect 302785 152219 302851 152222
rect 172329 152146 172395 152149
rect 371693 152146 371759 152149
rect 169924 152144 172395 152146
rect 169924 152088 172334 152144
rect 172390 152088 172395 152144
rect 169924 152086 172395 152088
rect 369932 152144 371759 152146
rect 369932 152088 371698 152144
rect 371754 152088 371759 152144
rect 369932 152086 371759 152088
rect 172329 152083 172395 152086
rect 371693 152083 371759 152086
rect 172421 151602 172487 151605
rect 371693 151602 371759 151605
rect 169924 151600 172487 151602
rect 169924 151544 172426 151600
rect 172482 151544 172487 151600
rect 169924 151542 172487 151544
rect 369932 151600 371759 151602
rect 369932 151544 371698 151600
rect 371754 151544 371759 151600
rect 369932 151542 371759 151544
rect 172421 151539 172487 151542
rect 371693 151539 371759 151542
rect 444833 151194 444899 151197
rect 441876 151192 444899 151194
rect 441876 151136 444838 151192
rect 444894 151136 444899 151192
rect 441876 151134 444899 151136
rect 444833 151131 444899 151134
rect 172329 151058 172395 151061
rect 371693 151058 371759 151061
rect 169924 151056 172395 151058
rect 169924 151000 172334 151056
rect 172390 151000 172395 151056
rect 169924 150998 172395 151000
rect 369932 151056 371759 151058
rect 369932 151000 371698 151056
rect 371754 151000 371759 151056
rect 369932 150998 371759 151000
rect 172329 150995 172395 150998
rect 371693 150995 371759 150998
rect 198365 150922 198431 150925
rect 198365 150920 200100 150922
rect 198365 150864 198370 150920
rect 198426 150864 200100 150920
rect 198365 150862 200100 150864
rect 198365 150859 198431 150862
rect 171869 150514 171935 150517
rect 371509 150514 371575 150517
rect 169924 150512 171935 150514
rect 169924 150456 171874 150512
rect 171930 150456 171935 150512
rect 169924 150454 171935 150456
rect 369932 150512 371575 150514
rect 369932 150456 371514 150512
rect 371570 150456 371575 150512
rect 369932 150454 371575 150456
rect 171869 150451 171935 150454
rect 371509 150451 371575 150454
rect 444925 150106 444991 150109
rect 441876 150104 444991 150106
rect 441876 150048 444930 150104
rect 444986 150048 444991 150104
rect 441876 150046 444991 150048
rect 444925 150043 444991 150046
rect 171501 149970 171567 149973
rect 371693 149970 371759 149973
rect 169924 149968 171567 149970
rect -960 149834 480 149924
rect 169924 149912 171506 149968
rect 171562 149912 171567 149968
rect 169924 149910 171567 149912
rect 369932 149968 371759 149970
rect 369932 149912 371698 149968
rect 371754 149912 371759 149968
rect 369932 149910 371759 149912
rect 171501 149907 171567 149910
rect 371693 149907 371759 149910
rect 3417 149834 3483 149837
rect -960 149832 3483 149834
rect -960 149776 3422 149832
rect 3478 149776 3483 149832
rect -960 149774 3483 149776
rect -960 149684 480 149774
rect 3417 149771 3483 149774
rect 171685 149426 171751 149429
rect 371509 149426 371575 149429
rect 169924 149424 171751 149426
rect 169924 149368 171690 149424
rect 171746 149368 171751 149424
rect 169924 149366 171751 149368
rect 369932 149424 371575 149426
rect 369932 149368 371514 149424
rect 371570 149368 371575 149424
rect 369932 149366 371575 149368
rect 171685 149363 171751 149366
rect 371509 149363 371575 149366
rect 302785 149154 302851 149157
rect 299828 149152 302851 149154
rect 299828 149096 302790 149152
rect 302846 149096 302851 149152
rect 299828 149094 302851 149096
rect 302785 149091 302851 149094
rect 171869 148882 171935 148885
rect 371693 148882 371759 148885
rect 445293 148882 445359 148885
rect 169924 148880 171935 148882
rect 169924 148824 171874 148880
rect 171930 148824 171935 148880
rect 169924 148822 171935 148824
rect 369932 148880 371759 148882
rect 369932 148824 371698 148880
rect 371754 148824 371759 148880
rect 369932 148822 371759 148824
rect 441876 148880 445359 148882
rect 441876 148824 445298 148880
rect 445354 148824 445359 148880
rect 441876 148822 445359 148824
rect 171869 148819 171935 148822
rect 371693 148819 371759 148822
rect 445293 148819 445359 148822
rect 198273 148746 198339 148749
rect 198273 148744 200100 148746
rect 198273 148688 198278 148744
rect 198334 148688 200100 148744
rect 198273 148686 200100 148688
rect 198273 148683 198339 148686
rect 171685 148338 171751 148341
rect 371693 148338 371759 148341
rect 169924 148336 171751 148338
rect 169924 148280 171690 148336
rect 171746 148280 171751 148336
rect 169924 148278 171751 148280
rect 369932 148336 371759 148338
rect 369932 148280 371698 148336
rect 371754 148280 371759 148336
rect 369932 148278 371759 148280
rect 171685 148275 171751 148278
rect 371693 148275 371759 148278
rect 171685 147794 171751 147797
rect 371693 147794 371759 147797
rect 445569 147794 445635 147797
rect 169924 147792 171751 147794
rect 169924 147736 171690 147792
rect 171746 147736 171751 147792
rect 169924 147734 171751 147736
rect 369932 147792 371759 147794
rect 369932 147736 371698 147792
rect 371754 147736 371759 147792
rect 369932 147734 371759 147736
rect 441876 147792 445635 147794
rect 441876 147736 445574 147792
rect 445630 147736 445635 147792
rect 441876 147734 445635 147736
rect 171685 147731 171751 147734
rect 371693 147731 371759 147734
rect 445569 147731 445635 147734
rect 172421 147250 172487 147253
rect 371233 147250 371299 147253
rect 169924 147248 172487 147250
rect 169924 147192 172426 147248
rect 172482 147192 172487 147248
rect 169924 147190 172487 147192
rect 369932 147248 371299 147250
rect 369932 147192 371238 147248
rect 371294 147192 371299 147248
rect 369932 147190 371299 147192
rect 172421 147187 172487 147190
rect 371233 147187 371299 147190
rect 171869 146706 171935 146709
rect 371233 146706 371299 146709
rect 169924 146704 171935 146706
rect 169924 146648 171874 146704
rect 171930 146648 171935 146704
rect 169924 146646 171935 146648
rect 369932 146704 371299 146706
rect 369932 146648 371238 146704
rect 371294 146648 371299 146704
rect 369932 146646 371299 146648
rect 171869 146643 171935 146646
rect 371233 146643 371299 146646
rect 197721 146570 197787 146573
rect 444833 146570 444899 146573
rect 197721 146568 200100 146570
rect 197721 146512 197726 146568
rect 197782 146512 200100 146568
rect 197721 146510 200100 146512
rect 441876 146568 444899 146570
rect 441876 146512 444838 146568
rect 444894 146512 444899 146568
rect 441876 146510 444899 146512
rect 197721 146507 197787 146510
rect 444833 146507 444899 146510
rect 172237 146162 172303 146165
rect 371693 146162 371759 146165
rect 169924 146160 172303 146162
rect 169924 146104 172242 146160
rect 172298 146104 172303 146160
rect 169924 146102 172303 146104
rect 369932 146160 371759 146162
rect 369932 146104 371698 146160
rect 371754 146104 371759 146160
rect 369932 146102 371759 146104
rect 172237 146099 172303 146102
rect 371693 146099 371759 146102
rect 302785 145890 302851 145893
rect 299828 145888 302851 145890
rect 299828 145832 302790 145888
rect 302846 145832 302851 145888
rect 299828 145830 302851 145832
rect 302785 145827 302851 145830
rect 172421 145618 172487 145621
rect 371509 145618 371575 145621
rect 169924 145616 172487 145618
rect 169924 145560 172426 145616
rect 172482 145560 172487 145616
rect 169924 145558 172487 145560
rect 369932 145616 371575 145618
rect 369932 145560 371514 145616
rect 371570 145560 371575 145616
rect 369932 145558 371575 145560
rect 172421 145555 172487 145558
rect 371509 145555 371575 145558
rect 445477 145482 445543 145485
rect 441876 145480 445543 145482
rect 441876 145424 445482 145480
rect 445538 145424 445543 145480
rect 441876 145422 445543 145424
rect 445477 145419 445543 145422
rect 172329 145074 172395 145077
rect 371693 145074 371759 145077
rect 169924 145072 172395 145074
rect 169924 145016 172334 145072
rect 172390 145016 172395 145072
rect 169924 145014 172395 145016
rect 369932 145072 371759 145074
rect 369932 145016 371698 145072
rect 371754 145016 371759 145072
rect 369932 145014 371759 145016
rect 172329 145011 172395 145014
rect 371693 145011 371759 145014
rect 172421 144530 172487 144533
rect 371693 144530 371759 144533
rect 169924 144528 172487 144530
rect 169924 144472 172426 144528
rect 172482 144472 172487 144528
rect 169924 144470 172487 144472
rect 369932 144528 371759 144530
rect 369932 144472 371698 144528
rect 371754 144472 371759 144528
rect 369932 144470 371759 144472
rect 172421 144467 172487 144470
rect 371693 144467 371759 144470
rect 197353 144394 197419 144397
rect 197353 144392 200100 144394
rect 197353 144336 197358 144392
rect 197414 144336 200100 144392
rect 197353 144334 200100 144336
rect 197353 144331 197419 144334
rect 445109 144258 445175 144261
rect 441876 144256 445175 144258
rect 441876 144200 445114 144256
rect 445170 144200 445175 144256
rect 441876 144198 445175 144200
rect 445109 144195 445175 144198
rect 172145 144122 172211 144125
rect 371509 144122 371575 144125
rect 169924 144120 172211 144122
rect 169924 144064 172150 144120
rect 172206 144064 172211 144120
rect 169924 144062 172211 144064
rect 369932 144120 371575 144122
rect 369932 144064 371514 144120
rect 371570 144064 371575 144120
rect 369932 144062 371575 144064
rect 172145 144059 172211 144062
rect 371509 144059 371575 144062
rect 171777 143578 171843 143581
rect 372061 143578 372127 143581
rect 169924 143576 171843 143578
rect 169924 143520 171782 143576
rect 171838 143520 171843 143576
rect 169924 143518 171843 143520
rect 369932 143576 372127 143578
rect 369932 143520 372066 143576
rect 372122 143520 372127 143576
rect 369932 143518 372127 143520
rect 171777 143515 171843 143518
rect 372061 143515 372127 143518
rect 445109 143170 445175 143173
rect 441876 143168 445175 143170
rect 441876 143112 445114 143168
rect 445170 143112 445175 143168
rect 441876 143110 445175 143112
rect 445109 143107 445175 143110
rect 171869 143034 171935 143037
rect 371693 143034 371759 143037
rect 169924 143032 171935 143034
rect 169924 142976 171874 143032
rect 171930 142976 171935 143032
rect 169924 142974 171935 142976
rect 369932 143032 371759 143034
rect 369932 142976 371698 143032
rect 371754 142976 371759 143032
rect 369932 142974 371759 142976
rect 171869 142971 171935 142974
rect 371693 142971 371759 142974
rect 302785 142762 302851 142765
rect 299828 142760 302851 142762
rect 299828 142704 302790 142760
rect 302846 142704 302851 142760
rect 299828 142702 302851 142704
rect 302785 142699 302851 142702
rect 171685 142490 171751 142493
rect 371233 142490 371299 142493
rect 169924 142488 171751 142490
rect 169924 142432 171690 142488
rect 171746 142432 171751 142488
rect 169924 142430 171751 142432
rect 369932 142488 371299 142490
rect 369932 142432 371238 142488
rect 371294 142432 371299 142488
rect 369932 142430 371299 142432
rect 171685 142427 171751 142430
rect 371233 142427 371299 142430
rect 197353 142218 197419 142221
rect 197353 142216 200100 142218
rect 197353 142160 197358 142216
rect 197414 142160 200100 142216
rect 197353 142158 200100 142160
rect 197353 142155 197419 142158
rect 171501 141946 171567 141949
rect 371693 141946 371759 141949
rect 444373 141946 444439 141949
rect 169924 141944 171567 141946
rect 169924 141888 171506 141944
rect 171562 141888 171567 141944
rect 169924 141886 171567 141888
rect 369932 141944 371759 141946
rect 369932 141888 371698 141944
rect 371754 141888 371759 141944
rect 369932 141886 371759 141888
rect 441876 141944 444439 141946
rect 441876 141888 444378 141944
rect 444434 141888 444439 141944
rect 441876 141886 444439 141888
rect 171501 141883 171567 141886
rect 371693 141883 371759 141886
rect 444373 141883 444439 141886
rect 171777 141402 171843 141405
rect 371509 141402 371575 141405
rect 169924 141400 171843 141402
rect 169924 141344 171782 141400
rect 171838 141344 171843 141400
rect 169924 141342 171843 141344
rect 369932 141400 371575 141402
rect 369932 141344 371514 141400
rect 371570 141344 371575 141400
rect 369932 141342 371575 141344
rect 171777 141339 171843 141342
rect 371509 141339 371575 141342
rect 172421 140858 172487 140861
rect 371233 140858 371299 140861
rect 444741 140858 444807 140861
rect 169924 140856 172487 140858
rect 169924 140800 172426 140856
rect 172482 140800 172487 140856
rect 169924 140798 172487 140800
rect 369932 140856 371299 140858
rect 369932 140800 371238 140856
rect 371294 140800 371299 140856
rect 369932 140798 371299 140800
rect 441876 140856 444807 140858
rect 441876 140800 444746 140856
rect 444802 140800 444807 140856
rect 441876 140798 444807 140800
rect 172421 140795 172487 140798
rect 371233 140795 371299 140798
rect 444741 140795 444807 140798
rect 171685 140314 171751 140317
rect 371693 140314 371759 140317
rect 169924 140312 171751 140314
rect 169924 140256 171690 140312
rect 171746 140256 171751 140312
rect 169924 140254 171751 140256
rect 369932 140312 371759 140314
rect 369932 140256 371698 140312
rect 371754 140256 371759 140312
rect 369932 140254 371759 140256
rect 171685 140251 171751 140254
rect 371693 140251 371759 140254
rect 198273 140042 198339 140045
rect 198273 140040 200100 140042
rect 198273 139984 198278 140040
rect 198334 139984 200100 140040
rect 198273 139982 200100 139984
rect 198273 139979 198339 139982
rect 171685 139770 171751 139773
rect 372705 139770 372771 139773
rect 169924 139768 171751 139770
rect 169924 139712 171690 139768
rect 171746 139712 171751 139768
rect 169924 139710 171751 139712
rect 369932 139768 372771 139770
rect 369932 139712 372710 139768
rect 372766 139712 372771 139768
rect 369932 139710 372771 139712
rect 171685 139707 171751 139710
rect 372705 139707 372771 139710
rect 302877 139634 302943 139637
rect 444373 139634 444439 139637
rect 299828 139632 302943 139634
rect 299828 139576 302882 139632
rect 302938 139576 302943 139632
rect 299828 139574 302943 139576
rect 441876 139632 444439 139634
rect 441876 139576 444378 139632
rect 444434 139576 444439 139632
rect 441876 139574 444439 139576
rect 302877 139571 302943 139574
rect 444373 139571 444439 139574
rect 580165 139362 580231 139365
rect 583520 139362 584960 139452
rect 580165 139360 584960 139362
rect 580165 139304 580170 139360
rect 580226 139304 584960 139360
rect 580165 139302 584960 139304
rect 580165 139299 580231 139302
rect 172421 139226 172487 139229
rect 371693 139226 371759 139229
rect 169924 139224 172487 139226
rect 169924 139168 172426 139224
rect 172482 139168 172487 139224
rect 169924 139166 172487 139168
rect 369932 139224 371759 139226
rect 369932 139168 371698 139224
rect 371754 139168 371759 139224
rect 583520 139212 584960 139302
rect 369932 139166 371759 139168
rect 172421 139163 172487 139166
rect 371693 139163 371759 139166
rect 171593 138682 171659 138685
rect 371693 138682 371759 138685
rect 169924 138680 171659 138682
rect 169924 138624 171598 138680
rect 171654 138624 171659 138680
rect 169924 138622 171659 138624
rect 369932 138680 371759 138682
rect 369932 138624 371698 138680
rect 371754 138624 371759 138680
rect 369932 138622 371759 138624
rect 171593 138619 171659 138622
rect 371693 138619 371759 138622
rect 444373 138546 444439 138549
rect 441876 138544 444439 138546
rect 441876 138488 444378 138544
rect 444434 138488 444439 138544
rect 441876 138486 444439 138488
rect 444373 138483 444439 138486
rect 171501 138138 171567 138141
rect 371509 138138 371575 138141
rect 169924 138136 171567 138138
rect 169924 138080 171506 138136
rect 171562 138080 171567 138136
rect 169924 138078 171567 138080
rect 369932 138136 371575 138138
rect 369932 138080 371514 138136
rect 371570 138080 371575 138136
rect 369932 138078 371575 138080
rect 171501 138075 171567 138078
rect 371509 138075 371575 138078
rect 197537 137866 197603 137869
rect 197537 137864 200100 137866
rect 197537 137808 197542 137864
rect 197598 137808 200100 137864
rect 197537 137806 200100 137808
rect 197537 137803 197603 137806
rect 172053 137594 172119 137597
rect 371366 137594 371372 137596
rect 169924 137592 172119 137594
rect 169924 137536 172058 137592
rect 172114 137536 172119 137592
rect 169924 137534 172119 137536
rect 369932 137534 371372 137594
rect 172053 137531 172119 137534
rect 371366 137532 371372 137534
rect 371436 137532 371442 137596
rect 444373 137322 444439 137325
rect 441876 137320 444439 137322
rect 441876 137264 444378 137320
rect 444434 137264 444439 137320
rect 441876 137262 444439 137264
rect 444373 137259 444439 137262
rect 172329 137050 172395 137053
rect 372470 137050 372476 137052
rect 169924 137048 172395 137050
rect 169924 136992 172334 137048
rect 172390 136992 172395 137048
rect 169924 136990 172395 136992
rect 369932 136990 372476 137050
rect 172329 136987 172395 136990
rect 372470 136988 372476 136990
rect 372540 136988 372546 137052
rect -960 136778 480 136868
rect 3233 136778 3299 136781
rect -960 136776 3299 136778
rect -960 136720 3238 136776
rect 3294 136720 3299 136776
rect -960 136718 3299 136720
rect -960 136628 480 136718
rect 3233 136715 3299 136718
rect 172421 136506 172487 136509
rect 371734 136506 371740 136508
rect 169924 136504 172487 136506
rect 169924 136448 172426 136504
rect 172482 136448 172487 136504
rect 169924 136446 172487 136448
rect 369932 136446 371740 136506
rect 172421 136443 172487 136446
rect 371734 136444 371740 136446
rect 371804 136444 371810 136508
rect 302969 136370 303035 136373
rect 299828 136368 303035 136370
rect 299828 136312 302974 136368
rect 303030 136312 303035 136368
rect 299828 136310 303035 136312
rect 302969 136307 303035 136310
rect 444741 136234 444807 136237
rect 445937 136234 446003 136237
rect 441876 136232 446003 136234
rect 441876 136176 444746 136232
rect 444802 136176 445942 136232
rect 445998 136176 446003 136232
rect 441876 136174 446003 136176
rect 444741 136171 444807 136174
rect 445937 136171 446003 136174
rect 172237 135962 172303 135965
rect 370129 135962 370195 135965
rect 169924 135960 172303 135962
rect 169924 135904 172242 135960
rect 172298 135904 172303 135960
rect 169924 135902 172303 135904
rect 369932 135960 370195 135962
rect 369932 135904 370134 135960
rect 370190 135904 370195 135960
rect 369932 135902 370195 135904
rect 172237 135899 172303 135902
rect 370129 135899 370195 135902
rect 198089 135690 198155 135693
rect 198089 135688 200100 135690
rect 198089 135632 198094 135688
rect 198150 135632 200100 135688
rect 198089 135630 200100 135632
rect 198089 135627 198155 135630
rect 171685 135418 171751 135421
rect 370221 135418 370287 135421
rect 169924 135416 171751 135418
rect 169924 135360 171690 135416
rect 171746 135360 171751 135416
rect 169924 135358 171751 135360
rect 369932 135416 370287 135418
rect 369932 135360 370226 135416
rect 370282 135360 370287 135416
rect 369932 135358 370287 135360
rect 171685 135355 171751 135358
rect 370221 135355 370287 135358
rect 369393 135146 369459 135149
rect 369350 135144 369459 135146
rect 369350 135088 369398 135144
rect 369454 135088 369459 135144
rect 369350 135083 369459 135088
rect 172421 134874 172487 134877
rect 169924 134872 172487 134874
rect 169924 134816 172426 134872
rect 172482 134816 172487 134872
rect 369350 134844 369410 135083
rect 444833 135010 444899 135013
rect 441876 135008 444899 135010
rect 441876 134952 444838 135008
rect 444894 134952 444899 135008
rect 441876 134950 444899 134952
rect 444833 134947 444899 134950
rect 169924 134814 172487 134816
rect 172421 134811 172487 134814
rect 369853 134602 369919 134605
rect 369853 134600 369962 134602
rect 369853 134544 369858 134600
rect 369914 134544 369962 134600
rect 369853 134539 369962 134544
rect 172237 134330 172303 134333
rect 169924 134328 172303 134330
rect 169924 134272 172242 134328
rect 172298 134272 172303 134328
rect 369902 134300 369962 134539
rect 169924 134270 172303 134272
rect 172237 134267 172303 134270
rect 370037 134058 370103 134061
rect 369902 134056 370103 134058
rect 369902 134000 370042 134056
rect 370098 134000 370103 134056
rect 369902 133998 370103 134000
rect 171225 133922 171291 133925
rect 169924 133920 171291 133922
rect 169924 133864 171230 133920
rect 171286 133864 171291 133920
rect 369902 133892 369962 133998
rect 370037 133995 370103 133998
rect 444649 133922 444715 133925
rect 441876 133920 444715 133922
rect 169924 133862 171291 133864
rect 441876 133864 444654 133920
rect 444710 133864 444715 133920
rect 441876 133862 444715 133864
rect 171225 133859 171291 133862
rect 444649 133859 444715 133862
rect 369945 133650 370011 133653
rect 369902 133648 370011 133650
rect 369902 133592 369950 133648
rect 370006 133592 370011 133648
rect 369902 133587 370011 133592
rect 197537 133514 197603 133517
rect 197537 133512 200100 133514
rect 197537 133456 197542 133512
rect 197598 133456 200100 133512
rect 197537 133454 200100 133456
rect 197537 133451 197603 133454
rect 172421 133378 172487 133381
rect 169924 133376 172487 133378
rect 169924 133320 172426 133376
rect 172482 133320 172487 133376
rect 369902 133348 369962 133587
rect 169924 133318 172487 133320
rect 172421 133315 172487 133318
rect 303061 133242 303127 133245
rect 299828 133240 303127 133242
rect 299828 133184 303066 133240
rect 303122 133184 303127 133240
rect 299828 133182 303127 133184
rect 303061 133179 303127 133182
rect 172329 132834 172395 132837
rect 370313 132834 370379 132837
rect 169924 132832 172395 132834
rect 169924 132776 172334 132832
rect 172390 132776 172395 132832
rect 169924 132774 172395 132776
rect 369932 132832 370379 132834
rect 369932 132776 370318 132832
rect 370374 132776 370379 132832
rect 369932 132774 370379 132776
rect 172329 132771 172395 132774
rect 370313 132771 370379 132774
rect 444557 132698 444623 132701
rect 441876 132696 444623 132698
rect 441876 132640 444562 132696
rect 444618 132640 444623 132696
rect 441876 132638 444623 132640
rect 444557 132635 444623 132638
rect 369301 132426 369367 132429
rect 369301 132424 369410 132426
rect 369301 132368 369306 132424
rect 369362 132368 369410 132424
rect 369301 132363 369410 132368
rect 171133 132290 171199 132293
rect 169924 132288 171199 132290
rect 169924 132232 171138 132288
rect 171194 132232 171199 132288
rect 369350 132260 369410 132363
rect 169924 132230 171199 132232
rect 171133 132227 171199 132230
rect 369485 132018 369551 132021
rect 369485 132016 369594 132018
rect 369485 131960 369490 132016
rect 369546 131960 369594 132016
rect 369485 131955 369594 131960
rect 172421 131746 172487 131749
rect 169924 131744 172487 131746
rect 169924 131688 172426 131744
rect 172482 131688 172487 131744
rect 369534 131716 369594 131955
rect 169924 131686 172487 131688
rect 172421 131683 172487 131686
rect 444465 131610 444531 131613
rect 441876 131608 444531 131610
rect 441876 131552 444470 131608
rect 444526 131552 444531 131608
rect 441876 131550 444531 131552
rect 444465 131547 444531 131550
rect 369301 131474 369367 131477
rect 369301 131472 369410 131474
rect 369301 131416 369306 131472
rect 369362 131416 369410 131472
rect 369301 131411 369410 131416
rect 197905 131338 197971 131341
rect 197905 131336 200100 131338
rect 197905 131280 197910 131336
rect 197966 131280 200100 131336
rect 197905 131278 200100 131280
rect 197905 131275 197971 131278
rect 171501 131202 171567 131205
rect 169924 131200 171567 131202
rect 169924 131144 171506 131200
rect 171562 131144 171567 131200
rect 369350 131172 369410 131411
rect 169924 131142 171567 131144
rect 171501 131139 171567 131142
rect 172329 130658 172395 130661
rect 370221 130658 370287 130661
rect 169924 130656 172395 130658
rect 169924 130600 172334 130656
rect 172390 130600 172395 130656
rect 169924 130598 172395 130600
rect 369932 130656 370287 130658
rect 369932 130600 370226 130656
rect 370282 130600 370287 130656
rect 369932 130598 370287 130600
rect 172329 130595 172395 130598
rect 370221 130595 370287 130598
rect 442993 130386 443059 130389
rect 443913 130386 443979 130389
rect 441876 130384 443979 130386
rect 441876 130328 442998 130384
rect 443054 130328 443918 130384
rect 443974 130328 443979 130384
rect 441876 130326 443979 130328
rect 442993 130323 443059 130326
rect 443913 130323 443979 130326
rect 171869 130114 171935 130117
rect 302785 130114 302851 130117
rect 370497 130114 370563 130117
rect 169924 130112 171935 130114
rect 169924 130056 171874 130112
rect 171930 130056 171935 130112
rect 169924 130054 171935 130056
rect 299828 130112 302851 130114
rect 299828 130056 302790 130112
rect 302846 130056 302851 130112
rect 369932 130112 370563 130114
rect 369932 130084 370502 130112
rect 299828 130054 302851 130056
rect 171869 130051 171935 130054
rect 302785 130051 302851 130054
rect 369902 130056 370502 130084
rect 370558 130056 370563 130112
rect 369902 130054 370563 130056
rect 369902 129845 369962 130054
rect 370497 130051 370563 130054
rect 369902 129840 370011 129845
rect 369902 129784 369950 129840
rect 370006 129784 370011 129840
rect 369902 129782 370011 129784
rect 369945 129779 370011 129782
rect 172421 129570 172487 129573
rect 169924 129568 172487 129570
rect 169924 129512 172426 129568
rect 172482 129512 172487 129568
rect 169924 129510 172487 129512
rect 172421 129507 172487 129510
rect 369902 129165 369962 129540
rect 443637 129298 443703 129301
rect 441876 129296 443703 129298
rect 441876 129240 443642 129296
rect 443698 129240 443703 129296
rect 441876 129238 443703 129240
rect 443637 129235 443703 129238
rect 197353 129162 197419 129165
rect 197353 129160 200100 129162
rect 197353 129104 197358 129160
rect 197414 129104 200100 129160
rect 197353 129102 200100 129104
rect 369853 129160 369962 129165
rect 369853 129104 369858 129160
rect 369914 129104 369962 129160
rect 369853 129102 369962 129104
rect 197353 129099 197419 129102
rect 369853 129099 369919 129102
rect 172053 129026 172119 129029
rect 370313 129026 370379 129029
rect 169924 129024 172119 129026
rect 169924 128968 172058 129024
rect 172114 128968 172119 129024
rect 169924 128966 172119 128968
rect 369932 129024 370379 129026
rect 369932 128968 370318 129024
rect 370374 128968 370379 129024
rect 369932 128966 370379 128968
rect 172053 128963 172119 128966
rect 370313 128963 370379 128966
rect 370037 128618 370103 128621
rect 371969 128618 372035 128621
rect 369902 128616 372035 128618
rect 369902 128560 370042 128616
rect 370098 128560 371974 128616
rect 372030 128560 372035 128616
rect 369902 128558 372035 128560
rect 171869 128482 171935 128485
rect 169924 128480 171935 128482
rect 169924 128424 171874 128480
rect 171930 128424 171935 128480
rect 369902 128452 369962 128558
rect 370037 128555 370103 128558
rect 371969 128555 372035 128558
rect 169924 128422 171935 128424
rect 171869 128419 171935 128422
rect 443085 128074 443151 128077
rect 444373 128074 444439 128077
rect 441876 128072 444439 128074
rect 441876 128016 443090 128072
rect 443146 128016 444378 128072
rect 444434 128016 444439 128072
rect 441876 128014 444439 128016
rect 443085 128011 443151 128014
rect 444373 128011 444439 128014
rect 171961 127938 172027 127941
rect 371233 127938 371299 127941
rect 372061 127938 372127 127941
rect 169924 127936 172027 127938
rect 169924 127880 171966 127936
rect 172022 127880 172027 127936
rect 169924 127878 172027 127880
rect 369932 127936 372127 127938
rect 369932 127880 371238 127936
rect 371294 127880 372066 127936
rect 372122 127880 372127 127936
rect 369932 127878 372127 127880
rect 171961 127875 172027 127878
rect 371233 127875 371299 127878
rect 372061 127875 372127 127878
rect 171777 127394 171843 127397
rect 370129 127394 370195 127397
rect 371877 127394 371943 127397
rect 169924 127392 171843 127394
rect 169924 127336 171782 127392
rect 171838 127336 171843 127392
rect 169924 127334 171843 127336
rect 369932 127392 371943 127394
rect 369932 127336 370134 127392
rect 370190 127336 371882 127392
rect 371938 127336 371943 127392
rect 369932 127334 371943 127336
rect 171777 127331 171843 127334
rect 370129 127331 370195 127334
rect 371877 127331 371943 127334
rect 197353 126986 197419 126989
rect 445661 126986 445727 126989
rect 197353 126984 200100 126986
rect 197353 126928 197358 126984
rect 197414 126928 200100 126984
rect 441876 126984 445727 126986
rect 441876 126956 445666 126984
rect 197353 126926 200100 126928
rect 441846 126928 445666 126956
rect 445722 126928 445727 126984
rect 441846 126926 445727 126928
rect 197353 126923 197419 126926
rect 172237 126850 172303 126853
rect 302601 126850 302667 126853
rect 371785 126850 371851 126853
rect 169924 126848 172303 126850
rect 169924 126792 172242 126848
rect 172298 126792 172303 126848
rect 169924 126790 172303 126792
rect 299828 126848 302667 126850
rect 299828 126792 302606 126848
rect 302662 126792 302667 126848
rect 299828 126790 302667 126792
rect 369932 126848 371851 126850
rect 369932 126792 371790 126848
rect 371846 126792 371851 126848
rect 369932 126790 371851 126792
rect 172237 126787 172303 126790
rect 302601 126787 302667 126790
rect 371785 126787 371851 126790
rect 441846 126445 441906 126926
rect 445661 126923 445727 126926
rect 441846 126440 441955 126445
rect 441846 126384 441894 126440
rect 441950 126384 441955 126440
rect 441846 126382 441955 126384
rect 441889 126379 441955 126382
rect 172329 126306 172395 126309
rect 370405 126306 370471 126309
rect 169924 126304 172395 126306
rect 169924 126248 172334 126304
rect 172390 126248 172395 126304
rect 169924 126246 172395 126248
rect 369932 126304 370471 126306
rect 369932 126248 370410 126304
rect 370466 126248 370471 126304
rect 369932 126246 370471 126248
rect 172329 126243 172395 126246
rect 370405 126243 370471 126246
rect 580165 126034 580231 126037
rect 583520 126034 584960 126124
rect 580165 126032 584960 126034
rect 580165 125976 580170 126032
rect 580226 125976 584960 126032
rect 580165 125974 584960 125976
rect 580165 125971 580231 125974
rect 583520 125884 584960 125974
rect 172421 125762 172487 125765
rect 370589 125762 370655 125765
rect 372429 125762 372495 125765
rect 444373 125762 444439 125765
rect 169924 125760 172487 125762
rect 169924 125704 172426 125760
rect 172482 125704 172487 125760
rect 169924 125702 172487 125704
rect 369932 125760 372495 125762
rect 369932 125704 370594 125760
rect 370650 125704 372434 125760
rect 372490 125704 372495 125760
rect 441692 125760 444439 125762
rect 441692 125732 444378 125760
rect 369932 125702 372495 125704
rect 172421 125699 172487 125702
rect 370589 125699 370655 125702
rect 372429 125699 372495 125702
rect 441662 125704 444378 125732
rect 444434 125704 444439 125760
rect 441662 125702 444439 125704
rect 441662 125493 441722 125702
rect 444373 125699 444439 125702
rect 441613 125488 441722 125493
rect 441613 125432 441618 125488
rect 441674 125432 441722 125488
rect 441613 125430 441722 125432
rect 441613 125427 441679 125430
rect 172421 125218 172487 125221
rect 371325 125218 371391 125221
rect 169924 125216 172487 125218
rect 169924 125160 172426 125216
rect 172482 125160 172487 125216
rect 169924 125158 172487 125160
rect 369932 125216 371391 125218
rect 369932 125160 371330 125216
rect 371386 125160 371391 125216
rect 369932 125158 371391 125160
rect 172421 125155 172487 125158
rect 371325 125155 371391 125158
rect 441889 124946 441955 124949
rect 441846 124944 441955 124946
rect 441846 124888 441894 124944
rect 441950 124888 441955 124944
rect 441846 124883 441955 124888
rect 198549 124810 198615 124813
rect 369945 124810 370011 124813
rect 370497 124810 370563 124813
rect 198549 124808 200100 124810
rect 198549 124752 198554 124808
rect 198610 124752 200100 124808
rect 198549 124750 200100 124752
rect 369902 124808 370563 124810
rect 369902 124752 369950 124808
rect 370006 124752 370502 124808
rect 370558 124752 370563 124808
rect 369902 124750 370563 124752
rect 198549 124747 198615 124750
rect 369902 124747 370011 124750
rect 370497 124747 370563 124750
rect 171685 124674 171751 124677
rect 169924 124672 171751 124674
rect 169924 124616 171690 124672
rect 171746 124616 171751 124672
rect 369902 124644 369962 124747
rect 441846 124644 441906 124883
rect 169924 124614 171751 124616
rect 171685 124611 171751 124614
rect 369853 124402 369919 124405
rect 369853 124400 369962 124402
rect 369853 124344 369858 124400
rect 369914 124344 369962 124400
rect 369853 124339 369962 124344
rect 172145 124266 172211 124269
rect 169924 124264 172211 124266
rect 169924 124208 172150 124264
rect 172206 124208 172211 124264
rect 369902 124266 369962 124339
rect 370773 124266 370839 124269
rect 369902 124264 370839 124266
rect 369902 124236 370778 124264
rect 169924 124206 172211 124208
rect 369932 124208 370778 124236
rect 370834 124208 370839 124264
rect 369932 124206 370839 124208
rect 172145 124203 172211 124206
rect 370773 124203 370839 124206
rect 362769 123996 362835 123997
rect 362718 123932 362724 123996
rect 362788 123994 362835 123996
rect 365161 123994 365227 123997
rect 365294 123994 365300 123996
rect 362788 123992 362880 123994
rect 362830 123936 362880 123992
rect 362788 123934 362880 123936
rect 365161 123992 365300 123994
rect 365161 123936 365166 123992
rect 365222 123936 365300 123992
rect 365161 123934 365300 123936
rect 362788 123932 362835 123934
rect 362769 123931 362835 123932
rect 365161 123931 365227 123934
rect 365294 123932 365300 123934
rect 365364 123932 365370 123996
rect -960 123572 480 123812
rect 302693 123722 302759 123725
rect 299828 123720 302759 123722
rect 299828 123664 302698 123720
rect 302754 123664 302759 123720
rect 299828 123662 302759 123664
rect 302693 123659 302759 123662
rect 197997 122634 198063 122637
rect 197997 122632 200100 122634
rect 197997 122576 198002 122632
rect 198058 122576 200100 122632
rect 197997 122574 200100 122576
rect 197997 122571 198063 122574
rect 302785 120594 302851 120597
rect 299828 120592 302851 120594
rect 299828 120536 302790 120592
rect 302846 120536 302851 120592
rect 299828 120534 302851 120536
rect 302785 120531 302851 120534
rect 197537 120458 197603 120461
rect 197537 120456 200100 120458
rect 197537 120400 197542 120456
rect 197598 120400 200100 120456
rect 197537 120398 200100 120400
rect 197537 120395 197603 120398
rect 198089 118282 198155 118285
rect 198089 118280 200100 118282
rect 198089 118224 198094 118280
rect 198150 118224 200100 118280
rect 198089 118222 200100 118224
rect 198089 118219 198155 118222
rect 302785 117330 302851 117333
rect 299828 117328 302851 117330
rect 299828 117272 302790 117328
rect 302846 117272 302851 117328
rect 299828 117270 302851 117272
rect 302785 117267 302851 117270
rect 197537 116106 197603 116109
rect 197537 116104 200100 116106
rect 197537 116048 197542 116104
rect 197598 116048 200100 116104
rect 197537 116046 200100 116048
rect 197537 116043 197603 116046
rect 302969 114202 303035 114205
rect 299828 114200 303035 114202
rect 299828 114144 302974 114200
rect 303030 114144 303035 114200
rect 299828 114142 303035 114144
rect 302969 114139 303035 114142
rect 197353 113930 197419 113933
rect 197353 113928 200100 113930
rect 197353 113872 197358 113928
rect 197414 113872 200100 113928
rect 197353 113870 200100 113872
rect 197353 113867 197419 113870
rect 579797 112842 579863 112845
rect 583520 112842 584960 112932
rect 579797 112840 584960 112842
rect 579797 112784 579802 112840
rect 579858 112784 584960 112840
rect 579797 112782 584960 112784
rect 579797 112779 579863 112782
rect 583520 112692 584960 112782
rect 197353 111754 197419 111757
rect 197353 111752 200100 111754
rect 197353 111696 197358 111752
rect 197414 111696 200100 111752
rect 197353 111694 200100 111696
rect 197353 111691 197419 111694
rect 302325 111074 302391 111077
rect 299828 111072 302391 111074
rect 299828 111016 302330 111072
rect 302386 111016 302391 111072
rect 299828 111014 302391 111016
rect 302325 111011 302391 111014
rect -960 110666 480 110756
rect 3417 110666 3483 110669
rect -960 110664 3483 110666
rect -960 110608 3422 110664
rect 3478 110608 3483 110664
rect -960 110606 3483 110608
rect -960 110516 480 110606
rect 3417 110603 3483 110606
rect 197997 109578 198063 109581
rect 197997 109576 200100 109578
rect 197997 109520 198002 109576
rect 198058 109520 200100 109576
rect 197997 109518 200100 109520
rect 197997 109515 198063 109518
rect 302785 107810 302851 107813
rect 299828 107808 302851 107810
rect 299828 107752 302790 107808
rect 302846 107752 302851 107808
rect 299828 107750 302851 107752
rect 302785 107747 302851 107750
rect 198549 107402 198615 107405
rect 198549 107400 200100 107402
rect 198549 107344 198554 107400
rect 198610 107344 200100 107400
rect 198549 107342 200100 107344
rect 198549 107339 198615 107342
rect 197537 105226 197603 105229
rect 197537 105224 200100 105226
rect 197537 105168 197542 105224
rect 197598 105168 200100 105224
rect 197537 105166 200100 105168
rect 197537 105163 197603 105166
rect 302877 104682 302943 104685
rect 299828 104680 302943 104682
rect 299828 104624 302882 104680
rect 302938 104624 302943 104680
rect 299828 104622 302943 104624
rect 302877 104619 302943 104622
rect 197905 103050 197971 103053
rect 197905 103048 200100 103050
rect 197905 102992 197910 103048
rect 197966 102992 200100 103048
rect 197905 102990 200100 102992
rect 197905 102987 197971 102990
rect 302785 101554 302851 101557
rect 299828 101552 302851 101554
rect 299828 101496 302790 101552
rect 302846 101496 302851 101552
rect 299828 101494 302851 101496
rect 302785 101491 302851 101494
rect 197537 101010 197603 101013
rect 197537 101008 200100 101010
rect 197537 100952 197542 101008
rect 197598 100952 200100 101008
rect 197537 100950 200100 100952
rect 197537 100947 197603 100950
rect 580165 99514 580231 99517
rect 583520 99514 584960 99604
rect 580165 99512 584960 99514
rect 580165 99456 580170 99512
rect 580226 99456 584960 99512
rect 580165 99454 584960 99456
rect 580165 99451 580231 99454
rect 583520 99364 584960 99454
rect -960 97610 480 97700
rect 3417 97610 3483 97613
rect -960 97608 3483 97610
rect -960 97552 3422 97608
rect 3478 97552 3483 97608
rect -960 97550 3483 97552
rect -960 97460 480 97550
rect 3417 97547 3483 97550
rect 50337 97610 50403 97613
rect 206093 97610 206159 97613
rect 50337 97608 206159 97610
rect 50337 97552 50342 97608
rect 50398 97552 206098 97608
rect 206154 97552 206159 97608
rect 50337 97550 206159 97552
rect 50337 97547 50403 97550
rect 206093 97547 206159 97550
rect 39297 97474 39363 97477
rect 203517 97474 203583 97477
rect 39297 97472 203583 97474
rect 39297 97416 39302 97472
rect 39358 97416 203522 97472
rect 203578 97416 203583 97472
rect 39297 97414 203583 97416
rect 39297 97411 39363 97414
rect 203517 97411 203583 97414
rect 279325 97474 279391 97477
rect 436737 97474 436803 97477
rect 279325 97472 436803 97474
rect 279325 97416 279330 97472
rect 279386 97416 436742 97472
rect 436798 97416 436803 97472
rect 279325 97414 436803 97416
rect 279325 97411 279391 97414
rect 436737 97411 436803 97414
rect 38561 97338 38627 97341
rect 206553 97338 206619 97341
rect 38561 97336 206619 97338
rect 38561 97280 38566 97336
rect 38622 97280 206558 97336
rect 206614 97280 206619 97336
rect 38561 97278 206619 97280
rect 38561 97275 38627 97278
rect 206553 97275 206619 97278
rect 280521 97338 280587 97341
rect 443637 97338 443703 97341
rect 280521 97336 443703 97338
rect 280521 97280 280526 97336
rect 280582 97280 443642 97336
rect 443698 97280 443703 97336
rect 280521 97278 443703 97280
rect 280521 97275 280587 97278
rect 443637 97275 443703 97278
rect 32397 97202 32463 97205
rect 204897 97202 204963 97205
rect 32397 97200 204963 97202
rect 32397 97144 32402 97200
rect 32458 97144 204902 97200
rect 204958 97144 204963 97200
rect 32397 97142 204963 97144
rect 32397 97139 32463 97142
rect 204897 97139 204963 97142
rect 282637 97202 282703 97205
rect 283005 97202 283071 97205
rect 282637 97200 283071 97202
rect 282637 97144 282642 97200
rect 282698 97144 283010 97200
rect 283066 97144 283071 97200
rect 282637 97142 283071 97144
rect 282637 97139 282703 97142
rect 283005 97139 283071 97142
rect 299105 97202 299171 97205
rect 580257 97202 580323 97205
rect 299105 97200 580323 97202
rect 299105 97144 299110 97200
rect 299166 97144 580262 97200
rect 580318 97144 580323 97200
rect 299105 97142 580323 97144
rect 299105 97139 299171 97142
rect 580257 97139 580323 97142
rect 274173 97066 274239 97069
rect 278681 97066 278747 97069
rect 274173 97064 278747 97066
rect 274173 97008 274178 97064
rect 274234 97008 278686 97064
rect 278742 97008 278747 97064
rect 274173 97006 278747 97008
rect 274173 97003 274239 97006
rect 278681 97003 278747 97006
rect 289813 95978 289879 95981
rect 525793 95978 525859 95981
rect 289813 95976 525859 95978
rect 289813 95920 289818 95976
rect 289874 95920 525798 95976
rect 525854 95920 525859 95976
rect 289813 95918 525859 95920
rect 289813 95915 289879 95918
rect 525793 95915 525859 95918
rect 294045 95842 294111 95845
rect 550633 95842 550699 95845
rect 294045 95840 550699 95842
rect 294045 95784 294050 95840
rect 294106 95784 550638 95840
rect 550694 95784 550699 95840
rect 294045 95782 550699 95784
rect 294045 95779 294111 95782
rect 550633 95779 550699 95782
rect 580165 86186 580231 86189
rect 583520 86186 584960 86276
rect 580165 86184 584960 86186
rect 580165 86128 580170 86184
rect 580226 86128 584960 86184
rect 580165 86126 584960 86128
rect 580165 86123 580231 86126
rect 583520 86036 584960 86126
rect -960 84690 480 84780
rect 3141 84690 3207 84693
rect -960 84688 3207 84690
rect -960 84632 3146 84688
rect 3202 84632 3207 84688
rect -960 84630 3207 84632
rect -960 84540 480 84630
rect 3141 84627 3207 84630
rect 579981 72994 580047 72997
rect 583520 72994 584960 73084
rect 579981 72992 584960 72994
rect 579981 72936 579986 72992
rect 580042 72936 584960 72992
rect 579981 72934 584960 72936
rect 579981 72931 580047 72934
rect 583520 72844 584960 72934
rect -960 71634 480 71724
rect 2773 71634 2839 71637
rect -960 71632 2839 71634
rect -960 71576 2778 71632
rect 2834 71576 2839 71632
rect -960 71574 2839 71576
rect -960 71484 480 71574
rect 2773 71571 2839 71574
rect 580165 59666 580231 59669
rect 583520 59666 584960 59756
rect 580165 59664 584960 59666
rect 580165 59608 580170 59664
rect 580226 59608 584960 59664
rect 580165 59606 584960 59608
rect 580165 59603 580231 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 3049 58578 3115 58581
rect -960 58576 3115 58578
rect -960 58520 3054 58576
rect 3110 58520 3115 58576
rect -960 58518 3115 58520
rect -960 58428 480 58518
rect 3049 58515 3115 58518
rect 582465 46338 582531 46341
rect 583520 46338 584960 46428
rect 582465 46336 584960 46338
rect 582465 46280 582470 46336
rect 582526 46280 584960 46336
rect 582465 46278 584960 46280
rect 582465 46275 582531 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 3417 45522 3483 45525
rect -960 45520 3483 45522
rect -960 45464 3422 45520
rect 3478 45464 3483 45520
rect -960 45462 3483 45464
rect -960 45372 480 45462
rect 3417 45459 3483 45462
rect 580165 33146 580231 33149
rect 583520 33146 584960 33236
rect 580165 33144 584960 33146
rect 580165 33088 580170 33144
rect 580226 33088 584960 33144
rect 580165 33086 584960 33088
rect 580165 33083 580231 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 3141 32466 3207 32469
rect -960 32464 3207 32466
rect -960 32408 3146 32464
rect 3202 32408 3207 32464
rect -960 32406 3207 32408
rect -960 32316 480 32406
rect 3141 32403 3207 32406
rect 580165 19818 580231 19821
rect 583520 19818 584960 19908
rect 580165 19816 584960 19818
rect 580165 19760 580170 19816
rect 580226 19760 584960 19816
rect 580165 19758 584960 19760
rect 580165 19755 580231 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3417 19410 3483 19413
rect -960 19408 3483 19410
rect -960 19352 3422 19408
rect 3478 19352 3483 19408
rect -960 19350 3483 19352
rect -960 19260 480 19350
rect 3417 19347 3483 19350
rect 582373 6626 582439 6629
rect 583520 6626 584960 6716
rect 582373 6624 584960 6626
rect -960 6490 480 6580
rect 582373 6568 582378 6624
rect 582434 6568 584960 6624
rect 582373 6566 584960 6568
rect 582373 6563 582439 6566
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect 583520 6476 584960 6566
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
<< via3 >>
rect 371924 353500 371988 353564
rect 371740 352956 371804 353020
rect 372108 352412 372172 352476
rect 371556 351324 371620 351388
rect 371188 350780 371252 350844
rect 361620 337724 361684 337788
rect 364380 337724 364444 337788
rect 371372 281556 371436 281620
rect 371924 281556 371988 281620
rect 371740 281012 371804 281076
rect 372108 280468 372172 280532
rect 371556 279380 371620 279444
rect 371188 278836 371252 278900
rect 370084 276932 370148 276996
rect 370268 275300 370332 275364
rect 361620 267820 361684 267884
rect 364380 266188 364444 266252
rect 361620 266052 361684 266116
rect 371372 224980 371436 225044
rect 371740 223892 371804 223956
rect 371372 209476 371436 209540
rect 371740 208932 371804 208996
rect 371924 208388 371988 208452
rect 371556 207300 371620 207364
rect 371924 207300 371988 207364
rect 371188 206756 371252 206820
rect 372292 206756 372356 206820
rect 370084 205260 370148 205324
rect 370268 203628 370332 203692
rect 364380 196012 364444 196076
rect 371372 196012 371436 196076
rect 372476 195196 372540 195260
rect 361620 194516 361684 194580
rect 362724 194516 362788 194580
rect 365300 194516 365364 194580
rect 371740 175612 371804 175676
rect 372292 175204 372356 175268
rect 371924 174932 371988 174996
rect 372292 173164 372356 173228
rect 371924 171668 371988 171732
rect 372292 162692 372356 162756
rect 371924 152900 371988 152964
rect 371372 137532 371436 137596
rect 372476 136988 372540 137052
rect 371740 136444 371804 136508
rect 362724 123992 362788 123996
rect 362724 123936 362774 123992
rect 362774 123936 362788 123992
rect 362724 123932 362788 123936
rect 365300 123932 365364 123996
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 680614 -8106 711002
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 -8106 680614
rect -8726 680294 -8106 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 -8106 680294
rect -8726 644614 -8106 680058
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 -8106 644614
rect -8726 644294 -8106 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 -8106 644294
rect -8726 608614 -8106 644058
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 -8106 608614
rect -8726 608294 -8106 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 -8106 608294
rect -8726 572614 -8106 608058
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 -8106 572614
rect -8726 572294 -8106 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 -8106 572294
rect -8726 536614 -8106 572058
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 -8106 536614
rect -8726 536294 -8106 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 -8106 536294
rect -8726 500614 -8106 536058
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 -8106 500614
rect -8726 500294 -8106 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 -8106 500294
rect -8726 464614 -8106 500058
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 -8106 464614
rect -8726 464294 -8106 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 -8106 464294
rect -8726 428614 -8106 464058
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 -8106 428614
rect -8726 428294 -8106 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 -8106 428294
rect -8726 392614 -8106 428058
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 -8106 392614
rect -8726 392294 -8106 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 -8106 392294
rect -8726 356614 -8106 392058
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 -8106 356614
rect -8726 356294 -8106 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 -8106 356294
rect -8726 320614 -8106 356058
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 -8106 320614
rect -8726 320294 -8106 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 -8106 320294
rect -8726 284614 -8106 320058
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 -8106 284614
rect -8726 284294 -8106 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 -8106 284294
rect -8726 248614 -8106 284058
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 -8106 248614
rect -8726 248294 -8106 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 -8106 248294
rect -8726 212614 -8106 248058
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 -8106 212614
rect -8726 212294 -8106 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 -8106 212294
rect -8726 176614 -8106 212058
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 -8106 176614
rect -8726 176294 -8106 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 -8106 176294
rect -8726 140614 -8106 176058
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 -8106 140614
rect -8726 140294 -8106 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 -8106 140294
rect -8726 104614 -8106 140058
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 -8106 104614
rect -8726 104294 -8106 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 -8106 104294
rect -8726 68614 -8106 104058
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 -8106 68614
rect -8726 68294 -8106 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 -8106 68294
rect -8726 32614 -8106 68058
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 -8106 32614
rect -8726 32294 -8106 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 -8106 32294
rect -8726 -7066 -8106 32058
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 698614 -7146 710042
rect 12954 710598 13574 711590
rect 12954 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 13574 710598
rect 12954 710278 13574 710362
rect 12954 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 13574 710278
rect -7766 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 -7146 698614
rect -7766 698294 -7146 698378
rect -7766 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 -7146 698294
rect -7766 662614 -7146 698058
rect -7766 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 -7146 662614
rect -7766 662294 -7146 662378
rect -7766 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 -7146 662294
rect -7766 626614 -7146 662058
rect -7766 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 -7146 626614
rect -7766 626294 -7146 626378
rect -7766 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 -7146 626294
rect -7766 590614 -7146 626058
rect -7766 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 -7146 590614
rect -7766 590294 -7146 590378
rect -7766 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 -7146 590294
rect -7766 554614 -7146 590058
rect -7766 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 -7146 554614
rect -7766 554294 -7146 554378
rect -7766 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 -7146 554294
rect -7766 518614 -7146 554058
rect -7766 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 -7146 518614
rect -7766 518294 -7146 518378
rect -7766 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 -7146 518294
rect -7766 482614 -7146 518058
rect -7766 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 -7146 482614
rect -7766 482294 -7146 482378
rect -7766 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 -7146 482294
rect -7766 446614 -7146 482058
rect -7766 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 -7146 446614
rect -7766 446294 -7146 446378
rect -7766 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 -7146 446294
rect -7766 410614 -7146 446058
rect -7766 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 -7146 410614
rect -7766 410294 -7146 410378
rect -7766 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 -7146 410294
rect -7766 374614 -7146 410058
rect -7766 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 -7146 374614
rect -7766 374294 -7146 374378
rect -7766 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 -7146 374294
rect -7766 338614 -7146 374058
rect -7766 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 -7146 338614
rect -7766 338294 -7146 338378
rect -7766 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 -7146 338294
rect -7766 302614 -7146 338058
rect -7766 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 -7146 302614
rect -7766 302294 -7146 302378
rect -7766 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 -7146 302294
rect -7766 266614 -7146 302058
rect -7766 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 -7146 266614
rect -7766 266294 -7146 266378
rect -7766 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 -7146 266294
rect -7766 230614 -7146 266058
rect -7766 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 -7146 230614
rect -7766 230294 -7146 230378
rect -7766 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 -7146 230294
rect -7766 194614 -7146 230058
rect -7766 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 -7146 194614
rect -7766 194294 -7146 194378
rect -7766 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 -7146 194294
rect -7766 158614 -7146 194058
rect -7766 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 -7146 158614
rect -7766 158294 -7146 158378
rect -7766 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 -7146 158294
rect -7766 122614 -7146 158058
rect -7766 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 -7146 122614
rect -7766 122294 -7146 122378
rect -7766 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 -7146 122294
rect -7766 86614 -7146 122058
rect -7766 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 -7146 86614
rect -7766 86294 -7146 86378
rect -7766 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 -7146 86294
rect -7766 50614 -7146 86058
rect -7766 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 -7146 50614
rect -7766 50294 -7146 50378
rect -7766 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 -7146 50294
rect -7766 14614 -7146 50058
rect -7766 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 -7146 14614
rect -7766 14294 -7146 14378
rect -7766 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 -7146 14294
rect -7766 -6106 -7146 14058
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 676894 -6186 709082
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 -6186 676894
rect -6806 676574 -6186 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 -6186 676574
rect -6806 640894 -6186 676338
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 -6186 640894
rect -6806 640574 -6186 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 -6186 640574
rect -6806 604894 -6186 640338
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 -6186 604894
rect -6806 604574 -6186 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 -6186 604574
rect -6806 568894 -6186 604338
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 -6186 568894
rect -6806 568574 -6186 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 -6186 568574
rect -6806 532894 -6186 568338
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 -6186 532894
rect -6806 532574 -6186 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 -6186 532574
rect -6806 496894 -6186 532338
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 -6186 496894
rect -6806 496574 -6186 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 -6186 496574
rect -6806 460894 -6186 496338
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 -6186 460894
rect -6806 460574 -6186 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 -6186 460574
rect -6806 424894 -6186 460338
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 -6186 424894
rect -6806 424574 -6186 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 -6186 424574
rect -6806 388894 -6186 424338
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 -6186 388894
rect -6806 388574 -6186 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 -6186 388574
rect -6806 352894 -6186 388338
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 -6186 352894
rect -6806 352574 -6186 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 -6186 352574
rect -6806 316894 -6186 352338
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 -6186 316894
rect -6806 316574 -6186 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 -6186 316574
rect -6806 280894 -6186 316338
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 -6186 280894
rect -6806 280574 -6186 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 -6186 280574
rect -6806 244894 -6186 280338
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 -6186 244894
rect -6806 244574 -6186 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 -6186 244574
rect -6806 208894 -6186 244338
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 -6186 208894
rect -6806 208574 -6186 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 -6186 208574
rect -6806 172894 -6186 208338
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 -6186 172894
rect -6806 172574 -6186 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 -6186 172574
rect -6806 136894 -6186 172338
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 -6186 136894
rect -6806 136574 -6186 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 -6186 136574
rect -6806 100894 -6186 136338
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 -6186 100894
rect -6806 100574 -6186 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 -6186 100574
rect -6806 64894 -6186 100338
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 -6186 64894
rect -6806 64574 -6186 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 -6186 64574
rect -6806 28894 -6186 64338
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 -6186 28894
rect -6806 28574 -6186 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 -6186 28574
rect -6806 -5146 -6186 28338
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 694894 -5226 708122
rect 9234 708678 9854 709670
rect 9234 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 9854 708678
rect 9234 708358 9854 708442
rect 9234 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 9854 708358
rect -5846 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 -5226 694894
rect -5846 694574 -5226 694658
rect -5846 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 -5226 694574
rect -5846 658894 -5226 694338
rect -5846 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 -5226 658894
rect -5846 658574 -5226 658658
rect -5846 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 -5226 658574
rect -5846 622894 -5226 658338
rect -5846 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 -5226 622894
rect -5846 622574 -5226 622658
rect -5846 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 -5226 622574
rect -5846 586894 -5226 622338
rect -5846 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 -5226 586894
rect -5846 586574 -5226 586658
rect -5846 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 -5226 586574
rect -5846 550894 -5226 586338
rect -5846 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 -5226 550894
rect -5846 550574 -5226 550658
rect -5846 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 -5226 550574
rect -5846 514894 -5226 550338
rect -5846 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 -5226 514894
rect -5846 514574 -5226 514658
rect -5846 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 -5226 514574
rect -5846 478894 -5226 514338
rect -5846 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 -5226 478894
rect -5846 478574 -5226 478658
rect -5846 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 -5226 478574
rect -5846 442894 -5226 478338
rect -5846 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 -5226 442894
rect -5846 442574 -5226 442658
rect -5846 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 -5226 442574
rect -5846 406894 -5226 442338
rect -5846 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 -5226 406894
rect -5846 406574 -5226 406658
rect -5846 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 -5226 406574
rect -5846 370894 -5226 406338
rect -5846 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 -5226 370894
rect -5846 370574 -5226 370658
rect -5846 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 -5226 370574
rect -5846 334894 -5226 370338
rect -5846 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 -5226 334894
rect -5846 334574 -5226 334658
rect -5846 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 -5226 334574
rect -5846 298894 -5226 334338
rect -5846 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 -5226 298894
rect -5846 298574 -5226 298658
rect -5846 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 -5226 298574
rect -5846 262894 -5226 298338
rect -5846 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 -5226 262894
rect -5846 262574 -5226 262658
rect -5846 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 -5226 262574
rect -5846 226894 -5226 262338
rect -5846 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 -5226 226894
rect -5846 226574 -5226 226658
rect -5846 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 -5226 226574
rect -5846 190894 -5226 226338
rect -5846 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 -5226 190894
rect -5846 190574 -5226 190658
rect -5846 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 -5226 190574
rect -5846 154894 -5226 190338
rect -5846 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 -5226 154894
rect -5846 154574 -5226 154658
rect -5846 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 -5226 154574
rect -5846 118894 -5226 154338
rect -5846 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 -5226 118894
rect -5846 118574 -5226 118658
rect -5846 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 -5226 118574
rect -5846 82894 -5226 118338
rect -5846 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 -5226 82894
rect -5846 82574 -5226 82658
rect -5846 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 -5226 82574
rect -5846 46894 -5226 82338
rect -5846 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 -5226 46894
rect -5846 46574 -5226 46658
rect -5846 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 -5226 46574
rect -5846 10894 -5226 46338
rect -5846 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 -5226 10894
rect -5846 10574 -5226 10658
rect -5846 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 -5226 10574
rect -5846 -4186 -5226 10338
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 673174 -4266 707162
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 -4266 673174
rect -4886 672854 -4266 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 -4266 672854
rect -4886 637174 -4266 672618
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 -4266 637174
rect -4886 636854 -4266 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 -4266 636854
rect -4886 601174 -4266 636618
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 -4266 601174
rect -4886 600854 -4266 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 -4266 600854
rect -4886 565174 -4266 600618
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 -4266 565174
rect -4886 564854 -4266 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 -4266 564854
rect -4886 529174 -4266 564618
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 -4266 529174
rect -4886 528854 -4266 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 -4266 528854
rect -4886 493174 -4266 528618
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 -4266 493174
rect -4886 492854 -4266 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 -4266 492854
rect -4886 457174 -4266 492618
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 -4266 457174
rect -4886 456854 -4266 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 -4266 456854
rect -4886 421174 -4266 456618
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 -4266 421174
rect -4886 420854 -4266 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 -4266 420854
rect -4886 385174 -4266 420618
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 -4266 385174
rect -4886 384854 -4266 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 -4266 384854
rect -4886 349174 -4266 384618
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 -4266 349174
rect -4886 348854 -4266 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 -4266 348854
rect -4886 313174 -4266 348618
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 -4266 313174
rect -4886 312854 -4266 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 -4266 312854
rect -4886 277174 -4266 312618
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 -4266 277174
rect -4886 276854 -4266 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 -4266 276854
rect -4886 241174 -4266 276618
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 -4266 241174
rect -4886 240854 -4266 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 -4266 240854
rect -4886 205174 -4266 240618
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 -4266 205174
rect -4886 204854 -4266 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 -4266 204854
rect -4886 169174 -4266 204618
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 -4266 169174
rect -4886 168854 -4266 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 -4266 168854
rect -4886 133174 -4266 168618
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 -4266 133174
rect -4886 132854 -4266 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 -4266 132854
rect -4886 97174 -4266 132618
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 -4266 97174
rect -4886 96854 -4266 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 -4266 96854
rect -4886 61174 -4266 96618
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 -4266 61174
rect -4886 60854 -4266 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 -4266 60854
rect -4886 25174 -4266 60618
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 -4266 25174
rect -4886 24854 -4266 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 -4266 24854
rect -4886 -3226 -4266 24618
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 691174 -3306 706202
rect 5514 706758 6134 707750
rect 5514 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 6134 706758
rect 5514 706438 6134 706522
rect 5514 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 6134 706438
rect -3926 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 -3306 691174
rect -3926 690854 -3306 690938
rect -3926 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 -3306 690854
rect -3926 655174 -3306 690618
rect -3926 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 -3306 655174
rect -3926 654854 -3306 654938
rect -3926 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 -3306 654854
rect -3926 619174 -3306 654618
rect -3926 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 -3306 619174
rect -3926 618854 -3306 618938
rect -3926 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 -3306 618854
rect -3926 583174 -3306 618618
rect -3926 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 -3306 583174
rect -3926 582854 -3306 582938
rect -3926 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 -3306 582854
rect -3926 547174 -3306 582618
rect -3926 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 -3306 547174
rect -3926 546854 -3306 546938
rect -3926 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 -3306 546854
rect -3926 511174 -3306 546618
rect -3926 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 -3306 511174
rect -3926 510854 -3306 510938
rect -3926 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 -3306 510854
rect -3926 475174 -3306 510618
rect -3926 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 -3306 475174
rect -3926 474854 -3306 474938
rect -3926 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 -3306 474854
rect -3926 439174 -3306 474618
rect -3926 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 -3306 439174
rect -3926 438854 -3306 438938
rect -3926 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 -3306 438854
rect -3926 403174 -3306 438618
rect -3926 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 -3306 403174
rect -3926 402854 -3306 402938
rect -3926 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 -3306 402854
rect -3926 367174 -3306 402618
rect -3926 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 -3306 367174
rect -3926 366854 -3306 366938
rect -3926 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 -3306 366854
rect -3926 331174 -3306 366618
rect -3926 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 -3306 331174
rect -3926 330854 -3306 330938
rect -3926 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 -3306 330854
rect -3926 295174 -3306 330618
rect -3926 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 -3306 295174
rect -3926 294854 -3306 294938
rect -3926 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 -3306 294854
rect -3926 259174 -3306 294618
rect -3926 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 -3306 259174
rect -3926 258854 -3306 258938
rect -3926 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 -3306 258854
rect -3926 223174 -3306 258618
rect -3926 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 -3306 223174
rect -3926 222854 -3306 222938
rect -3926 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 -3306 222854
rect -3926 187174 -3306 222618
rect -3926 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 -3306 187174
rect -3926 186854 -3306 186938
rect -3926 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 -3306 186854
rect -3926 151174 -3306 186618
rect -3926 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 -3306 151174
rect -3926 150854 -3306 150938
rect -3926 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 -3306 150854
rect -3926 115174 -3306 150618
rect -3926 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 -3306 115174
rect -3926 114854 -3306 114938
rect -3926 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 -3306 114854
rect -3926 79174 -3306 114618
rect -3926 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 -3306 79174
rect -3926 78854 -3306 78938
rect -3926 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 -3306 78854
rect -3926 43174 -3306 78618
rect -3926 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 -3306 43174
rect -3926 42854 -3306 42938
rect -3926 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 -3306 42854
rect -3926 7174 -3306 42618
rect -3926 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 -3306 7174
rect -3926 6854 -3306 6938
rect -3926 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 -3306 6854
rect -3926 -2266 -3306 6618
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 669454 -2346 705242
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 -2346 669454
rect -2966 669134 -2346 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 -2346 669134
rect -2966 633454 -2346 668898
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 -2346 633454
rect -2966 633134 -2346 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 -2346 633134
rect -2966 597454 -2346 632898
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 -2346 597454
rect -2966 597134 -2346 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 -2346 597134
rect -2966 561454 -2346 596898
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 -2346 561454
rect -2966 561134 -2346 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 -2346 561134
rect -2966 525454 -2346 560898
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 -2346 525454
rect -2966 525134 -2346 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 -2346 525134
rect -2966 489454 -2346 524898
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 -2346 489454
rect -2966 489134 -2346 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 -2346 489134
rect -2966 453454 -2346 488898
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 -2346 453454
rect -2966 453134 -2346 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 -2346 453134
rect -2966 417454 -2346 452898
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 -2346 417454
rect -2966 417134 -2346 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 -2346 417134
rect -2966 381454 -2346 416898
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 -2346 381454
rect -2966 381134 -2346 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 -2346 381134
rect -2966 345454 -2346 380898
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 -2346 345454
rect -2966 345134 -2346 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 -2346 345134
rect -2966 309454 -2346 344898
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 -2346 309454
rect -2966 309134 -2346 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 -2346 309134
rect -2966 273454 -2346 308898
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 -2346 273454
rect -2966 273134 -2346 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 -2346 273134
rect -2966 237454 -2346 272898
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 -2346 237454
rect -2966 237134 -2346 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 -2346 237134
rect -2966 201454 -2346 236898
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 -2346 201454
rect -2966 201134 -2346 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 -2346 201134
rect -2966 165454 -2346 200898
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 -2346 165454
rect -2966 165134 -2346 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 -2346 165134
rect -2966 129454 -2346 164898
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 -2346 129454
rect -2966 129134 -2346 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 -2346 129134
rect -2966 93454 -2346 128898
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 -2346 93454
rect -2966 93134 -2346 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 -2346 93134
rect -2966 57454 -2346 92898
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 -2346 57454
rect -2966 57134 -2346 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 -2346 57134
rect -2966 21454 -2346 56898
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 -2346 21454
rect -2966 21134 -2346 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 -2346 21134
rect -2966 -1306 -2346 20898
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 705830
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 1794 -1894 2414 -902
rect 5514 691174 6134 706202
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 5514 619174 6134 654618
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 5514 259174 6134 294618
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 5514 223174 6134 258618
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 5514 187174 6134 222618
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 5514 151174 6134 186618
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 5514 115174 6134 150618
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 5514 79174 6134 114618
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 5514 43174 6134 78618
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 5514 7174 6134 42618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect 5514 -2266 6134 6618
rect 5514 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 6134 -2266
rect 5514 -2586 6134 -2502
rect 5514 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 6134 -2586
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect 5514 -3814 6134 -2822
rect 9234 694894 9854 708122
rect 9234 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 9854 694894
rect 9234 694574 9854 694658
rect 9234 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 9854 694574
rect 9234 658894 9854 694338
rect 9234 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 9854 658894
rect 9234 658574 9854 658658
rect 9234 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 9854 658574
rect 9234 622894 9854 658338
rect 9234 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 9854 622894
rect 9234 622574 9854 622658
rect 9234 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 9854 622574
rect 9234 586894 9854 622338
rect 9234 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 9854 586894
rect 9234 586574 9854 586658
rect 9234 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 9854 586574
rect 9234 550894 9854 586338
rect 9234 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 9854 550894
rect 9234 550574 9854 550658
rect 9234 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 9854 550574
rect 9234 514894 9854 550338
rect 9234 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 9854 514894
rect 9234 514574 9854 514658
rect 9234 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 9854 514574
rect 9234 478894 9854 514338
rect 9234 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 9854 478894
rect 9234 478574 9854 478658
rect 9234 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 9854 478574
rect 9234 442894 9854 478338
rect 9234 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 9854 442894
rect 9234 442574 9854 442658
rect 9234 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 9854 442574
rect 9234 406894 9854 442338
rect 9234 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 9854 406894
rect 9234 406574 9854 406658
rect 9234 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 9854 406574
rect 9234 370894 9854 406338
rect 9234 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 9854 370894
rect 9234 370574 9854 370658
rect 9234 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 9854 370574
rect 9234 334894 9854 370338
rect 9234 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 9854 334894
rect 9234 334574 9854 334658
rect 9234 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 9854 334574
rect 9234 298894 9854 334338
rect 9234 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 9854 298894
rect 9234 298574 9854 298658
rect 9234 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 9854 298574
rect 9234 262894 9854 298338
rect 9234 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 9854 262894
rect 9234 262574 9854 262658
rect 9234 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 9854 262574
rect 9234 226894 9854 262338
rect 9234 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 9854 226894
rect 9234 226574 9854 226658
rect 9234 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 9854 226574
rect 9234 190894 9854 226338
rect 9234 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 9854 190894
rect 9234 190574 9854 190658
rect 9234 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 9854 190574
rect 9234 154894 9854 190338
rect 9234 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 9854 154894
rect 9234 154574 9854 154658
rect 9234 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 9854 154574
rect 9234 118894 9854 154338
rect 9234 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 9854 118894
rect 9234 118574 9854 118658
rect 9234 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 9854 118574
rect 9234 82894 9854 118338
rect 9234 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 9854 82894
rect 9234 82574 9854 82658
rect 9234 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 9854 82574
rect 9234 46894 9854 82338
rect 9234 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 9854 46894
rect 9234 46574 9854 46658
rect 9234 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 9854 46574
rect 9234 10894 9854 46338
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect 9234 -4186 9854 10338
rect 9234 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 9854 -4186
rect 9234 -4506 9854 -4422
rect 9234 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 9854 -4506
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect 9234 -5734 9854 -4742
rect 12954 698614 13574 710042
rect 30954 711558 31574 711590
rect 30954 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 31574 711558
rect 30954 711238 31574 711322
rect 30954 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 31574 711238
rect 27234 709638 27854 709670
rect 27234 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 27854 709638
rect 27234 709318 27854 709402
rect 27234 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 27854 709318
rect 23514 707718 24134 707750
rect 23514 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 24134 707718
rect 23514 707398 24134 707482
rect 23514 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 24134 707398
rect 12954 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 13574 698614
rect 12954 698294 13574 698378
rect 12954 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 13574 698294
rect 12954 662614 13574 698058
rect 12954 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 13574 662614
rect 12954 662294 13574 662378
rect 12954 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 13574 662294
rect 12954 626614 13574 662058
rect 12954 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 13574 626614
rect 12954 626294 13574 626378
rect 12954 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 13574 626294
rect 12954 590614 13574 626058
rect 12954 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 13574 590614
rect 12954 590294 13574 590378
rect 12954 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 13574 590294
rect 12954 554614 13574 590058
rect 12954 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 13574 554614
rect 12954 554294 13574 554378
rect 12954 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 13574 554294
rect 12954 518614 13574 554058
rect 12954 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 13574 518614
rect 12954 518294 13574 518378
rect 12954 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 13574 518294
rect 12954 482614 13574 518058
rect 12954 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 13574 482614
rect 12954 482294 13574 482378
rect 12954 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 13574 482294
rect 12954 446614 13574 482058
rect 12954 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 13574 446614
rect 12954 446294 13574 446378
rect 12954 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 13574 446294
rect 12954 410614 13574 446058
rect 12954 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 13574 410614
rect 12954 410294 13574 410378
rect 12954 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 13574 410294
rect 12954 374614 13574 410058
rect 12954 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 13574 374614
rect 12954 374294 13574 374378
rect 12954 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 13574 374294
rect 12954 338614 13574 374058
rect 12954 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 13574 338614
rect 12954 338294 13574 338378
rect 12954 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 13574 338294
rect 12954 302614 13574 338058
rect 12954 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 13574 302614
rect 12954 302294 13574 302378
rect 12954 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 13574 302294
rect 12954 266614 13574 302058
rect 12954 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 13574 266614
rect 12954 266294 13574 266378
rect 12954 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 13574 266294
rect 12954 230614 13574 266058
rect 12954 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 13574 230614
rect 12954 230294 13574 230378
rect 12954 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 13574 230294
rect 12954 194614 13574 230058
rect 12954 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 13574 194614
rect 12954 194294 13574 194378
rect 12954 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 13574 194294
rect 12954 158614 13574 194058
rect 12954 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 13574 158614
rect 12954 158294 13574 158378
rect 12954 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 13574 158294
rect 12954 122614 13574 158058
rect 12954 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 13574 122614
rect 12954 122294 13574 122378
rect 12954 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 13574 122294
rect 12954 86614 13574 122058
rect 12954 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 13574 86614
rect 12954 86294 13574 86378
rect 12954 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 13574 86294
rect 12954 50614 13574 86058
rect 12954 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 13574 50614
rect 12954 50294 13574 50378
rect 12954 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 13574 50294
rect 12954 14614 13574 50058
rect 12954 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 13574 14614
rect 12954 14294 13574 14378
rect 12954 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 13574 14294
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect 12954 -6106 13574 14058
rect 19794 705798 20414 705830
rect 19794 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 20414 705798
rect 19794 705478 20414 705562
rect 19794 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 20414 705478
rect 19794 669454 20414 705242
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -1306 20414 20898
rect 19794 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 20414 -1306
rect 19794 -1626 20414 -1542
rect 19794 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 20414 -1626
rect 19794 -1894 20414 -1862
rect 23514 673174 24134 707162
rect 23514 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 24134 673174
rect 23514 672854 24134 672938
rect 23514 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 24134 672854
rect 23514 637174 24134 672618
rect 23514 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 24134 637174
rect 23514 636854 24134 636938
rect 23514 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 24134 636854
rect 23514 601174 24134 636618
rect 23514 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 24134 601174
rect 23514 600854 24134 600938
rect 23514 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 24134 600854
rect 23514 565174 24134 600618
rect 23514 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 24134 565174
rect 23514 564854 24134 564938
rect 23514 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 24134 564854
rect 23514 529174 24134 564618
rect 23514 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 24134 529174
rect 23514 528854 24134 528938
rect 23514 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 24134 528854
rect 23514 493174 24134 528618
rect 23514 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 24134 493174
rect 23514 492854 24134 492938
rect 23514 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 24134 492854
rect 23514 457174 24134 492618
rect 23514 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 24134 457174
rect 23514 456854 24134 456938
rect 23514 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 24134 456854
rect 23514 421174 24134 456618
rect 23514 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 24134 421174
rect 23514 420854 24134 420938
rect 23514 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 24134 420854
rect 23514 385174 24134 420618
rect 23514 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 24134 385174
rect 23514 384854 24134 384938
rect 23514 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 24134 384854
rect 23514 349174 24134 384618
rect 23514 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 24134 349174
rect 23514 348854 24134 348938
rect 23514 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 24134 348854
rect 23514 313174 24134 348618
rect 23514 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 24134 313174
rect 23514 312854 24134 312938
rect 23514 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 24134 312854
rect 23514 277174 24134 312618
rect 23514 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 24134 277174
rect 23514 276854 24134 276938
rect 23514 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 24134 276854
rect 23514 241174 24134 276618
rect 23514 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 24134 241174
rect 23514 240854 24134 240938
rect 23514 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 24134 240854
rect 23514 205174 24134 240618
rect 23514 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 24134 205174
rect 23514 204854 24134 204938
rect 23514 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 24134 204854
rect 23514 169174 24134 204618
rect 23514 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 24134 169174
rect 23514 168854 24134 168938
rect 23514 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 24134 168854
rect 23514 133174 24134 168618
rect 23514 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 24134 133174
rect 23514 132854 24134 132938
rect 23514 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 24134 132854
rect 23514 97174 24134 132618
rect 23514 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 24134 97174
rect 23514 96854 24134 96938
rect 23514 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 24134 96854
rect 23514 61174 24134 96618
rect 23514 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 24134 61174
rect 23514 60854 24134 60938
rect 23514 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 24134 60854
rect 23514 25174 24134 60618
rect 23514 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 24134 25174
rect 23514 24854 24134 24938
rect 23514 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 24134 24854
rect 23514 -3226 24134 24618
rect 23514 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 24134 -3226
rect 23514 -3546 24134 -3462
rect 23514 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 24134 -3546
rect 23514 -3814 24134 -3782
rect 27234 676894 27854 709082
rect 27234 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 27854 676894
rect 27234 676574 27854 676658
rect 27234 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 27854 676574
rect 27234 640894 27854 676338
rect 27234 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 27854 640894
rect 27234 640574 27854 640658
rect 27234 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 27854 640574
rect 27234 604894 27854 640338
rect 27234 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 27854 604894
rect 27234 604574 27854 604658
rect 27234 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 27854 604574
rect 27234 568894 27854 604338
rect 27234 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 27854 568894
rect 27234 568574 27854 568658
rect 27234 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 27854 568574
rect 27234 532894 27854 568338
rect 27234 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 27854 532894
rect 27234 532574 27854 532658
rect 27234 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 27854 532574
rect 27234 496894 27854 532338
rect 27234 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 27854 496894
rect 27234 496574 27854 496658
rect 27234 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 27854 496574
rect 27234 460894 27854 496338
rect 27234 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 27854 460894
rect 27234 460574 27854 460658
rect 27234 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 27854 460574
rect 27234 424894 27854 460338
rect 27234 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 27854 424894
rect 27234 424574 27854 424658
rect 27234 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 27854 424574
rect 27234 388894 27854 424338
rect 27234 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 27854 388894
rect 27234 388574 27854 388658
rect 27234 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 27854 388574
rect 27234 352894 27854 388338
rect 27234 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 27854 352894
rect 27234 352574 27854 352658
rect 27234 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 27854 352574
rect 27234 316894 27854 352338
rect 27234 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 27854 316894
rect 27234 316574 27854 316658
rect 27234 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 27854 316574
rect 27234 280894 27854 316338
rect 27234 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 27854 280894
rect 27234 280574 27854 280658
rect 27234 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 27854 280574
rect 27234 244894 27854 280338
rect 27234 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 27854 244894
rect 27234 244574 27854 244658
rect 27234 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 27854 244574
rect 27234 208894 27854 244338
rect 27234 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 27854 208894
rect 27234 208574 27854 208658
rect 27234 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 27854 208574
rect 27234 172894 27854 208338
rect 27234 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 27854 172894
rect 27234 172574 27854 172658
rect 27234 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 27854 172574
rect 27234 136894 27854 172338
rect 27234 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 27854 136894
rect 27234 136574 27854 136658
rect 27234 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 27854 136574
rect 27234 100894 27854 136338
rect 27234 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 27854 100894
rect 27234 100574 27854 100658
rect 27234 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 27854 100574
rect 27234 64894 27854 100338
rect 27234 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 27854 64894
rect 27234 64574 27854 64658
rect 27234 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 27854 64574
rect 27234 28894 27854 64338
rect 27234 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 27854 28894
rect 27234 28574 27854 28658
rect 27234 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 27854 28574
rect 27234 -5146 27854 28338
rect 27234 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 27854 -5146
rect 27234 -5466 27854 -5382
rect 27234 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 27854 -5466
rect 27234 -5734 27854 -5702
rect 30954 680614 31574 711002
rect 48954 710598 49574 711590
rect 48954 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 49574 710598
rect 48954 710278 49574 710362
rect 48954 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 49574 710278
rect 45234 708678 45854 709670
rect 45234 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 45854 708678
rect 45234 708358 45854 708442
rect 45234 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 45854 708358
rect 41514 706758 42134 707750
rect 41514 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 42134 706758
rect 41514 706438 42134 706522
rect 41514 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 42134 706438
rect 30954 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 31574 680614
rect 30954 680294 31574 680378
rect 30954 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 31574 680294
rect 30954 644614 31574 680058
rect 30954 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 31574 644614
rect 30954 644294 31574 644378
rect 30954 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 31574 644294
rect 30954 608614 31574 644058
rect 30954 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 31574 608614
rect 30954 608294 31574 608378
rect 30954 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 31574 608294
rect 30954 572614 31574 608058
rect 30954 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 31574 572614
rect 30954 572294 31574 572378
rect 30954 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 31574 572294
rect 30954 536614 31574 572058
rect 30954 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 31574 536614
rect 30954 536294 31574 536378
rect 30954 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 31574 536294
rect 30954 500614 31574 536058
rect 30954 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 31574 500614
rect 30954 500294 31574 500378
rect 30954 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 31574 500294
rect 30954 464614 31574 500058
rect 30954 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 31574 464614
rect 30954 464294 31574 464378
rect 30954 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 31574 464294
rect 30954 428614 31574 464058
rect 30954 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 31574 428614
rect 30954 428294 31574 428378
rect 30954 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 31574 428294
rect 30954 392614 31574 428058
rect 30954 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 31574 392614
rect 30954 392294 31574 392378
rect 30954 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 31574 392294
rect 30954 356614 31574 392058
rect 30954 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 31574 356614
rect 30954 356294 31574 356378
rect 30954 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 31574 356294
rect 30954 320614 31574 356058
rect 30954 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 31574 320614
rect 30954 320294 31574 320378
rect 30954 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 31574 320294
rect 30954 284614 31574 320058
rect 30954 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 31574 284614
rect 30954 284294 31574 284378
rect 30954 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 31574 284294
rect 30954 248614 31574 284058
rect 30954 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 31574 248614
rect 30954 248294 31574 248378
rect 30954 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 31574 248294
rect 30954 212614 31574 248058
rect 30954 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 31574 212614
rect 30954 212294 31574 212378
rect 30954 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 31574 212294
rect 30954 176614 31574 212058
rect 30954 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 31574 176614
rect 30954 176294 31574 176378
rect 30954 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 31574 176294
rect 30954 140614 31574 176058
rect 30954 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 31574 140614
rect 30954 140294 31574 140378
rect 30954 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 31574 140294
rect 30954 104614 31574 140058
rect 30954 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 31574 104614
rect 30954 104294 31574 104378
rect 30954 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 31574 104294
rect 30954 68614 31574 104058
rect 30954 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 31574 68614
rect 30954 68294 31574 68378
rect 30954 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 31574 68294
rect 30954 32614 31574 68058
rect 30954 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 31574 32614
rect 30954 32294 31574 32378
rect 30954 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 31574 32294
rect 12954 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 13574 -6106
rect 12954 -6426 13574 -6342
rect 12954 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 13574 -6426
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 12954 -7654 13574 -6662
rect 30954 -7066 31574 32058
rect 37794 704838 38414 705830
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -1894 38414 -902
rect 41514 691174 42134 706202
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 41514 655174 42134 690618
rect 41514 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 42134 655174
rect 41514 654854 42134 654938
rect 41514 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 42134 654854
rect 41514 619174 42134 654618
rect 41514 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 42134 619174
rect 41514 618854 42134 618938
rect 41514 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 42134 618854
rect 41514 583174 42134 618618
rect 41514 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 42134 583174
rect 41514 582854 42134 582938
rect 41514 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 42134 582854
rect 41514 547174 42134 582618
rect 41514 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 42134 547174
rect 41514 546854 42134 546938
rect 41514 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 42134 546854
rect 41514 511174 42134 546618
rect 41514 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 42134 511174
rect 41514 510854 42134 510938
rect 41514 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 42134 510854
rect 41514 475174 42134 510618
rect 41514 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 42134 475174
rect 41514 474854 42134 474938
rect 41514 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 42134 474854
rect 41514 439174 42134 474618
rect 41514 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 42134 439174
rect 41514 438854 42134 438938
rect 41514 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 42134 438854
rect 41514 403174 42134 438618
rect 41514 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 42134 403174
rect 41514 402854 42134 402938
rect 41514 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 42134 402854
rect 41514 367174 42134 402618
rect 41514 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 42134 367174
rect 41514 366854 42134 366938
rect 41514 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 42134 366854
rect 41514 331174 42134 366618
rect 41514 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 42134 331174
rect 41514 330854 42134 330938
rect 41514 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 42134 330854
rect 41514 295174 42134 330618
rect 41514 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 42134 295174
rect 41514 294854 42134 294938
rect 41514 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 42134 294854
rect 41514 259174 42134 294618
rect 41514 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 42134 259174
rect 41514 258854 42134 258938
rect 41514 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 42134 258854
rect 41514 223174 42134 258618
rect 41514 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 42134 223174
rect 41514 222854 42134 222938
rect 41514 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 42134 222854
rect 41514 187174 42134 222618
rect 41514 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 42134 187174
rect 41514 186854 42134 186938
rect 41514 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 42134 186854
rect 41514 151174 42134 186618
rect 41514 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 42134 151174
rect 41514 150854 42134 150938
rect 41514 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 42134 150854
rect 41514 115174 42134 150618
rect 41514 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 42134 115174
rect 41514 114854 42134 114938
rect 41514 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 42134 114854
rect 41514 79174 42134 114618
rect 41514 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 42134 79174
rect 41514 78854 42134 78938
rect 41514 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 42134 78854
rect 41514 43174 42134 78618
rect 41514 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 42134 43174
rect 41514 42854 42134 42938
rect 41514 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 42134 42854
rect 41514 7174 42134 42618
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -2266 42134 6618
rect 41514 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 42134 -2266
rect 41514 -2586 42134 -2502
rect 41514 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 42134 -2586
rect 41514 -3814 42134 -2822
rect 45234 694894 45854 708122
rect 45234 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 45854 694894
rect 45234 694574 45854 694658
rect 45234 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 45854 694574
rect 45234 658894 45854 694338
rect 45234 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 45854 658894
rect 45234 658574 45854 658658
rect 45234 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 45854 658574
rect 45234 622894 45854 658338
rect 45234 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 45854 622894
rect 45234 622574 45854 622658
rect 45234 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 45854 622574
rect 45234 586894 45854 622338
rect 45234 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 45854 586894
rect 45234 586574 45854 586658
rect 45234 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 45854 586574
rect 45234 550894 45854 586338
rect 45234 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 45854 550894
rect 45234 550574 45854 550658
rect 45234 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 45854 550574
rect 45234 514894 45854 550338
rect 45234 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 45854 514894
rect 45234 514574 45854 514658
rect 45234 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 45854 514574
rect 45234 478894 45854 514338
rect 45234 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 45854 478894
rect 45234 478574 45854 478658
rect 45234 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 45854 478574
rect 45234 442894 45854 478338
rect 45234 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 45854 442894
rect 45234 442574 45854 442658
rect 45234 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 45854 442574
rect 45234 406894 45854 442338
rect 45234 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 45854 406894
rect 45234 406574 45854 406658
rect 45234 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 45854 406574
rect 45234 370894 45854 406338
rect 45234 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 45854 370894
rect 45234 370574 45854 370658
rect 45234 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 45854 370574
rect 45234 334894 45854 370338
rect 45234 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 45854 334894
rect 45234 334574 45854 334658
rect 45234 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 45854 334574
rect 45234 298894 45854 334338
rect 45234 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 45854 298894
rect 45234 298574 45854 298658
rect 45234 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 45854 298574
rect 45234 262894 45854 298338
rect 45234 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 45854 262894
rect 45234 262574 45854 262658
rect 45234 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 45854 262574
rect 45234 226894 45854 262338
rect 45234 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 45854 226894
rect 45234 226574 45854 226658
rect 45234 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 45854 226574
rect 45234 190894 45854 226338
rect 45234 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 45854 190894
rect 45234 190574 45854 190658
rect 45234 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 45854 190574
rect 45234 154894 45854 190338
rect 45234 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 45854 154894
rect 45234 154574 45854 154658
rect 45234 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 45854 154574
rect 45234 118894 45854 154338
rect 45234 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 45854 118894
rect 45234 118574 45854 118658
rect 45234 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 45854 118574
rect 45234 82894 45854 118338
rect 45234 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 45854 82894
rect 45234 82574 45854 82658
rect 45234 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 45854 82574
rect 45234 46894 45854 82338
rect 45234 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 45854 46894
rect 45234 46574 45854 46658
rect 45234 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 45854 46574
rect 45234 10894 45854 46338
rect 45234 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 45854 10894
rect 45234 10574 45854 10658
rect 45234 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 45854 10574
rect 45234 -4186 45854 10338
rect 45234 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 45854 -4186
rect 45234 -4506 45854 -4422
rect 45234 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 45854 -4506
rect 45234 -5734 45854 -4742
rect 48954 698614 49574 710042
rect 66954 711558 67574 711590
rect 66954 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 67574 711558
rect 66954 711238 67574 711322
rect 66954 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 67574 711238
rect 63234 709638 63854 709670
rect 63234 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 63854 709638
rect 63234 709318 63854 709402
rect 63234 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 63854 709318
rect 59514 707718 60134 707750
rect 59514 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 60134 707718
rect 59514 707398 60134 707482
rect 59514 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 60134 707398
rect 48954 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 49574 698614
rect 48954 698294 49574 698378
rect 48954 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 49574 698294
rect 48954 662614 49574 698058
rect 48954 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 49574 662614
rect 48954 662294 49574 662378
rect 48954 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 49574 662294
rect 48954 626614 49574 662058
rect 48954 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 49574 626614
rect 48954 626294 49574 626378
rect 48954 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 49574 626294
rect 48954 590614 49574 626058
rect 48954 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 49574 590614
rect 48954 590294 49574 590378
rect 48954 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 49574 590294
rect 48954 554614 49574 590058
rect 48954 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 49574 554614
rect 48954 554294 49574 554378
rect 48954 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 49574 554294
rect 48954 518614 49574 554058
rect 48954 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 49574 518614
rect 48954 518294 49574 518378
rect 48954 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 49574 518294
rect 48954 482614 49574 518058
rect 48954 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 49574 482614
rect 48954 482294 49574 482378
rect 48954 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 49574 482294
rect 48954 446614 49574 482058
rect 48954 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 49574 446614
rect 48954 446294 49574 446378
rect 48954 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 49574 446294
rect 48954 410614 49574 446058
rect 48954 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 49574 410614
rect 48954 410294 49574 410378
rect 48954 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 49574 410294
rect 48954 374614 49574 410058
rect 48954 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 49574 374614
rect 48954 374294 49574 374378
rect 48954 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 49574 374294
rect 48954 338614 49574 374058
rect 48954 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 49574 338614
rect 48954 338294 49574 338378
rect 48954 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 49574 338294
rect 48954 302614 49574 338058
rect 48954 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 49574 302614
rect 48954 302294 49574 302378
rect 48954 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 49574 302294
rect 48954 266614 49574 302058
rect 48954 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 49574 266614
rect 48954 266294 49574 266378
rect 48954 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 49574 266294
rect 48954 230614 49574 266058
rect 48954 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 49574 230614
rect 48954 230294 49574 230378
rect 48954 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 49574 230294
rect 48954 194614 49574 230058
rect 48954 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 49574 194614
rect 48954 194294 49574 194378
rect 48954 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 49574 194294
rect 48954 158614 49574 194058
rect 48954 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 49574 158614
rect 48954 158294 49574 158378
rect 48954 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 49574 158294
rect 48954 122614 49574 158058
rect 48954 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 49574 122614
rect 48954 122294 49574 122378
rect 48954 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 49574 122294
rect 48954 86614 49574 122058
rect 48954 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 49574 86614
rect 48954 86294 49574 86378
rect 48954 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 49574 86294
rect 48954 50614 49574 86058
rect 48954 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 49574 50614
rect 48954 50294 49574 50378
rect 48954 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 49574 50294
rect 48954 14614 49574 50058
rect 48954 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 49574 14614
rect 48954 14294 49574 14378
rect 48954 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 49574 14294
rect 30954 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 31574 -7066
rect 30954 -7386 31574 -7302
rect 30954 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 31574 -7386
rect 30954 -7654 31574 -7622
rect 48954 -6106 49574 14058
rect 55794 705798 56414 705830
rect 55794 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 56414 705798
rect 55794 705478 56414 705562
rect 55794 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 56414 705478
rect 55794 669454 56414 705242
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 273454 56414 308898
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 237454 56414 272898
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55794 201454 56414 236898
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -1306 56414 20898
rect 55794 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 56414 -1306
rect 55794 -1626 56414 -1542
rect 55794 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 56414 -1626
rect 55794 -1894 56414 -1862
rect 59514 673174 60134 707162
rect 59514 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 60134 673174
rect 59514 672854 60134 672938
rect 59514 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 60134 672854
rect 59514 637174 60134 672618
rect 59514 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 60134 637174
rect 59514 636854 60134 636938
rect 59514 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 60134 636854
rect 59514 601174 60134 636618
rect 59514 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 60134 601174
rect 59514 600854 60134 600938
rect 59514 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 60134 600854
rect 59514 565174 60134 600618
rect 59514 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 60134 565174
rect 59514 564854 60134 564938
rect 59514 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 60134 564854
rect 59514 529174 60134 564618
rect 59514 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 60134 529174
rect 59514 528854 60134 528938
rect 59514 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 60134 528854
rect 59514 493174 60134 528618
rect 59514 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 60134 493174
rect 59514 492854 60134 492938
rect 59514 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 60134 492854
rect 59514 457174 60134 492618
rect 59514 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 60134 457174
rect 59514 456854 60134 456938
rect 59514 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 60134 456854
rect 59514 421174 60134 456618
rect 59514 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 60134 421174
rect 59514 420854 60134 420938
rect 59514 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 60134 420854
rect 59514 385174 60134 420618
rect 59514 384938 59546 385174
rect 59782 384938 59866 385174
rect 60102 384938 60134 385174
rect 59514 384854 60134 384938
rect 59514 384618 59546 384854
rect 59782 384618 59866 384854
rect 60102 384618 60134 384854
rect 59514 349174 60134 384618
rect 59514 348938 59546 349174
rect 59782 348938 59866 349174
rect 60102 348938 60134 349174
rect 59514 348854 60134 348938
rect 59514 348618 59546 348854
rect 59782 348618 59866 348854
rect 60102 348618 60134 348854
rect 59514 313174 60134 348618
rect 59514 312938 59546 313174
rect 59782 312938 59866 313174
rect 60102 312938 60134 313174
rect 59514 312854 60134 312938
rect 59514 312618 59546 312854
rect 59782 312618 59866 312854
rect 60102 312618 60134 312854
rect 59514 277174 60134 312618
rect 59514 276938 59546 277174
rect 59782 276938 59866 277174
rect 60102 276938 60134 277174
rect 59514 276854 60134 276938
rect 59514 276618 59546 276854
rect 59782 276618 59866 276854
rect 60102 276618 60134 276854
rect 59514 241174 60134 276618
rect 59514 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 60134 241174
rect 59514 240854 60134 240938
rect 59514 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 60134 240854
rect 59514 205174 60134 240618
rect 59514 204938 59546 205174
rect 59782 204938 59866 205174
rect 60102 204938 60134 205174
rect 59514 204854 60134 204938
rect 59514 204618 59546 204854
rect 59782 204618 59866 204854
rect 60102 204618 60134 204854
rect 59514 169174 60134 204618
rect 59514 168938 59546 169174
rect 59782 168938 59866 169174
rect 60102 168938 60134 169174
rect 59514 168854 60134 168938
rect 59514 168618 59546 168854
rect 59782 168618 59866 168854
rect 60102 168618 60134 168854
rect 59514 133174 60134 168618
rect 59514 132938 59546 133174
rect 59782 132938 59866 133174
rect 60102 132938 60134 133174
rect 59514 132854 60134 132938
rect 59514 132618 59546 132854
rect 59782 132618 59866 132854
rect 60102 132618 60134 132854
rect 59514 97174 60134 132618
rect 59514 96938 59546 97174
rect 59782 96938 59866 97174
rect 60102 96938 60134 97174
rect 59514 96854 60134 96938
rect 59514 96618 59546 96854
rect 59782 96618 59866 96854
rect 60102 96618 60134 96854
rect 59514 61174 60134 96618
rect 59514 60938 59546 61174
rect 59782 60938 59866 61174
rect 60102 60938 60134 61174
rect 59514 60854 60134 60938
rect 59514 60618 59546 60854
rect 59782 60618 59866 60854
rect 60102 60618 60134 60854
rect 59514 25174 60134 60618
rect 59514 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 60134 25174
rect 59514 24854 60134 24938
rect 59514 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 60134 24854
rect 59514 -3226 60134 24618
rect 59514 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 60134 -3226
rect 59514 -3546 60134 -3462
rect 59514 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 60134 -3546
rect 59514 -3814 60134 -3782
rect 63234 676894 63854 709082
rect 63234 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 63854 676894
rect 63234 676574 63854 676658
rect 63234 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 63854 676574
rect 63234 640894 63854 676338
rect 63234 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 63854 640894
rect 63234 640574 63854 640658
rect 63234 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 63854 640574
rect 63234 604894 63854 640338
rect 63234 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 63854 604894
rect 63234 604574 63854 604658
rect 63234 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 63854 604574
rect 63234 568894 63854 604338
rect 63234 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 63854 568894
rect 63234 568574 63854 568658
rect 63234 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 63854 568574
rect 63234 532894 63854 568338
rect 63234 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 63854 532894
rect 63234 532574 63854 532658
rect 63234 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 63854 532574
rect 63234 496894 63854 532338
rect 63234 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 63854 496894
rect 63234 496574 63854 496658
rect 63234 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 63854 496574
rect 63234 460894 63854 496338
rect 63234 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 63854 460894
rect 63234 460574 63854 460658
rect 63234 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 63854 460574
rect 63234 424894 63854 460338
rect 63234 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 63854 424894
rect 63234 424574 63854 424658
rect 63234 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 63854 424574
rect 63234 388894 63854 424338
rect 63234 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 63854 388894
rect 63234 388574 63854 388658
rect 63234 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 63854 388574
rect 63234 352894 63854 388338
rect 63234 352658 63266 352894
rect 63502 352658 63586 352894
rect 63822 352658 63854 352894
rect 63234 352574 63854 352658
rect 63234 352338 63266 352574
rect 63502 352338 63586 352574
rect 63822 352338 63854 352574
rect 63234 316894 63854 352338
rect 63234 316658 63266 316894
rect 63502 316658 63586 316894
rect 63822 316658 63854 316894
rect 63234 316574 63854 316658
rect 63234 316338 63266 316574
rect 63502 316338 63586 316574
rect 63822 316338 63854 316574
rect 63234 280894 63854 316338
rect 63234 280658 63266 280894
rect 63502 280658 63586 280894
rect 63822 280658 63854 280894
rect 63234 280574 63854 280658
rect 63234 280338 63266 280574
rect 63502 280338 63586 280574
rect 63822 280338 63854 280574
rect 63234 244894 63854 280338
rect 63234 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 63854 244894
rect 63234 244574 63854 244658
rect 63234 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 63854 244574
rect 63234 208894 63854 244338
rect 63234 208658 63266 208894
rect 63502 208658 63586 208894
rect 63822 208658 63854 208894
rect 63234 208574 63854 208658
rect 63234 208338 63266 208574
rect 63502 208338 63586 208574
rect 63822 208338 63854 208574
rect 63234 172894 63854 208338
rect 63234 172658 63266 172894
rect 63502 172658 63586 172894
rect 63822 172658 63854 172894
rect 63234 172574 63854 172658
rect 63234 172338 63266 172574
rect 63502 172338 63586 172574
rect 63822 172338 63854 172574
rect 63234 136894 63854 172338
rect 63234 136658 63266 136894
rect 63502 136658 63586 136894
rect 63822 136658 63854 136894
rect 63234 136574 63854 136658
rect 63234 136338 63266 136574
rect 63502 136338 63586 136574
rect 63822 136338 63854 136574
rect 63234 100894 63854 136338
rect 63234 100658 63266 100894
rect 63502 100658 63586 100894
rect 63822 100658 63854 100894
rect 63234 100574 63854 100658
rect 63234 100338 63266 100574
rect 63502 100338 63586 100574
rect 63822 100338 63854 100574
rect 63234 64894 63854 100338
rect 63234 64658 63266 64894
rect 63502 64658 63586 64894
rect 63822 64658 63854 64894
rect 63234 64574 63854 64658
rect 63234 64338 63266 64574
rect 63502 64338 63586 64574
rect 63822 64338 63854 64574
rect 63234 28894 63854 64338
rect 63234 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 63854 28894
rect 63234 28574 63854 28658
rect 63234 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 63854 28574
rect 63234 -5146 63854 28338
rect 63234 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 63854 -5146
rect 63234 -5466 63854 -5382
rect 63234 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 63854 -5466
rect 63234 -5734 63854 -5702
rect 66954 680614 67574 711002
rect 84954 710598 85574 711590
rect 84954 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 85574 710598
rect 84954 710278 85574 710362
rect 84954 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 85574 710278
rect 81234 708678 81854 709670
rect 81234 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 81854 708678
rect 81234 708358 81854 708442
rect 81234 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 81854 708358
rect 77514 706758 78134 707750
rect 77514 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 78134 706758
rect 77514 706438 78134 706522
rect 77514 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 78134 706438
rect 66954 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 67574 680614
rect 66954 680294 67574 680378
rect 66954 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 67574 680294
rect 66954 644614 67574 680058
rect 66954 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 67574 644614
rect 66954 644294 67574 644378
rect 66954 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 67574 644294
rect 66954 608614 67574 644058
rect 66954 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 67574 608614
rect 66954 608294 67574 608378
rect 66954 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 67574 608294
rect 66954 572614 67574 608058
rect 66954 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 67574 572614
rect 66954 572294 67574 572378
rect 66954 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 67574 572294
rect 66954 536614 67574 572058
rect 66954 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 67574 536614
rect 66954 536294 67574 536378
rect 66954 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 67574 536294
rect 66954 500614 67574 536058
rect 66954 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 67574 500614
rect 66954 500294 67574 500378
rect 66954 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 67574 500294
rect 66954 464614 67574 500058
rect 66954 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 67574 464614
rect 66954 464294 67574 464378
rect 66954 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 67574 464294
rect 66954 428614 67574 464058
rect 66954 428378 66986 428614
rect 67222 428378 67306 428614
rect 67542 428378 67574 428614
rect 66954 428294 67574 428378
rect 66954 428058 66986 428294
rect 67222 428058 67306 428294
rect 67542 428058 67574 428294
rect 66954 392614 67574 428058
rect 66954 392378 66986 392614
rect 67222 392378 67306 392614
rect 67542 392378 67574 392614
rect 66954 392294 67574 392378
rect 66954 392058 66986 392294
rect 67222 392058 67306 392294
rect 67542 392058 67574 392294
rect 66954 356614 67574 392058
rect 66954 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 67574 356614
rect 66954 356294 67574 356378
rect 66954 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 67574 356294
rect 66954 320614 67574 356058
rect 66954 320378 66986 320614
rect 67222 320378 67306 320614
rect 67542 320378 67574 320614
rect 66954 320294 67574 320378
rect 66954 320058 66986 320294
rect 67222 320058 67306 320294
rect 67542 320058 67574 320294
rect 66954 284614 67574 320058
rect 66954 284378 66986 284614
rect 67222 284378 67306 284614
rect 67542 284378 67574 284614
rect 66954 284294 67574 284378
rect 66954 284058 66986 284294
rect 67222 284058 67306 284294
rect 67542 284058 67574 284294
rect 66954 248614 67574 284058
rect 66954 248378 66986 248614
rect 67222 248378 67306 248614
rect 67542 248378 67574 248614
rect 66954 248294 67574 248378
rect 66954 248058 66986 248294
rect 67222 248058 67306 248294
rect 67542 248058 67574 248294
rect 66954 212614 67574 248058
rect 66954 212378 66986 212614
rect 67222 212378 67306 212614
rect 67542 212378 67574 212614
rect 66954 212294 67574 212378
rect 66954 212058 66986 212294
rect 67222 212058 67306 212294
rect 67542 212058 67574 212294
rect 66954 176614 67574 212058
rect 66954 176378 66986 176614
rect 67222 176378 67306 176614
rect 67542 176378 67574 176614
rect 66954 176294 67574 176378
rect 66954 176058 66986 176294
rect 67222 176058 67306 176294
rect 67542 176058 67574 176294
rect 66954 140614 67574 176058
rect 66954 140378 66986 140614
rect 67222 140378 67306 140614
rect 67542 140378 67574 140614
rect 66954 140294 67574 140378
rect 66954 140058 66986 140294
rect 67222 140058 67306 140294
rect 67542 140058 67574 140294
rect 66954 104614 67574 140058
rect 66954 104378 66986 104614
rect 67222 104378 67306 104614
rect 67542 104378 67574 104614
rect 66954 104294 67574 104378
rect 66954 104058 66986 104294
rect 67222 104058 67306 104294
rect 67542 104058 67574 104294
rect 66954 68614 67574 104058
rect 66954 68378 66986 68614
rect 67222 68378 67306 68614
rect 67542 68378 67574 68614
rect 66954 68294 67574 68378
rect 66954 68058 66986 68294
rect 67222 68058 67306 68294
rect 67542 68058 67574 68294
rect 66954 32614 67574 68058
rect 66954 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 67574 32614
rect 66954 32294 67574 32378
rect 66954 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 67574 32294
rect 48954 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 49574 -6106
rect 48954 -6426 49574 -6342
rect 48954 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 49574 -6426
rect 48954 -7654 49574 -6662
rect 66954 -7066 67574 32058
rect 73794 704838 74414 705830
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 579454 74414 614898
rect 73794 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 74414 579454
rect 73794 579134 74414 579218
rect 73794 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 74414 579134
rect 73794 543454 74414 578898
rect 73794 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 74414 543454
rect 73794 543134 74414 543218
rect 73794 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 74414 543134
rect 73794 507454 74414 542898
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 471454 74414 506898
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73794 435454 74414 470898
rect 73794 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 74414 435454
rect 73794 435134 74414 435218
rect 73794 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 74414 435134
rect 73794 399454 74414 434898
rect 73794 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 74414 399454
rect 73794 399134 74414 399218
rect 73794 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 74414 399134
rect 73794 363454 74414 398898
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 73794 327454 74414 362898
rect 73794 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 74414 327454
rect 73794 327134 74414 327218
rect 73794 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 74414 327134
rect 73794 291454 74414 326898
rect 73794 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 74414 291454
rect 73794 291134 74414 291218
rect 73794 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 74414 291134
rect 73794 255454 74414 290898
rect 73794 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 74414 255454
rect 73794 255134 74414 255218
rect 73794 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 74414 255134
rect 73794 219454 74414 254898
rect 73794 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 74414 219454
rect 73794 219134 74414 219218
rect 73794 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 74414 219134
rect 73794 183454 74414 218898
rect 73794 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 74414 183454
rect 73794 183134 74414 183218
rect 73794 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 74414 183134
rect 73794 147454 74414 182898
rect 73794 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 74414 147454
rect 73794 147134 74414 147218
rect 73794 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 74414 147134
rect 73794 111454 74414 146898
rect 73794 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 74414 111454
rect 73794 111134 74414 111218
rect 73794 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 74414 111134
rect 73794 75454 74414 110898
rect 73794 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 74414 75454
rect 73794 75134 74414 75218
rect 73794 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 74414 75134
rect 73794 39454 74414 74898
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -1894 74414 -902
rect 77514 691174 78134 706202
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 655174 78134 690618
rect 77514 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 78134 655174
rect 77514 654854 78134 654938
rect 77514 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 78134 654854
rect 77514 619174 78134 654618
rect 77514 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 78134 619174
rect 77514 618854 78134 618938
rect 77514 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 78134 618854
rect 77514 583174 78134 618618
rect 77514 582938 77546 583174
rect 77782 582938 77866 583174
rect 78102 582938 78134 583174
rect 77514 582854 78134 582938
rect 77514 582618 77546 582854
rect 77782 582618 77866 582854
rect 78102 582618 78134 582854
rect 77514 547174 78134 582618
rect 77514 546938 77546 547174
rect 77782 546938 77866 547174
rect 78102 546938 78134 547174
rect 77514 546854 78134 546938
rect 77514 546618 77546 546854
rect 77782 546618 77866 546854
rect 78102 546618 78134 546854
rect 77514 511174 78134 546618
rect 77514 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 78134 511174
rect 77514 510854 78134 510938
rect 77514 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 78134 510854
rect 77514 475174 78134 510618
rect 77514 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 78134 475174
rect 77514 474854 78134 474938
rect 77514 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 78134 474854
rect 77514 439174 78134 474618
rect 77514 438938 77546 439174
rect 77782 438938 77866 439174
rect 78102 438938 78134 439174
rect 77514 438854 78134 438938
rect 77514 438618 77546 438854
rect 77782 438618 77866 438854
rect 78102 438618 78134 438854
rect 77514 403174 78134 438618
rect 77514 402938 77546 403174
rect 77782 402938 77866 403174
rect 78102 402938 78134 403174
rect 77514 402854 78134 402938
rect 77514 402618 77546 402854
rect 77782 402618 77866 402854
rect 78102 402618 78134 402854
rect 77514 367174 78134 402618
rect 77514 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 78134 367174
rect 77514 366854 78134 366938
rect 77514 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 78134 366854
rect 77514 331174 78134 366618
rect 77514 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 78134 331174
rect 77514 330854 78134 330938
rect 77514 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 78134 330854
rect 77514 295174 78134 330618
rect 77514 294938 77546 295174
rect 77782 294938 77866 295174
rect 78102 294938 78134 295174
rect 77514 294854 78134 294938
rect 77514 294618 77546 294854
rect 77782 294618 77866 294854
rect 78102 294618 78134 294854
rect 77514 259174 78134 294618
rect 77514 258938 77546 259174
rect 77782 258938 77866 259174
rect 78102 258938 78134 259174
rect 77514 258854 78134 258938
rect 77514 258618 77546 258854
rect 77782 258618 77866 258854
rect 78102 258618 78134 258854
rect 77514 223174 78134 258618
rect 77514 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 78134 223174
rect 77514 222854 78134 222938
rect 77514 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 78134 222854
rect 77514 187174 78134 222618
rect 77514 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 78134 187174
rect 77514 186854 78134 186938
rect 77514 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 78134 186854
rect 77514 151174 78134 186618
rect 77514 150938 77546 151174
rect 77782 150938 77866 151174
rect 78102 150938 78134 151174
rect 77514 150854 78134 150938
rect 77514 150618 77546 150854
rect 77782 150618 77866 150854
rect 78102 150618 78134 150854
rect 77514 115174 78134 150618
rect 77514 114938 77546 115174
rect 77782 114938 77866 115174
rect 78102 114938 78134 115174
rect 77514 114854 78134 114938
rect 77514 114618 77546 114854
rect 77782 114618 77866 114854
rect 78102 114618 78134 114854
rect 77514 79174 78134 114618
rect 77514 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 78134 79174
rect 77514 78854 78134 78938
rect 77514 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 78134 78854
rect 77514 43174 78134 78618
rect 77514 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 78134 43174
rect 77514 42854 78134 42938
rect 77514 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 78134 42854
rect 77514 7174 78134 42618
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 77514 -2266 78134 6618
rect 77514 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 78134 -2266
rect 77514 -2586 78134 -2502
rect 77514 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 78134 -2586
rect 77514 -3814 78134 -2822
rect 81234 694894 81854 708122
rect 81234 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 81854 694894
rect 81234 694574 81854 694658
rect 81234 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 81854 694574
rect 81234 658894 81854 694338
rect 81234 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 81854 658894
rect 81234 658574 81854 658658
rect 81234 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 81854 658574
rect 81234 622894 81854 658338
rect 81234 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 81854 622894
rect 81234 622574 81854 622658
rect 81234 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 81854 622574
rect 81234 586894 81854 622338
rect 81234 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 81854 586894
rect 81234 586574 81854 586658
rect 81234 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 81854 586574
rect 81234 550894 81854 586338
rect 81234 550658 81266 550894
rect 81502 550658 81586 550894
rect 81822 550658 81854 550894
rect 81234 550574 81854 550658
rect 81234 550338 81266 550574
rect 81502 550338 81586 550574
rect 81822 550338 81854 550574
rect 81234 514894 81854 550338
rect 81234 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 81854 514894
rect 81234 514574 81854 514658
rect 81234 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 81854 514574
rect 81234 478894 81854 514338
rect 81234 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 81854 478894
rect 81234 478574 81854 478658
rect 81234 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 81854 478574
rect 81234 442894 81854 478338
rect 81234 442658 81266 442894
rect 81502 442658 81586 442894
rect 81822 442658 81854 442894
rect 81234 442574 81854 442658
rect 81234 442338 81266 442574
rect 81502 442338 81586 442574
rect 81822 442338 81854 442574
rect 81234 406894 81854 442338
rect 81234 406658 81266 406894
rect 81502 406658 81586 406894
rect 81822 406658 81854 406894
rect 81234 406574 81854 406658
rect 81234 406338 81266 406574
rect 81502 406338 81586 406574
rect 81822 406338 81854 406574
rect 81234 370894 81854 406338
rect 81234 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 81854 370894
rect 81234 370574 81854 370658
rect 81234 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 81854 370574
rect 81234 334894 81854 370338
rect 81234 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 81854 334894
rect 81234 334574 81854 334658
rect 81234 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 81854 334574
rect 81234 298894 81854 334338
rect 81234 298658 81266 298894
rect 81502 298658 81586 298894
rect 81822 298658 81854 298894
rect 81234 298574 81854 298658
rect 81234 298338 81266 298574
rect 81502 298338 81586 298574
rect 81822 298338 81854 298574
rect 81234 262894 81854 298338
rect 81234 262658 81266 262894
rect 81502 262658 81586 262894
rect 81822 262658 81854 262894
rect 81234 262574 81854 262658
rect 81234 262338 81266 262574
rect 81502 262338 81586 262574
rect 81822 262338 81854 262574
rect 81234 226894 81854 262338
rect 81234 226658 81266 226894
rect 81502 226658 81586 226894
rect 81822 226658 81854 226894
rect 81234 226574 81854 226658
rect 81234 226338 81266 226574
rect 81502 226338 81586 226574
rect 81822 226338 81854 226574
rect 81234 190894 81854 226338
rect 81234 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 81854 190894
rect 81234 190574 81854 190658
rect 81234 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 81854 190574
rect 81234 154894 81854 190338
rect 81234 154658 81266 154894
rect 81502 154658 81586 154894
rect 81822 154658 81854 154894
rect 81234 154574 81854 154658
rect 81234 154338 81266 154574
rect 81502 154338 81586 154574
rect 81822 154338 81854 154574
rect 81234 118894 81854 154338
rect 81234 118658 81266 118894
rect 81502 118658 81586 118894
rect 81822 118658 81854 118894
rect 81234 118574 81854 118658
rect 81234 118338 81266 118574
rect 81502 118338 81586 118574
rect 81822 118338 81854 118574
rect 81234 82894 81854 118338
rect 81234 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 81854 82894
rect 81234 82574 81854 82658
rect 81234 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 81854 82574
rect 81234 46894 81854 82338
rect 81234 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 81854 46894
rect 81234 46574 81854 46658
rect 81234 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 81854 46574
rect 81234 10894 81854 46338
rect 81234 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 81854 10894
rect 81234 10574 81854 10658
rect 81234 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 81854 10574
rect 81234 -4186 81854 10338
rect 81234 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 81854 -4186
rect 81234 -4506 81854 -4422
rect 81234 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 81854 -4506
rect 81234 -5734 81854 -4742
rect 84954 698614 85574 710042
rect 102954 711558 103574 711590
rect 102954 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 103574 711558
rect 102954 711238 103574 711322
rect 102954 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 103574 711238
rect 99234 709638 99854 709670
rect 99234 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 99854 709638
rect 99234 709318 99854 709402
rect 99234 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 99854 709318
rect 95514 707718 96134 707750
rect 95514 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 96134 707718
rect 95514 707398 96134 707482
rect 95514 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 96134 707398
rect 84954 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 85574 698614
rect 84954 698294 85574 698378
rect 84954 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 85574 698294
rect 84954 662614 85574 698058
rect 84954 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 85574 662614
rect 84954 662294 85574 662378
rect 84954 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 85574 662294
rect 84954 626614 85574 662058
rect 84954 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 85574 626614
rect 84954 626294 85574 626378
rect 84954 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 85574 626294
rect 84954 590614 85574 626058
rect 84954 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 85574 590614
rect 84954 590294 85574 590378
rect 84954 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 85574 590294
rect 84954 554614 85574 590058
rect 84954 554378 84986 554614
rect 85222 554378 85306 554614
rect 85542 554378 85574 554614
rect 84954 554294 85574 554378
rect 84954 554058 84986 554294
rect 85222 554058 85306 554294
rect 85542 554058 85574 554294
rect 84954 518614 85574 554058
rect 84954 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 85574 518614
rect 84954 518294 85574 518378
rect 84954 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 85574 518294
rect 84954 482614 85574 518058
rect 84954 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 85574 482614
rect 84954 482294 85574 482378
rect 84954 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 85574 482294
rect 84954 446614 85574 482058
rect 84954 446378 84986 446614
rect 85222 446378 85306 446614
rect 85542 446378 85574 446614
rect 84954 446294 85574 446378
rect 84954 446058 84986 446294
rect 85222 446058 85306 446294
rect 85542 446058 85574 446294
rect 84954 410614 85574 446058
rect 84954 410378 84986 410614
rect 85222 410378 85306 410614
rect 85542 410378 85574 410614
rect 84954 410294 85574 410378
rect 84954 410058 84986 410294
rect 85222 410058 85306 410294
rect 85542 410058 85574 410294
rect 84954 374614 85574 410058
rect 84954 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 85574 374614
rect 84954 374294 85574 374378
rect 84954 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 85574 374294
rect 84954 338614 85574 374058
rect 84954 338378 84986 338614
rect 85222 338378 85306 338614
rect 85542 338378 85574 338614
rect 84954 338294 85574 338378
rect 84954 338058 84986 338294
rect 85222 338058 85306 338294
rect 85542 338058 85574 338294
rect 84954 302614 85574 338058
rect 84954 302378 84986 302614
rect 85222 302378 85306 302614
rect 85542 302378 85574 302614
rect 84954 302294 85574 302378
rect 84954 302058 84986 302294
rect 85222 302058 85306 302294
rect 85542 302058 85574 302294
rect 84954 266614 85574 302058
rect 84954 266378 84986 266614
rect 85222 266378 85306 266614
rect 85542 266378 85574 266614
rect 84954 266294 85574 266378
rect 84954 266058 84986 266294
rect 85222 266058 85306 266294
rect 85542 266058 85574 266294
rect 84954 230614 85574 266058
rect 84954 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 85574 230614
rect 84954 230294 85574 230378
rect 84954 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 85574 230294
rect 84954 194614 85574 230058
rect 84954 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 85574 194614
rect 84954 194294 85574 194378
rect 84954 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 85574 194294
rect 84954 158614 85574 194058
rect 84954 158378 84986 158614
rect 85222 158378 85306 158614
rect 85542 158378 85574 158614
rect 84954 158294 85574 158378
rect 84954 158058 84986 158294
rect 85222 158058 85306 158294
rect 85542 158058 85574 158294
rect 84954 122614 85574 158058
rect 84954 122378 84986 122614
rect 85222 122378 85306 122614
rect 85542 122378 85574 122614
rect 84954 122294 85574 122378
rect 84954 122058 84986 122294
rect 85222 122058 85306 122294
rect 85542 122058 85574 122294
rect 84954 86614 85574 122058
rect 84954 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 85574 86614
rect 84954 86294 85574 86378
rect 84954 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 85574 86294
rect 84954 50614 85574 86058
rect 84954 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 85574 50614
rect 84954 50294 85574 50378
rect 84954 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 85574 50294
rect 84954 14614 85574 50058
rect 84954 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 85574 14614
rect 84954 14294 85574 14378
rect 84954 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 85574 14294
rect 66954 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 67574 -7066
rect 66954 -7386 67574 -7302
rect 66954 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 67574 -7386
rect 66954 -7654 67574 -7622
rect 84954 -6106 85574 14058
rect 91794 705798 92414 705830
rect 91794 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 92414 705798
rect 91794 705478 92414 705562
rect 91794 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 92414 705478
rect 91794 669454 92414 705242
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 91794 561454 92414 596898
rect 91794 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 92414 561454
rect 91794 561134 92414 561218
rect 91794 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 92414 561134
rect 91794 525454 92414 560898
rect 91794 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 92414 525454
rect 91794 525134 92414 525218
rect 91794 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 92414 525134
rect 91794 489454 92414 524898
rect 91794 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 92414 489454
rect 91794 489134 92414 489218
rect 91794 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 92414 489134
rect 91794 453454 92414 488898
rect 91794 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 92414 453454
rect 91794 453134 92414 453218
rect 91794 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 92414 453134
rect 91794 417454 92414 452898
rect 91794 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 92414 417454
rect 91794 417134 92414 417218
rect 91794 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 92414 417134
rect 91794 381454 92414 416898
rect 91794 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 92414 381454
rect 91794 381134 92414 381218
rect 91794 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 92414 381134
rect 91794 345454 92414 380898
rect 91794 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 92414 345454
rect 91794 345134 92414 345218
rect 91794 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 92414 345134
rect 91794 309454 92414 344898
rect 91794 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 92414 309454
rect 91794 309134 92414 309218
rect 91794 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 92414 309134
rect 91794 273454 92414 308898
rect 91794 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 92414 273454
rect 91794 273134 92414 273218
rect 91794 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 92414 273134
rect 91794 237454 92414 272898
rect 91794 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 92414 237454
rect 91794 237134 92414 237218
rect 91794 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 92414 237134
rect 91794 201454 92414 236898
rect 91794 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 92414 201454
rect 91794 201134 92414 201218
rect 91794 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 92414 201134
rect 91794 165454 92414 200898
rect 91794 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 92414 165454
rect 91794 165134 92414 165218
rect 91794 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 92414 165134
rect 91794 129454 92414 164898
rect 91794 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 92414 129454
rect 91794 129134 92414 129218
rect 91794 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 92414 129134
rect 91794 93454 92414 128898
rect 91794 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 92414 93454
rect 91794 93134 92414 93218
rect 91794 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 92414 93134
rect 91794 57454 92414 92898
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -1306 92414 20898
rect 91794 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 92414 -1306
rect 91794 -1626 92414 -1542
rect 91794 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 92414 -1626
rect 91794 -1894 92414 -1862
rect 95514 673174 96134 707162
rect 95514 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 96134 673174
rect 95514 672854 96134 672938
rect 95514 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 96134 672854
rect 95514 637174 96134 672618
rect 95514 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 96134 637174
rect 95514 636854 96134 636938
rect 95514 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 96134 636854
rect 95514 601174 96134 636618
rect 95514 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 96134 601174
rect 95514 600854 96134 600938
rect 95514 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 96134 600854
rect 95514 565174 96134 600618
rect 95514 564938 95546 565174
rect 95782 564938 95866 565174
rect 96102 564938 96134 565174
rect 95514 564854 96134 564938
rect 95514 564618 95546 564854
rect 95782 564618 95866 564854
rect 96102 564618 96134 564854
rect 95514 529174 96134 564618
rect 95514 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 96134 529174
rect 95514 528854 96134 528938
rect 95514 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 96134 528854
rect 95514 493174 96134 528618
rect 95514 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 96134 493174
rect 95514 492854 96134 492938
rect 95514 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 96134 492854
rect 95514 457174 96134 492618
rect 95514 456938 95546 457174
rect 95782 456938 95866 457174
rect 96102 456938 96134 457174
rect 95514 456854 96134 456938
rect 95514 456618 95546 456854
rect 95782 456618 95866 456854
rect 96102 456618 96134 456854
rect 95514 421174 96134 456618
rect 95514 420938 95546 421174
rect 95782 420938 95866 421174
rect 96102 420938 96134 421174
rect 95514 420854 96134 420938
rect 95514 420618 95546 420854
rect 95782 420618 95866 420854
rect 96102 420618 96134 420854
rect 95514 385174 96134 420618
rect 95514 384938 95546 385174
rect 95782 384938 95866 385174
rect 96102 384938 96134 385174
rect 95514 384854 96134 384938
rect 95514 384618 95546 384854
rect 95782 384618 95866 384854
rect 96102 384618 96134 384854
rect 95514 349174 96134 384618
rect 95514 348938 95546 349174
rect 95782 348938 95866 349174
rect 96102 348938 96134 349174
rect 95514 348854 96134 348938
rect 95514 348618 95546 348854
rect 95782 348618 95866 348854
rect 96102 348618 96134 348854
rect 95514 313174 96134 348618
rect 95514 312938 95546 313174
rect 95782 312938 95866 313174
rect 96102 312938 96134 313174
rect 95514 312854 96134 312938
rect 95514 312618 95546 312854
rect 95782 312618 95866 312854
rect 96102 312618 96134 312854
rect 95514 277174 96134 312618
rect 95514 276938 95546 277174
rect 95782 276938 95866 277174
rect 96102 276938 96134 277174
rect 95514 276854 96134 276938
rect 95514 276618 95546 276854
rect 95782 276618 95866 276854
rect 96102 276618 96134 276854
rect 95514 241174 96134 276618
rect 95514 240938 95546 241174
rect 95782 240938 95866 241174
rect 96102 240938 96134 241174
rect 95514 240854 96134 240938
rect 95514 240618 95546 240854
rect 95782 240618 95866 240854
rect 96102 240618 96134 240854
rect 95514 205174 96134 240618
rect 95514 204938 95546 205174
rect 95782 204938 95866 205174
rect 96102 204938 96134 205174
rect 95514 204854 96134 204938
rect 95514 204618 95546 204854
rect 95782 204618 95866 204854
rect 96102 204618 96134 204854
rect 95514 169174 96134 204618
rect 95514 168938 95546 169174
rect 95782 168938 95866 169174
rect 96102 168938 96134 169174
rect 95514 168854 96134 168938
rect 95514 168618 95546 168854
rect 95782 168618 95866 168854
rect 96102 168618 96134 168854
rect 95514 133174 96134 168618
rect 95514 132938 95546 133174
rect 95782 132938 95866 133174
rect 96102 132938 96134 133174
rect 95514 132854 96134 132938
rect 95514 132618 95546 132854
rect 95782 132618 95866 132854
rect 96102 132618 96134 132854
rect 95514 97174 96134 132618
rect 95514 96938 95546 97174
rect 95782 96938 95866 97174
rect 96102 96938 96134 97174
rect 95514 96854 96134 96938
rect 95514 96618 95546 96854
rect 95782 96618 95866 96854
rect 96102 96618 96134 96854
rect 95514 61174 96134 96618
rect 95514 60938 95546 61174
rect 95782 60938 95866 61174
rect 96102 60938 96134 61174
rect 95514 60854 96134 60938
rect 95514 60618 95546 60854
rect 95782 60618 95866 60854
rect 96102 60618 96134 60854
rect 95514 25174 96134 60618
rect 95514 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 96134 25174
rect 95514 24854 96134 24938
rect 95514 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 96134 24854
rect 95514 -3226 96134 24618
rect 95514 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 96134 -3226
rect 95514 -3546 96134 -3462
rect 95514 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 96134 -3546
rect 95514 -3814 96134 -3782
rect 99234 676894 99854 709082
rect 99234 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 99854 676894
rect 99234 676574 99854 676658
rect 99234 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 99854 676574
rect 99234 640894 99854 676338
rect 99234 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 99854 640894
rect 99234 640574 99854 640658
rect 99234 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 99854 640574
rect 99234 604894 99854 640338
rect 99234 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 99854 604894
rect 99234 604574 99854 604658
rect 99234 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 99854 604574
rect 99234 568894 99854 604338
rect 99234 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 99854 568894
rect 99234 568574 99854 568658
rect 99234 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 99854 568574
rect 99234 532894 99854 568338
rect 99234 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 99854 532894
rect 99234 532574 99854 532658
rect 99234 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 99854 532574
rect 99234 496894 99854 532338
rect 99234 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 99854 496894
rect 99234 496574 99854 496658
rect 99234 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 99854 496574
rect 99234 460894 99854 496338
rect 99234 460658 99266 460894
rect 99502 460658 99586 460894
rect 99822 460658 99854 460894
rect 99234 460574 99854 460658
rect 99234 460338 99266 460574
rect 99502 460338 99586 460574
rect 99822 460338 99854 460574
rect 99234 424894 99854 460338
rect 99234 424658 99266 424894
rect 99502 424658 99586 424894
rect 99822 424658 99854 424894
rect 99234 424574 99854 424658
rect 99234 424338 99266 424574
rect 99502 424338 99586 424574
rect 99822 424338 99854 424574
rect 99234 388894 99854 424338
rect 99234 388658 99266 388894
rect 99502 388658 99586 388894
rect 99822 388658 99854 388894
rect 99234 388574 99854 388658
rect 99234 388338 99266 388574
rect 99502 388338 99586 388574
rect 99822 388338 99854 388574
rect 99234 352894 99854 388338
rect 99234 352658 99266 352894
rect 99502 352658 99586 352894
rect 99822 352658 99854 352894
rect 99234 352574 99854 352658
rect 99234 352338 99266 352574
rect 99502 352338 99586 352574
rect 99822 352338 99854 352574
rect 99234 316894 99854 352338
rect 99234 316658 99266 316894
rect 99502 316658 99586 316894
rect 99822 316658 99854 316894
rect 99234 316574 99854 316658
rect 99234 316338 99266 316574
rect 99502 316338 99586 316574
rect 99822 316338 99854 316574
rect 99234 280894 99854 316338
rect 99234 280658 99266 280894
rect 99502 280658 99586 280894
rect 99822 280658 99854 280894
rect 99234 280574 99854 280658
rect 99234 280338 99266 280574
rect 99502 280338 99586 280574
rect 99822 280338 99854 280574
rect 99234 244894 99854 280338
rect 99234 244658 99266 244894
rect 99502 244658 99586 244894
rect 99822 244658 99854 244894
rect 99234 244574 99854 244658
rect 99234 244338 99266 244574
rect 99502 244338 99586 244574
rect 99822 244338 99854 244574
rect 99234 208894 99854 244338
rect 99234 208658 99266 208894
rect 99502 208658 99586 208894
rect 99822 208658 99854 208894
rect 99234 208574 99854 208658
rect 99234 208338 99266 208574
rect 99502 208338 99586 208574
rect 99822 208338 99854 208574
rect 99234 172894 99854 208338
rect 99234 172658 99266 172894
rect 99502 172658 99586 172894
rect 99822 172658 99854 172894
rect 99234 172574 99854 172658
rect 99234 172338 99266 172574
rect 99502 172338 99586 172574
rect 99822 172338 99854 172574
rect 99234 136894 99854 172338
rect 99234 136658 99266 136894
rect 99502 136658 99586 136894
rect 99822 136658 99854 136894
rect 99234 136574 99854 136658
rect 99234 136338 99266 136574
rect 99502 136338 99586 136574
rect 99822 136338 99854 136574
rect 99234 100894 99854 136338
rect 99234 100658 99266 100894
rect 99502 100658 99586 100894
rect 99822 100658 99854 100894
rect 99234 100574 99854 100658
rect 99234 100338 99266 100574
rect 99502 100338 99586 100574
rect 99822 100338 99854 100574
rect 99234 64894 99854 100338
rect 99234 64658 99266 64894
rect 99502 64658 99586 64894
rect 99822 64658 99854 64894
rect 99234 64574 99854 64658
rect 99234 64338 99266 64574
rect 99502 64338 99586 64574
rect 99822 64338 99854 64574
rect 99234 28894 99854 64338
rect 99234 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 99854 28894
rect 99234 28574 99854 28658
rect 99234 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 99854 28574
rect 99234 -5146 99854 28338
rect 99234 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 99854 -5146
rect 99234 -5466 99854 -5382
rect 99234 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 99854 -5466
rect 99234 -5734 99854 -5702
rect 102954 680614 103574 711002
rect 120954 710598 121574 711590
rect 120954 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 121574 710598
rect 120954 710278 121574 710362
rect 120954 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 121574 710278
rect 117234 708678 117854 709670
rect 117234 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 117854 708678
rect 117234 708358 117854 708442
rect 117234 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 117854 708358
rect 113514 706758 114134 707750
rect 113514 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 114134 706758
rect 113514 706438 114134 706522
rect 113514 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 114134 706438
rect 102954 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 103574 680614
rect 102954 680294 103574 680378
rect 102954 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 103574 680294
rect 102954 644614 103574 680058
rect 102954 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 103574 644614
rect 102954 644294 103574 644378
rect 102954 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 103574 644294
rect 102954 608614 103574 644058
rect 102954 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 103574 608614
rect 102954 608294 103574 608378
rect 102954 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 103574 608294
rect 102954 572614 103574 608058
rect 102954 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 103574 572614
rect 102954 572294 103574 572378
rect 102954 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 103574 572294
rect 102954 536614 103574 572058
rect 102954 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 103574 536614
rect 102954 536294 103574 536378
rect 102954 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 103574 536294
rect 102954 500614 103574 536058
rect 102954 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 103574 500614
rect 102954 500294 103574 500378
rect 102954 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 103574 500294
rect 102954 464614 103574 500058
rect 102954 464378 102986 464614
rect 103222 464378 103306 464614
rect 103542 464378 103574 464614
rect 102954 464294 103574 464378
rect 102954 464058 102986 464294
rect 103222 464058 103306 464294
rect 103542 464058 103574 464294
rect 102954 428614 103574 464058
rect 102954 428378 102986 428614
rect 103222 428378 103306 428614
rect 103542 428378 103574 428614
rect 102954 428294 103574 428378
rect 102954 428058 102986 428294
rect 103222 428058 103306 428294
rect 103542 428058 103574 428294
rect 102954 392614 103574 428058
rect 102954 392378 102986 392614
rect 103222 392378 103306 392614
rect 103542 392378 103574 392614
rect 102954 392294 103574 392378
rect 102954 392058 102986 392294
rect 103222 392058 103306 392294
rect 103542 392058 103574 392294
rect 102954 356614 103574 392058
rect 102954 356378 102986 356614
rect 103222 356378 103306 356614
rect 103542 356378 103574 356614
rect 102954 356294 103574 356378
rect 102954 356058 102986 356294
rect 103222 356058 103306 356294
rect 103542 356058 103574 356294
rect 102954 320614 103574 356058
rect 102954 320378 102986 320614
rect 103222 320378 103306 320614
rect 103542 320378 103574 320614
rect 102954 320294 103574 320378
rect 102954 320058 102986 320294
rect 103222 320058 103306 320294
rect 103542 320058 103574 320294
rect 102954 284614 103574 320058
rect 102954 284378 102986 284614
rect 103222 284378 103306 284614
rect 103542 284378 103574 284614
rect 102954 284294 103574 284378
rect 102954 284058 102986 284294
rect 103222 284058 103306 284294
rect 103542 284058 103574 284294
rect 102954 248614 103574 284058
rect 102954 248378 102986 248614
rect 103222 248378 103306 248614
rect 103542 248378 103574 248614
rect 102954 248294 103574 248378
rect 102954 248058 102986 248294
rect 103222 248058 103306 248294
rect 103542 248058 103574 248294
rect 102954 212614 103574 248058
rect 102954 212378 102986 212614
rect 103222 212378 103306 212614
rect 103542 212378 103574 212614
rect 102954 212294 103574 212378
rect 102954 212058 102986 212294
rect 103222 212058 103306 212294
rect 103542 212058 103574 212294
rect 102954 176614 103574 212058
rect 102954 176378 102986 176614
rect 103222 176378 103306 176614
rect 103542 176378 103574 176614
rect 102954 176294 103574 176378
rect 102954 176058 102986 176294
rect 103222 176058 103306 176294
rect 103542 176058 103574 176294
rect 102954 140614 103574 176058
rect 102954 140378 102986 140614
rect 103222 140378 103306 140614
rect 103542 140378 103574 140614
rect 102954 140294 103574 140378
rect 102954 140058 102986 140294
rect 103222 140058 103306 140294
rect 103542 140058 103574 140294
rect 102954 104614 103574 140058
rect 102954 104378 102986 104614
rect 103222 104378 103306 104614
rect 103542 104378 103574 104614
rect 102954 104294 103574 104378
rect 102954 104058 102986 104294
rect 103222 104058 103306 104294
rect 103542 104058 103574 104294
rect 102954 68614 103574 104058
rect 102954 68378 102986 68614
rect 103222 68378 103306 68614
rect 103542 68378 103574 68614
rect 102954 68294 103574 68378
rect 102954 68058 102986 68294
rect 103222 68058 103306 68294
rect 103542 68058 103574 68294
rect 102954 32614 103574 68058
rect 102954 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 103574 32614
rect 102954 32294 103574 32378
rect 102954 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 103574 32294
rect 84954 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 85574 -6106
rect 84954 -6426 85574 -6342
rect 84954 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 85574 -6426
rect 84954 -7654 85574 -6662
rect 102954 -7066 103574 32058
rect 109794 704838 110414 705830
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 109794 543454 110414 578898
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 109794 507454 110414 542898
rect 109794 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 110414 507454
rect 109794 507134 110414 507218
rect 109794 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 110414 507134
rect 109794 471454 110414 506898
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 109794 435454 110414 470898
rect 109794 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 110414 435454
rect 109794 435134 110414 435218
rect 109794 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 110414 435134
rect 109794 399454 110414 434898
rect 109794 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 110414 399454
rect 109794 399134 110414 399218
rect 109794 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 110414 399134
rect 109794 363454 110414 398898
rect 109794 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 110414 363454
rect 109794 363134 110414 363218
rect 109794 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 110414 363134
rect 109794 327454 110414 362898
rect 109794 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 110414 327454
rect 109794 327134 110414 327218
rect 109794 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 110414 327134
rect 109794 291454 110414 326898
rect 109794 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 110414 291454
rect 109794 291134 110414 291218
rect 109794 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 110414 291134
rect 109794 255454 110414 290898
rect 109794 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 110414 255454
rect 109794 255134 110414 255218
rect 109794 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 110414 255134
rect 109794 219454 110414 254898
rect 109794 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 110414 219454
rect 109794 219134 110414 219218
rect 109794 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 110414 219134
rect 109794 183454 110414 218898
rect 109794 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 110414 183454
rect 109794 183134 110414 183218
rect 109794 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 110414 183134
rect 109794 147454 110414 182898
rect 109794 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 110414 147454
rect 109794 147134 110414 147218
rect 109794 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 110414 147134
rect 109794 111454 110414 146898
rect 109794 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 110414 111454
rect 109794 111134 110414 111218
rect 109794 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 110414 111134
rect 109794 75454 110414 110898
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 109794 75134 110414 75218
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 109794 39454 110414 74898
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -1894 110414 -902
rect 113514 691174 114134 706202
rect 113514 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 114134 691174
rect 113514 690854 114134 690938
rect 113514 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 114134 690854
rect 113514 655174 114134 690618
rect 113514 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 114134 655174
rect 113514 654854 114134 654938
rect 113514 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 114134 654854
rect 113514 619174 114134 654618
rect 113514 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 114134 619174
rect 113514 618854 114134 618938
rect 113514 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 114134 618854
rect 113514 583174 114134 618618
rect 113514 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 114134 583174
rect 113514 582854 114134 582938
rect 113514 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 114134 582854
rect 113514 547174 114134 582618
rect 113514 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 114134 547174
rect 113514 546854 114134 546938
rect 113514 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 114134 546854
rect 113514 511174 114134 546618
rect 113514 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 114134 511174
rect 113514 510854 114134 510938
rect 113514 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 114134 510854
rect 113514 475174 114134 510618
rect 113514 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 114134 475174
rect 113514 474854 114134 474938
rect 113514 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 114134 474854
rect 113514 439174 114134 474618
rect 113514 438938 113546 439174
rect 113782 438938 113866 439174
rect 114102 438938 114134 439174
rect 113514 438854 114134 438938
rect 113514 438618 113546 438854
rect 113782 438618 113866 438854
rect 114102 438618 114134 438854
rect 113514 403174 114134 438618
rect 113514 402938 113546 403174
rect 113782 402938 113866 403174
rect 114102 402938 114134 403174
rect 113514 402854 114134 402938
rect 113514 402618 113546 402854
rect 113782 402618 113866 402854
rect 114102 402618 114134 402854
rect 113514 367174 114134 402618
rect 113514 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 114134 367174
rect 113514 366854 114134 366938
rect 113514 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 114134 366854
rect 113514 331174 114134 366618
rect 113514 330938 113546 331174
rect 113782 330938 113866 331174
rect 114102 330938 114134 331174
rect 113514 330854 114134 330938
rect 113514 330618 113546 330854
rect 113782 330618 113866 330854
rect 114102 330618 114134 330854
rect 113514 295174 114134 330618
rect 113514 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 114134 295174
rect 113514 294854 114134 294938
rect 113514 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 114134 294854
rect 113514 259174 114134 294618
rect 113514 258938 113546 259174
rect 113782 258938 113866 259174
rect 114102 258938 114134 259174
rect 113514 258854 114134 258938
rect 113514 258618 113546 258854
rect 113782 258618 113866 258854
rect 114102 258618 114134 258854
rect 113514 223174 114134 258618
rect 113514 222938 113546 223174
rect 113782 222938 113866 223174
rect 114102 222938 114134 223174
rect 113514 222854 114134 222938
rect 113514 222618 113546 222854
rect 113782 222618 113866 222854
rect 114102 222618 114134 222854
rect 113514 187174 114134 222618
rect 113514 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 114134 187174
rect 113514 186854 114134 186938
rect 113514 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 114134 186854
rect 113514 151174 114134 186618
rect 113514 150938 113546 151174
rect 113782 150938 113866 151174
rect 114102 150938 114134 151174
rect 113514 150854 114134 150938
rect 113514 150618 113546 150854
rect 113782 150618 113866 150854
rect 114102 150618 114134 150854
rect 113514 115174 114134 150618
rect 113514 114938 113546 115174
rect 113782 114938 113866 115174
rect 114102 114938 114134 115174
rect 113514 114854 114134 114938
rect 113514 114618 113546 114854
rect 113782 114618 113866 114854
rect 114102 114618 114134 114854
rect 113514 79174 114134 114618
rect 113514 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 114134 79174
rect 113514 78854 114134 78938
rect 113514 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 114134 78854
rect 113514 43174 114134 78618
rect 113514 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 114134 43174
rect 113514 42854 114134 42938
rect 113514 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 114134 42854
rect 113514 7174 114134 42618
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 113514 -2266 114134 6618
rect 113514 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 114134 -2266
rect 113514 -2586 114134 -2502
rect 113514 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 114134 -2586
rect 113514 -3814 114134 -2822
rect 117234 694894 117854 708122
rect 117234 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 117854 694894
rect 117234 694574 117854 694658
rect 117234 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 117854 694574
rect 117234 658894 117854 694338
rect 117234 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 117854 658894
rect 117234 658574 117854 658658
rect 117234 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 117854 658574
rect 117234 622894 117854 658338
rect 117234 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 117854 622894
rect 117234 622574 117854 622658
rect 117234 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 117854 622574
rect 117234 586894 117854 622338
rect 117234 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 117854 586894
rect 117234 586574 117854 586658
rect 117234 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 117854 586574
rect 117234 550894 117854 586338
rect 117234 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 117854 550894
rect 117234 550574 117854 550658
rect 117234 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 117854 550574
rect 117234 514894 117854 550338
rect 117234 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 117854 514894
rect 117234 514574 117854 514658
rect 117234 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 117854 514574
rect 117234 478894 117854 514338
rect 117234 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 117854 478894
rect 117234 478574 117854 478658
rect 117234 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 117854 478574
rect 117234 442894 117854 478338
rect 117234 442658 117266 442894
rect 117502 442658 117586 442894
rect 117822 442658 117854 442894
rect 117234 442574 117854 442658
rect 117234 442338 117266 442574
rect 117502 442338 117586 442574
rect 117822 442338 117854 442574
rect 117234 406894 117854 442338
rect 117234 406658 117266 406894
rect 117502 406658 117586 406894
rect 117822 406658 117854 406894
rect 117234 406574 117854 406658
rect 117234 406338 117266 406574
rect 117502 406338 117586 406574
rect 117822 406338 117854 406574
rect 117234 370894 117854 406338
rect 117234 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 117854 370894
rect 117234 370574 117854 370658
rect 117234 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 117854 370574
rect 117234 334894 117854 370338
rect 117234 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 117854 334894
rect 117234 334574 117854 334658
rect 117234 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 117854 334574
rect 117234 298894 117854 334338
rect 117234 298658 117266 298894
rect 117502 298658 117586 298894
rect 117822 298658 117854 298894
rect 117234 298574 117854 298658
rect 117234 298338 117266 298574
rect 117502 298338 117586 298574
rect 117822 298338 117854 298574
rect 117234 262894 117854 298338
rect 117234 262658 117266 262894
rect 117502 262658 117586 262894
rect 117822 262658 117854 262894
rect 117234 262574 117854 262658
rect 117234 262338 117266 262574
rect 117502 262338 117586 262574
rect 117822 262338 117854 262574
rect 117234 226894 117854 262338
rect 117234 226658 117266 226894
rect 117502 226658 117586 226894
rect 117822 226658 117854 226894
rect 117234 226574 117854 226658
rect 117234 226338 117266 226574
rect 117502 226338 117586 226574
rect 117822 226338 117854 226574
rect 117234 190894 117854 226338
rect 117234 190658 117266 190894
rect 117502 190658 117586 190894
rect 117822 190658 117854 190894
rect 117234 190574 117854 190658
rect 117234 190338 117266 190574
rect 117502 190338 117586 190574
rect 117822 190338 117854 190574
rect 117234 154894 117854 190338
rect 117234 154658 117266 154894
rect 117502 154658 117586 154894
rect 117822 154658 117854 154894
rect 117234 154574 117854 154658
rect 117234 154338 117266 154574
rect 117502 154338 117586 154574
rect 117822 154338 117854 154574
rect 117234 118894 117854 154338
rect 117234 118658 117266 118894
rect 117502 118658 117586 118894
rect 117822 118658 117854 118894
rect 117234 118574 117854 118658
rect 117234 118338 117266 118574
rect 117502 118338 117586 118574
rect 117822 118338 117854 118574
rect 117234 82894 117854 118338
rect 117234 82658 117266 82894
rect 117502 82658 117586 82894
rect 117822 82658 117854 82894
rect 117234 82574 117854 82658
rect 117234 82338 117266 82574
rect 117502 82338 117586 82574
rect 117822 82338 117854 82574
rect 117234 46894 117854 82338
rect 117234 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 117854 46894
rect 117234 46574 117854 46658
rect 117234 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 117854 46574
rect 117234 10894 117854 46338
rect 117234 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 117854 10894
rect 117234 10574 117854 10658
rect 117234 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 117854 10574
rect 117234 -4186 117854 10338
rect 117234 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 117854 -4186
rect 117234 -4506 117854 -4422
rect 117234 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 117854 -4506
rect 117234 -5734 117854 -4742
rect 120954 698614 121574 710042
rect 138954 711558 139574 711590
rect 138954 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 139574 711558
rect 138954 711238 139574 711322
rect 138954 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 139574 711238
rect 135234 709638 135854 709670
rect 135234 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 135854 709638
rect 135234 709318 135854 709402
rect 135234 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 135854 709318
rect 131514 707718 132134 707750
rect 131514 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 132134 707718
rect 131514 707398 132134 707482
rect 131514 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 132134 707398
rect 120954 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 121574 698614
rect 120954 698294 121574 698378
rect 120954 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 121574 698294
rect 120954 662614 121574 698058
rect 120954 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 121574 662614
rect 120954 662294 121574 662378
rect 120954 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 121574 662294
rect 120954 626614 121574 662058
rect 120954 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 121574 626614
rect 120954 626294 121574 626378
rect 120954 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 121574 626294
rect 120954 590614 121574 626058
rect 120954 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 121574 590614
rect 120954 590294 121574 590378
rect 120954 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 121574 590294
rect 120954 554614 121574 590058
rect 120954 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 121574 554614
rect 120954 554294 121574 554378
rect 120954 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 121574 554294
rect 120954 518614 121574 554058
rect 120954 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 121574 518614
rect 120954 518294 121574 518378
rect 120954 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 121574 518294
rect 120954 482614 121574 518058
rect 120954 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 121574 482614
rect 120954 482294 121574 482378
rect 120954 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 121574 482294
rect 120954 446614 121574 482058
rect 120954 446378 120986 446614
rect 121222 446378 121306 446614
rect 121542 446378 121574 446614
rect 120954 446294 121574 446378
rect 120954 446058 120986 446294
rect 121222 446058 121306 446294
rect 121542 446058 121574 446294
rect 120954 410614 121574 446058
rect 120954 410378 120986 410614
rect 121222 410378 121306 410614
rect 121542 410378 121574 410614
rect 120954 410294 121574 410378
rect 120954 410058 120986 410294
rect 121222 410058 121306 410294
rect 121542 410058 121574 410294
rect 120954 374614 121574 410058
rect 120954 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 121574 374614
rect 120954 374294 121574 374378
rect 120954 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 121574 374294
rect 120954 338614 121574 374058
rect 120954 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 121574 338614
rect 120954 338294 121574 338378
rect 120954 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 121574 338294
rect 120954 302614 121574 338058
rect 120954 302378 120986 302614
rect 121222 302378 121306 302614
rect 121542 302378 121574 302614
rect 120954 302294 121574 302378
rect 120954 302058 120986 302294
rect 121222 302058 121306 302294
rect 121542 302058 121574 302294
rect 120954 266614 121574 302058
rect 120954 266378 120986 266614
rect 121222 266378 121306 266614
rect 121542 266378 121574 266614
rect 120954 266294 121574 266378
rect 120954 266058 120986 266294
rect 121222 266058 121306 266294
rect 121542 266058 121574 266294
rect 120954 230614 121574 266058
rect 120954 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 121574 230614
rect 120954 230294 121574 230378
rect 120954 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 121574 230294
rect 120954 194614 121574 230058
rect 120954 194378 120986 194614
rect 121222 194378 121306 194614
rect 121542 194378 121574 194614
rect 120954 194294 121574 194378
rect 120954 194058 120986 194294
rect 121222 194058 121306 194294
rect 121542 194058 121574 194294
rect 120954 158614 121574 194058
rect 120954 158378 120986 158614
rect 121222 158378 121306 158614
rect 121542 158378 121574 158614
rect 120954 158294 121574 158378
rect 120954 158058 120986 158294
rect 121222 158058 121306 158294
rect 121542 158058 121574 158294
rect 120954 122614 121574 158058
rect 120954 122378 120986 122614
rect 121222 122378 121306 122614
rect 121542 122378 121574 122614
rect 120954 122294 121574 122378
rect 120954 122058 120986 122294
rect 121222 122058 121306 122294
rect 121542 122058 121574 122294
rect 120954 86614 121574 122058
rect 120954 86378 120986 86614
rect 121222 86378 121306 86614
rect 121542 86378 121574 86614
rect 120954 86294 121574 86378
rect 120954 86058 120986 86294
rect 121222 86058 121306 86294
rect 121542 86058 121574 86294
rect 120954 50614 121574 86058
rect 120954 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 121574 50614
rect 120954 50294 121574 50378
rect 120954 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 121574 50294
rect 120954 14614 121574 50058
rect 120954 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 121574 14614
rect 120954 14294 121574 14378
rect 120954 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 121574 14294
rect 102954 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 103574 -7066
rect 102954 -7386 103574 -7302
rect 102954 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 103574 -7386
rect 102954 -7654 103574 -7622
rect 120954 -6106 121574 14058
rect 127794 705798 128414 705830
rect 127794 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 128414 705798
rect 127794 705478 128414 705562
rect 127794 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 128414 705478
rect 127794 669454 128414 705242
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 127794 561454 128414 596898
rect 127794 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 128414 561454
rect 127794 561134 128414 561218
rect 127794 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 128414 561134
rect 127794 525454 128414 560898
rect 127794 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 128414 525454
rect 127794 525134 128414 525218
rect 127794 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 128414 525134
rect 127794 489454 128414 524898
rect 127794 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 128414 489454
rect 127794 489134 128414 489218
rect 127794 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 128414 489134
rect 127794 453454 128414 488898
rect 127794 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 128414 453454
rect 127794 453134 128414 453218
rect 127794 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 128414 453134
rect 127794 417454 128414 452898
rect 127794 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 128414 417454
rect 127794 417134 128414 417218
rect 127794 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 128414 417134
rect 127794 381454 128414 416898
rect 127794 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 128414 381454
rect 127794 381134 128414 381218
rect 127794 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 128414 381134
rect 127794 345454 128414 380898
rect 127794 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 128414 345454
rect 127794 345134 128414 345218
rect 127794 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 128414 345134
rect 127794 309454 128414 344898
rect 127794 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 128414 309454
rect 127794 309134 128414 309218
rect 127794 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 128414 309134
rect 127794 273454 128414 308898
rect 127794 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 128414 273454
rect 127794 273134 128414 273218
rect 127794 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 128414 273134
rect 127794 237454 128414 272898
rect 127794 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 128414 237454
rect 127794 237134 128414 237218
rect 127794 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 128414 237134
rect 127794 201454 128414 236898
rect 127794 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 128414 201454
rect 127794 201134 128414 201218
rect 127794 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 128414 201134
rect 127794 165454 128414 200898
rect 127794 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 128414 165454
rect 127794 165134 128414 165218
rect 127794 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 128414 165134
rect 127794 129454 128414 164898
rect 127794 129218 127826 129454
rect 128062 129218 128146 129454
rect 128382 129218 128414 129454
rect 127794 129134 128414 129218
rect 127794 128898 127826 129134
rect 128062 128898 128146 129134
rect 128382 128898 128414 129134
rect 127794 93454 128414 128898
rect 127794 93218 127826 93454
rect 128062 93218 128146 93454
rect 128382 93218 128414 93454
rect 127794 93134 128414 93218
rect 127794 92898 127826 93134
rect 128062 92898 128146 93134
rect 128382 92898 128414 93134
rect 127794 57454 128414 92898
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -1306 128414 20898
rect 127794 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 128414 -1306
rect 127794 -1626 128414 -1542
rect 127794 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 128414 -1626
rect 127794 -1894 128414 -1862
rect 131514 673174 132134 707162
rect 131514 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 132134 673174
rect 131514 672854 132134 672938
rect 131514 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 132134 672854
rect 131514 637174 132134 672618
rect 131514 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 132134 637174
rect 131514 636854 132134 636938
rect 131514 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 132134 636854
rect 131514 601174 132134 636618
rect 131514 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 132134 601174
rect 131514 600854 132134 600938
rect 131514 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 132134 600854
rect 131514 565174 132134 600618
rect 131514 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 132134 565174
rect 131514 564854 132134 564938
rect 131514 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 132134 564854
rect 131514 529174 132134 564618
rect 131514 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 132134 529174
rect 131514 528854 132134 528938
rect 131514 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 132134 528854
rect 131514 493174 132134 528618
rect 131514 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 132134 493174
rect 131514 492854 132134 492938
rect 131514 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 132134 492854
rect 131514 457174 132134 492618
rect 131514 456938 131546 457174
rect 131782 456938 131866 457174
rect 132102 456938 132134 457174
rect 131514 456854 132134 456938
rect 131514 456618 131546 456854
rect 131782 456618 131866 456854
rect 132102 456618 132134 456854
rect 131514 421174 132134 456618
rect 131514 420938 131546 421174
rect 131782 420938 131866 421174
rect 132102 420938 132134 421174
rect 131514 420854 132134 420938
rect 131514 420618 131546 420854
rect 131782 420618 131866 420854
rect 132102 420618 132134 420854
rect 131514 385174 132134 420618
rect 131514 384938 131546 385174
rect 131782 384938 131866 385174
rect 132102 384938 132134 385174
rect 131514 384854 132134 384938
rect 131514 384618 131546 384854
rect 131782 384618 131866 384854
rect 132102 384618 132134 384854
rect 131514 349174 132134 384618
rect 131514 348938 131546 349174
rect 131782 348938 131866 349174
rect 132102 348938 132134 349174
rect 131514 348854 132134 348938
rect 131514 348618 131546 348854
rect 131782 348618 131866 348854
rect 132102 348618 132134 348854
rect 131514 313174 132134 348618
rect 131514 312938 131546 313174
rect 131782 312938 131866 313174
rect 132102 312938 132134 313174
rect 131514 312854 132134 312938
rect 131514 312618 131546 312854
rect 131782 312618 131866 312854
rect 132102 312618 132134 312854
rect 131514 277174 132134 312618
rect 131514 276938 131546 277174
rect 131782 276938 131866 277174
rect 132102 276938 132134 277174
rect 131514 276854 132134 276938
rect 131514 276618 131546 276854
rect 131782 276618 131866 276854
rect 132102 276618 132134 276854
rect 131514 241174 132134 276618
rect 131514 240938 131546 241174
rect 131782 240938 131866 241174
rect 132102 240938 132134 241174
rect 131514 240854 132134 240938
rect 131514 240618 131546 240854
rect 131782 240618 131866 240854
rect 132102 240618 132134 240854
rect 131514 205174 132134 240618
rect 131514 204938 131546 205174
rect 131782 204938 131866 205174
rect 132102 204938 132134 205174
rect 131514 204854 132134 204938
rect 131514 204618 131546 204854
rect 131782 204618 131866 204854
rect 132102 204618 132134 204854
rect 131514 169174 132134 204618
rect 131514 168938 131546 169174
rect 131782 168938 131866 169174
rect 132102 168938 132134 169174
rect 131514 168854 132134 168938
rect 131514 168618 131546 168854
rect 131782 168618 131866 168854
rect 132102 168618 132134 168854
rect 131514 133174 132134 168618
rect 131514 132938 131546 133174
rect 131782 132938 131866 133174
rect 132102 132938 132134 133174
rect 131514 132854 132134 132938
rect 131514 132618 131546 132854
rect 131782 132618 131866 132854
rect 132102 132618 132134 132854
rect 131514 97174 132134 132618
rect 131514 96938 131546 97174
rect 131782 96938 131866 97174
rect 132102 96938 132134 97174
rect 131514 96854 132134 96938
rect 131514 96618 131546 96854
rect 131782 96618 131866 96854
rect 132102 96618 132134 96854
rect 131514 61174 132134 96618
rect 131514 60938 131546 61174
rect 131782 60938 131866 61174
rect 132102 60938 132134 61174
rect 131514 60854 132134 60938
rect 131514 60618 131546 60854
rect 131782 60618 131866 60854
rect 132102 60618 132134 60854
rect 131514 25174 132134 60618
rect 131514 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 132134 25174
rect 131514 24854 132134 24938
rect 131514 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 132134 24854
rect 131514 -3226 132134 24618
rect 131514 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 132134 -3226
rect 131514 -3546 132134 -3462
rect 131514 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 132134 -3546
rect 131514 -3814 132134 -3782
rect 135234 676894 135854 709082
rect 135234 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 135854 676894
rect 135234 676574 135854 676658
rect 135234 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 135854 676574
rect 135234 640894 135854 676338
rect 135234 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 135854 640894
rect 135234 640574 135854 640658
rect 135234 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 135854 640574
rect 135234 604894 135854 640338
rect 135234 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 135854 604894
rect 135234 604574 135854 604658
rect 135234 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 135854 604574
rect 135234 568894 135854 604338
rect 135234 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 135854 568894
rect 135234 568574 135854 568658
rect 135234 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 135854 568574
rect 135234 532894 135854 568338
rect 135234 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 135854 532894
rect 135234 532574 135854 532658
rect 135234 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 135854 532574
rect 135234 496894 135854 532338
rect 135234 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 135854 496894
rect 135234 496574 135854 496658
rect 135234 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 135854 496574
rect 135234 460894 135854 496338
rect 135234 460658 135266 460894
rect 135502 460658 135586 460894
rect 135822 460658 135854 460894
rect 135234 460574 135854 460658
rect 135234 460338 135266 460574
rect 135502 460338 135586 460574
rect 135822 460338 135854 460574
rect 135234 424894 135854 460338
rect 135234 424658 135266 424894
rect 135502 424658 135586 424894
rect 135822 424658 135854 424894
rect 135234 424574 135854 424658
rect 135234 424338 135266 424574
rect 135502 424338 135586 424574
rect 135822 424338 135854 424574
rect 135234 388894 135854 424338
rect 135234 388658 135266 388894
rect 135502 388658 135586 388894
rect 135822 388658 135854 388894
rect 135234 388574 135854 388658
rect 135234 388338 135266 388574
rect 135502 388338 135586 388574
rect 135822 388338 135854 388574
rect 135234 352894 135854 388338
rect 135234 352658 135266 352894
rect 135502 352658 135586 352894
rect 135822 352658 135854 352894
rect 135234 352574 135854 352658
rect 135234 352338 135266 352574
rect 135502 352338 135586 352574
rect 135822 352338 135854 352574
rect 135234 316894 135854 352338
rect 135234 316658 135266 316894
rect 135502 316658 135586 316894
rect 135822 316658 135854 316894
rect 135234 316574 135854 316658
rect 135234 316338 135266 316574
rect 135502 316338 135586 316574
rect 135822 316338 135854 316574
rect 135234 280894 135854 316338
rect 135234 280658 135266 280894
rect 135502 280658 135586 280894
rect 135822 280658 135854 280894
rect 135234 280574 135854 280658
rect 135234 280338 135266 280574
rect 135502 280338 135586 280574
rect 135822 280338 135854 280574
rect 135234 244894 135854 280338
rect 135234 244658 135266 244894
rect 135502 244658 135586 244894
rect 135822 244658 135854 244894
rect 135234 244574 135854 244658
rect 135234 244338 135266 244574
rect 135502 244338 135586 244574
rect 135822 244338 135854 244574
rect 135234 208894 135854 244338
rect 135234 208658 135266 208894
rect 135502 208658 135586 208894
rect 135822 208658 135854 208894
rect 135234 208574 135854 208658
rect 135234 208338 135266 208574
rect 135502 208338 135586 208574
rect 135822 208338 135854 208574
rect 135234 172894 135854 208338
rect 135234 172658 135266 172894
rect 135502 172658 135586 172894
rect 135822 172658 135854 172894
rect 135234 172574 135854 172658
rect 135234 172338 135266 172574
rect 135502 172338 135586 172574
rect 135822 172338 135854 172574
rect 135234 136894 135854 172338
rect 135234 136658 135266 136894
rect 135502 136658 135586 136894
rect 135822 136658 135854 136894
rect 135234 136574 135854 136658
rect 135234 136338 135266 136574
rect 135502 136338 135586 136574
rect 135822 136338 135854 136574
rect 135234 100894 135854 136338
rect 135234 100658 135266 100894
rect 135502 100658 135586 100894
rect 135822 100658 135854 100894
rect 135234 100574 135854 100658
rect 135234 100338 135266 100574
rect 135502 100338 135586 100574
rect 135822 100338 135854 100574
rect 135234 64894 135854 100338
rect 135234 64658 135266 64894
rect 135502 64658 135586 64894
rect 135822 64658 135854 64894
rect 135234 64574 135854 64658
rect 135234 64338 135266 64574
rect 135502 64338 135586 64574
rect 135822 64338 135854 64574
rect 135234 28894 135854 64338
rect 135234 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 135854 28894
rect 135234 28574 135854 28658
rect 135234 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 135854 28574
rect 135234 -5146 135854 28338
rect 135234 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 135854 -5146
rect 135234 -5466 135854 -5382
rect 135234 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 135854 -5466
rect 135234 -5734 135854 -5702
rect 138954 680614 139574 711002
rect 156954 710598 157574 711590
rect 156954 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 157574 710598
rect 156954 710278 157574 710362
rect 156954 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 157574 710278
rect 153234 708678 153854 709670
rect 153234 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 153854 708678
rect 153234 708358 153854 708442
rect 153234 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 153854 708358
rect 149514 706758 150134 707750
rect 149514 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 150134 706758
rect 149514 706438 150134 706522
rect 149514 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 150134 706438
rect 138954 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 139574 680614
rect 138954 680294 139574 680378
rect 138954 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 139574 680294
rect 138954 644614 139574 680058
rect 138954 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 139574 644614
rect 138954 644294 139574 644378
rect 138954 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 139574 644294
rect 138954 608614 139574 644058
rect 138954 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 139574 608614
rect 138954 608294 139574 608378
rect 138954 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 139574 608294
rect 138954 572614 139574 608058
rect 138954 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 139574 572614
rect 138954 572294 139574 572378
rect 138954 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 139574 572294
rect 138954 536614 139574 572058
rect 138954 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 139574 536614
rect 138954 536294 139574 536378
rect 138954 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 139574 536294
rect 138954 500614 139574 536058
rect 138954 500378 138986 500614
rect 139222 500378 139306 500614
rect 139542 500378 139574 500614
rect 138954 500294 139574 500378
rect 138954 500058 138986 500294
rect 139222 500058 139306 500294
rect 139542 500058 139574 500294
rect 138954 464614 139574 500058
rect 138954 464378 138986 464614
rect 139222 464378 139306 464614
rect 139542 464378 139574 464614
rect 138954 464294 139574 464378
rect 138954 464058 138986 464294
rect 139222 464058 139306 464294
rect 139542 464058 139574 464294
rect 138954 428614 139574 464058
rect 138954 428378 138986 428614
rect 139222 428378 139306 428614
rect 139542 428378 139574 428614
rect 138954 428294 139574 428378
rect 138954 428058 138986 428294
rect 139222 428058 139306 428294
rect 139542 428058 139574 428294
rect 138954 392614 139574 428058
rect 138954 392378 138986 392614
rect 139222 392378 139306 392614
rect 139542 392378 139574 392614
rect 138954 392294 139574 392378
rect 138954 392058 138986 392294
rect 139222 392058 139306 392294
rect 139542 392058 139574 392294
rect 138954 356614 139574 392058
rect 138954 356378 138986 356614
rect 139222 356378 139306 356614
rect 139542 356378 139574 356614
rect 138954 356294 139574 356378
rect 138954 356058 138986 356294
rect 139222 356058 139306 356294
rect 139542 356058 139574 356294
rect 138954 320614 139574 356058
rect 138954 320378 138986 320614
rect 139222 320378 139306 320614
rect 139542 320378 139574 320614
rect 138954 320294 139574 320378
rect 138954 320058 138986 320294
rect 139222 320058 139306 320294
rect 139542 320058 139574 320294
rect 138954 284614 139574 320058
rect 138954 284378 138986 284614
rect 139222 284378 139306 284614
rect 139542 284378 139574 284614
rect 138954 284294 139574 284378
rect 138954 284058 138986 284294
rect 139222 284058 139306 284294
rect 139542 284058 139574 284294
rect 138954 248614 139574 284058
rect 138954 248378 138986 248614
rect 139222 248378 139306 248614
rect 139542 248378 139574 248614
rect 138954 248294 139574 248378
rect 138954 248058 138986 248294
rect 139222 248058 139306 248294
rect 139542 248058 139574 248294
rect 138954 212614 139574 248058
rect 138954 212378 138986 212614
rect 139222 212378 139306 212614
rect 139542 212378 139574 212614
rect 138954 212294 139574 212378
rect 138954 212058 138986 212294
rect 139222 212058 139306 212294
rect 139542 212058 139574 212294
rect 138954 176614 139574 212058
rect 138954 176378 138986 176614
rect 139222 176378 139306 176614
rect 139542 176378 139574 176614
rect 138954 176294 139574 176378
rect 138954 176058 138986 176294
rect 139222 176058 139306 176294
rect 139542 176058 139574 176294
rect 138954 140614 139574 176058
rect 138954 140378 138986 140614
rect 139222 140378 139306 140614
rect 139542 140378 139574 140614
rect 138954 140294 139574 140378
rect 138954 140058 138986 140294
rect 139222 140058 139306 140294
rect 139542 140058 139574 140294
rect 138954 104614 139574 140058
rect 138954 104378 138986 104614
rect 139222 104378 139306 104614
rect 139542 104378 139574 104614
rect 138954 104294 139574 104378
rect 138954 104058 138986 104294
rect 139222 104058 139306 104294
rect 139542 104058 139574 104294
rect 138954 68614 139574 104058
rect 138954 68378 138986 68614
rect 139222 68378 139306 68614
rect 139542 68378 139574 68614
rect 138954 68294 139574 68378
rect 138954 68058 138986 68294
rect 139222 68058 139306 68294
rect 139542 68058 139574 68294
rect 138954 32614 139574 68058
rect 138954 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 139574 32614
rect 138954 32294 139574 32378
rect 138954 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 139574 32294
rect 120954 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 121574 -6106
rect 120954 -6426 121574 -6342
rect 120954 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 121574 -6426
rect 120954 -7654 121574 -6662
rect 138954 -7066 139574 32058
rect 145794 704838 146414 705830
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 543454 146414 578898
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 507454 146414 542898
rect 145794 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 146414 507454
rect 145794 507134 146414 507218
rect 145794 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 146414 507134
rect 145794 471454 146414 506898
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 435454 146414 470898
rect 145794 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 146414 435454
rect 145794 435134 146414 435218
rect 145794 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 146414 435134
rect 145794 399454 146414 434898
rect 145794 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 146414 399454
rect 145794 399134 146414 399218
rect 145794 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 146414 399134
rect 145794 363454 146414 398898
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 145794 327454 146414 362898
rect 145794 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 146414 327454
rect 145794 327134 146414 327218
rect 145794 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 146414 327134
rect 145794 291454 146414 326898
rect 145794 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 146414 291454
rect 145794 291134 146414 291218
rect 145794 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 146414 291134
rect 145794 255454 146414 290898
rect 145794 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 146414 255454
rect 145794 255134 146414 255218
rect 145794 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 146414 255134
rect 145794 219454 146414 254898
rect 145794 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 146414 219454
rect 145794 219134 146414 219218
rect 145794 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 146414 219134
rect 145794 183454 146414 218898
rect 145794 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 146414 183454
rect 145794 183134 146414 183218
rect 145794 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 146414 183134
rect 145794 147454 146414 182898
rect 145794 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 146414 147454
rect 145794 147134 146414 147218
rect 145794 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 146414 147134
rect 145794 111454 146414 146898
rect 145794 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 146414 111454
rect 145794 111134 146414 111218
rect 145794 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 146414 111134
rect 145794 75454 146414 110898
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145794 75134 146414 75218
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 145794 39454 146414 74898
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -1894 146414 -902
rect 149514 691174 150134 706202
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 655174 150134 690618
rect 149514 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 150134 655174
rect 149514 654854 150134 654938
rect 149514 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 150134 654854
rect 149514 619174 150134 654618
rect 149514 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 150134 619174
rect 149514 618854 150134 618938
rect 149514 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 150134 618854
rect 149514 583174 150134 618618
rect 149514 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 150134 583174
rect 149514 582854 150134 582938
rect 149514 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 150134 582854
rect 149514 547174 150134 582618
rect 149514 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 150134 547174
rect 149514 546854 150134 546938
rect 149514 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 150134 546854
rect 149514 511174 150134 546618
rect 149514 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 150134 511174
rect 149514 510854 150134 510938
rect 149514 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 150134 510854
rect 149514 475174 150134 510618
rect 149514 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 150134 475174
rect 149514 474854 150134 474938
rect 149514 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 150134 474854
rect 149514 439174 150134 474618
rect 149514 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 150134 439174
rect 149514 438854 150134 438938
rect 149514 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 150134 438854
rect 149514 403174 150134 438618
rect 149514 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 150134 403174
rect 149514 402854 150134 402938
rect 149514 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 150134 402854
rect 149514 367174 150134 402618
rect 149514 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 150134 367174
rect 149514 366854 150134 366938
rect 149514 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 150134 366854
rect 149514 331174 150134 366618
rect 149514 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 150134 331174
rect 149514 330854 150134 330938
rect 149514 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 150134 330854
rect 149514 295174 150134 330618
rect 149514 294938 149546 295174
rect 149782 294938 149866 295174
rect 150102 294938 150134 295174
rect 149514 294854 150134 294938
rect 149514 294618 149546 294854
rect 149782 294618 149866 294854
rect 150102 294618 150134 294854
rect 149514 259174 150134 294618
rect 149514 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 150134 259174
rect 149514 258854 150134 258938
rect 149514 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 150134 258854
rect 149514 223174 150134 258618
rect 149514 222938 149546 223174
rect 149782 222938 149866 223174
rect 150102 222938 150134 223174
rect 149514 222854 150134 222938
rect 149514 222618 149546 222854
rect 149782 222618 149866 222854
rect 150102 222618 150134 222854
rect 149514 187174 150134 222618
rect 149514 186938 149546 187174
rect 149782 186938 149866 187174
rect 150102 186938 150134 187174
rect 149514 186854 150134 186938
rect 149514 186618 149546 186854
rect 149782 186618 149866 186854
rect 150102 186618 150134 186854
rect 149514 151174 150134 186618
rect 149514 150938 149546 151174
rect 149782 150938 149866 151174
rect 150102 150938 150134 151174
rect 149514 150854 150134 150938
rect 149514 150618 149546 150854
rect 149782 150618 149866 150854
rect 150102 150618 150134 150854
rect 149514 115174 150134 150618
rect 149514 114938 149546 115174
rect 149782 114938 149866 115174
rect 150102 114938 150134 115174
rect 149514 114854 150134 114938
rect 149514 114618 149546 114854
rect 149782 114618 149866 114854
rect 150102 114618 150134 114854
rect 149514 79174 150134 114618
rect 149514 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 150134 79174
rect 149514 78854 150134 78938
rect 149514 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 150134 78854
rect 149514 43174 150134 78618
rect 149514 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 150134 43174
rect 149514 42854 150134 42938
rect 149514 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 150134 42854
rect 149514 7174 150134 42618
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 149514 -2266 150134 6618
rect 149514 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 150134 -2266
rect 149514 -2586 150134 -2502
rect 149514 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 150134 -2586
rect 149514 -3814 150134 -2822
rect 153234 694894 153854 708122
rect 153234 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 153854 694894
rect 153234 694574 153854 694658
rect 153234 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 153854 694574
rect 153234 658894 153854 694338
rect 153234 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 153854 658894
rect 153234 658574 153854 658658
rect 153234 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 153854 658574
rect 153234 622894 153854 658338
rect 153234 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 153854 622894
rect 153234 622574 153854 622658
rect 153234 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 153854 622574
rect 153234 586894 153854 622338
rect 153234 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 153854 586894
rect 153234 586574 153854 586658
rect 153234 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 153854 586574
rect 153234 550894 153854 586338
rect 153234 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 153854 550894
rect 153234 550574 153854 550658
rect 153234 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 153854 550574
rect 153234 514894 153854 550338
rect 153234 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 153854 514894
rect 153234 514574 153854 514658
rect 153234 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 153854 514574
rect 153234 478894 153854 514338
rect 153234 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 153854 478894
rect 153234 478574 153854 478658
rect 153234 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 153854 478574
rect 153234 442894 153854 478338
rect 153234 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 153854 442894
rect 153234 442574 153854 442658
rect 153234 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 153854 442574
rect 153234 406894 153854 442338
rect 153234 406658 153266 406894
rect 153502 406658 153586 406894
rect 153822 406658 153854 406894
rect 153234 406574 153854 406658
rect 153234 406338 153266 406574
rect 153502 406338 153586 406574
rect 153822 406338 153854 406574
rect 153234 370894 153854 406338
rect 153234 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 153854 370894
rect 153234 370574 153854 370658
rect 153234 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 153854 370574
rect 153234 334894 153854 370338
rect 153234 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 153854 334894
rect 153234 334574 153854 334658
rect 153234 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 153854 334574
rect 153234 298894 153854 334338
rect 153234 298658 153266 298894
rect 153502 298658 153586 298894
rect 153822 298658 153854 298894
rect 153234 298574 153854 298658
rect 153234 298338 153266 298574
rect 153502 298338 153586 298574
rect 153822 298338 153854 298574
rect 153234 262894 153854 298338
rect 153234 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 153854 262894
rect 153234 262574 153854 262658
rect 153234 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 153854 262574
rect 153234 226894 153854 262338
rect 153234 226658 153266 226894
rect 153502 226658 153586 226894
rect 153822 226658 153854 226894
rect 153234 226574 153854 226658
rect 153234 226338 153266 226574
rect 153502 226338 153586 226574
rect 153822 226338 153854 226574
rect 153234 190894 153854 226338
rect 153234 190658 153266 190894
rect 153502 190658 153586 190894
rect 153822 190658 153854 190894
rect 153234 190574 153854 190658
rect 153234 190338 153266 190574
rect 153502 190338 153586 190574
rect 153822 190338 153854 190574
rect 153234 154894 153854 190338
rect 153234 154658 153266 154894
rect 153502 154658 153586 154894
rect 153822 154658 153854 154894
rect 153234 154574 153854 154658
rect 153234 154338 153266 154574
rect 153502 154338 153586 154574
rect 153822 154338 153854 154574
rect 153234 118894 153854 154338
rect 153234 118658 153266 118894
rect 153502 118658 153586 118894
rect 153822 118658 153854 118894
rect 153234 118574 153854 118658
rect 153234 118338 153266 118574
rect 153502 118338 153586 118574
rect 153822 118338 153854 118574
rect 153234 82894 153854 118338
rect 153234 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 153854 82894
rect 153234 82574 153854 82658
rect 153234 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 153854 82574
rect 153234 46894 153854 82338
rect 153234 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 153854 46894
rect 153234 46574 153854 46658
rect 153234 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 153854 46574
rect 153234 10894 153854 46338
rect 153234 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 153854 10894
rect 153234 10574 153854 10658
rect 153234 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 153854 10574
rect 153234 -4186 153854 10338
rect 153234 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 153854 -4186
rect 153234 -4506 153854 -4422
rect 153234 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 153854 -4506
rect 153234 -5734 153854 -4742
rect 156954 698614 157574 710042
rect 174954 711558 175574 711590
rect 174954 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 175574 711558
rect 174954 711238 175574 711322
rect 174954 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 175574 711238
rect 171234 709638 171854 709670
rect 171234 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 171854 709638
rect 171234 709318 171854 709402
rect 171234 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 171854 709318
rect 167514 707718 168134 707750
rect 167514 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 168134 707718
rect 167514 707398 168134 707482
rect 167514 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 168134 707398
rect 156954 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 157574 698614
rect 156954 698294 157574 698378
rect 156954 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 157574 698294
rect 156954 662614 157574 698058
rect 156954 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 157574 662614
rect 156954 662294 157574 662378
rect 156954 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 157574 662294
rect 156954 626614 157574 662058
rect 156954 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 157574 626614
rect 156954 626294 157574 626378
rect 156954 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 157574 626294
rect 156954 590614 157574 626058
rect 156954 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 157574 590614
rect 156954 590294 157574 590378
rect 156954 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 157574 590294
rect 156954 554614 157574 590058
rect 156954 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 157574 554614
rect 156954 554294 157574 554378
rect 156954 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 157574 554294
rect 156954 518614 157574 554058
rect 156954 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 157574 518614
rect 156954 518294 157574 518378
rect 156954 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 157574 518294
rect 156954 482614 157574 518058
rect 156954 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 157574 482614
rect 156954 482294 157574 482378
rect 156954 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 157574 482294
rect 156954 446614 157574 482058
rect 156954 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 157574 446614
rect 156954 446294 157574 446378
rect 156954 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 157574 446294
rect 156954 410614 157574 446058
rect 156954 410378 156986 410614
rect 157222 410378 157306 410614
rect 157542 410378 157574 410614
rect 156954 410294 157574 410378
rect 156954 410058 156986 410294
rect 157222 410058 157306 410294
rect 157542 410058 157574 410294
rect 156954 374614 157574 410058
rect 156954 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 157574 374614
rect 156954 374294 157574 374378
rect 156954 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 157574 374294
rect 156954 338614 157574 374058
rect 156954 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 157574 338614
rect 156954 338294 157574 338378
rect 156954 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 157574 338294
rect 156954 302614 157574 338058
rect 156954 302378 156986 302614
rect 157222 302378 157306 302614
rect 157542 302378 157574 302614
rect 156954 302294 157574 302378
rect 156954 302058 156986 302294
rect 157222 302058 157306 302294
rect 157542 302058 157574 302294
rect 156954 266614 157574 302058
rect 156954 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 157574 266614
rect 156954 266294 157574 266378
rect 156954 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 157574 266294
rect 156954 230614 157574 266058
rect 156954 230378 156986 230614
rect 157222 230378 157306 230614
rect 157542 230378 157574 230614
rect 156954 230294 157574 230378
rect 156954 230058 156986 230294
rect 157222 230058 157306 230294
rect 157542 230058 157574 230294
rect 156954 194614 157574 230058
rect 156954 194378 156986 194614
rect 157222 194378 157306 194614
rect 157542 194378 157574 194614
rect 156954 194294 157574 194378
rect 156954 194058 156986 194294
rect 157222 194058 157306 194294
rect 157542 194058 157574 194294
rect 156954 158614 157574 194058
rect 163794 705798 164414 705830
rect 163794 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 164414 705798
rect 163794 705478 164414 705562
rect 163794 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 164414 705478
rect 163794 669454 164414 705242
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 163794 561454 164414 596898
rect 163794 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 164414 561454
rect 163794 561134 164414 561218
rect 163794 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 164414 561134
rect 163794 525454 164414 560898
rect 163794 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 164414 525454
rect 163794 525134 164414 525218
rect 163794 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 164414 525134
rect 163794 489454 164414 524898
rect 163794 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 164414 489454
rect 163794 489134 164414 489218
rect 163794 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 164414 489134
rect 163794 453454 164414 488898
rect 163794 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 164414 453454
rect 163794 453134 164414 453218
rect 163794 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 164414 453134
rect 163794 417454 164414 452898
rect 163794 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 164414 417454
rect 163794 417134 164414 417218
rect 163794 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 164414 417134
rect 163794 381454 164414 416898
rect 163794 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 164414 381454
rect 163794 381134 164414 381218
rect 163794 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 164414 381134
rect 163794 345454 164414 380898
rect 163794 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 164414 345454
rect 163794 345134 164414 345218
rect 163794 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 164414 345134
rect 163794 309454 164414 344898
rect 163794 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 164414 309454
rect 163794 309134 164414 309218
rect 163794 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 164414 309134
rect 163794 273454 164414 308898
rect 163794 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 164414 273454
rect 163794 273134 164414 273218
rect 163794 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 164414 273134
rect 163794 237454 164414 272898
rect 163794 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 164414 237454
rect 163794 237134 164414 237218
rect 163794 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 164414 237134
rect 163794 201454 164414 236898
rect 163794 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 164414 201454
rect 163794 201134 164414 201218
rect 163794 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 164414 201134
rect 163794 192000 164414 200898
rect 167514 673174 168134 707162
rect 167514 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 168134 673174
rect 167514 672854 168134 672938
rect 167514 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 168134 672854
rect 167514 637174 168134 672618
rect 167514 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 168134 637174
rect 167514 636854 168134 636938
rect 167514 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 168134 636854
rect 167514 601174 168134 636618
rect 167514 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 168134 601174
rect 167514 600854 168134 600938
rect 167514 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 168134 600854
rect 167514 565174 168134 600618
rect 167514 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 168134 565174
rect 167514 564854 168134 564938
rect 167514 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 168134 564854
rect 167514 529174 168134 564618
rect 167514 528938 167546 529174
rect 167782 528938 167866 529174
rect 168102 528938 168134 529174
rect 167514 528854 168134 528938
rect 167514 528618 167546 528854
rect 167782 528618 167866 528854
rect 168102 528618 168134 528854
rect 167514 493174 168134 528618
rect 167514 492938 167546 493174
rect 167782 492938 167866 493174
rect 168102 492938 168134 493174
rect 167514 492854 168134 492938
rect 167514 492618 167546 492854
rect 167782 492618 167866 492854
rect 168102 492618 168134 492854
rect 167514 457174 168134 492618
rect 167514 456938 167546 457174
rect 167782 456938 167866 457174
rect 168102 456938 168134 457174
rect 167514 456854 168134 456938
rect 167514 456618 167546 456854
rect 167782 456618 167866 456854
rect 168102 456618 168134 456854
rect 167514 421174 168134 456618
rect 167514 420938 167546 421174
rect 167782 420938 167866 421174
rect 168102 420938 168134 421174
rect 167514 420854 168134 420938
rect 167514 420618 167546 420854
rect 167782 420618 167866 420854
rect 168102 420618 168134 420854
rect 167514 385174 168134 420618
rect 167514 384938 167546 385174
rect 167782 384938 167866 385174
rect 168102 384938 168134 385174
rect 167514 384854 168134 384938
rect 167514 384618 167546 384854
rect 167782 384618 167866 384854
rect 168102 384618 168134 384854
rect 167514 349174 168134 384618
rect 167514 348938 167546 349174
rect 167782 348938 167866 349174
rect 168102 348938 168134 349174
rect 167514 348854 168134 348938
rect 167514 348618 167546 348854
rect 167782 348618 167866 348854
rect 168102 348618 168134 348854
rect 167514 313174 168134 348618
rect 167514 312938 167546 313174
rect 167782 312938 167866 313174
rect 168102 312938 168134 313174
rect 167514 312854 168134 312938
rect 167514 312618 167546 312854
rect 167782 312618 167866 312854
rect 168102 312618 168134 312854
rect 167514 277174 168134 312618
rect 167514 276938 167546 277174
rect 167782 276938 167866 277174
rect 168102 276938 168134 277174
rect 167514 276854 168134 276938
rect 167514 276618 167546 276854
rect 167782 276618 167866 276854
rect 168102 276618 168134 276854
rect 167514 241174 168134 276618
rect 167514 240938 167546 241174
rect 167782 240938 167866 241174
rect 168102 240938 168134 241174
rect 167514 240854 168134 240938
rect 167514 240618 167546 240854
rect 167782 240618 167866 240854
rect 168102 240618 168134 240854
rect 167514 205174 168134 240618
rect 167514 204938 167546 205174
rect 167782 204938 167866 205174
rect 168102 204938 168134 205174
rect 167514 204854 168134 204938
rect 167514 204618 167546 204854
rect 167782 204618 167866 204854
rect 168102 204618 168134 204854
rect 167514 192000 168134 204618
rect 171234 676894 171854 709082
rect 171234 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 171854 676894
rect 171234 676574 171854 676658
rect 171234 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 171854 676574
rect 171234 640894 171854 676338
rect 171234 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 171854 640894
rect 171234 640574 171854 640658
rect 171234 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 171854 640574
rect 171234 604894 171854 640338
rect 171234 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 171854 604894
rect 171234 604574 171854 604658
rect 171234 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 171854 604574
rect 171234 568894 171854 604338
rect 171234 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 171854 568894
rect 171234 568574 171854 568658
rect 171234 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 171854 568574
rect 171234 532894 171854 568338
rect 171234 532658 171266 532894
rect 171502 532658 171586 532894
rect 171822 532658 171854 532894
rect 171234 532574 171854 532658
rect 171234 532338 171266 532574
rect 171502 532338 171586 532574
rect 171822 532338 171854 532574
rect 171234 496894 171854 532338
rect 171234 496658 171266 496894
rect 171502 496658 171586 496894
rect 171822 496658 171854 496894
rect 171234 496574 171854 496658
rect 171234 496338 171266 496574
rect 171502 496338 171586 496574
rect 171822 496338 171854 496574
rect 171234 460894 171854 496338
rect 171234 460658 171266 460894
rect 171502 460658 171586 460894
rect 171822 460658 171854 460894
rect 171234 460574 171854 460658
rect 171234 460338 171266 460574
rect 171502 460338 171586 460574
rect 171822 460338 171854 460574
rect 171234 424894 171854 460338
rect 171234 424658 171266 424894
rect 171502 424658 171586 424894
rect 171822 424658 171854 424894
rect 171234 424574 171854 424658
rect 171234 424338 171266 424574
rect 171502 424338 171586 424574
rect 171822 424338 171854 424574
rect 171234 388894 171854 424338
rect 171234 388658 171266 388894
rect 171502 388658 171586 388894
rect 171822 388658 171854 388894
rect 171234 388574 171854 388658
rect 171234 388338 171266 388574
rect 171502 388338 171586 388574
rect 171822 388338 171854 388574
rect 171234 352894 171854 388338
rect 171234 352658 171266 352894
rect 171502 352658 171586 352894
rect 171822 352658 171854 352894
rect 171234 352574 171854 352658
rect 171234 352338 171266 352574
rect 171502 352338 171586 352574
rect 171822 352338 171854 352574
rect 171234 316894 171854 352338
rect 171234 316658 171266 316894
rect 171502 316658 171586 316894
rect 171822 316658 171854 316894
rect 171234 316574 171854 316658
rect 171234 316338 171266 316574
rect 171502 316338 171586 316574
rect 171822 316338 171854 316574
rect 171234 280894 171854 316338
rect 171234 280658 171266 280894
rect 171502 280658 171586 280894
rect 171822 280658 171854 280894
rect 171234 280574 171854 280658
rect 171234 280338 171266 280574
rect 171502 280338 171586 280574
rect 171822 280338 171854 280574
rect 171234 244894 171854 280338
rect 171234 244658 171266 244894
rect 171502 244658 171586 244894
rect 171822 244658 171854 244894
rect 171234 244574 171854 244658
rect 171234 244338 171266 244574
rect 171502 244338 171586 244574
rect 171822 244338 171854 244574
rect 171234 208894 171854 244338
rect 171234 208658 171266 208894
rect 171502 208658 171586 208894
rect 171822 208658 171854 208894
rect 171234 208574 171854 208658
rect 171234 208338 171266 208574
rect 171502 208338 171586 208574
rect 171822 208338 171854 208574
rect 171234 192000 171854 208338
rect 174954 680614 175574 711002
rect 192954 710598 193574 711590
rect 192954 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 193574 710598
rect 192954 710278 193574 710362
rect 192954 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 193574 710278
rect 189234 708678 189854 709670
rect 189234 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 189854 708678
rect 189234 708358 189854 708442
rect 189234 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 189854 708358
rect 185514 706758 186134 707750
rect 185514 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 186134 706758
rect 185514 706438 186134 706522
rect 185514 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 186134 706438
rect 174954 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 175574 680614
rect 174954 680294 175574 680378
rect 174954 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 175574 680294
rect 174954 644614 175574 680058
rect 174954 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 175574 644614
rect 174954 644294 175574 644378
rect 174954 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 175574 644294
rect 174954 608614 175574 644058
rect 174954 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 175574 608614
rect 174954 608294 175574 608378
rect 174954 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 175574 608294
rect 174954 572614 175574 608058
rect 174954 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 175574 572614
rect 174954 572294 175574 572378
rect 174954 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 175574 572294
rect 174954 536614 175574 572058
rect 174954 536378 174986 536614
rect 175222 536378 175306 536614
rect 175542 536378 175574 536614
rect 174954 536294 175574 536378
rect 174954 536058 174986 536294
rect 175222 536058 175306 536294
rect 175542 536058 175574 536294
rect 174954 500614 175574 536058
rect 174954 500378 174986 500614
rect 175222 500378 175306 500614
rect 175542 500378 175574 500614
rect 174954 500294 175574 500378
rect 174954 500058 174986 500294
rect 175222 500058 175306 500294
rect 175542 500058 175574 500294
rect 174954 464614 175574 500058
rect 174954 464378 174986 464614
rect 175222 464378 175306 464614
rect 175542 464378 175574 464614
rect 174954 464294 175574 464378
rect 174954 464058 174986 464294
rect 175222 464058 175306 464294
rect 175542 464058 175574 464294
rect 174954 428614 175574 464058
rect 174954 428378 174986 428614
rect 175222 428378 175306 428614
rect 175542 428378 175574 428614
rect 174954 428294 175574 428378
rect 174954 428058 174986 428294
rect 175222 428058 175306 428294
rect 175542 428058 175574 428294
rect 174954 392614 175574 428058
rect 174954 392378 174986 392614
rect 175222 392378 175306 392614
rect 175542 392378 175574 392614
rect 174954 392294 175574 392378
rect 174954 392058 174986 392294
rect 175222 392058 175306 392294
rect 175542 392058 175574 392294
rect 174954 356614 175574 392058
rect 174954 356378 174986 356614
rect 175222 356378 175306 356614
rect 175542 356378 175574 356614
rect 174954 356294 175574 356378
rect 174954 356058 174986 356294
rect 175222 356058 175306 356294
rect 175542 356058 175574 356294
rect 174954 320614 175574 356058
rect 174954 320378 174986 320614
rect 175222 320378 175306 320614
rect 175542 320378 175574 320614
rect 174954 320294 175574 320378
rect 174954 320058 174986 320294
rect 175222 320058 175306 320294
rect 175542 320058 175574 320294
rect 174954 284614 175574 320058
rect 174954 284378 174986 284614
rect 175222 284378 175306 284614
rect 175542 284378 175574 284614
rect 174954 284294 175574 284378
rect 174954 284058 174986 284294
rect 175222 284058 175306 284294
rect 175542 284058 175574 284294
rect 174954 248614 175574 284058
rect 174954 248378 174986 248614
rect 175222 248378 175306 248614
rect 175542 248378 175574 248614
rect 174954 248294 175574 248378
rect 174954 248058 174986 248294
rect 175222 248058 175306 248294
rect 175542 248058 175574 248294
rect 174954 212614 175574 248058
rect 174954 212378 174986 212614
rect 175222 212378 175306 212614
rect 175542 212378 175574 212614
rect 174954 212294 175574 212378
rect 174954 212058 174986 212294
rect 175222 212058 175306 212294
rect 175542 212058 175574 212294
rect 162243 183454 162563 183486
rect 162243 183218 162285 183454
rect 162521 183218 162563 183454
rect 162243 183134 162563 183218
rect 162243 182898 162285 183134
rect 162521 182898 162563 183134
rect 162243 182866 162563 182898
rect 164840 183454 165160 183486
rect 164840 183218 164882 183454
rect 165118 183218 165160 183454
rect 164840 183134 165160 183218
rect 164840 182898 164882 183134
rect 165118 182898 165160 183134
rect 164840 182866 165160 182898
rect 167437 183454 167757 183486
rect 167437 183218 167479 183454
rect 167715 183218 167757 183454
rect 167437 183134 167757 183218
rect 167437 182898 167479 183134
rect 167715 182898 167757 183134
rect 167437 182866 167757 182898
rect 174954 176614 175574 212058
rect 174954 176378 174986 176614
rect 175222 176378 175306 176614
rect 175542 176378 175574 176614
rect 174954 176294 175574 176378
rect 174954 176058 174986 176294
rect 175222 176058 175306 176294
rect 175542 176058 175574 176294
rect 163541 165454 163861 165486
rect 163541 165218 163583 165454
rect 163819 165218 163861 165454
rect 163541 165134 163861 165218
rect 163541 164898 163583 165134
rect 163819 164898 163861 165134
rect 163541 164866 163861 164898
rect 166138 165454 166458 165486
rect 166138 165218 166180 165454
rect 166416 165218 166458 165454
rect 166138 165134 166458 165218
rect 166138 164898 166180 165134
rect 166416 164898 166458 165134
rect 166138 164866 166458 164898
rect 156954 158378 156986 158614
rect 157222 158378 157306 158614
rect 157542 158378 157574 158614
rect 156954 158294 157574 158378
rect 156954 158058 156986 158294
rect 157222 158058 157306 158294
rect 157542 158058 157574 158294
rect 156954 122614 157574 158058
rect 163794 156000 164414 158000
rect 167514 156000 168134 158000
rect 171234 156000 171854 158000
rect 162243 147454 162563 147486
rect 162243 147218 162285 147454
rect 162521 147218 162563 147454
rect 162243 147134 162563 147218
rect 162243 146898 162285 147134
rect 162521 146898 162563 147134
rect 162243 146866 162563 146898
rect 164840 147454 165160 147486
rect 164840 147218 164882 147454
rect 165118 147218 165160 147454
rect 164840 147134 165160 147218
rect 164840 146898 164882 147134
rect 165118 146898 165160 147134
rect 164840 146866 165160 146898
rect 167437 147454 167757 147486
rect 167437 147218 167479 147454
rect 167715 147218 167757 147454
rect 167437 147134 167757 147218
rect 167437 146898 167479 147134
rect 167715 146898 167757 147134
rect 167437 146866 167757 146898
rect 174954 140614 175574 176058
rect 174954 140378 174986 140614
rect 175222 140378 175306 140614
rect 175542 140378 175574 140614
rect 174954 140294 175574 140378
rect 174954 140058 174986 140294
rect 175222 140058 175306 140294
rect 175542 140058 175574 140294
rect 163541 129454 163861 129486
rect 163541 129218 163583 129454
rect 163819 129218 163861 129454
rect 163541 129134 163861 129218
rect 163541 128898 163583 129134
rect 163819 128898 163861 129134
rect 163541 128866 163861 128898
rect 166138 129454 166458 129486
rect 166138 129218 166180 129454
rect 166416 129218 166458 129454
rect 166138 129134 166458 129218
rect 166138 128898 166180 129134
rect 166416 128898 166458 129134
rect 166138 128866 166458 128898
rect 156954 122378 156986 122614
rect 157222 122378 157306 122614
rect 157542 122378 157574 122614
rect 156954 122294 157574 122378
rect 156954 122058 156986 122294
rect 157222 122058 157306 122294
rect 157542 122058 157574 122294
rect 156954 86614 157574 122058
rect 156954 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 157574 86614
rect 156954 86294 157574 86378
rect 156954 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 157574 86294
rect 156954 50614 157574 86058
rect 156954 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 157574 50614
rect 156954 50294 157574 50378
rect 156954 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 157574 50294
rect 156954 14614 157574 50058
rect 156954 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 157574 14614
rect 156954 14294 157574 14378
rect 156954 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 157574 14294
rect 138954 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 139574 -7066
rect 138954 -7386 139574 -7302
rect 138954 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 139574 -7386
rect 138954 -7654 139574 -7622
rect 156954 -6106 157574 14058
rect 163794 93454 164414 122000
rect 163794 93218 163826 93454
rect 164062 93218 164146 93454
rect 164382 93218 164414 93454
rect 163794 93134 164414 93218
rect 163794 92898 163826 93134
rect 164062 92898 164146 93134
rect 164382 92898 164414 93134
rect 163794 57454 164414 92898
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -1306 164414 20898
rect 163794 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 164414 -1306
rect 163794 -1626 164414 -1542
rect 163794 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 164414 -1626
rect 163794 -1894 164414 -1862
rect 167514 97174 168134 122000
rect 167514 96938 167546 97174
rect 167782 96938 167866 97174
rect 168102 96938 168134 97174
rect 167514 96854 168134 96938
rect 167514 96618 167546 96854
rect 167782 96618 167866 96854
rect 168102 96618 168134 96854
rect 167514 61174 168134 96618
rect 167514 60938 167546 61174
rect 167782 60938 167866 61174
rect 168102 60938 168134 61174
rect 167514 60854 168134 60938
rect 167514 60618 167546 60854
rect 167782 60618 167866 60854
rect 168102 60618 168134 60854
rect 167514 25174 168134 60618
rect 167514 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 168134 25174
rect 167514 24854 168134 24938
rect 167514 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 168134 24854
rect 167514 -3226 168134 24618
rect 167514 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 168134 -3226
rect 167514 -3546 168134 -3462
rect 167514 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 168134 -3546
rect 167514 -3814 168134 -3782
rect 171234 100894 171854 122000
rect 171234 100658 171266 100894
rect 171502 100658 171586 100894
rect 171822 100658 171854 100894
rect 171234 100574 171854 100658
rect 171234 100338 171266 100574
rect 171502 100338 171586 100574
rect 171822 100338 171854 100574
rect 171234 64894 171854 100338
rect 171234 64658 171266 64894
rect 171502 64658 171586 64894
rect 171822 64658 171854 64894
rect 171234 64574 171854 64658
rect 171234 64338 171266 64574
rect 171502 64338 171586 64574
rect 171822 64338 171854 64574
rect 171234 28894 171854 64338
rect 171234 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 171854 28894
rect 171234 28574 171854 28658
rect 171234 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 171854 28574
rect 171234 -5146 171854 28338
rect 171234 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 171854 -5146
rect 171234 -5466 171854 -5382
rect 171234 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 171854 -5466
rect 171234 -5734 171854 -5702
rect 174954 104614 175574 140058
rect 174954 104378 174986 104614
rect 175222 104378 175306 104614
rect 175542 104378 175574 104614
rect 174954 104294 175574 104378
rect 174954 104058 174986 104294
rect 175222 104058 175306 104294
rect 175542 104058 175574 104294
rect 174954 68614 175574 104058
rect 174954 68378 174986 68614
rect 175222 68378 175306 68614
rect 175542 68378 175574 68614
rect 174954 68294 175574 68378
rect 174954 68058 174986 68294
rect 175222 68058 175306 68294
rect 175542 68058 175574 68294
rect 174954 32614 175574 68058
rect 174954 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 175574 32614
rect 174954 32294 175574 32378
rect 174954 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 175574 32294
rect 156954 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 157574 -6106
rect 156954 -6426 157574 -6342
rect 156954 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 157574 -6426
rect 156954 -7654 157574 -6662
rect 174954 -7066 175574 32058
rect 181794 704838 182414 705830
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 543454 182414 578898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 507454 182414 542898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 181794 471454 182414 506898
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 181794 435454 182414 470898
rect 181794 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 182414 435454
rect 181794 435134 182414 435218
rect 181794 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 182414 435134
rect 181794 399454 182414 434898
rect 181794 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 182414 399454
rect 181794 399134 182414 399218
rect 181794 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 182414 399134
rect 181794 363454 182414 398898
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 181794 327454 182414 362898
rect 181794 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 182414 327454
rect 181794 327134 182414 327218
rect 181794 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 182414 327134
rect 181794 291454 182414 326898
rect 181794 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 182414 291454
rect 181794 291134 182414 291218
rect 181794 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 182414 291134
rect 181794 255454 182414 290898
rect 181794 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 182414 255454
rect 181794 255134 182414 255218
rect 181794 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 182414 255134
rect 181794 219454 182414 254898
rect 181794 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 182414 219454
rect 181794 219134 182414 219218
rect 181794 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 182414 219134
rect 181794 183454 182414 218898
rect 181794 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 182414 183454
rect 181794 183134 182414 183218
rect 181794 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 182414 183134
rect 181794 147454 182414 182898
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 111454 182414 146898
rect 181794 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 182414 111454
rect 181794 111134 182414 111218
rect 181794 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 182414 111134
rect 181794 75454 182414 110898
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 181794 39454 182414 74898
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -1894 182414 -902
rect 185514 691174 186134 706202
rect 185514 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 186134 691174
rect 185514 690854 186134 690938
rect 185514 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 186134 690854
rect 185514 655174 186134 690618
rect 185514 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 186134 655174
rect 185514 654854 186134 654938
rect 185514 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 186134 654854
rect 185514 619174 186134 654618
rect 185514 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 186134 619174
rect 185514 618854 186134 618938
rect 185514 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 186134 618854
rect 185514 583174 186134 618618
rect 185514 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 186134 583174
rect 185514 582854 186134 582938
rect 185514 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 186134 582854
rect 185514 547174 186134 582618
rect 185514 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 186134 547174
rect 185514 546854 186134 546938
rect 185514 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 186134 546854
rect 185514 511174 186134 546618
rect 185514 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 186134 511174
rect 185514 510854 186134 510938
rect 185514 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 186134 510854
rect 185514 475174 186134 510618
rect 185514 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 186134 475174
rect 185514 474854 186134 474938
rect 185514 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 186134 474854
rect 185514 439174 186134 474618
rect 185514 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 186134 439174
rect 185514 438854 186134 438938
rect 185514 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 186134 438854
rect 185514 403174 186134 438618
rect 185514 402938 185546 403174
rect 185782 402938 185866 403174
rect 186102 402938 186134 403174
rect 185514 402854 186134 402938
rect 185514 402618 185546 402854
rect 185782 402618 185866 402854
rect 186102 402618 186134 402854
rect 185514 367174 186134 402618
rect 185514 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 186134 367174
rect 185514 366854 186134 366938
rect 185514 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 186134 366854
rect 185514 331174 186134 366618
rect 185514 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 186134 331174
rect 185514 330854 186134 330938
rect 185514 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 186134 330854
rect 185514 295174 186134 330618
rect 185514 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 186134 295174
rect 185514 294854 186134 294938
rect 185514 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 186134 294854
rect 185514 259174 186134 294618
rect 185514 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 186134 259174
rect 185514 258854 186134 258938
rect 185514 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 186134 258854
rect 185514 223174 186134 258618
rect 185514 222938 185546 223174
rect 185782 222938 185866 223174
rect 186102 222938 186134 223174
rect 185514 222854 186134 222938
rect 185514 222618 185546 222854
rect 185782 222618 185866 222854
rect 186102 222618 186134 222854
rect 185514 187174 186134 222618
rect 185514 186938 185546 187174
rect 185782 186938 185866 187174
rect 186102 186938 186134 187174
rect 185514 186854 186134 186938
rect 185514 186618 185546 186854
rect 185782 186618 185866 186854
rect 186102 186618 186134 186854
rect 185514 151174 186134 186618
rect 185514 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 186134 151174
rect 185514 150854 186134 150938
rect 185514 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 186134 150854
rect 185514 115174 186134 150618
rect 185514 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 186134 115174
rect 185514 114854 186134 114938
rect 185514 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 186134 114854
rect 185514 79174 186134 114618
rect 185514 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 186134 79174
rect 185514 78854 186134 78938
rect 185514 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 186134 78854
rect 185514 43174 186134 78618
rect 185514 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 186134 43174
rect 185514 42854 186134 42938
rect 185514 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 186134 42854
rect 185514 7174 186134 42618
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 185514 -2266 186134 6618
rect 185514 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 186134 -2266
rect 185514 -2586 186134 -2502
rect 185514 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 186134 -2586
rect 185514 -3814 186134 -2822
rect 189234 694894 189854 708122
rect 189234 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 189854 694894
rect 189234 694574 189854 694658
rect 189234 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 189854 694574
rect 189234 658894 189854 694338
rect 189234 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 189854 658894
rect 189234 658574 189854 658658
rect 189234 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 189854 658574
rect 189234 622894 189854 658338
rect 189234 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 189854 622894
rect 189234 622574 189854 622658
rect 189234 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 189854 622574
rect 189234 586894 189854 622338
rect 189234 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 189854 586894
rect 189234 586574 189854 586658
rect 189234 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 189854 586574
rect 189234 550894 189854 586338
rect 189234 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 189854 550894
rect 189234 550574 189854 550658
rect 189234 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 189854 550574
rect 189234 514894 189854 550338
rect 189234 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 189854 514894
rect 189234 514574 189854 514658
rect 189234 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 189854 514574
rect 189234 478894 189854 514338
rect 189234 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 189854 478894
rect 189234 478574 189854 478658
rect 189234 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 189854 478574
rect 189234 442894 189854 478338
rect 189234 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 189854 442894
rect 189234 442574 189854 442658
rect 189234 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 189854 442574
rect 189234 406894 189854 442338
rect 189234 406658 189266 406894
rect 189502 406658 189586 406894
rect 189822 406658 189854 406894
rect 189234 406574 189854 406658
rect 189234 406338 189266 406574
rect 189502 406338 189586 406574
rect 189822 406338 189854 406574
rect 189234 370894 189854 406338
rect 189234 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 189854 370894
rect 189234 370574 189854 370658
rect 189234 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 189854 370574
rect 189234 334894 189854 370338
rect 189234 334658 189266 334894
rect 189502 334658 189586 334894
rect 189822 334658 189854 334894
rect 189234 334574 189854 334658
rect 189234 334338 189266 334574
rect 189502 334338 189586 334574
rect 189822 334338 189854 334574
rect 189234 298894 189854 334338
rect 189234 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 189854 298894
rect 189234 298574 189854 298658
rect 189234 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 189854 298574
rect 189234 262894 189854 298338
rect 189234 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 189854 262894
rect 189234 262574 189854 262658
rect 189234 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 189854 262574
rect 189234 226894 189854 262338
rect 189234 226658 189266 226894
rect 189502 226658 189586 226894
rect 189822 226658 189854 226894
rect 189234 226574 189854 226658
rect 189234 226338 189266 226574
rect 189502 226338 189586 226574
rect 189822 226338 189854 226574
rect 189234 190894 189854 226338
rect 189234 190658 189266 190894
rect 189502 190658 189586 190894
rect 189822 190658 189854 190894
rect 189234 190574 189854 190658
rect 189234 190338 189266 190574
rect 189502 190338 189586 190574
rect 189822 190338 189854 190574
rect 189234 154894 189854 190338
rect 189234 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 189854 154894
rect 189234 154574 189854 154658
rect 189234 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 189854 154574
rect 189234 118894 189854 154338
rect 189234 118658 189266 118894
rect 189502 118658 189586 118894
rect 189822 118658 189854 118894
rect 189234 118574 189854 118658
rect 189234 118338 189266 118574
rect 189502 118338 189586 118574
rect 189822 118338 189854 118574
rect 189234 82894 189854 118338
rect 189234 82658 189266 82894
rect 189502 82658 189586 82894
rect 189822 82658 189854 82894
rect 189234 82574 189854 82658
rect 189234 82338 189266 82574
rect 189502 82338 189586 82574
rect 189822 82338 189854 82574
rect 189234 46894 189854 82338
rect 189234 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 189854 46894
rect 189234 46574 189854 46658
rect 189234 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 189854 46574
rect 189234 10894 189854 46338
rect 189234 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 189854 10894
rect 189234 10574 189854 10658
rect 189234 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 189854 10574
rect 189234 -4186 189854 10338
rect 189234 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 189854 -4186
rect 189234 -4506 189854 -4422
rect 189234 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 189854 -4506
rect 189234 -5734 189854 -4742
rect 192954 698614 193574 710042
rect 210954 711558 211574 711590
rect 210954 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 211574 711558
rect 210954 711238 211574 711322
rect 210954 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 211574 711238
rect 207234 709638 207854 709670
rect 207234 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 207854 709638
rect 207234 709318 207854 709402
rect 207234 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 207854 709318
rect 203514 707718 204134 707750
rect 203514 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 204134 707718
rect 203514 707398 204134 707482
rect 203514 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 204134 707398
rect 192954 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 193574 698614
rect 192954 698294 193574 698378
rect 192954 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 193574 698294
rect 192954 662614 193574 698058
rect 192954 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 193574 662614
rect 192954 662294 193574 662378
rect 192954 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 193574 662294
rect 192954 626614 193574 662058
rect 192954 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 193574 626614
rect 192954 626294 193574 626378
rect 192954 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 193574 626294
rect 192954 590614 193574 626058
rect 192954 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 193574 590614
rect 192954 590294 193574 590378
rect 192954 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 193574 590294
rect 192954 554614 193574 590058
rect 192954 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 193574 554614
rect 192954 554294 193574 554378
rect 192954 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 193574 554294
rect 192954 518614 193574 554058
rect 192954 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 193574 518614
rect 192954 518294 193574 518378
rect 192954 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 193574 518294
rect 192954 482614 193574 518058
rect 192954 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 193574 482614
rect 192954 482294 193574 482378
rect 192954 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 193574 482294
rect 192954 446614 193574 482058
rect 192954 446378 192986 446614
rect 193222 446378 193306 446614
rect 193542 446378 193574 446614
rect 192954 446294 193574 446378
rect 192954 446058 192986 446294
rect 193222 446058 193306 446294
rect 193542 446058 193574 446294
rect 192954 410614 193574 446058
rect 192954 410378 192986 410614
rect 193222 410378 193306 410614
rect 193542 410378 193574 410614
rect 192954 410294 193574 410378
rect 192954 410058 192986 410294
rect 193222 410058 193306 410294
rect 193542 410058 193574 410294
rect 192954 374614 193574 410058
rect 192954 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 193574 374614
rect 192954 374294 193574 374378
rect 192954 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 193574 374294
rect 192954 338614 193574 374058
rect 192954 338378 192986 338614
rect 193222 338378 193306 338614
rect 193542 338378 193574 338614
rect 192954 338294 193574 338378
rect 192954 338058 192986 338294
rect 193222 338058 193306 338294
rect 193542 338058 193574 338294
rect 192954 302614 193574 338058
rect 192954 302378 192986 302614
rect 193222 302378 193306 302614
rect 193542 302378 193574 302614
rect 192954 302294 193574 302378
rect 192954 302058 192986 302294
rect 193222 302058 193306 302294
rect 193542 302058 193574 302294
rect 192954 266614 193574 302058
rect 199794 705798 200414 705830
rect 199794 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 200414 705798
rect 199794 705478 200414 705562
rect 199794 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 200414 705478
rect 199794 669454 200414 705242
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 561454 200414 596898
rect 199794 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 200414 561454
rect 199794 561134 200414 561218
rect 199794 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 200414 561134
rect 199794 525454 200414 560898
rect 199794 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 200414 525454
rect 199794 525134 200414 525218
rect 199794 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 200414 525134
rect 199794 489454 200414 524898
rect 199794 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 200414 489454
rect 199794 489134 200414 489218
rect 199794 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 200414 489134
rect 199794 453454 200414 488898
rect 199794 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 200414 453454
rect 199794 453134 200414 453218
rect 199794 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 200414 453134
rect 199794 417454 200414 452898
rect 199794 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 200414 417454
rect 199794 417134 200414 417218
rect 199794 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 200414 417134
rect 199794 381454 200414 416898
rect 199794 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 200414 381454
rect 199794 381134 200414 381218
rect 199794 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 200414 381134
rect 199794 345454 200414 380898
rect 199794 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 200414 345454
rect 199794 345134 200414 345218
rect 199794 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 200414 345134
rect 199794 309454 200414 344898
rect 199794 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 200414 309454
rect 199794 309134 200414 309218
rect 199794 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 200414 309134
rect 199794 302000 200414 308898
rect 203514 673174 204134 707162
rect 203514 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 204134 673174
rect 203514 672854 204134 672938
rect 203514 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 204134 672854
rect 203514 637174 204134 672618
rect 203514 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 204134 637174
rect 203514 636854 204134 636938
rect 203514 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 204134 636854
rect 203514 601174 204134 636618
rect 203514 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 204134 601174
rect 203514 600854 204134 600938
rect 203514 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 204134 600854
rect 203514 565174 204134 600618
rect 203514 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 204134 565174
rect 203514 564854 204134 564938
rect 203514 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 204134 564854
rect 203514 529174 204134 564618
rect 203514 528938 203546 529174
rect 203782 528938 203866 529174
rect 204102 528938 204134 529174
rect 203514 528854 204134 528938
rect 203514 528618 203546 528854
rect 203782 528618 203866 528854
rect 204102 528618 204134 528854
rect 203514 493174 204134 528618
rect 203514 492938 203546 493174
rect 203782 492938 203866 493174
rect 204102 492938 204134 493174
rect 203514 492854 204134 492938
rect 203514 492618 203546 492854
rect 203782 492618 203866 492854
rect 204102 492618 204134 492854
rect 203514 457174 204134 492618
rect 203514 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 204134 457174
rect 203514 456854 204134 456938
rect 203514 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 204134 456854
rect 203514 421174 204134 456618
rect 203514 420938 203546 421174
rect 203782 420938 203866 421174
rect 204102 420938 204134 421174
rect 203514 420854 204134 420938
rect 203514 420618 203546 420854
rect 203782 420618 203866 420854
rect 204102 420618 204134 420854
rect 203514 385174 204134 420618
rect 203514 384938 203546 385174
rect 203782 384938 203866 385174
rect 204102 384938 204134 385174
rect 203514 384854 204134 384938
rect 203514 384618 203546 384854
rect 203782 384618 203866 384854
rect 204102 384618 204134 384854
rect 203514 349174 204134 384618
rect 203514 348938 203546 349174
rect 203782 348938 203866 349174
rect 204102 348938 204134 349174
rect 203514 348854 204134 348938
rect 203514 348618 203546 348854
rect 203782 348618 203866 348854
rect 204102 348618 204134 348854
rect 203514 313174 204134 348618
rect 203514 312938 203546 313174
rect 203782 312938 203866 313174
rect 204102 312938 204134 313174
rect 203514 312854 204134 312938
rect 203514 312618 203546 312854
rect 203782 312618 203866 312854
rect 204102 312618 204134 312854
rect 203514 302000 204134 312618
rect 207234 676894 207854 709082
rect 207234 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 207854 676894
rect 207234 676574 207854 676658
rect 207234 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 207854 676574
rect 207234 640894 207854 676338
rect 207234 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 207854 640894
rect 207234 640574 207854 640658
rect 207234 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 207854 640574
rect 207234 604894 207854 640338
rect 207234 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 207854 604894
rect 207234 604574 207854 604658
rect 207234 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 207854 604574
rect 207234 568894 207854 604338
rect 207234 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 207854 568894
rect 207234 568574 207854 568658
rect 207234 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 207854 568574
rect 207234 532894 207854 568338
rect 207234 532658 207266 532894
rect 207502 532658 207586 532894
rect 207822 532658 207854 532894
rect 207234 532574 207854 532658
rect 207234 532338 207266 532574
rect 207502 532338 207586 532574
rect 207822 532338 207854 532574
rect 207234 496894 207854 532338
rect 207234 496658 207266 496894
rect 207502 496658 207586 496894
rect 207822 496658 207854 496894
rect 207234 496574 207854 496658
rect 207234 496338 207266 496574
rect 207502 496338 207586 496574
rect 207822 496338 207854 496574
rect 207234 460894 207854 496338
rect 207234 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 207854 460894
rect 207234 460574 207854 460658
rect 207234 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 207854 460574
rect 207234 424894 207854 460338
rect 207234 424658 207266 424894
rect 207502 424658 207586 424894
rect 207822 424658 207854 424894
rect 207234 424574 207854 424658
rect 207234 424338 207266 424574
rect 207502 424338 207586 424574
rect 207822 424338 207854 424574
rect 207234 388894 207854 424338
rect 207234 388658 207266 388894
rect 207502 388658 207586 388894
rect 207822 388658 207854 388894
rect 207234 388574 207854 388658
rect 207234 388338 207266 388574
rect 207502 388338 207586 388574
rect 207822 388338 207854 388574
rect 207234 352894 207854 388338
rect 207234 352658 207266 352894
rect 207502 352658 207586 352894
rect 207822 352658 207854 352894
rect 207234 352574 207854 352658
rect 207234 352338 207266 352574
rect 207502 352338 207586 352574
rect 207822 352338 207854 352574
rect 207234 316894 207854 352338
rect 207234 316658 207266 316894
rect 207502 316658 207586 316894
rect 207822 316658 207854 316894
rect 207234 316574 207854 316658
rect 207234 316338 207266 316574
rect 207502 316338 207586 316574
rect 207822 316338 207854 316574
rect 207234 302000 207854 316338
rect 210954 680614 211574 711002
rect 228954 710598 229574 711590
rect 228954 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 229574 710598
rect 228954 710278 229574 710362
rect 228954 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 229574 710278
rect 225234 708678 225854 709670
rect 225234 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 225854 708678
rect 225234 708358 225854 708442
rect 225234 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 225854 708358
rect 221514 706758 222134 707750
rect 221514 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 222134 706758
rect 221514 706438 222134 706522
rect 221514 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 222134 706438
rect 210954 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 211574 680614
rect 210954 680294 211574 680378
rect 210954 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 211574 680294
rect 210954 644614 211574 680058
rect 210954 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 211574 644614
rect 210954 644294 211574 644378
rect 210954 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 211574 644294
rect 210954 608614 211574 644058
rect 210954 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 211574 608614
rect 210954 608294 211574 608378
rect 210954 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 211574 608294
rect 210954 572614 211574 608058
rect 210954 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 211574 572614
rect 210954 572294 211574 572378
rect 210954 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 211574 572294
rect 210954 536614 211574 572058
rect 210954 536378 210986 536614
rect 211222 536378 211306 536614
rect 211542 536378 211574 536614
rect 210954 536294 211574 536378
rect 210954 536058 210986 536294
rect 211222 536058 211306 536294
rect 211542 536058 211574 536294
rect 210954 500614 211574 536058
rect 210954 500378 210986 500614
rect 211222 500378 211306 500614
rect 211542 500378 211574 500614
rect 210954 500294 211574 500378
rect 210954 500058 210986 500294
rect 211222 500058 211306 500294
rect 211542 500058 211574 500294
rect 210954 464614 211574 500058
rect 210954 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 211574 464614
rect 210954 464294 211574 464378
rect 210954 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 211574 464294
rect 210954 428614 211574 464058
rect 210954 428378 210986 428614
rect 211222 428378 211306 428614
rect 211542 428378 211574 428614
rect 210954 428294 211574 428378
rect 210954 428058 210986 428294
rect 211222 428058 211306 428294
rect 211542 428058 211574 428294
rect 210954 392614 211574 428058
rect 210954 392378 210986 392614
rect 211222 392378 211306 392614
rect 211542 392378 211574 392614
rect 210954 392294 211574 392378
rect 210954 392058 210986 392294
rect 211222 392058 211306 392294
rect 211542 392058 211574 392294
rect 210954 356614 211574 392058
rect 210954 356378 210986 356614
rect 211222 356378 211306 356614
rect 211542 356378 211574 356614
rect 210954 356294 211574 356378
rect 210954 356058 210986 356294
rect 211222 356058 211306 356294
rect 211542 356058 211574 356294
rect 210954 320614 211574 356058
rect 210954 320378 210986 320614
rect 211222 320378 211306 320614
rect 211542 320378 211574 320614
rect 210954 320294 211574 320378
rect 210954 320058 210986 320294
rect 211222 320058 211306 320294
rect 211542 320058 211574 320294
rect 210954 302000 211574 320058
rect 217794 704838 218414 705830
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 543454 218414 578898
rect 217794 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 218414 543454
rect 217794 543134 218414 543218
rect 217794 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 218414 543134
rect 217794 507454 218414 542898
rect 217794 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 218414 507454
rect 217794 507134 218414 507218
rect 217794 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 218414 507134
rect 217794 471454 218414 506898
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 217794 435454 218414 470898
rect 217794 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 218414 435454
rect 217794 435134 218414 435218
rect 217794 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 218414 435134
rect 217794 399454 218414 434898
rect 217794 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 218414 399454
rect 217794 399134 218414 399218
rect 217794 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 218414 399134
rect 217794 363454 218414 398898
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 217794 327454 218414 362898
rect 217794 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 218414 327454
rect 217794 327134 218414 327218
rect 217794 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 218414 327134
rect 217794 302000 218414 326898
rect 221514 691174 222134 706202
rect 221514 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 222134 691174
rect 221514 690854 222134 690938
rect 221514 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 222134 690854
rect 221514 655174 222134 690618
rect 221514 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 222134 655174
rect 221514 654854 222134 654938
rect 221514 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 222134 654854
rect 221514 619174 222134 654618
rect 221514 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 222134 619174
rect 221514 618854 222134 618938
rect 221514 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 222134 618854
rect 221514 583174 222134 618618
rect 221514 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 222134 583174
rect 221514 582854 222134 582938
rect 221514 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 222134 582854
rect 221514 547174 222134 582618
rect 221514 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 222134 547174
rect 221514 546854 222134 546938
rect 221514 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 222134 546854
rect 221514 511174 222134 546618
rect 221514 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 222134 511174
rect 221514 510854 222134 510938
rect 221514 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 222134 510854
rect 221514 475174 222134 510618
rect 221514 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 222134 475174
rect 221514 474854 222134 474938
rect 221514 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 222134 474854
rect 221514 439174 222134 474618
rect 221514 438938 221546 439174
rect 221782 438938 221866 439174
rect 222102 438938 222134 439174
rect 221514 438854 222134 438938
rect 221514 438618 221546 438854
rect 221782 438618 221866 438854
rect 222102 438618 222134 438854
rect 221514 403174 222134 438618
rect 221514 402938 221546 403174
rect 221782 402938 221866 403174
rect 222102 402938 222134 403174
rect 221514 402854 222134 402938
rect 221514 402618 221546 402854
rect 221782 402618 221866 402854
rect 222102 402618 222134 402854
rect 221514 367174 222134 402618
rect 221514 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 222134 367174
rect 221514 366854 222134 366938
rect 221514 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 222134 366854
rect 221514 331174 222134 366618
rect 221514 330938 221546 331174
rect 221782 330938 221866 331174
rect 222102 330938 222134 331174
rect 221514 330854 222134 330938
rect 221514 330618 221546 330854
rect 221782 330618 221866 330854
rect 222102 330618 222134 330854
rect 221514 302000 222134 330618
rect 225234 694894 225854 708122
rect 225234 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 225854 694894
rect 225234 694574 225854 694658
rect 225234 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 225854 694574
rect 225234 658894 225854 694338
rect 225234 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 225854 658894
rect 225234 658574 225854 658658
rect 225234 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 225854 658574
rect 225234 622894 225854 658338
rect 225234 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 225854 622894
rect 225234 622574 225854 622658
rect 225234 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 225854 622574
rect 225234 586894 225854 622338
rect 225234 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 225854 586894
rect 225234 586574 225854 586658
rect 225234 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 225854 586574
rect 225234 550894 225854 586338
rect 225234 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 225854 550894
rect 225234 550574 225854 550658
rect 225234 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 225854 550574
rect 225234 514894 225854 550338
rect 225234 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 225854 514894
rect 225234 514574 225854 514658
rect 225234 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 225854 514574
rect 225234 478894 225854 514338
rect 225234 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 225854 478894
rect 225234 478574 225854 478658
rect 225234 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 225854 478574
rect 225234 442894 225854 478338
rect 225234 442658 225266 442894
rect 225502 442658 225586 442894
rect 225822 442658 225854 442894
rect 225234 442574 225854 442658
rect 225234 442338 225266 442574
rect 225502 442338 225586 442574
rect 225822 442338 225854 442574
rect 225234 406894 225854 442338
rect 225234 406658 225266 406894
rect 225502 406658 225586 406894
rect 225822 406658 225854 406894
rect 225234 406574 225854 406658
rect 225234 406338 225266 406574
rect 225502 406338 225586 406574
rect 225822 406338 225854 406574
rect 225234 370894 225854 406338
rect 225234 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 225854 370894
rect 225234 370574 225854 370658
rect 225234 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 225854 370574
rect 225234 334894 225854 370338
rect 225234 334658 225266 334894
rect 225502 334658 225586 334894
rect 225822 334658 225854 334894
rect 225234 334574 225854 334658
rect 225234 334338 225266 334574
rect 225502 334338 225586 334574
rect 225822 334338 225854 334574
rect 225234 302000 225854 334338
rect 228954 698614 229574 710042
rect 246954 711558 247574 711590
rect 246954 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 247574 711558
rect 246954 711238 247574 711322
rect 246954 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 247574 711238
rect 243234 709638 243854 709670
rect 243234 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 243854 709638
rect 243234 709318 243854 709402
rect 243234 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 243854 709318
rect 239514 707718 240134 707750
rect 239514 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 240134 707718
rect 239514 707398 240134 707482
rect 239514 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 240134 707398
rect 228954 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 229574 698614
rect 228954 698294 229574 698378
rect 228954 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 229574 698294
rect 228954 662614 229574 698058
rect 228954 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 229574 662614
rect 228954 662294 229574 662378
rect 228954 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 229574 662294
rect 228954 626614 229574 662058
rect 228954 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 229574 626614
rect 228954 626294 229574 626378
rect 228954 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 229574 626294
rect 228954 590614 229574 626058
rect 228954 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 229574 590614
rect 228954 590294 229574 590378
rect 228954 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 229574 590294
rect 228954 554614 229574 590058
rect 228954 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 229574 554614
rect 228954 554294 229574 554378
rect 228954 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 229574 554294
rect 228954 518614 229574 554058
rect 228954 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 229574 518614
rect 228954 518294 229574 518378
rect 228954 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 229574 518294
rect 228954 482614 229574 518058
rect 228954 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 229574 482614
rect 228954 482294 229574 482378
rect 228954 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 229574 482294
rect 228954 446614 229574 482058
rect 228954 446378 228986 446614
rect 229222 446378 229306 446614
rect 229542 446378 229574 446614
rect 228954 446294 229574 446378
rect 228954 446058 228986 446294
rect 229222 446058 229306 446294
rect 229542 446058 229574 446294
rect 228954 410614 229574 446058
rect 228954 410378 228986 410614
rect 229222 410378 229306 410614
rect 229542 410378 229574 410614
rect 228954 410294 229574 410378
rect 228954 410058 228986 410294
rect 229222 410058 229306 410294
rect 229542 410058 229574 410294
rect 228954 374614 229574 410058
rect 228954 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 229574 374614
rect 228954 374294 229574 374378
rect 228954 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 229574 374294
rect 228954 338614 229574 374058
rect 228954 338378 228986 338614
rect 229222 338378 229306 338614
rect 229542 338378 229574 338614
rect 228954 338294 229574 338378
rect 228954 338058 228986 338294
rect 229222 338058 229306 338294
rect 229542 338058 229574 338294
rect 228954 302614 229574 338058
rect 228954 302378 228986 302614
rect 229222 302378 229306 302614
rect 229542 302378 229574 302614
rect 228954 302294 229574 302378
rect 228954 302058 228986 302294
rect 229222 302058 229306 302294
rect 229542 302058 229574 302294
rect 228954 302000 229574 302058
rect 235794 705798 236414 705830
rect 235794 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 236414 705798
rect 235794 705478 236414 705562
rect 235794 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 236414 705478
rect 235794 669454 236414 705242
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 597454 236414 632898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 561454 236414 596898
rect 235794 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 236414 561454
rect 235794 561134 236414 561218
rect 235794 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 236414 561134
rect 235794 525454 236414 560898
rect 235794 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 236414 525454
rect 235794 525134 236414 525218
rect 235794 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 236414 525134
rect 235794 489454 236414 524898
rect 235794 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 236414 489454
rect 235794 489134 236414 489218
rect 235794 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 236414 489134
rect 235794 453454 236414 488898
rect 235794 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 236414 453454
rect 235794 453134 236414 453218
rect 235794 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 236414 453134
rect 235794 417454 236414 452898
rect 235794 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 236414 417454
rect 235794 417134 236414 417218
rect 235794 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 236414 417134
rect 235794 381454 236414 416898
rect 235794 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 236414 381454
rect 235794 381134 236414 381218
rect 235794 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 236414 381134
rect 235794 345454 236414 380898
rect 235794 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 236414 345454
rect 235794 345134 236414 345218
rect 235794 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 236414 345134
rect 235794 309454 236414 344898
rect 235794 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 236414 309454
rect 235794 309134 236414 309218
rect 235794 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 236414 309134
rect 235794 302000 236414 308898
rect 239514 673174 240134 707162
rect 239514 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 240134 673174
rect 239514 672854 240134 672938
rect 239514 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 240134 672854
rect 239514 637174 240134 672618
rect 239514 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 240134 637174
rect 239514 636854 240134 636938
rect 239514 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 240134 636854
rect 239514 601174 240134 636618
rect 239514 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 240134 601174
rect 239514 600854 240134 600938
rect 239514 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 240134 600854
rect 239514 565174 240134 600618
rect 239514 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 240134 565174
rect 239514 564854 240134 564938
rect 239514 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 240134 564854
rect 239514 529174 240134 564618
rect 239514 528938 239546 529174
rect 239782 528938 239866 529174
rect 240102 528938 240134 529174
rect 239514 528854 240134 528938
rect 239514 528618 239546 528854
rect 239782 528618 239866 528854
rect 240102 528618 240134 528854
rect 239514 493174 240134 528618
rect 239514 492938 239546 493174
rect 239782 492938 239866 493174
rect 240102 492938 240134 493174
rect 239514 492854 240134 492938
rect 239514 492618 239546 492854
rect 239782 492618 239866 492854
rect 240102 492618 240134 492854
rect 239514 457174 240134 492618
rect 239514 456938 239546 457174
rect 239782 456938 239866 457174
rect 240102 456938 240134 457174
rect 239514 456854 240134 456938
rect 239514 456618 239546 456854
rect 239782 456618 239866 456854
rect 240102 456618 240134 456854
rect 239514 421174 240134 456618
rect 239514 420938 239546 421174
rect 239782 420938 239866 421174
rect 240102 420938 240134 421174
rect 239514 420854 240134 420938
rect 239514 420618 239546 420854
rect 239782 420618 239866 420854
rect 240102 420618 240134 420854
rect 239514 385174 240134 420618
rect 239514 384938 239546 385174
rect 239782 384938 239866 385174
rect 240102 384938 240134 385174
rect 239514 384854 240134 384938
rect 239514 384618 239546 384854
rect 239782 384618 239866 384854
rect 240102 384618 240134 384854
rect 239514 349174 240134 384618
rect 239514 348938 239546 349174
rect 239782 348938 239866 349174
rect 240102 348938 240134 349174
rect 239514 348854 240134 348938
rect 239514 348618 239546 348854
rect 239782 348618 239866 348854
rect 240102 348618 240134 348854
rect 239514 313174 240134 348618
rect 239514 312938 239546 313174
rect 239782 312938 239866 313174
rect 240102 312938 240134 313174
rect 239514 312854 240134 312938
rect 239514 312618 239546 312854
rect 239782 312618 239866 312854
rect 240102 312618 240134 312854
rect 239514 302000 240134 312618
rect 243234 676894 243854 709082
rect 243234 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 243854 676894
rect 243234 676574 243854 676658
rect 243234 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 243854 676574
rect 243234 640894 243854 676338
rect 243234 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 243854 640894
rect 243234 640574 243854 640658
rect 243234 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 243854 640574
rect 243234 604894 243854 640338
rect 243234 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 243854 604894
rect 243234 604574 243854 604658
rect 243234 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 243854 604574
rect 243234 568894 243854 604338
rect 243234 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 243854 568894
rect 243234 568574 243854 568658
rect 243234 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 243854 568574
rect 243234 532894 243854 568338
rect 243234 532658 243266 532894
rect 243502 532658 243586 532894
rect 243822 532658 243854 532894
rect 243234 532574 243854 532658
rect 243234 532338 243266 532574
rect 243502 532338 243586 532574
rect 243822 532338 243854 532574
rect 243234 496894 243854 532338
rect 243234 496658 243266 496894
rect 243502 496658 243586 496894
rect 243822 496658 243854 496894
rect 243234 496574 243854 496658
rect 243234 496338 243266 496574
rect 243502 496338 243586 496574
rect 243822 496338 243854 496574
rect 243234 460894 243854 496338
rect 243234 460658 243266 460894
rect 243502 460658 243586 460894
rect 243822 460658 243854 460894
rect 243234 460574 243854 460658
rect 243234 460338 243266 460574
rect 243502 460338 243586 460574
rect 243822 460338 243854 460574
rect 243234 424894 243854 460338
rect 243234 424658 243266 424894
rect 243502 424658 243586 424894
rect 243822 424658 243854 424894
rect 243234 424574 243854 424658
rect 243234 424338 243266 424574
rect 243502 424338 243586 424574
rect 243822 424338 243854 424574
rect 243234 388894 243854 424338
rect 243234 388658 243266 388894
rect 243502 388658 243586 388894
rect 243822 388658 243854 388894
rect 243234 388574 243854 388658
rect 243234 388338 243266 388574
rect 243502 388338 243586 388574
rect 243822 388338 243854 388574
rect 243234 352894 243854 388338
rect 243234 352658 243266 352894
rect 243502 352658 243586 352894
rect 243822 352658 243854 352894
rect 243234 352574 243854 352658
rect 243234 352338 243266 352574
rect 243502 352338 243586 352574
rect 243822 352338 243854 352574
rect 243234 316894 243854 352338
rect 243234 316658 243266 316894
rect 243502 316658 243586 316894
rect 243822 316658 243854 316894
rect 243234 316574 243854 316658
rect 243234 316338 243266 316574
rect 243502 316338 243586 316574
rect 243822 316338 243854 316574
rect 243234 302000 243854 316338
rect 246954 680614 247574 711002
rect 264954 710598 265574 711590
rect 264954 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 265574 710598
rect 264954 710278 265574 710362
rect 264954 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 265574 710278
rect 261234 708678 261854 709670
rect 261234 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 261854 708678
rect 261234 708358 261854 708442
rect 261234 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 261854 708358
rect 257514 706758 258134 707750
rect 257514 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 258134 706758
rect 257514 706438 258134 706522
rect 257514 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 258134 706438
rect 246954 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 247574 680614
rect 246954 680294 247574 680378
rect 246954 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 247574 680294
rect 246954 644614 247574 680058
rect 246954 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 247574 644614
rect 246954 644294 247574 644378
rect 246954 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 247574 644294
rect 246954 608614 247574 644058
rect 246954 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 247574 608614
rect 246954 608294 247574 608378
rect 246954 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 247574 608294
rect 246954 572614 247574 608058
rect 246954 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 247574 572614
rect 246954 572294 247574 572378
rect 246954 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 247574 572294
rect 246954 536614 247574 572058
rect 246954 536378 246986 536614
rect 247222 536378 247306 536614
rect 247542 536378 247574 536614
rect 246954 536294 247574 536378
rect 246954 536058 246986 536294
rect 247222 536058 247306 536294
rect 247542 536058 247574 536294
rect 246954 500614 247574 536058
rect 246954 500378 246986 500614
rect 247222 500378 247306 500614
rect 247542 500378 247574 500614
rect 246954 500294 247574 500378
rect 246954 500058 246986 500294
rect 247222 500058 247306 500294
rect 247542 500058 247574 500294
rect 246954 464614 247574 500058
rect 246954 464378 246986 464614
rect 247222 464378 247306 464614
rect 247542 464378 247574 464614
rect 246954 464294 247574 464378
rect 246954 464058 246986 464294
rect 247222 464058 247306 464294
rect 247542 464058 247574 464294
rect 246954 428614 247574 464058
rect 246954 428378 246986 428614
rect 247222 428378 247306 428614
rect 247542 428378 247574 428614
rect 246954 428294 247574 428378
rect 246954 428058 246986 428294
rect 247222 428058 247306 428294
rect 247542 428058 247574 428294
rect 246954 392614 247574 428058
rect 246954 392378 246986 392614
rect 247222 392378 247306 392614
rect 247542 392378 247574 392614
rect 246954 392294 247574 392378
rect 246954 392058 246986 392294
rect 247222 392058 247306 392294
rect 247542 392058 247574 392294
rect 246954 356614 247574 392058
rect 246954 356378 246986 356614
rect 247222 356378 247306 356614
rect 247542 356378 247574 356614
rect 246954 356294 247574 356378
rect 246954 356058 246986 356294
rect 247222 356058 247306 356294
rect 247542 356058 247574 356294
rect 246954 320614 247574 356058
rect 246954 320378 246986 320614
rect 247222 320378 247306 320614
rect 247542 320378 247574 320614
rect 246954 320294 247574 320378
rect 246954 320058 246986 320294
rect 247222 320058 247306 320294
rect 247542 320058 247574 320294
rect 246954 302000 247574 320058
rect 253794 704838 254414 705830
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 543454 254414 578898
rect 253794 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 254414 543454
rect 253794 543134 254414 543218
rect 253794 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 254414 543134
rect 253794 507454 254414 542898
rect 253794 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 254414 507454
rect 253794 507134 254414 507218
rect 253794 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 254414 507134
rect 253794 471454 254414 506898
rect 253794 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 254414 471454
rect 253794 471134 254414 471218
rect 253794 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 254414 471134
rect 253794 435454 254414 470898
rect 253794 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 254414 435454
rect 253794 435134 254414 435218
rect 253794 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 254414 435134
rect 253794 399454 254414 434898
rect 253794 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 254414 399454
rect 253794 399134 254414 399218
rect 253794 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 254414 399134
rect 253794 363454 254414 398898
rect 253794 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 254414 363454
rect 253794 363134 254414 363218
rect 253794 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 254414 363134
rect 253794 327454 254414 362898
rect 253794 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 254414 327454
rect 253794 327134 254414 327218
rect 253794 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 254414 327134
rect 253794 302000 254414 326898
rect 257514 691174 258134 706202
rect 257514 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 258134 691174
rect 257514 690854 258134 690938
rect 257514 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 258134 690854
rect 257514 655174 258134 690618
rect 257514 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 258134 655174
rect 257514 654854 258134 654938
rect 257514 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 258134 654854
rect 257514 619174 258134 654618
rect 257514 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 258134 619174
rect 257514 618854 258134 618938
rect 257514 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 258134 618854
rect 257514 583174 258134 618618
rect 257514 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 258134 583174
rect 257514 582854 258134 582938
rect 257514 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 258134 582854
rect 257514 547174 258134 582618
rect 257514 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 258134 547174
rect 257514 546854 258134 546938
rect 257514 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 258134 546854
rect 257514 511174 258134 546618
rect 257514 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 258134 511174
rect 257514 510854 258134 510938
rect 257514 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 258134 510854
rect 257514 475174 258134 510618
rect 257514 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 258134 475174
rect 257514 474854 258134 474938
rect 257514 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 258134 474854
rect 257514 439174 258134 474618
rect 257514 438938 257546 439174
rect 257782 438938 257866 439174
rect 258102 438938 258134 439174
rect 257514 438854 258134 438938
rect 257514 438618 257546 438854
rect 257782 438618 257866 438854
rect 258102 438618 258134 438854
rect 257514 403174 258134 438618
rect 257514 402938 257546 403174
rect 257782 402938 257866 403174
rect 258102 402938 258134 403174
rect 257514 402854 258134 402938
rect 257514 402618 257546 402854
rect 257782 402618 257866 402854
rect 258102 402618 258134 402854
rect 257514 367174 258134 402618
rect 257514 366938 257546 367174
rect 257782 366938 257866 367174
rect 258102 366938 258134 367174
rect 257514 366854 258134 366938
rect 257514 366618 257546 366854
rect 257782 366618 257866 366854
rect 258102 366618 258134 366854
rect 257514 331174 258134 366618
rect 257514 330938 257546 331174
rect 257782 330938 257866 331174
rect 258102 330938 258134 331174
rect 257514 330854 258134 330938
rect 257514 330618 257546 330854
rect 257782 330618 257866 330854
rect 258102 330618 258134 330854
rect 257514 302000 258134 330618
rect 261234 694894 261854 708122
rect 261234 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 261854 694894
rect 261234 694574 261854 694658
rect 261234 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 261854 694574
rect 261234 658894 261854 694338
rect 261234 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 261854 658894
rect 261234 658574 261854 658658
rect 261234 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 261854 658574
rect 261234 622894 261854 658338
rect 261234 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 261854 622894
rect 261234 622574 261854 622658
rect 261234 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 261854 622574
rect 261234 586894 261854 622338
rect 261234 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 261854 586894
rect 261234 586574 261854 586658
rect 261234 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 261854 586574
rect 261234 550894 261854 586338
rect 261234 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 261854 550894
rect 261234 550574 261854 550658
rect 261234 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 261854 550574
rect 261234 514894 261854 550338
rect 261234 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 261854 514894
rect 261234 514574 261854 514658
rect 261234 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 261854 514574
rect 261234 478894 261854 514338
rect 261234 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 261854 478894
rect 261234 478574 261854 478658
rect 261234 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 261854 478574
rect 261234 442894 261854 478338
rect 261234 442658 261266 442894
rect 261502 442658 261586 442894
rect 261822 442658 261854 442894
rect 261234 442574 261854 442658
rect 261234 442338 261266 442574
rect 261502 442338 261586 442574
rect 261822 442338 261854 442574
rect 261234 406894 261854 442338
rect 261234 406658 261266 406894
rect 261502 406658 261586 406894
rect 261822 406658 261854 406894
rect 261234 406574 261854 406658
rect 261234 406338 261266 406574
rect 261502 406338 261586 406574
rect 261822 406338 261854 406574
rect 261234 370894 261854 406338
rect 261234 370658 261266 370894
rect 261502 370658 261586 370894
rect 261822 370658 261854 370894
rect 261234 370574 261854 370658
rect 261234 370338 261266 370574
rect 261502 370338 261586 370574
rect 261822 370338 261854 370574
rect 261234 334894 261854 370338
rect 261234 334658 261266 334894
rect 261502 334658 261586 334894
rect 261822 334658 261854 334894
rect 261234 334574 261854 334658
rect 261234 334338 261266 334574
rect 261502 334338 261586 334574
rect 261822 334338 261854 334574
rect 261234 302000 261854 334338
rect 264954 698614 265574 710042
rect 282954 711558 283574 711590
rect 282954 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 283574 711558
rect 282954 711238 283574 711322
rect 282954 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 283574 711238
rect 279234 709638 279854 709670
rect 279234 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 279854 709638
rect 279234 709318 279854 709402
rect 279234 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 279854 709318
rect 275514 707718 276134 707750
rect 275514 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 276134 707718
rect 275514 707398 276134 707482
rect 275514 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 276134 707398
rect 264954 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 265574 698614
rect 264954 698294 265574 698378
rect 264954 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 265574 698294
rect 264954 662614 265574 698058
rect 264954 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 265574 662614
rect 264954 662294 265574 662378
rect 264954 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 265574 662294
rect 264954 626614 265574 662058
rect 264954 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 265574 626614
rect 264954 626294 265574 626378
rect 264954 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 265574 626294
rect 264954 590614 265574 626058
rect 264954 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 265574 590614
rect 264954 590294 265574 590378
rect 264954 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 265574 590294
rect 264954 554614 265574 590058
rect 264954 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 265574 554614
rect 264954 554294 265574 554378
rect 264954 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 265574 554294
rect 264954 518614 265574 554058
rect 264954 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 265574 518614
rect 264954 518294 265574 518378
rect 264954 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 265574 518294
rect 264954 482614 265574 518058
rect 264954 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 265574 482614
rect 264954 482294 265574 482378
rect 264954 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 265574 482294
rect 264954 446614 265574 482058
rect 264954 446378 264986 446614
rect 265222 446378 265306 446614
rect 265542 446378 265574 446614
rect 264954 446294 265574 446378
rect 264954 446058 264986 446294
rect 265222 446058 265306 446294
rect 265542 446058 265574 446294
rect 264954 410614 265574 446058
rect 264954 410378 264986 410614
rect 265222 410378 265306 410614
rect 265542 410378 265574 410614
rect 264954 410294 265574 410378
rect 264954 410058 264986 410294
rect 265222 410058 265306 410294
rect 265542 410058 265574 410294
rect 264954 374614 265574 410058
rect 264954 374378 264986 374614
rect 265222 374378 265306 374614
rect 265542 374378 265574 374614
rect 264954 374294 265574 374378
rect 264954 374058 264986 374294
rect 265222 374058 265306 374294
rect 265542 374058 265574 374294
rect 264954 338614 265574 374058
rect 264954 338378 264986 338614
rect 265222 338378 265306 338614
rect 265542 338378 265574 338614
rect 264954 338294 265574 338378
rect 264954 338058 264986 338294
rect 265222 338058 265306 338294
rect 265542 338058 265574 338294
rect 264954 302614 265574 338058
rect 264954 302378 264986 302614
rect 265222 302378 265306 302614
rect 265542 302378 265574 302614
rect 264954 302294 265574 302378
rect 264954 302058 264986 302294
rect 265222 302058 265306 302294
rect 265542 302058 265574 302294
rect 264954 302000 265574 302058
rect 271794 705798 272414 705830
rect 271794 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 272414 705798
rect 271794 705478 272414 705562
rect 271794 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 272414 705478
rect 271794 669454 272414 705242
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 561454 272414 596898
rect 271794 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 272414 561454
rect 271794 561134 272414 561218
rect 271794 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 272414 561134
rect 271794 525454 272414 560898
rect 271794 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 272414 525454
rect 271794 525134 272414 525218
rect 271794 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 272414 525134
rect 271794 489454 272414 524898
rect 271794 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 272414 489454
rect 271794 489134 272414 489218
rect 271794 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 272414 489134
rect 271794 453454 272414 488898
rect 271794 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 272414 453454
rect 271794 453134 272414 453218
rect 271794 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 272414 453134
rect 271794 417454 272414 452898
rect 271794 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 272414 417454
rect 271794 417134 272414 417218
rect 271794 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 272414 417134
rect 271794 381454 272414 416898
rect 271794 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 272414 381454
rect 271794 381134 272414 381218
rect 271794 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 272414 381134
rect 271794 345454 272414 380898
rect 271794 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 272414 345454
rect 271794 345134 272414 345218
rect 271794 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 272414 345134
rect 271794 309454 272414 344898
rect 271794 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 272414 309454
rect 271794 309134 272414 309218
rect 271794 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 272414 309134
rect 271794 302000 272414 308898
rect 275514 673174 276134 707162
rect 275514 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 276134 673174
rect 275514 672854 276134 672938
rect 275514 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 276134 672854
rect 275514 637174 276134 672618
rect 275514 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 276134 637174
rect 275514 636854 276134 636938
rect 275514 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 276134 636854
rect 275514 601174 276134 636618
rect 275514 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 276134 601174
rect 275514 600854 276134 600938
rect 275514 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 276134 600854
rect 275514 565174 276134 600618
rect 275514 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 276134 565174
rect 275514 564854 276134 564938
rect 275514 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 276134 564854
rect 275514 529174 276134 564618
rect 275514 528938 275546 529174
rect 275782 528938 275866 529174
rect 276102 528938 276134 529174
rect 275514 528854 276134 528938
rect 275514 528618 275546 528854
rect 275782 528618 275866 528854
rect 276102 528618 276134 528854
rect 275514 493174 276134 528618
rect 275514 492938 275546 493174
rect 275782 492938 275866 493174
rect 276102 492938 276134 493174
rect 275514 492854 276134 492938
rect 275514 492618 275546 492854
rect 275782 492618 275866 492854
rect 276102 492618 276134 492854
rect 275514 457174 276134 492618
rect 275514 456938 275546 457174
rect 275782 456938 275866 457174
rect 276102 456938 276134 457174
rect 275514 456854 276134 456938
rect 275514 456618 275546 456854
rect 275782 456618 275866 456854
rect 276102 456618 276134 456854
rect 275514 421174 276134 456618
rect 275514 420938 275546 421174
rect 275782 420938 275866 421174
rect 276102 420938 276134 421174
rect 275514 420854 276134 420938
rect 275514 420618 275546 420854
rect 275782 420618 275866 420854
rect 276102 420618 276134 420854
rect 275514 385174 276134 420618
rect 275514 384938 275546 385174
rect 275782 384938 275866 385174
rect 276102 384938 276134 385174
rect 275514 384854 276134 384938
rect 275514 384618 275546 384854
rect 275782 384618 275866 384854
rect 276102 384618 276134 384854
rect 275514 349174 276134 384618
rect 275514 348938 275546 349174
rect 275782 348938 275866 349174
rect 276102 348938 276134 349174
rect 275514 348854 276134 348938
rect 275514 348618 275546 348854
rect 275782 348618 275866 348854
rect 276102 348618 276134 348854
rect 275514 313174 276134 348618
rect 275514 312938 275546 313174
rect 275782 312938 275866 313174
rect 276102 312938 276134 313174
rect 275514 312854 276134 312938
rect 275514 312618 275546 312854
rect 275782 312618 275866 312854
rect 276102 312618 276134 312854
rect 275514 302000 276134 312618
rect 279234 676894 279854 709082
rect 279234 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 279854 676894
rect 279234 676574 279854 676658
rect 279234 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 279854 676574
rect 279234 640894 279854 676338
rect 279234 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 279854 640894
rect 279234 640574 279854 640658
rect 279234 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 279854 640574
rect 279234 604894 279854 640338
rect 279234 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 279854 604894
rect 279234 604574 279854 604658
rect 279234 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 279854 604574
rect 279234 568894 279854 604338
rect 279234 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 279854 568894
rect 279234 568574 279854 568658
rect 279234 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 279854 568574
rect 279234 532894 279854 568338
rect 279234 532658 279266 532894
rect 279502 532658 279586 532894
rect 279822 532658 279854 532894
rect 279234 532574 279854 532658
rect 279234 532338 279266 532574
rect 279502 532338 279586 532574
rect 279822 532338 279854 532574
rect 279234 496894 279854 532338
rect 279234 496658 279266 496894
rect 279502 496658 279586 496894
rect 279822 496658 279854 496894
rect 279234 496574 279854 496658
rect 279234 496338 279266 496574
rect 279502 496338 279586 496574
rect 279822 496338 279854 496574
rect 279234 460894 279854 496338
rect 279234 460658 279266 460894
rect 279502 460658 279586 460894
rect 279822 460658 279854 460894
rect 279234 460574 279854 460658
rect 279234 460338 279266 460574
rect 279502 460338 279586 460574
rect 279822 460338 279854 460574
rect 279234 424894 279854 460338
rect 279234 424658 279266 424894
rect 279502 424658 279586 424894
rect 279822 424658 279854 424894
rect 279234 424574 279854 424658
rect 279234 424338 279266 424574
rect 279502 424338 279586 424574
rect 279822 424338 279854 424574
rect 279234 388894 279854 424338
rect 279234 388658 279266 388894
rect 279502 388658 279586 388894
rect 279822 388658 279854 388894
rect 279234 388574 279854 388658
rect 279234 388338 279266 388574
rect 279502 388338 279586 388574
rect 279822 388338 279854 388574
rect 279234 352894 279854 388338
rect 279234 352658 279266 352894
rect 279502 352658 279586 352894
rect 279822 352658 279854 352894
rect 279234 352574 279854 352658
rect 279234 352338 279266 352574
rect 279502 352338 279586 352574
rect 279822 352338 279854 352574
rect 279234 316894 279854 352338
rect 279234 316658 279266 316894
rect 279502 316658 279586 316894
rect 279822 316658 279854 316894
rect 279234 316574 279854 316658
rect 279234 316338 279266 316574
rect 279502 316338 279586 316574
rect 279822 316338 279854 316574
rect 279234 302000 279854 316338
rect 282954 680614 283574 711002
rect 300954 710598 301574 711590
rect 300954 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 301574 710598
rect 300954 710278 301574 710362
rect 300954 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 301574 710278
rect 297234 708678 297854 709670
rect 297234 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 297854 708678
rect 297234 708358 297854 708442
rect 297234 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 297854 708358
rect 293514 706758 294134 707750
rect 293514 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 294134 706758
rect 293514 706438 294134 706522
rect 293514 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 294134 706438
rect 282954 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 283574 680614
rect 282954 680294 283574 680378
rect 282954 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 283574 680294
rect 282954 644614 283574 680058
rect 282954 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 283574 644614
rect 282954 644294 283574 644378
rect 282954 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 283574 644294
rect 282954 608614 283574 644058
rect 282954 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 283574 608614
rect 282954 608294 283574 608378
rect 282954 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 283574 608294
rect 282954 572614 283574 608058
rect 282954 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 283574 572614
rect 282954 572294 283574 572378
rect 282954 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 283574 572294
rect 282954 536614 283574 572058
rect 282954 536378 282986 536614
rect 283222 536378 283306 536614
rect 283542 536378 283574 536614
rect 282954 536294 283574 536378
rect 282954 536058 282986 536294
rect 283222 536058 283306 536294
rect 283542 536058 283574 536294
rect 282954 500614 283574 536058
rect 282954 500378 282986 500614
rect 283222 500378 283306 500614
rect 283542 500378 283574 500614
rect 282954 500294 283574 500378
rect 282954 500058 282986 500294
rect 283222 500058 283306 500294
rect 283542 500058 283574 500294
rect 282954 464614 283574 500058
rect 282954 464378 282986 464614
rect 283222 464378 283306 464614
rect 283542 464378 283574 464614
rect 282954 464294 283574 464378
rect 282954 464058 282986 464294
rect 283222 464058 283306 464294
rect 283542 464058 283574 464294
rect 282954 428614 283574 464058
rect 282954 428378 282986 428614
rect 283222 428378 283306 428614
rect 283542 428378 283574 428614
rect 282954 428294 283574 428378
rect 282954 428058 282986 428294
rect 283222 428058 283306 428294
rect 283542 428058 283574 428294
rect 282954 392614 283574 428058
rect 282954 392378 282986 392614
rect 283222 392378 283306 392614
rect 283542 392378 283574 392614
rect 282954 392294 283574 392378
rect 282954 392058 282986 392294
rect 283222 392058 283306 392294
rect 283542 392058 283574 392294
rect 282954 356614 283574 392058
rect 282954 356378 282986 356614
rect 283222 356378 283306 356614
rect 283542 356378 283574 356614
rect 282954 356294 283574 356378
rect 282954 356058 282986 356294
rect 283222 356058 283306 356294
rect 283542 356058 283574 356294
rect 282954 320614 283574 356058
rect 282954 320378 282986 320614
rect 283222 320378 283306 320614
rect 283542 320378 283574 320614
rect 282954 320294 283574 320378
rect 282954 320058 282986 320294
rect 283222 320058 283306 320294
rect 283542 320058 283574 320294
rect 282954 302000 283574 320058
rect 289794 704838 290414 705830
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 543454 290414 578898
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289794 507454 290414 542898
rect 289794 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 290414 507454
rect 289794 507134 290414 507218
rect 289794 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 290414 507134
rect 289794 471454 290414 506898
rect 289794 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 290414 471454
rect 289794 471134 290414 471218
rect 289794 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 290414 471134
rect 289794 435454 290414 470898
rect 289794 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 290414 435454
rect 289794 435134 290414 435218
rect 289794 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 290414 435134
rect 289794 399454 290414 434898
rect 289794 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 290414 399454
rect 289794 399134 290414 399218
rect 289794 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 290414 399134
rect 289794 363454 290414 398898
rect 289794 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 290414 363454
rect 289794 363134 290414 363218
rect 289794 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 290414 363134
rect 289794 327454 290414 362898
rect 289794 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 290414 327454
rect 289794 327134 290414 327218
rect 289794 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 290414 327134
rect 289794 302000 290414 326898
rect 293514 691174 294134 706202
rect 293514 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 294134 691174
rect 293514 690854 294134 690938
rect 293514 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 294134 690854
rect 293514 655174 294134 690618
rect 293514 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 294134 655174
rect 293514 654854 294134 654938
rect 293514 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 294134 654854
rect 293514 619174 294134 654618
rect 293514 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 294134 619174
rect 293514 618854 294134 618938
rect 293514 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 294134 618854
rect 293514 583174 294134 618618
rect 293514 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 294134 583174
rect 293514 582854 294134 582938
rect 293514 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 294134 582854
rect 293514 547174 294134 582618
rect 293514 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 294134 547174
rect 293514 546854 294134 546938
rect 293514 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 294134 546854
rect 293514 511174 294134 546618
rect 293514 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 294134 511174
rect 293514 510854 294134 510938
rect 293514 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 294134 510854
rect 293514 475174 294134 510618
rect 293514 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 294134 475174
rect 293514 474854 294134 474938
rect 293514 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 294134 474854
rect 293514 439174 294134 474618
rect 293514 438938 293546 439174
rect 293782 438938 293866 439174
rect 294102 438938 294134 439174
rect 293514 438854 294134 438938
rect 293514 438618 293546 438854
rect 293782 438618 293866 438854
rect 294102 438618 294134 438854
rect 293514 403174 294134 438618
rect 293514 402938 293546 403174
rect 293782 402938 293866 403174
rect 294102 402938 294134 403174
rect 293514 402854 294134 402938
rect 293514 402618 293546 402854
rect 293782 402618 293866 402854
rect 294102 402618 294134 402854
rect 293514 367174 294134 402618
rect 293514 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 294134 367174
rect 293514 366854 294134 366938
rect 293514 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 294134 366854
rect 293514 331174 294134 366618
rect 293514 330938 293546 331174
rect 293782 330938 293866 331174
rect 294102 330938 294134 331174
rect 293514 330854 294134 330938
rect 293514 330618 293546 330854
rect 293782 330618 293866 330854
rect 294102 330618 294134 330854
rect 293514 302000 294134 330618
rect 297234 694894 297854 708122
rect 297234 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 297854 694894
rect 297234 694574 297854 694658
rect 297234 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 297854 694574
rect 297234 658894 297854 694338
rect 297234 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 297854 658894
rect 297234 658574 297854 658658
rect 297234 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 297854 658574
rect 297234 622894 297854 658338
rect 297234 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 297854 622894
rect 297234 622574 297854 622658
rect 297234 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 297854 622574
rect 297234 586894 297854 622338
rect 297234 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 297854 586894
rect 297234 586574 297854 586658
rect 297234 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 297854 586574
rect 297234 550894 297854 586338
rect 297234 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 297854 550894
rect 297234 550574 297854 550658
rect 297234 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 297854 550574
rect 297234 514894 297854 550338
rect 297234 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 297854 514894
rect 297234 514574 297854 514658
rect 297234 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 297854 514574
rect 297234 478894 297854 514338
rect 297234 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 297854 478894
rect 297234 478574 297854 478658
rect 297234 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 297854 478574
rect 297234 442894 297854 478338
rect 297234 442658 297266 442894
rect 297502 442658 297586 442894
rect 297822 442658 297854 442894
rect 297234 442574 297854 442658
rect 297234 442338 297266 442574
rect 297502 442338 297586 442574
rect 297822 442338 297854 442574
rect 297234 406894 297854 442338
rect 297234 406658 297266 406894
rect 297502 406658 297586 406894
rect 297822 406658 297854 406894
rect 297234 406574 297854 406658
rect 297234 406338 297266 406574
rect 297502 406338 297586 406574
rect 297822 406338 297854 406574
rect 297234 370894 297854 406338
rect 297234 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 297854 370894
rect 297234 370574 297854 370658
rect 297234 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 297854 370574
rect 297234 334894 297854 370338
rect 297234 334658 297266 334894
rect 297502 334658 297586 334894
rect 297822 334658 297854 334894
rect 297234 334574 297854 334658
rect 297234 334338 297266 334574
rect 297502 334338 297586 334574
rect 297822 334338 297854 334574
rect 297234 302000 297854 334338
rect 300954 698614 301574 710042
rect 318954 711558 319574 711590
rect 318954 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 319574 711558
rect 318954 711238 319574 711322
rect 318954 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 319574 711238
rect 315234 709638 315854 709670
rect 315234 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 315854 709638
rect 315234 709318 315854 709402
rect 315234 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 315854 709318
rect 311514 707718 312134 707750
rect 311514 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 312134 707718
rect 311514 707398 312134 707482
rect 311514 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 312134 707398
rect 300954 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 301574 698614
rect 300954 698294 301574 698378
rect 300954 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 301574 698294
rect 300954 662614 301574 698058
rect 300954 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 301574 662614
rect 300954 662294 301574 662378
rect 300954 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 301574 662294
rect 300954 626614 301574 662058
rect 300954 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 301574 626614
rect 300954 626294 301574 626378
rect 300954 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 301574 626294
rect 300954 590614 301574 626058
rect 300954 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 301574 590614
rect 300954 590294 301574 590378
rect 300954 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 301574 590294
rect 300954 554614 301574 590058
rect 300954 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 301574 554614
rect 300954 554294 301574 554378
rect 300954 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 301574 554294
rect 300954 518614 301574 554058
rect 300954 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 301574 518614
rect 300954 518294 301574 518378
rect 300954 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 301574 518294
rect 300954 482614 301574 518058
rect 300954 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 301574 482614
rect 300954 482294 301574 482378
rect 300954 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 301574 482294
rect 300954 446614 301574 482058
rect 300954 446378 300986 446614
rect 301222 446378 301306 446614
rect 301542 446378 301574 446614
rect 300954 446294 301574 446378
rect 300954 446058 300986 446294
rect 301222 446058 301306 446294
rect 301542 446058 301574 446294
rect 300954 410614 301574 446058
rect 300954 410378 300986 410614
rect 301222 410378 301306 410614
rect 301542 410378 301574 410614
rect 300954 410294 301574 410378
rect 300954 410058 300986 410294
rect 301222 410058 301306 410294
rect 301542 410058 301574 410294
rect 300954 374614 301574 410058
rect 300954 374378 300986 374614
rect 301222 374378 301306 374614
rect 301542 374378 301574 374614
rect 300954 374294 301574 374378
rect 300954 374058 300986 374294
rect 301222 374058 301306 374294
rect 301542 374058 301574 374294
rect 300954 338614 301574 374058
rect 300954 338378 300986 338614
rect 301222 338378 301306 338614
rect 301542 338378 301574 338614
rect 300954 338294 301574 338378
rect 300954 338058 300986 338294
rect 301222 338058 301306 338294
rect 301542 338058 301574 338294
rect 300954 302614 301574 338058
rect 300954 302378 300986 302614
rect 301222 302378 301306 302614
rect 301542 302378 301574 302614
rect 300954 302294 301574 302378
rect 300954 302058 300986 302294
rect 301222 302058 301306 302294
rect 301542 302058 301574 302294
rect 300954 302000 301574 302058
rect 307794 705798 308414 705830
rect 307794 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 308414 705798
rect 307794 705478 308414 705562
rect 307794 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 308414 705478
rect 307794 669454 308414 705242
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 561454 308414 596898
rect 307794 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 308414 561454
rect 307794 561134 308414 561218
rect 307794 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 308414 561134
rect 307794 525454 308414 560898
rect 307794 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 308414 525454
rect 307794 525134 308414 525218
rect 307794 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 308414 525134
rect 307794 489454 308414 524898
rect 307794 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 308414 489454
rect 307794 489134 308414 489218
rect 307794 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 308414 489134
rect 307794 453454 308414 488898
rect 307794 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 308414 453454
rect 307794 453134 308414 453218
rect 307794 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 308414 453134
rect 307794 417454 308414 452898
rect 307794 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 308414 417454
rect 307794 417134 308414 417218
rect 307794 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 308414 417134
rect 307794 381454 308414 416898
rect 307794 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 308414 381454
rect 307794 381134 308414 381218
rect 307794 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 308414 381134
rect 307794 345454 308414 380898
rect 307794 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 308414 345454
rect 307794 345134 308414 345218
rect 307794 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 308414 345134
rect 307794 309454 308414 344898
rect 307794 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 308414 309454
rect 307794 309134 308414 309218
rect 307794 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 308414 309134
rect 204208 291454 204528 291486
rect 204208 291218 204250 291454
rect 204486 291218 204528 291454
rect 204208 291134 204528 291218
rect 204208 290898 204250 291134
rect 204486 290898 204528 291134
rect 204208 290866 204528 290898
rect 234928 291454 235248 291486
rect 234928 291218 234970 291454
rect 235206 291218 235248 291454
rect 234928 291134 235248 291218
rect 234928 290898 234970 291134
rect 235206 290898 235248 291134
rect 234928 290866 235248 290898
rect 265648 291454 265968 291486
rect 265648 291218 265690 291454
rect 265926 291218 265968 291454
rect 265648 291134 265968 291218
rect 265648 290898 265690 291134
rect 265926 290898 265968 291134
rect 265648 290866 265968 290898
rect 296368 291454 296688 291486
rect 296368 291218 296410 291454
rect 296646 291218 296688 291454
rect 296368 291134 296688 291218
rect 296368 290898 296410 291134
rect 296646 290898 296688 291134
rect 296368 290866 296688 290898
rect 219568 273454 219888 273486
rect 219568 273218 219610 273454
rect 219846 273218 219888 273454
rect 219568 273134 219888 273218
rect 219568 272898 219610 273134
rect 219846 272898 219888 273134
rect 219568 272866 219888 272898
rect 250288 273454 250608 273486
rect 250288 273218 250330 273454
rect 250566 273218 250608 273454
rect 250288 273134 250608 273218
rect 250288 272898 250330 273134
rect 250566 272898 250608 273134
rect 250288 272866 250608 272898
rect 281008 273454 281328 273486
rect 281008 273218 281050 273454
rect 281286 273218 281328 273454
rect 281008 273134 281328 273218
rect 281008 272898 281050 273134
rect 281286 272898 281328 273134
rect 281008 272866 281328 272898
rect 307794 273454 308414 308898
rect 307794 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 308414 273454
rect 307794 273134 308414 273218
rect 307794 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 308414 273134
rect 192954 266378 192986 266614
rect 193222 266378 193306 266614
rect 193542 266378 193574 266614
rect 192954 266294 193574 266378
rect 192954 266058 192986 266294
rect 193222 266058 193306 266294
rect 193542 266058 193574 266294
rect 192954 230614 193574 266058
rect 204208 255454 204528 255486
rect 204208 255218 204250 255454
rect 204486 255218 204528 255454
rect 204208 255134 204528 255218
rect 204208 254898 204250 255134
rect 204486 254898 204528 255134
rect 204208 254866 204528 254898
rect 234928 255454 235248 255486
rect 234928 255218 234970 255454
rect 235206 255218 235248 255454
rect 234928 255134 235248 255218
rect 234928 254898 234970 255134
rect 235206 254898 235248 255134
rect 234928 254866 235248 254898
rect 265648 255454 265968 255486
rect 265648 255218 265690 255454
rect 265926 255218 265968 255454
rect 265648 255134 265968 255218
rect 265648 254898 265690 255134
rect 265926 254898 265968 255134
rect 265648 254866 265968 254898
rect 296368 255454 296688 255486
rect 296368 255218 296410 255454
rect 296646 255218 296688 255454
rect 296368 255134 296688 255218
rect 296368 254898 296410 255134
rect 296646 254898 296688 255134
rect 296368 254866 296688 254898
rect 219568 237454 219888 237486
rect 219568 237218 219610 237454
rect 219846 237218 219888 237454
rect 219568 237134 219888 237218
rect 219568 236898 219610 237134
rect 219846 236898 219888 237134
rect 219568 236866 219888 236898
rect 250288 237454 250608 237486
rect 250288 237218 250330 237454
rect 250566 237218 250608 237454
rect 250288 237134 250608 237218
rect 250288 236898 250330 237134
rect 250566 236898 250608 237134
rect 250288 236866 250608 236898
rect 281008 237454 281328 237486
rect 281008 237218 281050 237454
rect 281286 237218 281328 237454
rect 281008 237134 281328 237218
rect 281008 236898 281050 237134
rect 281286 236898 281328 237134
rect 281008 236866 281328 236898
rect 307794 237454 308414 272898
rect 307794 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 308414 237454
rect 307794 237134 308414 237218
rect 307794 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 308414 237134
rect 192954 230378 192986 230614
rect 193222 230378 193306 230614
rect 193542 230378 193574 230614
rect 192954 230294 193574 230378
rect 192954 230058 192986 230294
rect 193222 230058 193306 230294
rect 193542 230058 193574 230294
rect 192954 194614 193574 230058
rect 204208 219454 204528 219486
rect 204208 219218 204250 219454
rect 204486 219218 204528 219454
rect 204208 219134 204528 219218
rect 204208 218898 204250 219134
rect 204486 218898 204528 219134
rect 204208 218866 204528 218898
rect 234928 219454 235248 219486
rect 234928 219218 234970 219454
rect 235206 219218 235248 219454
rect 234928 219134 235248 219218
rect 234928 218898 234970 219134
rect 235206 218898 235248 219134
rect 234928 218866 235248 218898
rect 265648 219454 265968 219486
rect 265648 219218 265690 219454
rect 265926 219218 265968 219454
rect 265648 219134 265968 219218
rect 265648 218898 265690 219134
rect 265926 218898 265968 219134
rect 265648 218866 265968 218898
rect 296368 219454 296688 219486
rect 296368 219218 296410 219454
rect 296646 219218 296688 219454
rect 296368 219134 296688 219218
rect 296368 218898 296410 219134
rect 296646 218898 296688 219134
rect 296368 218866 296688 218898
rect 219568 201454 219888 201486
rect 219568 201218 219610 201454
rect 219846 201218 219888 201454
rect 219568 201134 219888 201218
rect 219568 200898 219610 201134
rect 219846 200898 219888 201134
rect 219568 200866 219888 200898
rect 250288 201454 250608 201486
rect 250288 201218 250330 201454
rect 250566 201218 250608 201454
rect 250288 201134 250608 201218
rect 250288 200898 250330 201134
rect 250566 200898 250608 201134
rect 250288 200866 250608 200898
rect 281008 201454 281328 201486
rect 281008 201218 281050 201454
rect 281286 201218 281328 201454
rect 281008 201134 281328 201218
rect 281008 200898 281050 201134
rect 281286 200898 281328 201134
rect 281008 200866 281328 200898
rect 307794 201454 308414 236898
rect 307794 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 308414 201454
rect 307794 201134 308414 201218
rect 307794 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 308414 201134
rect 192954 194378 192986 194614
rect 193222 194378 193306 194614
rect 193542 194378 193574 194614
rect 192954 194294 193574 194378
rect 192954 194058 192986 194294
rect 193222 194058 193306 194294
rect 193542 194058 193574 194294
rect 192954 158614 193574 194058
rect 204208 183454 204528 183486
rect 204208 183218 204250 183454
rect 204486 183218 204528 183454
rect 204208 183134 204528 183218
rect 204208 182898 204250 183134
rect 204486 182898 204528 183134
rect 204208 182866 204528 182898
rect 234928 183454 235248 183486
rect 234928 183218 234970 183454
rect 235206 183218 235248 183454
rect 234928 183134 235248 183218
rect 234928 182898 234970 183134
rect 235206 182898 235248 183134
rect 234928 182866 235248 182898
rect 265648 183454 265968 183486
rect 265648 183218 265690 183454
rect 265926 183218 265968 183454
rect 265648 183134 265968 183218
rect 265648 182898 265690 183134
rect 265926 182898 265968 183134
rect 265648 182866 265968 182898
rect 296368 183454 296688 183486
rect 296368 183218 296410 183454
rect 296646 183218 296688 183454
rect 296368 183134 296688 183218
rect 296368 182898 296410 183134
rect 296646 182898 296688 183134
rect 296368 182866 296688 182898
rect 219568 165454 219888 165486
rect 219568 165218 219610 165454
rect 219846 165218 219888 165454
rect 219568 165134 219888 165218
rect 219568 164898 219610 165134
rect 219846 164898 219888 165134
rect 219568 164866 219888 164898
rect 250288 165454 250608 165486
rect 250288 165218 250330 165454
rect 250566 165218 250608 165454
rect 250288 165134 250608 165218
rect 250288 164898 250330 165134
rect 250566 164898 250608 165134
rect 250288 164866 250608 164898
rect 281008 165454 281328 165486
rect 281008 165218 281050 165454
rect 281286 165218 281328 165454
rect 281008 165134 281328 165218
rect 281008 164898 281050 165134
rect 281286 164898 281328 165134
rect 281008 164866 281328 164898
rect 307794 165454 308414 200898
rect 307794 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 308414 165454
rect 307794 165134 308414 165218
rect 307794 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 308414 165134
rect 192954 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 193574 158614
rect 192954 158294 193574 158378
rect 192954 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 193574 158294
rect 192954 122614 193574 158058
rect 204208 147454 204528 147486
rect 204208 147218 204250 147454
rect 204486 147218 204528 147454
rect 204208 147134 204528 147218
rect 204208 146898 204250 147134
rect 204486 146898 204528 147134
rect 204208 146866 204528 146898
rect 234928 147454 235248 147486
rect 234928 147218 234970 147454
rect 235206 147218 235248 147454
rect 234928 147134 235248 147218
rect 234928 146898 234970 147134
rect 235206 146898 235248 147134
rect 234928 146866 235248 146898
rect 265648 147454 265968 147486
rect 265648 147218 265690 147454
rect 265926 147218 265968 147454
rect 265648 147134 265968 147218
rect 265648 146898 265690 147134
rect 265926 146898 265968 147134
rect 265648 146866 265968 146898
rect 296368 147454 296688 147486
rect 296368 147218 296410 147454
rect 296646 147218 296688 147454
rect 296368 147134 296688 147218
rect 296368 146898 296410 147134
rect 296646 146898 296688 147134
rect 296368 146866 296688 146898
rect 219568 129454 219888 129486
rect 219568 129218 219610 129454
rect 219846 129218 219888 129454
rect 219568 129134 219888 129218
rect 219568 128898 219610 129134
rect 219846 128898 219888 129134
rect 219568 128866 219888 128898
rect 250288 129454 250608 129486
rect 250288 129218 250330 129454
rect 250566 129218 250608 129454
rect 250288 129134 250608 129218
rect 250288 128898 250330 129134
rect 250566 128898 250608 129134
rect 250288 128866 250608 128898
rect 281008 129454 281328 129486
rect 281008 129218 281050 129454
rect 281286 129218 281328 129454
rect 281008 129134 281328 129218
rect 281008 128898 281050 129134
rect 281286 128898 281328 129134
rect 281008 128866 281328 128898
rect 307794 129454 308414 164898
rect 307794 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 308414 129454
rect 307794 129134 308414 129218
rect 307794 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 308414 129134
rect 192954 122378 192986 122614
rect 193222 122378 193306 122614
rect 193542 122378 193574 122614
rect 192954 122294 193574 122378
rect 192954 122058 192986 122294
rect 193222 122058 193306 122294
rect 193542 122058 193574 122294
rect 192954 86614 193574 122058
rect 204208 111454 204528 111486
rect 204208 111218 204250 111454
rect 204486 111218 204528 111454
rect 204208 111134 204528 111218
rect 204208 110898 204250 111134
rect 204486 110898 204528 111134
rect 204208 110866 204528 110898
rect 234928 111454 235248 111486
rect 234928 111218 234970 111454
rect 235206 111218 235248 111454
rect 234928 111134 235248 111218
rect 234928 110898 234970 111134
rect 235206 110898 235248 111134
rect 234928 110866 235248 110898
rect 265648 111454 265968 111486
rect 265648 111218 265690 111454
rect 265926 111218 265968 111454
rect 265648 111134 265968 111218
rect 265648 110898 265690 111134
rect 265926 110898 265968 111134
rect 265648 110866 265968 110898
rect 296368 111454 296688 111486
rect 296368 111218 296410 111454
rect 296646 111218 296688 111454
rect 296368 111134 296688 111218
rect 296368 110898 296410 111134
rect 296646 110898 296688 111134
rect 296368 110866 296688 110898
rect 192954 86378 192986 86614
rect 193222 86378 193306 86614
rect 193542 86378 193574 86614
rect 192954 86294 193574 86378
rect 192954 86058 192986 86294
rect 193222 86058 193306 86294
rect 193542 86058 193574 86294
rect 192954 50614 193574 86058
rect 192954 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 193574 50614
rect 192954 50294 193574 50378
rect 192954 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 193574 50294
rect 192954 14614 193574 50058
rect 192954 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 193574 14614
rect 192954 14294 193574 14378
rect 192954 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 193574 14294
rect 174954 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 175574 -7066
rect 174954 -7386 175574 -7302
rect 174954 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 175574 -7386
rect 174954 -7654 175574 -7622
rect 192954 -6106 193574 14058
rect 199794 93454 200414 98000
rect 199794 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 200414 93454
rect 199794 93134 200414 93218
rect 199794 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 200414 93134
rect 199794 57454 200414 92898
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 21454 200414 56898
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -1306 200414 20898
rect 199794 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 200414 -1306
rect 199794 -1626 200414 -1542
rect 199794 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 200414 -1626
rect 199794 -1894 200414 -1862
rect 203514 97174 204134 98000
rect 203514 96938 203546 97174
rect 203782 96938 203866 97174
rect 204102 96938 204134 97174
rect 203514 96854 204134 96938
rect 203514 96618 203546 96854
rect 203782 96618 203866 96854
rect 204102 96618 204134 96854
rect 203514 61174 204134 96618
rect 203514 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 204134 61174
rect 203514 60854 204134 60938
rect 203514 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 204134 60854
rect 203514 25174 204134 60618
rect 203514 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 204134 25174
rect 203514 24854 204134 24938
rect 203514 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 204134 24854
rect 203514 -3226 204134 24618
rect 203514 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 204134 -3226
rect 203514 -3546 204134 -3462
rect 203514 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 204134 -3546
rect 203514 -3814 204134 -3782
rect 207234 64894 207854 98000
rect 207234 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 207854 64894
rect 207234 64574 207854 64658
rect 207234 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 207854 64574
rect 207234 28894 207854 64338
rect 207234 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 207854 28894
rect 207234 28574 207854 28658
rect 207234 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 207854 28574
rect 207234 -5146 207854 28338
rect 207234 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 207854 -5146
rect 207234 -5466 207854 -5382
rect 207234 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 207854 -5466
rect 207234 -5734 207854 -5702
rect 210954 68614 211574 98000
rect 210954 68378 210986 68614
rect 211222 68378 211306 68614
rect 211542 68378 211574 68614
rect 210954 68294 211574 68378
rect 210954 68058 210986 68294
rect 211222 68058 211306 68294
rect 211542 68058 211574 68294
rect 210954 32614 211574 68058
rect 210954 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 211574 32614
rect 210954 32294 211574 32378
rect 210954 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 211574 32294
rect 192954 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 193574 -6106
rect 192954 -6426 193574 -6342
rect 192954 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 193574 -6426
rect 192954 -7654 193574 -6662
rect 210954 -7066 211574 32058
rect 217794 75454 218414 98000
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 217794 39454 218414 74898
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -1894 218414 -902
rect 221514 79174 222134 98000
rect 221514 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 222134 79174
rect 221514 78854 222134 78938
rect 221514 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 222134 78854
rect 221514 43174 222134 78618
rect 221514 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 222134 43174
rect 221514 42854 222134 42938
rect 221514 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 222134 42854
rect 221514 7174 222134 42618
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -2266 222134 6618
rect 221514 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 222134 -2266
rect 221514 -2586 222134 -2502
rect 221514 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 222134 -2586
rect 221514 -3814 222134 -2822
rect 225234 82894 225854 98000
rect 225234 82658 225266 82894
rect 225502 82658 225586 82894
rect 225822 82658 225854 82894
rect 225234 82574 225854 82658
rect 225234 82338 225266 82574
rect 225502 82338 225586 82574
rect 225822 82338 225854 82574
rect 225234 46894 225854 82338
rect 225234 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 225854 46894
rect 225234 46574 225854 46658
rect 225234 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 225854 46574
rect 225234 10894 225854 46338
rect 225234 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 225854 10894
rect 225234 10574 225854 10658
rect 225234 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 225854 10574
rect 225234 -4186 225854 10338
rect 225234 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 225854 -4186
rect 225234 -4506 225854 -4422
rect 225234 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 225854 -4506
rect 225234 -5734 225854 -4742
rect 228954 86614 229574 98000
rect 228954 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 229574 86614
rect 228954 86294 229574 86378
rect 228954 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 229574 86294
rect 228954 50614 229574 86058
rect 228954 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 229574 50614
rect 228954 50294 229574 50378
rect 228954 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 229574 50294
rect 228954 14614 229574 50058
rect 228954 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 229574 14614
rect 228954 14294 229574 14378
rect 228954 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 229574 14294
rect 210954 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 211574 -7066
rect 210954 -7386 211574 -7302
rect 210954 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 211574 -7386
rect 210954 -7654 211574 -7622
rect 228954 -6106 229574 14058
rect 235794 93454 236414 98000
rect 235794 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 236414 93454
rect 235794 93134 236414 93218
rect 235794 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 236414 93134
rect 235794 57454 236414 92898
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -1306 236414 20898
rect 235794 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 236414 -1306
rect 235794 -1626 236414 -1542
rect 235794 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 236414 -1626
rect 235794 -1894 236414 -1862
rect 239514 97174 240134 98000
rect 239514 96938 239546 97174
rect 239782 96938 239866 97174
rect 240102 96938 240134 97174
rect 239514 96854 240134 96938
rect 239514 96618 239546 96854
rect 239782 96618 239866 96854
rect 240102 96618 240134 96854
rect 239514 61174 240134 96618
rect 239514 60938 239546 61174
rect 239782 60938 239866 61174
rect 240102 60938 240134 61174
rect 239514 60854 240134 60938
rect 239514 60618 239546 60854
rect 239782 60618 239866 60854
rect 240102 60618 240134 60854
rect 239514 25174 240134 60618
rect 239514 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 240134 25174
rect 239514 24854 240134 24938
rect 239514 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 240134 24854
rect 239514 -3226 240134 24618
rect 239514 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 240134 -3226
rect 239514 -3546 240134 -3462
rect 239514 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 240134 -3546
rect 239514 -3814 240134 -3782
rect 243234 64894 243854 98000
rect 243234 64658 243266 64894
rect 243502 64658 243586 64894
rect 243822 64658 243854 64894
rect 243234 64574 243854 64658
rect 243234 64338 243266 64574
rect 243502 64338 243586 64574
rect 243822 64338 243854 64574
rect 243234 28894 243854 64338
rect 243234 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 243854 28894
rect 243234 28574 243854 28658
rect 243234 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 243854 28574
rect 243234 -5146 243854 28338
rect 243234 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 243854 -5146
rect 243234 -5466 243854 -5382
rect 243234 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 243854 -5466
rect 243234 -5734 243854 -5702
rect 246954 68614 247574 98000
rect 246954 68378 246986 68614
rect 247222 68378 247306 68614
rect 247542 68378 247574 68614
rect 246954 68294 247574 68378
rect 246954 68058 246986 68294
rect 247222 68058 247306 68294
rect 247542 68058 247574 68294
rect 246954 32614 247574 68058
rect 246954 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 247574 32614
rect 246954 32294 247574 32378
rect 246954 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 247574 32294
rect 228954 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 229574 -6106
rect 228954 -6426 229574 -6342
rect 228954 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 229574 -6426
rect 228954 -7654 229574 -6662
rect 246954 -7066 247574 32058
rect 253794 75454 254414 98000
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253794 39454 254414 74898
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -1894 254414 -902
rect 257514 79174 258134 98000
rect 257514 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 258134 79174
rect 257514 78854 258134 78938
rect 257514 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 258134 78854
rect 257514 43174 258134 78618
rect 257514 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 258134 43174
rect 257514 42854 258134 42938
rect 257514 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 258134 42854
rect 257514 7174 258134 42618
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 257514 -2266 258134 6618
rect 257514 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 258134 -2266
rect 257514 -2586 258134 -2502
rect 257514 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 258134 -2586
rect 257514 -3814 258134 -2822
rect 261234 82894 261854 98000
rect 261234 82658 261266 82894
rect 261502 82658 261586 82894
rect 261822 82658 261854 82894
rect 261234 82574 261854 82658
rect 261234 82338 261266 82574
rect 261502 82338 261586 82574
rect 261822 82338 261854 82574
rect 261234 46894 261854 82338
rect 261234 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 261854 46894
rect 261234 46574 261854 46658
rect 261234 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 261854 46574
rect 261234 10894 261854 46338
rect 261234 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 261854 10894
rect 261234 10574 261854 10658
rect 261234 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 261854 10574
rect 261234 -4186 261854 10338
rect 261234 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 261854 -4186
rect 261234 -4506 261854 -4422
rect 261234 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 261854 -4506
rect 261234 -5734 261854 -4742
rect 264954 86614 265574 98000
rect 264954 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 265574 86614
rect 264954 86294 265574 86378
rect 264954 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 265574 86294
rect 264954 50614 265574 86058
rect 264954 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 265574 50614
rect 264954 50294 265574 50378
rect 264954 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 265574 50294
rect 264954 14614 265574 50058
rect 264954 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 265574 14614
rect 264954 14294 265574 14378
rect 264954 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 265574 14294
rect 246954 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 247574 -7066
rect 246954 -7386 247574 -7302
rect 246954 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 247574 -7386
rect 246954 -7654 247574 -7622
rect 264954 -6106 265574 14058
rect 271794 93454 272414 98000
rect 271794 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 272414 93454
rect 271794 93134 272414 93218
rect 271794 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 272414 93134
rect 271794 57454 272414 92898
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -1306 272414 20898
rect 271794 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 272414 -1306
rect 271794 -1626 272414 -1542
rect 271794 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 272414 -1626
rect 271794 -1894 272414 -1862
rect 275514 97174 276134 98000
rect 275514 96938 275546 97174
rect 275782 96938 275866 97174
rect 276102 96938 276134 97174
rect 275514 96854 276134 96938
rect 275514 96618 275546 96854
rect 275782 96618 275866 96854
rect 276102 96618 276134 96854
rect 275514 61174 276134 96618
rect 275514 60938 275546 61174
rect 275782 60938 275866 61174
rect 276102 60938 276134 61174
rect 275514 60854 276134 60938
rect 275514 60618 275546 60854
rect 275782 60618 275866 60854
rect 276102 60618 276134 60854
rect 275514 25174 276134 60618
rect 275514 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 276134 25174
rect 275514 24854 276134 24938
rect 275514 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 276134 24854
rect 275514 -3226 276134 24618
rect 275514 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 276134 -3226
rect 275514 -3546 276134 -3462
rect 275514 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 276134 -3546
rect 275514 -3814 276134 -3782
rect 279234 64894 279854 98000
rect 279234 64658 279266 64894
rect 279502 64658 279586 64894
rect 279822 64658 279854 64894
rect 279234 64574 279854 64658
rect 279234 64338 279266 64574
rect 279502 64338 279586 64574
rect 279822 64338 279854 64574
rect 279234 28894 279854 64338
rect 279234 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 279854 28894
rect 279234 28574 279854 28658
rect 279234 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 279854 28574
rect 279234 -5146 279854 28338
rect 279234 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 279854 -5146
rect 279234 -5466 279854 -5382
rect 279234 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 279854 -5466
rect 279234 -5734 279854 -5702
rect 282954 68614 283574 98000
rect 282954 68378 282986 68614
rect 283222 68378 283306 68614
rect 283542 68378 283574 68614
rect 282954 68294 283574 68378
rect 282954 68058 282986 68294
rect 283222 68058 283306 68294
rect 283542 68058 283574 68294
rect 282954 32614 283574 68058
rect 282954 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 283574 32614
rect 282954 32294 283574 32378
rect 282954 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 283574 32294
rect 264954 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 265574 -6106
rect 264954 -6426 265574 -6342
rect 264954 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 265574 -6426
rect 264954 -7654 265574 -6662
rect 282954 -7066 283574 32058
rect 289794 75454 290414 98000
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 289794 39454 290414 74898
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -1894 290414 -902
rect 293514 79174 294134 98000
rect 293514 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 294134 79174
rect 293514 78854 294134 78938
rect 293514 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 294134 78854
rect 293514 43174 294134 78618
rect 293514 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 294134 43174
rect 293514 42854 294134 42938
rect 293514 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 294134 42854
rect 293514 7174 294134 42618
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 293514 -2266 294134 6618
rect 293514 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 294134 -2266
rect 293514 -2586 294134 -2502
rect 293514 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 294134 -2586
rect 293514 -3814 294134 -2822
rect 297234 82894 297854 98000
rect 297234 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 297854 82894
rect 297234 82574 297854 82658
rect 297234 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 297854 82574
rect 297234 46894 297854 82338
rect 297234 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 297854 46894
rect 297234 46574 297854 46658
rect 297234 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 297854 46574
rect 297234 10894 297854 46338
rect 297234 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 297854 10894
rect 297234 10574 297854 10658
rect 297234 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 297854 10574
rect 297234 -4186 297854 10338
rect 297234 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 297854 -4186
rect 297234 -4506 297854 -4422
rect 297234 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 297854 -4506
rect 297234 -5734 297854 -4742
rect 300954 86614 301574 98000
rect 300954 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 301574 86614
rect 300954 86294 301574 86378
rect 300954 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 301574 86294
rect 300954 50614 301574 86058
rect 300954 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 301574 50614
rect 300954 50294 301574 50378
rect 300954 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 301574 50294
rect 300954 14614 301574 50058
rect 300954 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 301574 14614
rect 300954 14294 301574 14378
rect 300954 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 301574 14294
rect 282954 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 283574 -7066
rect 282954 -7386 283574 -7302
rect 282954 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 283574 -7386
rect 282954 -7654 283574 -7622
rect 300954 -6106 301574 14058
rect 307794 93454 308414 128898
rect 307794 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 308414 93454
rect 307794 93134 308414 93218
rect 307794 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 308414 93134
rect 307794 57454 308414 92898
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -1306 308414 20898
rect 307794 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 308414 -1306
rect 307794 -1626 308414 -1542
rect 307794 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 308414 -1626
rect 307794 -1894 308414 -1862
rect 311514 673174 312134 707162
rect 311514 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 312134 673174
rect 311514 672854 312134 672938
rect 311514 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 312134 672854
rect 311514 637174 312134 672618
rect 311514 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 312134 637174
rect 311514 636854 312134 636938
rect 311514 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 312134 636854
rect 311514 601174 312134 636618
rect 311514 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 312134 601174
rect 311514 600854 312134 600938
rect 311514 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 312134 600854
rect 311514 565174 312134 600618
rect 311514 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 312134 565174
rect 311514 564854 312134 564938
rect 311514 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 312134 564854
rect 311514 529174 312134 564618
rect 311514 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 312134 529174
rect 311514 528854 312134 528938
rect 311514 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 312134 528854
rect 311514 493174 312134 528618
rect 311514 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 312134 493174
rect 311514 492854 312134 492938
rect 311514 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 312134 492854
rect 311514 457174 312134 492618
rect 311514 456938 311546 457174
rect 311782 456938 311866 457174
rect 312102 456938 312134 457174
rect 311514 456854 312134 456938
rect 311514 456618 311546 456854
rect 311782 456618 311866 456854
rect 312102 456618 312134 456854
rect 311514 421174 312134 456618
rect 311514 420938 311546 421174
rect 311782 420938 311866 421174
rect 312102 420938 312134 421174
rect 311514 420854 312134 420938
rect 311514 420618 311546 420854
rect 311782 420618 311866 420854
rect 312102 420618 312134 420854
rect 311514 385174 312134 420618
rect 311514 384938 311546 385174
rect 311782 384938 311866 385174
rect 312102 384938 312134 385174
rect 311514 384854 312134 384938
rect 311514 384618 311546 384854
rect 311782 384618 311866 384854
rect 312102 384618 312134 384854
rect 311514 349174 312134 384618
rect 311514 348938 311546 349174
rect 311782 348938 311866 349174
rect 312102 348938 312134 349174
rect 311514 348854 312134 348938
rect 311514 348618 311546 348854
rect 311782 348618 311866 348854
rect 312102 348618 312134 348854
rect 311514 313174 312134 348618
rect 311514 312938 311546 313174
rect 311782 312938 311866 313174
rect 312102 312938 312134 313174
rect 311514 312854 312134 312938
rect 311514 312618 311546 312854
rect 311782 312618 311866 312854
rect 312102 312618 312134 312854
rect 311514 277174 312134 312618
rect 311514 276938 311546 277174
rect 311782 276938 311866 277174
rect 312102 276938 312134 277174
rect 311514 276854 312134 276938
rect 311514 276618 311546 276854
rect 311782 276618 311866 276854
rect 312102 276618 312134 276854
rect 311514 241174 312134 276618
rect 311514 240938 311546 241174
rect 311782 240938 311866 241174
rect 312102 240938 312134 241174
rect 311514 240854 312134 240938
rect 311514 240618 311546 240854
rect 311782 240618 311866 240854
rect 312102 240618 312134 240854
rect 311514 205174 312134 240618
rect 311514 204938 311546 205174
rect 311782 204938 311866 205174
rect 312102 204938 312134 205174
rect 311514 204854 312134 204938
rect 311514 204618 311546 204854
rect 311782 204618 311866 204854
rect 312102 204618 312134 204854
rect 311514 169174 312134 204618
rect 311514 168938 311546 169174
rect 311782 168938 311866 169174
rect 312102 168938 312134 169174
rect 311514 168854 312134 168938
rect 311514 168618 311546 168854
rect 311782 168618 311866 168854
rect 312102 168618 312134 168854
rect 311514 133174 312134 168618
rect 311514 132938 311546 133174
rect 311782 132938 311866 133174
rect 312102 132938 312134 133174
rect 311514 132854 312134 132938
rect 311514 132618 311546 132854
rect 311782 132618 311866 132854
rect 312102 132618 312134 132854
rect 311514 97174 312134 132618
rect 311514 96938 311546 97174
rect 311782 96938 311866 97174
rect 312102 96938 312134 97174
rect 311514 96854 312134 96938
rect 311514 96618 311546 96854
rect 311782 96618 311866 96854
rect 312102 96618 312134 96854
rect 311514 61174 312134 96618
rect 311514 60938 311546 61174
rect 311782 60938 311866 61174
rect 312102 60938 312134 61174
rect 311514 60854 312134 60938
rect 311514 60618 311546 60854
rect 311782 60618 311866 60854
rect 312102 60618 312134 60854
rect 311514 25174 312134 60618
rect 311514 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 312134 25174
rect 311514 24854 312134 24938
rect 311514 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 312134 24854
rect 311514 -3226 312134 24618
rect 311514 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 312134 -3226
rect 311514 -3546 312134 -3462
rect 311514 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 312134 -3546
rect 311514 -3814 312134 -3782
rect 315234 676894 315854 709082
rect 315234 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 315854 676894
rect 315234 676574 315854 676658
rect 315234 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 315854 676574
rect 315234 640894 315854 676338
rect 315234 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 315854 640894
rect 315234 640574 315854 640658
rect 315234 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 315854 640574
rect 315234 604894 315854 640338
rect 315234 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 315854 604894
rect 315234 604574 315854 604658
rect 315234 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 315854 604574
rect 315234 568894 315854 604338
rect 315234 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 315854 568894
rect 315234 568574 315854 568658
rect 315234 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 315854 568574
rect 315234 532894 315854 568338
rect 315234 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 315854 532894
rect 315234 532574 315854 532658
rect 315234 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 315854 532574
rect 315234 496894 315854 532338
rect 315234 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 315854 496894
rect 315234 496574 315854 496658
rect 315234 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 315854 496574
rect 315234 460894 315854 496338
rect 315234 460658 315266 460894
rect 315502 460658 315586 460894
rect 315822 460658 315854 460894
rect 315234 460574 315854 460658
rect 315234 460338 315266 460574
rect 315502 460338 315586 460574
rect 315822 460338 315854 460574
rect 315234 424894 315854 460338
rect 315234 424658 315266 424894
rect 315502 424658 315586 424894
rect 315822 424658 315854 424894
rect 315234 424574 315854 424658
rect 315234 424338 315266 424574
rect 315502 424338 315586 424574
rect 315822 424338 315854 424574
rect 315234 388894 315854 424338
rect 315234 388658 315266 388894
rect 315502 388658 315586 388894
rect 315822 388658 315854 388894
rect 315234 388574 315854 388658
rect 315234 388338 315266 388574
rect 315502 388338 315586 388574
rect 315822 388338 315854 388574
rect 315234 352894 315854 388338
rect 315234 352658 315266 352894
rect 315502 352658 315586 352894
rect 315822 352658 315854 352894
rect 315234 352574 315854 352658
rect 315234 352338 315266 352574
rect 315502 352338 315586 352574
rect 315822 352338 315854 352574
rect 315234 316894 315854 352338
rect 315234 316658 315266 316894
rect 315502 316658 315586 316894
rect 315822 316658 315854 316894
rect 315234 316574 315854 316658
rect 315234 316338 315266 316574
rect 315502 316338 315586 316574
rect 315822 316338 315854 316574
rect 315234 280894 315854 316338
rect 315234 280658 315266 280894
rect 315502 280658 315586 280894
rect 315822 280658 315854 280894
rect 315234 280574 315854 280658
rect 315234 280338 315266 280574
rect 315502 280338 315586 280574
rect 315822 280338 315854 280574
rect 315234 244894 315854 280338
rect 315234 244658 315266 244894
rect 315502 244658 315586 244894
rect 315822 244658 315854 244894
rect 315234 244574 315854 244658
rect 315234 244338 315266 244574
rect 315502 244338 315586 244574
rect 315822 244338 315854 244574
rect 315234 208894 315854 244338
rect 315234 208658 315266 208894
rect 315502 208658 315586 208894
rect 315822 208658 315854 208894
rect 315234 208574 315854 208658
rect 315234 208338 315266 208574
rect 315502 208338 315586 208574
rect 315822 208338 315854 208574
rect 315234 172894 315854 208338
rect 315234 172658 315266 172894
rect 315502 172658 315586 172894
rect 315822 172658 315854 172894
rect 315234 172574 315854 172658
rect 315234 172338 315266 172574
rect 315502 172338 315586 172574
rect 315822 172338 315854 172574
rect 315234 136894 315854 172338
rect 315234 136658 315266 136894
rect 315502 136658 315586 136894
rect 315822 136658 315854 136894
rect 315234 136574 315854 136658
rect 315234 136338 315266 136574
rect 315502 136338 315586 136574
rect 315822 136338 315854 136574
rect 315234 100894 315854 136338
rect 315234 100658 315266 100894
rect 315502 100658 315586 100894
rect 315822 100658 315854 100894
rect 315234 100574 315854 100658
rect 315234 100338 315266 100574
rect 315502 100338 315586 100574
rect 315822 100338 315854 100574
rect 315234 64894 315854 100338
rect 315234 64658 315266 64894
rect 315502 64658 315586 64894
rect 315822 64658 315854 64894
rect 315234 64574 315854 64658
rect 315234 64338 315266 64574
rect 315502 64338 315586 64574
rect 315822 64338 315854 64574
rect 315234 28894 315854 64338
rect 315234 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 315854 28894
rect 315234 28574 315854 28658
rect 315234 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 315854 28574
rect 315234 -5146 315854 28338
rect 315234 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 315854 -5146
rect 315234 -5466 315854 -5382
rect 315234 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 315854 -5466
rect 315234 -5734 315854 -5702
rect 318954 680614 319574 711002
rect 336954 710598 337574 711590
rect 336954 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 337574 710598
rect 336954 710278 337574 710362
rect 336954 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 337574 710278
rect 333234 708678 333854 709670
rect 333234 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 333854 708678
rect 333234 708358 333854 708442
rect 333234 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 333854 708358
rect 329514 706758 330134 707750
rect 329514 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 330134 706758
rect 329514 706438 330134 706522
rect 329514 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 330134 706438
rect 318954 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 319574 680614
rect 318954 680294 319574 680378
rect 318954 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 319574 680294
rect 318954 644614 319574 680058
rect 318954 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 319574 644614
rect 318954 644294 319574 644378
rect 318954 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 319574 644294
rect 318954 608614 319574 644058
rect 318954 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 319574 608614
rect 318954 608294 319574 608378
rect 318954 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 319574 608294
rect 318954 572614 319574 608058
rect 318954 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 319574 572614
rect 318954 572294 319574 572378
rect 318954 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 319574 572294
rect 318954 536614 319574 572058
rect 318954 536378 318986 536614
rect 319222 536378 319306 536614
rect 319542 536378 319574 536614
rect 318954 536294 319574 536378
rect 318954 536058 318986 536294
rect 319222 536058 319306 536294
rect 319542 536058 319574 536294
rect 318954 500614 319574 536058
rect 318954 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 319574 500614
rect 318954 500294 319574 500378
rect 318954 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 319574 500294
rect 318954 464614 319574 500058
rect 318954 464378 318986 464614
rect 319222 464378 319306 464614
rect 319542 464378 319574 464614
rect 318954 464294 319574 464378
rect 318954 464058 318986 464294
rect 319222 464058 319306 464294
rect 319542 464058 319574 464294
rect 318954 428614 319574 464058
rect 318954 428378 318986 428614
rect 319222 428378 319306 428614
rect 319542 428378 319574 428614
rect 318954 428294 319574 428378
rect 318954 428058 318986 428294
rect 319222 428058 319306 428294
rect 319542 428058 319574 428294
rect 318954 392614 319574 428058
rect 318954 392378 318986 392614
rect 319222 392378 319306 392614
rect 319542 392378 319574 392614
rect 318954 392294 319574 392378
rect 318954 392058 318986 392294
rect 319222 392058 319306 392294
rect 319542 392058 319574 392294
rect 318954 356614 319574 392058
rect 318954 356378 318986 356614
rect 319222 356378 319306 356614
rect 319542 356378 319574 356614
rect 318954 356294 319574 356378
rect 318954 356058 318986 356294
rect 319222 356058 319306 356294
rect 319542 356058 319574 356294
rect 318954 320614 319574 356058
rect 318954 320378 318986 320614
rect 319222 320378 319306 320614
rect 319542 320378 319574 320614
rect 318954 320294 319574 320378
rect 318954 320058 318986 320294
rect 319222 320058 319306 320294
rect 319542 320058 319574 320294
rect 318954 284614 319574 320058
rect 318954 284378 318986 284614
rect 319222 284378 319306 284614
rect 319542 284378 319574 284614
rect 318954 284294 319574 284378
rect 318954 284058 318986 284294
rect 319222 284058 319306 284294
rect 319542 284058 319574 284294
rect 318954 248614 319574 284058
rect 318954 248378 318986 248614
rect 319222 248378 319306 248614
rect 319542 248378 319574 248614
rect 318954 248294 319574 248378
rect 318954 248058 318986 248294
rect 319222 248058 319306 248294
rect 319542 248058 319574 248294
rect 318954 212614 319574 248058
rect 318954 212378 318986 212614
rect 319222 212378 319306 212614
rect 319542 212378 319574 212614
rect 318954 212294 319574 212378
rect 318954 212058 318986 212294
rect 319222 212058 319306 212294
rect 319542 212058 319574 212294
rect 318954 176614 319574 212058
rect 318954 176378 318986 176614
rect 319222 176378 319306 176614
rect 319542 176378 319574 176614
rect 318954 176294 319574 176378
rect 318954 176058 318986 176294
rect 319222 176058 319306 176294
rect 319542 176058 319574 176294
rect 318954 140614 319574 176058
rect 318954 140378 318986 140614
rect 319222 140378 319306 140614
rect 319542 140378 319574 140614
rect 318954 140294 319574 140378
rect 318954 140058 318986 140294
rect 319222 140058 319306 140294
rect 319542 140058 319574 140294
rect 318954 104614 319574 140058
rect 318954 104378 318986 104614
rect 319222 104378 319306 104614
rect 319542 104378 319574 104614
rect 318954 104294 319574 104378
rect 318954 104058 318986 104294
rect 319222 104058 319306 104294
rect 319542 104058 319574 104294
rect 318954 68614 319574 104058
rect 318954 68378 318986 68614
rect 319222 68378 319306 68614
rect 319542 68378 319574 68614
rect 318954 68294 319574 68378
rect 318954 68058 318986 68294
rect 319222 68058 319306 68294
rect 319542 68058 319574 68294
rect 318954 32614 319574 68058
rect 318954 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 319574 32614
rect 318954 32294 319574 32378
rect 318954 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 319574 32294
rect 300954 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 301574 -6106
rect 300954 -6426 301574 -6342
rect 300954 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 301574 -6426
rect 300954 -7654 301574 -6662
rect 318954 -7066 319574 32058
rect 325794 704838 326414 705830
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 543454 326414 578898
rect 325794 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 326414 543454
rect 325794 543134 326414 543218
rect 325794 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 326414 543134
rect 325794 507454 326414 542898
rect 325794 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 326414 507454
rect 325794 507134 326414 507218
rect 325794 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 326414 507134
rect 325794 471454 326414 506898
rect 325794 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 326414 471454
rect 325794 471134 326414 471218
rect 325794 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 326414 471134
rect 325794 435454 326414 470898
rect 325794 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 326414 435454
rect 325794 435134 326414 435218
rect 325794 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 326414 435134
rect 325794 399454 326414 434898
rect 325794 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 326414 399454
rect 325794 399134 326414 399218
rect 325794 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 326414 399134
rect 325794 363454 326414 398898
rect 325794 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 326414 363454
rect 325794 363134 326414 363218
rect 325794 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 326414 363134
rect 325794 327454 326414 362898
rect 325794 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 326414 327454
rect 325794 327134 326414 327218
rect 325794 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 326414 327134
rect 325794 291454 326414 326898
rect 325794 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 326414 291454
rect 325794 291134 326414 291218
rect 325794 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 326414 291134
rect 325794 255454 326414 290898
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 325794 219454 326414 254898
rect 325794 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 326414 219454
rect 325794 219134 326414 219218
rect 325794 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 326414 219134
rect 325794 183454 326414 218898
rect 325794 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 326414 183454
rect 325794 183134 326414 183218
rect 325794 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 326414 183134
rect 325794 147454 326414 182898
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 325794 111454 326414 146898
rect 325794 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 326414 111454
rect 325794 111134 326414 111218
rect 325794 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 326414 111134
rect 325794 75454 326414 110898
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -1894 326414 -902
rect 329514 691174 330134 706202
rect 329514 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 330134 691174
rect 329514 690854 330134 690938
rect 329514 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 330134 690854
rect 329514 655174 330134 690618
rect 329514 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 330134 655174
rect 329514 654854 330134 654938
rect 329514 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 330134 654854
rect 329514 619174 330134 654618
rect 329514 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 330134 619174
rect 329514 618854 330134 618938
rect 329514 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 330134 618854
rect 329514 583174 330134 618618
rect 329514 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 330134 583174
rect 329514 582854 330134 582938
rect 329514 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 330134 582854
rect 329514 547174 330134 582618
rect 329514 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 330134 547174
rect 329514 546854 330134 546938
rect 329514 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 330134 546854
rect 329514 511174 330134 546618
rect 329514 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 330134 511174
rect 329514 510854 330134 510938
rect 329514 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 330134 510854
rect 329514 475174 330134 510618
rect 329514 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 330134 475174
rect 329514 474854 330134 474938
rect 329514 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 330134 474854
rect 329514 439174 330134 474618
rect 329514 438938 329546 439174
rect 329782 438938 329866 439174
rect 330102 438938 330134 439174
rect 329514 438854 330134 438938
rect 329514 438618 329546 438854
rect 329782 438618 329866 438854
rect 330102 438618 330134 438854
rect 329514 403174 330134 438618
rect 329514 402938 329546 403174
rect 329782 402938 329866 403174
rect 330102 402938 330134 403174
rect 329514 402854 330134 402938
rect 329514 402618 329546 402854
rect 329782 402618 329866 402854
rect 330102 402618 330134 402854
rect 329514 367174 330134 402618
rect 329514 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 330134 367174
rect 329514 366854 330134 366938
rect 329514 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 330134 366854
rect 329514 331174 330134 366618
rect 329514 330938 329546 331174
rect 329782 330938 329866 331174
rect 330102 330938 330134 331174
rect 329514 330854 330134 330938
rect 329514 330618 329546 330854
rect 329782 330618 329866 330854
rect 330102 330618 330134 330854
rect 329514 295174 330134 330618
rect 329514 294938 329546 295174
rect 329782 294938 329866 295174
rect 330102 294938 330134 295174
rect 329514 294854 330134 294938
rect 329514 294618 329546 294854
rect 329782 294618 329866 294854
rect 330102 294618 330134 294854
rect 329514 259174 330134 294618
rect 329514 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 330134 259174
rect 329514 258854 330134 258938
rect 329514 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 330134 258854
rect 329514 223174 330134 258618
rect 329514 222938 329546 223174
rect 329782 222938 329866 223174
rect 330102 222938 330134 223174
rect 329514 222854 330134 222938
rect 329514 222618 329546 222854
rect 329782 222618 329866 222854
rect 330102 222618 330134 222854
rect 329514 187174 330134 222618
rect 329514 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 330134 187174
rect 329514 186854 330134 186938
rect 329514 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 330134 186854
rect 329514 151174 330134 186618
rect 329514 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 330134 151174
rect 329514 150854 330134 150938
rect 329514 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 330134 150854
rect 329514 115174 330134 150618
rect 329514 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 330134 115174
rect 329514 114854 330134 114938
rect 329514 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 330134 114854
rect 329514 79174 330134 114618
rect 329514 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 330134 79174
rect 329514 78854 330134 78938
rect 329514 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 330134 78854
rect 329514 43174 330134 78618
rect 329514 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 330134 43174
rect 329514 42854 330134 42938
rect 329514 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 330134 42854
rect 329514 7174 330134 42618
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 329514 -2266 330134 6618
rect 329514 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 330134 -2266
rect 329514 -2586 330134 -2502
rect 329514 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 330134 -2586
rect 329514 -3814 330134 -2822
rect 333234 694894 333854 708122
rect 333234 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 333854 694894
rect 333234 694574 333854 694658
rect 333234 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 333854 694574
rect 333234 658894 333854 694338
rect 333234 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 333854 658894
rect 333234 658574 333854 658658
rect 333234 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 333854 658574
rect 333234 622894 333854 658338
rect 333234 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 333854 622894
rect 333234 622574 333854 622658
rect 333234 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 333854 622574
rect 333234 586894 333854 622338
rect 333234 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 333854 586894
rect 333234 586574 333854 586658
rect 333234 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 333854 586574
rect 333234 550894 333854 586338
rect 333234 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 333854 550894
rect 333234 550574 333854 550658
rect 333234 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 333854 550574
rect 333234 514894 333854 550338
rect 333234 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 333854 514894
rect 333234 514574 333854 514658
rect 333234 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 333854 514574
rect 333234 478894 333854 514338
rect 333234 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 333854 478894
rect 333234 478574 333854 478658
rect 333234 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 333854 478574
rect 333234 442894 333854 478338
rect 333234 442658 333266 442894
rect 333502 442658 333586 442894
rect 333822 442658 333854 442894
rect 333234 442574 333854 442658
rect 333234 442338 333266 442574
rect 333502 442338 333586 442574
rect 333822 442338 333854 442574
rect 333234 406894 333854 442338
rect 333234 406658 333266 406894
rect 333502 406658 333586 406894
rect 333822 406658 333854 406894
rect 333234 406574 333854 406658
rect 333234 406338 333266 406574
rect 333502 406338 333586 406574
rect 333822 406338 333854 406574
rect 333234 370894 333854 406338
rect 333234 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 333854 370894
rect 333234 370574 333854 370658
rect 333234 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 333854 370574
rect 333234 334894 333854 370338
rect 333234 334658 333266 334894
rect 333502 334658 333586 334894
rect 333822 334658 333854 334894
rect 333234 334574 333854 334658
rect 333234 334338 333266 334574
rect 333502 334338 333586 334574
rect 333822 334338 333854 334574
rect 333234 298894 333854 334338
rect 333234 298658 333266 298894
rect 333502 298658 333586 298894
rect 333822 298658 333854 298894
rect 333234 298574 333854 298658
rect 333234 298338 333266 298574
rect 333502 298338 333586 298574
rect 333822 298338 333854 298574
rect 333234 262894 333854 298338
rect 333234 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 333854 262894
rect 333234 262574 333854 262658
rect 333234 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 333854 262574
rect 333234 226894 333854 262338
rect 333234 226658 333266 226894
rect 333502 226658 333586 226894
rect 333822 226658 333854 226894
rect 333234 226574 333854 226658
rect 333234 226338 333266 226574
rect 333502 226338 333586 226574
rect 333822 226338 333854 226574
rect 333234 190894 333854 226338
rect 333234 190658 333266 190894
rect 333502 190658 333586 190894
rect 333822 190658 333854 190894
rect 333234 190574 333854 190658
rect 333234 190338 333266 190574
rect 333502 190338 333586 190574
rect 333822 190338 333854 190574
rect 333234 154894 333854 190338
rect 333234 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 333854 154894
rect 333234 154574 333854 154658
rect 333234 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 333854 154574
rect 333234 118894 333854 154338
rect 333234 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 333854 118894
rect 333234 118574 333854 118658
rect 333234 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 333854 118574
rect 333234 82894 333854 118338
rect 333234 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 333854 82894
rect 333234 82574 333854 82658
rect 333234 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 333854 82574
rect 333234 46894 333854 82338
rect 333234 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 333854 46894
rect 333234 46574 333854 46658
rect 333234 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 333854 46574
rect 333234 10894 333854 46338
rect 333234 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 333854 10894
rect 333234 10574 333854 10658
rect 333234 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 333854 10574
rect 333234 -4186 333854 10338
rect 333234 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 333854 -4186
rect 333234 -4506 333854 -4422
rect 333234 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 333854 -4506
rect 333234 -5734 333854 -4742
rect 336954 698614 337574 710042
rect 354954 711558 355574 711590
rect 354954 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 355574 711558
rect 354954 711238 355574 711322
rect 354954 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 355574 711238
rect 351234 709638 351854 709670
rect 351234 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 351854 709638
rect 351234 709318 351854 709402
rect 351234 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 351854 709318
rect 347514 707718 348134 707750
rect 347514 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 348134 707718
rect 347514 707398 348134 707482
rect 347514 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 348134 707398
rect 336954 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 337574 698614
rect 336954 698294 337574 698378
rect 336954 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 337574 698294
rect 336954 662614 337574 698058
rect 336954 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 337574 662614
rect 336954 662294 337574 662378
rect 336954 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 337574 662294
rect 336954 626614 337574 662058
rect 336954 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 337574 626614
rect 336954 626294 337574 626378
rect 336954 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 337574 626294
rect 336954 590614 337574 626058
rect 336954 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 337574 590614
rect 336954 590294 337574 590378
rect 336954 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 337574 590294
rect 336954 554614 337574 590058
rect 336954 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 337574 554614
rect 336954 554294 337574 554378
rect 336954 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 337574 554294
rect 336954 518614 337574 554058
rect 336954 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 337574 518614
rect 336954 518294 337574 518378
rect 336954 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 337574 518294
rect 336954 482614 337574 518058
rect 336954 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 337574 482614
rect 336954 482294 337574 482378
rect 336954 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 337574 482294
rect 336954 446614 337574 482058
rect 336954 446378 336986 446614
rect 337222 446378 337306 446614
rect 337542 446378 337574 446614
rect 336954 446294 337574 446378
rect 336954 446058 336986 446294
rect 337222 446058 337306 446294
rect 337542 446058 337574 446294
rect 336954 410614 337574 446058
rect 336954 410378 336986 410614
rect 337222 410378 337306 410614
rect 337542 410378 337574 410614
rect 336954 410294 337574 410378
rect 336954 410058 336986 410294
rect 337222 410058 337306 410294
rect 337542 410058 337574 410294
rect 336954 374614 337574 410058
rect 336954 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 337574 374614
rect 336954 374294 337574 374378
rect 336954 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 337574 374294
rect 336954 338614 337574 374058
rect 336954 338378 336986 338614
rect 337222 338378 337306 338614
rect 337542 338378 337574 338614
rect 336954 338294 337574 338378
rect 336954 338058 336986 338294
rect 337222 338058 337306 338294
rect 337542 338058 337574 338294
rect 336954 302614 337574 338058
rect 336954 302378 336986 302614
rect 337222 302378 337306 302614
rect 337542 302378 337574 302614
rect 336954 302294 337574 302378
rect 336954 302058 336986 302294
rect 337222 302058 337306 302294
rect 337542 302058 337574 302294
rect 336954 266614 337574 302058
rect 336954 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 337574 266614
rect 336954 266294 337574 266378
rect 336954 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 337574 266294
rect 336954 230614 337574 266058
rect 336954 230378 336986 230614
rect 337222 230378 337306 230614
rect 337542 230378 337574 230614
rect 336954 230294 337574 230378
rect 336954 230058 336986 230294
rect 337222 230058 337306 230294
rect 337542 230058 337574 230294
rect 336954 194614 337574 230058
rect 336954 194378 336986 194614
rect 337222 194378 337306 194614
rect 337542 194378 337574 194614
rect 336954 194294 337574 194378
rect 336954 194058 336986 194294
rect 337222 194058 337306 194294
rect 337542 194058 337574 194294
rect 336954 158614 337574 194058
rect 336954 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 337574 158614
rect 336954 158294 337574 158378
rect 336954 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 337574 158294
rect 336954 122614 337574 158058
rect 336954 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 337574 122614
rect 336954 122294 337574 122378
rect 336954 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 337574 122294
rect 336954 86614 337574 122058
rect 336954 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 337574 86614
rect 336954 86294 337574 86378
rect 336954 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 337574 86294
rect 336954 50614 337574 86058
rect 336954 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 337574 50614
rect 336954 50294 337574 50378
rect 336954 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 337574 50294
rect 336954 14614 337574 50058
rect 336954 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 337574 14614
rect 336954 14294 337574 14378
rect 336954 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 337574 14294
rect 318954 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 319574 -7066
rect 318954 -7386 319574 -7302
rect 318954 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 319574 -7386
rect 318954 -7654 319574 -7622
rect 336954 -6106 337574 14058
rect 343794 705798 344414 705830
rect 343794 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 344414 705798
rect 343794 705478 344414 705562
rect 343794 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 344414 705478
rect 343794 669454 344414 705242
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 561454 344414 596898
rect 343794 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 344414 561454
rect 343794 561134 344414 561218
rect 343794 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 344414 561134
rect 343794 525454 344414 560898
rect 343794 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 344414 525454
rect 343794 525134 344414 525218
rect 343794 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 344414 525134
rect 343794 489454 344414 524898
rect 343794 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 344414 489454
rect 343794 489134 344414 489218
rect 343794 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 344414 489134
rect 343794 453454 344414 488898
rect 343794 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 344414 453454
rect 343794 453134 344414 453218
rect 343794 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 344414 453134
rect 343794 417454 344414 452898
rect 343794 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 344414 417454
rect 343794 417134 344414 417218
rect 343794 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 344414 417134
rect 343794 381454 344414 416898
rect 343794 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 344414 381454
rect 343794 381134 344414 381218
rect 343794 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 344414 381134
rect 343794 345454 344414 380898
rect 343794 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 344414 345454
rect 343794 345134 344414 345218
rect 343794 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 344414 345134
rect 343794 309454 344414 344898
rect 343794 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 344414 309454
rect 343794 309134 344414 309218
rect 343794 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 344414 309134
rect 343794 273454 344414 308898
rect 343794 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 344414 273454
rect 343794 273134 344414 273218
rect 343794 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 344414 273134
rect 343794 237454 344414 272898
rect 343794 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 344414 237454
rect 343794 237134 344414 237218
rect 343794 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 344414 237134
rect 343794 201454 344414 236898
rect 343794 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 344414 201454
rect 343794 201134 344414 201218
rect 343794 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 344414 201134
rect 343794 165454 344414 200898
rect 343794 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 344414 165454
rect 343794 165134 344414 165218
rect 343794 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 344414 165134
rect 343794 129454 344414 164898
rect 343794 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 344414 129454
rect 343794 129134 344414 129218
rect 343794 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 344414 129134
rect 343794 93454 344414 128898
rect 343794 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 344414 93454
rect 343794 93134 344414 93218
rect 343794 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 344414 93134
rect 343794 57454 344414 92898
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -1306 344414 20898
rect 343794 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 344414 -1306
rect 343794 -1626 344414 -1542
rect 343794 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 344414 -1626
rect 343794 -1894 344414 -1862
rect 347514 673174 348134 707162
rect 347514 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 348134 673174
rect 347514 672854 348134 672938
rect 347514 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 348134 672854
rect 347514 637174 348134 672618
rect 347514 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 348134 637174
rect 347514 636854 348134 636938
rect 347514 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 348134 636854
rect 347514 601174 348134 636618
rect 347514 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 348134 601174
rect 347514 600854 348134 600938
rect 347514 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 348134 600854
rect 347514 565174 348134 600618
rect 347514 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 348134 565174
rect 347514 564854 348134 564938
rect 347514 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 348134 564854
rect 347514 529174 348134 564618
rect 347514 528938 347546 529174
rect 347782 528938 347866 529174
rect 348102 528938 348134 529174
rect 347514 528854 348134 528938
rect 347514 528618 347546 528854
rect 347782 528618 347866 528854
rect 348102 528618 348134 528854
rect 347514 493174 348134 528618
rect 347514 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 348134 493174
rect 347514 492854 348134 492938
rect 347514 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 348134 492854
rect 347514 457174 348134 492618
rect 347514 456938 347546 457174
rect 347782 456938 347866 457174
rect 348102 456938 348134 457174
rect 347514 456854 348134 456938
rect 347514 456618 347546 456854
rect 347782 456618 347866 456854
rect 348102 456618 348134 456854
rect 347514 421174 348134 456618
rect 347514 420938 347546 421174
rect 347782 420938 347866 421174
rect 348102 420938 348134 421174
rect 347514 420854 348134 420938
rect 347514 420618 347546 420854
rect 347782 420618 347866 420854
rect 348102 420618 348134 420854
rect 347514 385174 348134 420618
rect 347514 384938 347546 385174
rect 347782 384938 347866 385174
rect 348102 384938 348134 385174
rect 347514 384854 348134 384938
rect 347514 384618 347546 384854
rect 347782 384618 347866 384854
rect 348102 384618 348134 384854
rect 347514 349174 348134 384618
rect 347514 348938 347546 349174
rect 347782 348938 347866 349174
rect 348102 348938 348134 349174
rect 347514 348854 348134 348938
rect 347514 348618 347546 348854
rect 347782 348618 347866 348854
rect 348102 348618 348134 348854
rect 347514 313174 348134 348618
rect 347514 312938 347546 313174
rect 347782 312938 347866 313174
rect 348102 312938 348134 313174
rect 347514 312854 348134 312938
rect 347514 312618 347546 312854
rect 347782 312618 347866 312854
rect 348102 312618 348134 312854
rect 347514 277174 348134 312618
rect 347514 276938 347546 277174
rect 347782 276938 347866 277174
rect 348102 276938 348134 277174
rect 347514 276854 348134 276938
rect 347514 276618 347546 276854
rect 347782 276618 347866 276854
rect 348102 276618 348134 276854
rect 347514 241174 348134 276618
rect 347514 240938 347546 241174
rect 347782 240938 347866 241174
rect 348102 240938 348134 241174
rect 347514 240854 348134 240938
rect 347514 240618 347546 240854
rect 347782 240618 347866 240854
rect 348102 240618 348134 240854
rect 347514 205174 348134 240618
rect 347514 204938 347546 205174
rect 347782 204938 347866 205174
rect 348102 204938 348134 205174
rect 347514 204854 348134 204938
rect 347514 204618 347546 204854
rect 347782 204618 347866 204854
rect 348102 204618 348134 204854
rect 347514 169174 348134 204618
rect 347514 168938 347546 169174
rect 347782 168938 347866 169174
rect 348102 168938 348134 169174
rect 347514 168854 348134 168938
rect 347514 168618 347546 168854
rect 347782 168618 347866 168854
rect 348102 168618 348134 168854
rect 347514 133174 348134 168618
rect 347514 132938 347546 133174
rect 347782 132938 347866 133174
rect 348102 132938 348134 133174
rect 347514 132854 348134 132938
rect 347514 132618 347546 132854
rect 347782 132618 347866 132854
rect 348102 132618 348134 132854
rect 347514 97174 348134 132618
rect 347514 96938 347546 97174
rect 347782 96938 347866 97174
rect 348102 96938 348134 97174
rect 347514 96854 348134 96938
rect 347514 96618 347546 96854
rect 347782 96618 347866 96854
rect 348102 96618 348134 96854
rect 347514 61174 348134 96618
rect 347514 60938 347546 61174
rect 347782 60938 347866 61174
rect 348102 60938 348134 61174
rect 347514 60854 348134 60938
rect 347514 60618 347546 60854
rect 347782 60618 347866 60854
rect 348102 60618 348134 60854
rect 347514 25174 348134 60618
rect 347514 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 348134 25174
rect 347514 24854 348134 24938
rect 347514 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 348134 24854
rect 347514 -3226 348134 24618
rect 347514 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 348134 -3226
rect 347514 -3546 348134 -3462
rect 347514 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 348134 -3546
rect 347514 -3814 348134 -3782
rect 351234 676894 351854 709082
rect 351234 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 351854 676894
rect 351234 676574 351854 676658
rect 351234 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 351854 676574
rect 351234 640894 351854 676338
rect 351234 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 351854 640894
rect 351234 640574 351854 640658
rect 351234 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 351854 640574
rect 351234 604894 351854 640338
rect 351234 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 351854 604894
rect 351234 604574 351854 604658
rect 351234 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 351854 604574
rect 351234 568894 351854 604338
rect 351234 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 351854 568894
rect 351234 568574 351854 568658
rect 351234 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 351854 568574
rect 351234 532894 351854 568338
rect 351234 532658 351266 532894
rect 351502 532658 351586 532894
rect 351822 532658 351854 532894
rect 351234 532574 351854 532658
rect 351234 532338 351266 532574
rect 351502 532338 351586 532574
rect 351822 532338 351854 532574
rect 351234 496894 351854 532338
rect 351234 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 351854 496894
rect 351234 496574 351854 496658
rect 351234 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 351854 496574
rect 351234 460894 351854 496338
rect 351234 460658 351266 460894
rect 351502 460658 351586 460894
rect 351822 460658 351854 460894
rect 351234 460574 351854 460658
rect 351234 460338 351266 460574
rect 351502 460338 351586 460574
rect 351822 460338 351854 460574
rect 351234 424894 351854 460338
rect 351234 424658 351266 424894
rect 351502 424658 351586 424894
rect 351822 424658 351854 424894
rect 351234 424574 351854 424658
rect 351234 424338 351266 424574
rect 351502 424338 351586 424574
rect 351822 424338 351854 424574
rect 351234 388894 351854 424338
rect 351234 388658 351266 388894
rect 351502 388658 351586 388894
rect 351822 388658 351854 388894
rect 351234 388574 351854 388658
rect 351234 388338 351266 388574
rect 351502 388338 351586 388574
rect 351822 388338 351854 388574
rect 351234 352894 351854 388338
rect 351234 352658 351266 352894
rect 351502 352658 351586 352894
rect 351822 352658 351854 352894
rect 351234 352574 351854 352658
rect 351234 352338 351266 352574
rect 351502 352338 351586 352574
rect 351822 352338 351854 352574
rect 351234 316894 351854 352338
rect 351234 316658 351266 316894
rect 351502 316658 351586 316894
rect 351822 316658 351854 316894
rect 351234 316574 351854 316658
rect 351234 316338 351266 316574
rect 351502 316338 351586 316574
rect 351822 316338 351854 316574
rect 351234 280894 351854 316338
rect 351234 280658 351266 280894
rect 351502 280658 351586 280894
rect 351822 280658 351854 280894
rect 351234 280574 351854 280658
rect 351234 280338 351266 280574
rect 351502 280338 351586 280574
rect 351822 280338 351854 280574
rect 351234 244894 351854 280338
rect 351234 244658 351266 244894
rect 351502 244658 351586 244894
rect 351822 244658 351854 244894
rect 351234 244574 351854 244658
rect 351234 244338 351266 244574
rect 351502 244338 351586 244574
rect 351822 244338 351854 244574
rect 351234 208894 351854 244338
rect 351234 208658 351266 208894
rect 351502 208658 351586 208894
rect 351822 208658 351854 208894
rect 351234 208574 351854 208658
rect 351234 208338 351266 208574
rect 351502 208338 351586 208574
rect 351822 208338 351854 208574
rect 351234 172894 351854 208338
rect 351234 172658 351266 172894
rect 351502 172658 351586 172894
rect 351822 172658 351854 172894
rect 351234 172574 351854 172658
rect 351234 172338 351266 172574
rect 351502 172338 351586 172574
rect 351822 172338 351854 172574
rect 351234 136894 351854 172338
rect 351234 136658 351266 136894
rect 351502 136658 351586 136894
rect 351822 136658 351854 136894
rect 351234 136574 351854 136658
rect 351234 136338 351266 136574
rect 351502 136338 351586 136574
rect 351822 136338 351854 136574
rect 351234 100894 351854 136338
rect 351234 100658 351266 100894
rect 351502 100658 351586 100894
rect 351822 100658 351854 100894
rect 351234 100574 351854 100658
rect 351234 100338 351266 100574
rect 351502 100338 351586 100574
rect 351822 100338 351854 100574
rect 351234 64894 351854 100338
rect 351234 64658 351266 64894
rect 351502 64658 351586 64894
rect 351822 64658 351854 64894
rect 351234 64574 351854 64658
rect 351234 64338 351266 64574
rect 351502 64338 351586 64574
rect 351822 64338 351854 64574
rect 351234 28894 351854 64338
rect 351234 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 351854 28894
rect 351234 28574 351854 28658
rect 351234 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 351854 28574
rect 351234 -5146 351854 28338
rect 351234 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 351854 -5146
rect 351234 -5466 351854 -5382
rect 351234 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 351854 -5466
rect 351234 -5734 351854 -5702
rect 354954 680614 355574 711002
rect 372954 710598 373574 711590
rect 372954 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 373574 710598
rect 372954 710278 373574 710362
rect 372954 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 373574 710278
rect 369234 708678 369854 709670
rect 369234 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 369854 708678
rect 369234 708358 369854 708442
rect 369234 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 369854 708358
rect 365514 706758 366134 707750
rect 365514 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 366134 706758
rect 365514 706438 366134 706522
rect 365514 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 366134 706438
rect 354954 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 355574 680614
rect 354954 680294 355574 680378
rect 354954 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 355574 680294
rect 354954 644614 355574 680058
rect 354954 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 355574 644614
rect 354954 644294 355574 644378
rect 354954 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 355574 644294
rect 354954 608614 355574 644058
rect 354954 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 355574 608614
rect 354954 608294 355574 608378
rect 354954 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 355574 608294
rect 354954 572614 355574 608058
rect 354954 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 355574 572614
rect 354954 572294 355574 572378
rect 354954 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 355574 572294
rect 354954 536614 355574 572058
rect 354954 536378 354986 536614
rect 355222 536378 355306 536614
rect 355542 536378 355574 536614
rect 354954 536294 355574 536378
rect 354954 536058 354986 536294
rect 355222 536058 355306 536294
rect 355542 536058 355574 536294
rect 354954 500614 355574 536058
rect 354954 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 355574 500614
rect 354954 500294 355574 500378
rect 354954 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 355574 500294
rect 354954 464614 355574 500058
rect 354954 464378 354986 464614
rect 355222 464378 355306 464614
rect 355542 464378 355574 464614
rect 354954 464294 355574 464378
rect 354954 464058 354986 464294
rect 355222 464058 355306 464294
rect 355542 464058 355574 464294
rect 354954 428614 355574 464058
rect 354954 428378 354986 428614
rect 355222 428378 355306 428614
rect 355542 428378 355574 428614
rect 354954 428294 355574 428378
rect 354954 428058 354986 428294
rect 355222 428058 355306 428294
rect 355542 428058 355574 428294
rect 354954 392614 355574 428058
rect 354954 392378 354986 392614
rect 355222 392378 355306 392614
rect 355542 392378 355574 392614
rect 354954 392294 355574 392378
rect 354954 392058 354986 392294
rect 355222 392058 355306 392294
rect 355542 392058 355574 392294
rect 354954 356614 355574 392058
rect 361794 704838 362414 705830
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 435454 362414 470898
rect 361794 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 362414 435454
rect 361794 435134 362414 435218
rect 361794 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 362414 435134
rect 361794 399454 362414 434898
rect 361794 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 362414 399454
rect 361794 399134 362414 399218
rect 361794 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 362414 399134
rect 361794 372000 362414 398898
rect 365514 691174 366134 706202
rect 365514 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 366134 691174
rect 365514 690854 366134 690938
rect 365514 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 366134 690854
rect 365514 655174 366134 690618
rect 365514 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 366134 655174
rect 365514 654854 366134 654938
rect 365514 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 366134 654854
rect 365514 619174 366134 654618
rect 365514 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 366134 619174
rect 365514 618854 366134 618938
rect 365514 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 366134 618854
rect 365514 583174 366134 618618
rect 365514 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 366134 583174
rect 365514 582854 366134 582938
rect 365514 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 366134 582854
rect 365514 547174 366134 582618
rect 365514 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 366134 547174
rect 365514 546854 366134 546938
rect 365514 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 366134 546854
rect 365514 511174 366134 546618
rect 365514 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 366134 511174
rect 365514 510854 366134 510938
rect 365514 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 366134 510854
rect 365514 475174 366134 510618
rect 365514 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 366134 475174
rect 365514 474854 366134 474938
rect 365514 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 366134 474854
rect 365514 439174 366134 474618
rect 365514 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 366134 439174
rect 365514 438854 366134 438938
rect 365514 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 366134 438854
rect 365514 403174 366134 438618
rect 365514 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 366134 403174
rect 365514 402854 366134 402938
rect 365514 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 366134 402854
rect 365514 372000 366134 402618
rect 369234 694894 369854 708122
rect 369234 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 369854 694894
rect 369234 694574 369854 694658
rect 369234 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 369854 694574
rect 369234 658894 369854 694338
rect 369234 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 369854 658894
rect 369234 658574 369854 658658
rect 369234 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 369854 658574
rect 369234 622894 369854 658338
rect 369234 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 369854 622894
rect 369234 622574 369854 622658
rect 369234 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 369854 622574
rect 369234 586894 369854 622338
rect 369234 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 369854 586894
rect 369234 586574 369854 586658
rect 369234 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 369854 586574
rect 369234 550894 369854 586338
rect 369234 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 369854 550894
rect 369234 550574 369854 550658
rect 369234 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 369854 550574
rect 369234 514894 369854 550338
rect 369234 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 369854 514894
rect 369234 514574 369854 514658
rect 369234 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 369854 514574
rect 369234 478894 369854 514338
rect 369234 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 369854 478894
rect 369234 478574 369854 478658
rect 369234 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 369854 478574
rect 369234 442894 369854 478338
rect 369234 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 369854 442894
rect 369234 442574 369854 442658
rect 369234 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 369854 442574
rect 369234 406894 369854 442338
rect 369234 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 369854 406894
rect 369234 406574 369854 406658
rect 369234 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 369854 406574
rect 369234 372000 369854 406338
rect 372954 698614 373574 710042
rect 390954 711558 391574 711590
rect 390954 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 391574 711558
rect 390954 711238 391574 711322
rect 390954 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 391574 711238
rect 387234 709638 387854 709670
rect 387234 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 387854 709638
rect 387234 709318 387854 709402
rect 387234 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 387854 709318
rect 383514 707718 384134 707750
rect 383514 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 384134 707718
rect 383514 707398 384134 707482
rect 383514 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 384134 707398
rect 372954 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 373574 698614
rect 372954 698294 373574 698378
rect 372954 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 373574 698294
rect 372954 662614 373574 698058
rect 372954 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 373574 662614
rect 372954 662294 373574 662378
rect 372954 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 373574 662294
rect 372954 626614 373574 662058
rect 372954 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 373574 626614
rect 372954 626294 373574 626378
rect 372954 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 373574 626294
rect 372954 590614 373574 626058
rect 372954 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 373574 590614
rect 372954 590294 373574 590378
rect 372954 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 373574 590294
rect 372954 554614 373574 590058
rect 372954 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 373574 554614
rect 372954 554294 373574 554378
rect 372954 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 373574 554294
rect 372954 518614 373574 554058
rect 372954 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 373574 518614
rect 372954 518294 373574 518378
rect 372954 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 373574 518294
rect 372954 482614 373574 518058
rect 372954 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 373574 482614
rect 372954 482294 373574 482378
rect 372954 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 373574 482294
rect 372954 446614 373574 482058
rect 372954 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 373574 446614
rect 372954 446294 373574 446378
rect 372954 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 373574 446294
rect 372954 410614 373574 446058
rect 372954 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 373574 410614
rect 372954 410294 373574 410378
rect 372954 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 373574 410294
rect 372954 374614 373574 410058
rect 372954 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 373574 374614
rect 372954 374294 373574 374378
rect 372954 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 373574 374294
rect 362243 363454 362563 363486
rect 362243 363218 362285 363454
rect 362521 363218 362563 363454
rect 362243 363134 362563 363218
rect 362243 362898 362285 363134
rect 362521 362898 362563 363134
rect 362243 362866 362563 362898
rect 364840 363454 365160 363486
rect 364840 363218 364882 363454
rect 365118 363218 365160 363454
rect 364840 363134 365160 363218
rect 364840 362898 364882 363134
rect 365118 362898 365160 363134
rect 364840 362866 365160 362898
rect 367437 363454 367757 363486
rect 367437 363218 367479 363454
rect 367715 363218 367757 363454
rect 367437 363134 367757 363218
rect 367437 362898 367479 363134
rect 367715 362898 367757 363134
rect 367437 362866 367757 362898
rect 354954 356378 354986 356614
rect 355222 356378 355306 356614
rect 355542 356378 355574 356614
rect 354954 356294 355574 356378
rect 354954 356058 354986 356294
rect 355222 356058 355306 356294
rect 355542 356058 355574 356294
rect 354954 320614 355574 356058
rect 371923 353564 371989 353565
rect 371923 353500 371924 353564
rect 371988 353500 371989 353564
rect 371923 353499 371989 353500
rect 371739 353020 371805 353021
rect 371739 352956 371740 353020
rect 371804 352956 371805 353020
rect 371739 352955 371805 352956
rect 371555 351388 371621 351389
rect 371555 351324 371556 351388
rect 371620 351324 371621 351388
rect 371555 351323 371621 351324
rect 371187 350844 371253 350845
rect 371187 350780 371188 350844
rect 371252 350780 371253 350844
rect 371187 350779 371253 350780
rect 363541 345454 363861 345486
rect 363541 345218 363583 345454
rect 363819 345218 363861 345454
rect 363541 345134 363861 345218
rect 363541 344898 363583 345134
rect 363819 344898 363861 345134
rect 363541 344866 363861 344898
rect 366138 345454 366458 345486
rect 366138 345218 366180 345454
rect 366416 345218 366458 345454
rect 366138 345134 366458 345218
rect 366138 344898 366180 345134
rect 366416 344898 366458 345134
rect 366138 344866 366458 344898
rect 361619 337788 361685 337789
rect 361619 337724 361620 337788
rect 361684 337724 361685 337788
rect 361619 337723 361685 337724
rect 354954 320378 354986 320614
rect 355222 320378 355306 320614
rect 355542 320378 355574 320614
rect 354954 320294 355574 320378
rect 354954 320058 354986 320294
rect 355222 320058 355306 320294
rect 355542 320058 355574 320294
rect 354954 284614 355574 320058
rect 354954 284378 354986 284614
rect 355222 284378 355306 284614
rect 355542 284378 355574 284614
rect 354954 284294 355574 284378
rect 354954 284058 354986 284294
rect 355222 284058 355306 284294
rect 355542 284058 355574 284294
rect 354954 248614 355574 284058
rect 361622 267885 361682 337723
rect 361794 327454 362414 338000
rect 364379 337788 364445 337789
rect 364379 337724 364380 337788
rect 364444 337724 364445 337788
rect 364379 337723 364445 337724
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 361794 300000 362414 326898
rect 362243 291454 362563 291486
rect 362243 291218 362285 291454
rect 362521 291218 362563 291454
rect 362243 291134 362563 291218
rect 362243 290898 362285 291134
rect 362521 290898 362563 291134
rect 362243 290866 362563 290898
rect 363541 273454 363861 273486
rect 363541 273218 363583 273454
rect 363819 273218 363861 273454
rect 363541 273134 363861 273218
rect 363541 272898 363583 273134
rect 363819 272898 363861 273134
rect 363541 272866 363861 272898
rect 361619 267884 361685 267885
rect 361619 267820 361620 267884
rect 361684 267820 361685 267884
rect 361619 267819 361685 267820
rect 361622 266117 361682 267819
rect 364382 266253 364442 337723
rect 365514 331174 366134 338000
rect 365514 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 366134 331174
rect 365514 330854 366134 330938
rect 365514 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 366134 330854
rect 365514 300000 366134 330618
rect 369234 334894 369854 338000
rect 369234 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 369854 334894
rect 369234 334574 369854 334658
rect 369234 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 369854 334574
rect 369234 300000 369854 334338
rect 364840 291454 365160 291486
rect 364840 291218 364882 291454
rect 365118 291218 365160 291454
rect 364840 291134 365160 291218
rect 364840 290898 364882 291134
rect 365118 290898 365160 291134
rect 364840 290866 365160 290898
rect 367437 291454 367757 291486
rect 367437 291218 367479 291454
rect 367715 291218 367757 291454
rect 367437 291134 367757 291218
rect 367437 290898 367479 291134
rect 367715 290898 367757 291134
rect 367437 290866 367757 290898
rect 371190 278901 371250 350779
rect 371371 281620 371437 281621
rect 371371 281556 371372 281620
rect 371436 281556 371437 281620
rect 371371 281555 371437 281556
rect 371187 278900 371253 278901
rect 371187 278836 371188 278900
rect 371252 278836 371253 278900
rect 371187 278835 371253 278836
rect 370083 276996 370149 276997
rect 370083 276932 370084 276996
rect 370148 276932 370149 276996
rect 370083 276931 370149 276932
rect 366138 273454 366458 273486
rect 366138 273218 366180 273454
rect 366416 273218 366458 273454
rect 366138 273134 366458 273218
rect 366138 272898 366180 273134
rect 366416 272898 366458 273134
rect 366138 272866 366458 272898
rect 364379 266252 364445 266253
rect 364379 266188 364380 266252
rect 364444 266188 364445 266252
rect 364379 266187 364445 266188
rect 361619 266116 361685 266117
rect 361619 266052 361620 266116
rect 361684 266052 361685 266116
rect 361619 266051 361685 266052
rect 354954 248378 354986 248614
rect 355222 248378 355306 248614
rect 355542 248378 355574 248614
rect 354954 248294 355574 248378
rect 354954 248058 354986 248294
rect 355222 248058 355306 248294
rect 355542 248058 355574 248294
rect 354954 212614 355574 248058
rect 354954 212378 354986 212614
rect 355222 212378 355306 212614
rect 355542 212378 355574 212614
rect 354954 212294 355574 212378
rect 354954 212058 354986 212294
rect 355222 212058 355306 212294
rect 355542 212058 355574 212294
rect 354954 176614 355574 212058
rect 361622 194581 361682 266051
rect 361794 255454 362414 266000
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 228000 362414 254898
rect 362243 219454 362563 219486
rect 362243 219218 362285 219454
rect 362521 219218 362563 219454
rect 362243 219134 362563 219218
rect 362243 218898 362285 219134
rect 362521 218898 362563 219134
rect 362243 218866 362563 218898
rect 363541 201454 363861 201486
rect 363541 201218 363583 201454
rect 363819 201218 363861 201454
rect 363541 201134 363861 201218
rect 363541 200898 363583 201134
rect 363819 200898 363861 201134
rect 363541 200866 363861 200898
rect 364382 196077 364442 266187
rect 365514 259174 366134 266000
rect 365514 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 366134 259174
rect 365514 258854 366134 258938
rect 365514 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 366134 258854
rect 365514 228000 366134 258618
rect 369234 262894 369854 266000
rect 369234 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 369854 262894
rect 369234 262574 369854 262658
rect 369234 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 369854 262574
rect 369234 228000 369854 262338
rect 364840 219454 365160 219486
rect 364840 219218 364882 219454
rect 365118 219218 365160 219454
rect 364840 219134 365160 219218
rect 364840 218898 364882 219134
rect 365118 218898 365160 219134
rect 364840 218866 365160 218898
rect 367437 219454 367757 219486
rect 367437 219218 367479 219454
rect 367715 219218 367757 219454
rect 367437 219134 367757 219218
rect 367437 218898 367479 219134
rect 367715 218898 367757 219134
rect 367437 218866 367757 218898
rect 370086 205325 370146 276931
rect 370267 275364 370333 275365
rect 370267 275300 370268 275364
rect 370332 275300 370333 275364
rect 370267 275299 370333 275300
rect 370083 205324 370149 205325
rect 370083 205260 370084 205324
rect 370148 205260 370149 205324
rect 370083 205259 370149 205260
rect 370270 203693 370330 275299
rect 371190 206821 371250 278835
rect 371374 225045 371434 281555
rect 371558 279445 371618 351323
rect 371742 281077 371802 352955
rect 371926 281621 371986 353499
rect 372107 352476 372173 352477
rect 372107 352412 372108 352476
rect 372172 352412 372173 352476
rect 372107 352411 372173 352412
rect 371923 281620 371989 281621
rect 371923 281556 371924 281620
rect 371988 281556 371989 281620
rect 371923 281555 371989 281556
rect 371739 281076 371805 281077
rect 371739 281012 371740 281076
rect 371804 281012 371805 281076
rect 371739 281011 371805 281012
rect 371555 279444 371621 279445
rect 371555 279380 371556 279444
rect 371620 279380 371621 279444
rect 371555 279379 371621 279380
rect 371371 225044 371437 225045
rect 371371 224980 371372 225044
rect 371436 224980 371437 225044
rect 371371 224979 371437 224980
rect 371374 209541 371434 224979
rect 371371 209540 371437 209541
rect 371371 209476 371372 209540
rect 371436 209476 371437 209540
rect 371371 209475 371437 209476
rect 371558 207365 371618 279379
rect 371742 223957 371802 281011
rect 372110 280533 372170 352411
rect 372954 338614 373574 374058
rect 372954 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 373574 338614
rect 372954 338294 373574 338378
rect 372954 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 373574 338294
rect 372954 302614 373574 338058
rect 372954 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 373574 302614
rect 372954 302294 373574 302378
rect 372954 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 373574 302294
rect 372107 280532 372173 280533
rect 372107 280468 372108 280532
rect 372172 280468 372173 280532
rect 372107 280467 372173 280468
rect 372110 277410 372170 280467
rect 371926 277350 372170 277410
rect 371739 223956 371805 223957
rect 371739 223892 371740 223956
rect 371804 223892 371805 223956
rect 371739 223891 371805 223892
rect 371742 208997 371802 223891
rect 371739 208996 371805 208997
rect 371739 208932 371740 208996
rect 371804 208932 371805 208996
rect 371739 208931 371805 208932
rect 371926 208453 371986 277350
rect 372954 266614 373574 302058
rect 372954 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 373574 266614
rect 372954 266294 373574 266378
rect 372954 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 373574 266294
rect 372954 230614 373574 266058
rect 372954 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 373574 230614
rect 372954 230294 373574 230378
rect 372954 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 373574 230294
rect 371923 208452 371989 208453
rect 371923 208388 371924 208452
rect 371988 208388 371989 208452
rect 371923 208387 371989 208388
rect 371555 207364 371621 207365
rect 371555 207300 371556 207364
rect 371620 207300 371621 207364
rect 371555 207299 371621 207300
rect 371923 207364 371989 207365
rect 371923 207300 371924 207364
rect 371988 207300 371989 207364
rect 371923 207299 371989 207300
rect 371187 206820 371253 206821
rect 371187 206756 371188 206820
rect 371252 206756 371253 206820
rect 371187 206755 371253 206756
rect 370267 203692 370333 203693
rect 370267 203628 370268 203692
rect 370332 203628 370333 203692
rect 370267 203627 370333 203628
rect 366138 201454 366458 201486
rect 366138 201218 366180 201454
rect 366416 201218 366458 201454
rect 366138 201134 366458 201218
rect 366138 200898 366180 201134
rect 366416 200898 366458 201134
rect 366138 200866 366458 200898
rect 364379 196076 364445 196077
rect 364379 196012 364380 196076
rect 364444 196012 364445 196076
rect 364379 196011 364445 196012
rect 371371 196076 371437 196077
rect 371371 196012 371372 196076
rect 371436 196012 371437 196076
rect 371371 196011 371437 196012
rect 361619 194580 361685 194581
rect 361619 194516 361620 194580
rect 361684 194516 361685 194580
rect 361619 194515 361685 194516
rect 362723 194580 362789 194581
rect 362723 194516 362724 194580
rect 362788 194516 362789 194580
rect 362723 194515 362789 194516
rect 365299 194580 365365 194581
rect 365299 194516 365300 194580
rect 365364 194516 365365 194580
rect 365299 194515 365365 194516
rect 354954 176378 354986 176614
rect 355222 176378 355306 176614
rect 355542 176378 355574 176614
rect 354954 176294 355574 176378
rect 354954 176058 354986 176294
rect 355222 176058 355306 176294
rect 355542 176058 355574 176294
rect 354954 140614 355574 176058
rect 361794 183454 362414 194000
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 361794 156000 362414 182898
rect 362243 147454 362563 147486
rect 362243 147218 362285 147454
rect 362521 147218 362563 147454
rect 362243 147134 362563 147218
rect 362243 146898 362285 147134
rect 362521 146898 362563 147134
rect 362243 146866 362563 146898
rect 354954 140378 354986 140614
rect 355222 140378 355306 140614
rect 355542 140378 355574 140614
rect 354954 140294 355574 140378
rect 354954 140058 354986 140294
rect 355222 140058 355306 140294
rect 355542 140058 355574 140294
rect 354954 104614 355574 140058
rect 362726 123997 362786 194515
rect 364840 147454 365160 147486
rect 364840 147218 364882 147454
rect 365118 147218 365160 147454
rect 364840 147134 365160 147218
rect 364840 146898 364882 147134
rect 365118 146898 365160 147134
rect 364840 146866 365160 146898
rect 363541 129454 363861 129486
rect 363541 129218 363583 129454
rect 363819 129218 363861 129454
rect 363541 129134 363861 129218
rect 363541 128898 363583 129134
rect 363819 128898 363861 129134
rect 363541 128866 363861 128898
rect 365302 123997 365362 194515
rect 365514 187174 366134 194000
rect 365514 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 366134 187174
rect 365514 186854 366134 186938
rect 365514 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 366134 186854
rect 365514 156000 366134 186618
rect 369234 190894 369854 194000
rect 369234 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 369854 190894
rect 369234 190574 369854 190658
rect 369234 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 369854 190574
rect 369234 156000 369854 190338
rect 367437 147454 367757 147486
rect 367437 147218 367479 147454
rect 367715 147218 367757 147454
rect 367437 147134 367757 147218
rect 367437 146898 367479 147134
rect 367715 146898 367757 147134
rect 367437 146866 367757 146898
rect 371374 137597 371434 196011
rect 371739 175676 371805 175677
rect 371739 175612 371740 175676
rect 371804 175612 371805 175676
rect 371739 175611 371805 175612
rect 371371 137596 371437 137597
rect 371371 137532 371372 137596
rect 371436 137532 371437 137596
rect 371371 137531 371437 137532
rect 371742 136509 371802 175611
rect 371926 175130 371986 207299
rect 372291 206820 372357 206821
rect 372291 206756 372292 206820
rect 372356 206756 372357 206820
rect 372291 206755 372357 206756
rect 372294 175269 372354 206755
rect 372475 195260 372541 195261
rect 372475 195196 372476 195260
rect 372540 195196 372541 195260
rect 372475 195195 372541 195196
rect 372291 175268 372357 175269
rect 372291 175204 372292 175268
rect 372356 175204 372357 175268
rect 372291 175203 372357 175204
rect 371926 175070 372354 175130
rect 371923 174996 371989 174997
rect 371923 174932 371924 174996
rect 371988 174932 371989 174996
rect 371923 174931 371989 174932
rect 371926 171733 371986 174931
rect 372294 173229 372354 175070
rect 372291 173228 372357 173229
rect 372291 173164 372292 173228
rect 372356 173164 372357 173228
rect 372291 173163 372357 173164
rect 371923 171732 371989 171733
rect 371923 171668 371924 171732
rect 371988 171668 371989 171732
rect 371923 171667 371989 171668
rect 371926 152965 371986 171667
rect 372294 162757 372354 173163
rect 372291 162756 372357 162757
rect 372291 162692 372292 162756
rect 372356 162692 372357 162756
rect 372291 162691 372357 162692
rect 371923 152964 371989 152965
rect 371923 152900 371924 152964
rect 371988 152900 371989 152964
rect 371923 152899 371989 152900
rect 372478 137053 372538 195195
rect 372954 194614 373574 230058
rect 372954 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 373574 194614
rect 372954 194294 373574 194378
rect 372954 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 373574 194294
rect 372954 158614 373574 194058
rect 372954 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 373574 158614
rect 372954 158294 373574 158378
rect 372954 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 373574 158294
rect 372475 137052 372541 137053
rect 372475 136988 372476 137052
rect 372540 136988 372541 137052
rect 372475 136987 372541 136988
rect 371739 136508 371805 136509
rect 371739 136444 371740 136508
rect 371804 136444 371805 136508
rect 371739 136443 371805 136444
rect 366138 129454 366458 129486
rect 366138 129218 366180 129454
rect 366416 129218 366458 129454
rect 366138 129134 366458 129218
rect 366138 128898 366180 129134
rect 366416 128898 366458 129134
rect 366138 128866 366458 128898
rect 362723 123996 362789 123997
rect 362723 123932 362724 123996
rect 362788 123932 362789 123996
rect 362723 123931 362789 123932
rect 365299 123996 365365 123997
rect 365299 123932 365300 123996
rect 365364 123932 365365 123996
rect 365299 123931 365365 123932
rect 372954 122614 373574 158058
rect 372954 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 373574 122614
rect 372954 122294 373574 122378
rect 372954 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 373574 122294
rect 354954 104378 354986 104614
rect 355222 104378 355306 104614
rect 355542 104378 355574 104614
rect 354954 104294 355574 104378
rect 354954 104058 354986 104294
rect 355222 104058 355306 104294
rect 355542 104058 355574 104294
rect 354954 68614 355574 104058
rect 354954 68378 354986 68614
rect 355222 68378 355306 68614
rect 355542 68378 355574 68614
rect 354954 68294 355574 68378
rect 354954 68058 354986 68294
rect 355222 68058 355306 68294
rect 355542 68058 355574 68294
rect 354954 32614 355574 68058
rect 354954 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 355574 32614
rect 354954 32294 355574 32378
rect 354954 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 355574 32294
rect 336954 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 337574 -6106
rect 336954 -6426 337574 -6342
rect 336954 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 337574 -6426
rect 336954 -7654 337574 -6662
rect 354954 -7066 355574 32058
rect 361794 111454 362414 122000
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -1894 362414 -902
rect 365514 115174 366134 122000
rect 365514 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 366134 115174
rect 365514 114854 366134 114938
rect 365514 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 366134 114854
rect 365514 79174 366134 114618
rect 365514 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 366134 79174
rect 365514 78854 366134 78938
rect 365514 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 366134 78854
rect 365514 43174 366134 78618
rect 365514 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 366134 43174
rect 365514 42854 366134 42938
rect 365514 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 366134 42854
rect 365514 7174 366134 42618
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 365514 -2266 366134 6618
rect 365514 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 366134 -2266
rect 365514 -2586 366134 -2502
rect 365514 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 366134 -2586
rect 365514 -3814 366134 -2822
rect 369234 118894 369854 122000
rect 369234 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 369854 118894
rect 369234 118574 369854 118658
rect 369234 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 369854 118574
rect 369234 82894 369854 118338
rect 369234 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 369854 82894
rect 369234 82574 369854 82658
rect 369234 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 369854 82574
rect 369234 46894 369854 82338
rect 369234 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 369854 46894
rect 369234 46574 369854 46658
rect 369234 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 369854 46574
rect 369234 10894 369854 46338
rect 369234 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 369854 10894
rect 369234 10574 369854 10658
rect 369234 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 369854 10574
rect 369234 -4186 369854 10338
rect 369234 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 369854 -4186
rect 369234 -4506 369854 -4422
rect 369234 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 369854 -4506
rect 369234 -5734 369854 -4742
rect 372954 86614 373574 122058
rect 372954 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 373574 86614
rect 372954 86294 373574 86378
rect 372954 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 373574 86294
rect 372954 50614 373574 86058
rect 372954 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 373574 50614
rect 372954 50294 373574 50378
rect 372954 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 373574 50294
rect 372954 14614 373574 50058
rect 372954 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 373574 14614
rect 372954 14294 373574 14378
rect 372954 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 373574 14294
rect 354954 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 355574 -7066
rect 354954 -7386 355574 -7302
rect 354954 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 355574 -7386
rect 354954 -7654 355574 -7622
rect 372954 -6106 373574 14058
rect 379794 705798 380414 705830
rect 379794 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 380414 705798
rect 379794 705478 380414 705562
rect 379794 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 380414 705478
rect 379794 669454 380414 705242
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 561454 380414 596898
rect 379794 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 380414 561454
rect 379794 561134 380414 561218
rect 379794 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 380414 561134
rect 379794 525454 380414 560898
rect 379794 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 380414 525454
rect 379794 525134 380414 525218
rect 379794 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 380414 525134
rect 379794 489454 380414 524898
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 379794 489134 380414 489218
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 379794 453454 380414 488898
rect 379794 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 380414 453454
rect 379794 453134 380414 453218
rect 379794 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 380414 453134
rect 379794 417454 380414 452898
rect 379794 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 380414 417454
rect 379794 417134 380414 417218
rect 379794 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 380414 417134
rect 379794 381454 380414 416898
rect 379794 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 380414 381454
rect 379794 381134 380414 381218
rect 379794 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 380414 381134
rect 379794 345454 380414 380898
rect 379794 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 380414 345454
rect 379794 345134 380414 345218
rect 379794 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 380414 345134
rect 379794 309454 380414 344898
rect 379794 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 380414 309454
rect 379794 309134 380414 309218
rect 379794 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 380414 309134
rect 379794 273454 380414 308898
rect 379794 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 380414 273454
rect 379794 273134 380414 273218
rect 379794 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 380414 273134
rect 379794 237454 380414 272898
rect 379794 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 380414 237454
rect 379794 237134 380414 237218
rect 379794 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 380414 237134
rect 379794 201454 380414 236898
rect 379794 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 380414 201454
rect 379794 201134 380414 201218
rect 379794 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 380414 201134
rect 379794 165454 380414 200898
rect 379794 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 380414 165454
rect 379794 165134 380414 165218
rect 379794 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 380414 165134
rect 379794 129454 380414 164898
rect 379794 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 380414 129454
rect 379794 129134 380414 129218
rect 379794 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 380414 129134
rect 379794 93454 380414 128898
rect 379794 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 380414 93454
rect 379794 93134 380414 93218
rect 379794 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 380414 93134
rect 379794 57454 380414 92898
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -1306 380414 20898
rect 379794 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 380414 -1306
rect 379794 -1626 380414 -1542
rect 379794 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 380414 -1626
rect 379794 -1894 380414 -1862
rect 383514 673174 384134 707162
rect 383514 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 384134 673174
rect 383514 672854 384134 672938
rect 383514 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 384134 672854
rect 383514 637174 384134 672618
rect 383514 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 384134 637174
rect 383514 636854 384134 636938
rect 383514 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 384134 636854
rect 383514 601174 384134 636618
rect 383514 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 384134 601174
rect 383514 600854 384134 600938
rect 383514 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 384134 600854
rect 383514 565174 384134 600618
rect 383514 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 384134 565174
rect 383514 564854 384134 564938
rect 383514 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 384134 564854
rect 383514 529174 384134 564618
rect 383514 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 384134 529174
rect 383514 528854 384134 528938
rect 383514 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 384134 528854
rect 383514 493174 384134 528618
rect 383514 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 384134 493174
rect 383514 492854 384134 492938
rect 383514 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 384134 492854
rect 383514 457174 384134 492618
rect 383514 456938 383546 457174
rect 383782 456938 383866 457174
rect 384102 456938 384134 457174
rect 383514 456854 384134 456938
rect 383514 456618 383546 456854
rect 383782 456618 383866 456854
rect 384102 456618 384134 456854
rect 383514 421174 384134 456618
rect 383514 420938 383546 421174
rect 383782 420938 383866 421174
rect 384102 420938 384134 421174
rect 383514 420854 384134 420938
rect 383514 420618 383546 420854
rect 383782 420618 383866 420854
rect 384102 420618 384134 420854
rect 383514 385174 384134 420618
rect 383514 384938 383546 385174
rect 383782 384938 383866 385174
rect 384102 384938 384134 385174
rect 383514 384854 384134 384938
rect 383514 384618 383546 384854
rect 383782 384618 383866 384854
rect 384102 384618 384134 384854
rect 383514 349174 384134 384618
rect 383514 348938 383546 349174
rect 383782 348938 383866 349174
rect 384102 348938 384134 349174
rect 383514 348854 384134 348938
rect 383514 348618 383546 348854
rect 383782 348618 383866 348854
rect 384102 348618 384134 348854
rect 383514 313174 384134 348618
rect 383514 312938 383546 313174
rect 383782 312938 383866 313174
rect 384102 312938 384134 313174
rect 383514 312854 384134 312938
rect 383514 312618 383546 312854
rect 383782 312618 383866 312854
rect 384102 312618 384134 312854
rect 383514 277174 384134 312618
rect 383514 276938 383546 277174
rect 383782 276938 383866 277174
rect 384102 276938 384134 277174
rect 383514 276854 384134 276938
rect 383514 276618 383546 276854
rect 383782 276618 383866 276854
rect 384102 276618 384134 276854
rect 383514 241174 384134 276618
rect 383514 240938 383546 241174
rect 383782 240938 383866 241174
rect 384102 240938 384134 241174
rect 383514 240854 384134 240938
rect 383514 240618 383546 240854
rect 383782 240618 383866 240854
rect 384102 240618 384134 240854
rect 383514 205174 384134 240618
rect 383514 204938 383546 205174
rect 383782 204938 383866 205174
rect 384102 204938 384134 205174
rect 383514 204854 384134 204938
rect 383514 204618 383546 204854
rect 383782 204618 383866 204854
rect 384102 204618 384134 204854
rect 383514 169174 384134 204618
rect 383514 168938 383546 169174
rect 383782 168938 383866 169174
rect 384102 168938 384134 169174
rect 383514 168854 384134 168938
rect 383514 168618 383546 168854
rect 383782 168618 383866 168854
rect 384102 168618 384134 168854
rect 383514 133174 384134 168618
rect 383514 132938 383546 133174
rect 383782 132938 383866 133174
rect 384102 132938 384134 133174
rect 383514 132854 384134 132938
rect 383514 132618 383546 132854
rect 383782 132618 383866 132854
rect 384102 132618 384134 132854
rect 383514 97174 384134 132618
rect 383514 96938 383546 97174
rect 383782 96938 383866 97174
rect 384102 96938 384134 97174
rect 383514 96854 384134 96938
rect 383514 96618 383546 96854
rect 383782 96618 383866 96854
rect 384102 96618 384134 96854
rect 383514 61174 384134 96618
rect 383514 60938 383546 61174
rect 383782 60938 383866 61174
rect 384102 60938 384134 61174
rect 383514 60854 384134 60938
rect 383514 60618 383546 60854
rect 383782 60618 383866 60854
rect 384102 60618 384134 60854
rect 383514 25174 384134 60618
rect 383514 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 384134 25174
rect 383514 24854 384134 24938
rect 383514 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 384134 24854
rect 383514 -3226 384134 24618
rect 383514 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 384134 -3226
rect 383514 -3546 384134 -3462
rect 383514 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 384134 -3546
rect 383514 -3814 384134 -3782
rect 387234 676894 387854 709082
rect 387234 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 387854 676894
rect 387234 676574 387854 676658
rect 387234 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 387854 676574
rect 387234 640894 387854 676338
rect 387234 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 387854 640894
rect 387234 640574 387854 640658
rect 387234 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 387854 640574
rect 387234 604894 387854 640338
rect 387234 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 387854 604894
rect 387234 604574 387854 604658
rect 387234 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 387854 604574
rect 387234 568894 387854 604338
rect 387234 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 387854 568894
rect 387234 568574 387854 568658
rect 387234 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 387854 568574
rect 387234 532894 387854 568338
rect 387234 532658 387266 532894
rect 387502 532658 387586 532894
rect 387822 532658 387854 532894
rect 387234 532574 387854 532658
rect 387234 532338 387266 532574
rect 387502 532338 387586 532574
rect 387822 532338 387854 532574
rect 387234 496894 387854 532338
rect 387234 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 387854 496894
rect 387234 496574 387854 496658
rect 387234 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 387854 496574
rect 387234 460894 387854 496338
rect 387234 460658 387266 460894
rect 387502 460658 387586 460894
rect 387822 460658 387854 460894
rect 387234 460574 387854 460658
rect 387234 460338 387266 460574
rect 387502 460338 387586 460574
rect 387822 460338 387854 460574
rect 387234 424894 387854 460338
rect 387234 424658 387266 424894
rect 387502 424658 387586 424894
rect 387822 424658 387854 424894
rect 387234 424574 387854 424658
rect 387234 424338 387266 424574
rect 387502 424338 387586 424574
rect 387822 424338 387854 424574
rect 387234 388894 387854 424338
rect 387234 388658 387266 388894
rect 387502 388658 387586 388894
rect 387822 388658 387854 388894
rect 387234 388574 387854 388658
rect 387234 388338 387266 388574
rect 387502 388338 387586 388574
rect 387822 388338 387854 388574
rect 387234 352894 387854 388338
rect 387234 352658 387266 352894
rect 387502 352658 387586 352894
rect 387822 352658 387854 352894
rect 387234 352574 387854 352658
rect 387234 352338 387266 352574
rect 387502 352338 387586 352574
rect 387822 352338 387854 352574
rect 387234 316894 387854 352338
rect 387234 316658 387266 316894
rect 387502 316658 387586 316894
rect 387822 316658 387854 316894
rect 387234 316574 387854 316658
rect 387234 316338 387266 316574
rect 387502 316338 387586 316574
rect 387822 316338 387854 316574
rect 387234 280894 387854 316338
rect 387234 280658 387266 280894
rect 387502 280658 387586 280894
rect 387822 280658 387854 280894
rect 387234 280574 387854 280658
rect 387234 280338 387266 280574
rect 387502 280338 387586 280574
rect 387822 280338 387854 280574
rect 387234 244894 387854 280338
rect 387234 244658 387266 244894
rect 387502 244658 387586 244894
rect 387822 244658 387854 244894
rect 387234 244574 387854 244658
rect 387234 244338 387266 244574
rect 387502 244338 387586 244574
rect 387822 244338 387854 244574
rect 387234 208894 387854 244338
rect 387234 208658 387266 208894
rect 387502 208658 387586 208894
rect 387822 208658 387854 208894
rect 387234 208574 387854 208658
rect 387234 208338 387266 208574
rect 387502 208338 387586 208574
rect 387822 208338 387854 208574
rect 387234 172894 387854 208338
rect 387234 172658 387266 172894
rect 387502 172658 387586 172894
rect 387822 172658 387854 172894
rect 387234 172574 387854 172658
rect 387234 172338 387266 172574
rect 387502 172338 387586 172574
rect 387822 172338 387854 172574
rect 387234 136894 387854 172338
rect 387234 136658 387266 136894
rect 387502 136658 387586 136894
rect 387822 136658 387854 136894
rect 387234 136574 387854 136658
rect 387234 136338 387266 136574
rect 387502 136338 387586 136574
rect 387822 136338 387854 136574
rect 387234 100894 387854 136338
rect 387234 100658 387266 100894
rect 387502 100658 387586 100894
rect 387822 100658 387854 100894
rect 387234 100574 387854 100658
rect 387234 100338 387266 100574
rect 387502 100338 387586 100574
rect 387822 100338 387854 100574
rect 387234 64894 387854 100338
rect 387234 64658 387266 64894
rect 387502 64658 387586 64894
rect 387822 64658 387854 64894
rect 387234 64574 387854 64658
rect 387234 64338 387266 64574
rect 387502 64338 387586 64574
rect 387822 64338 387854 64574
rect 387234 28894 387854 64338
rect 387234 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 387854 28894
rect 387234 28574 387854 28658
rect 387234 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 387854 28574
rect 387234 -5146 387854 28338
rect 387234 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 387854 -5146
rect 387234 -5466 387854 -5382
rect 387234 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 387854 -5466
rect 387234 -5734 387854 -5702
rect 390954 680614 391574 711002
rect 408954 710598 409574 711590
rect 408954 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 409574 710598
rect 408954 710278 409574 710362
rect 408954 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 409574 710278
rect 405234 708678 405854 709670
rect 405234 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 405854 708678
rect 405234 708358 405854 708442
rect 405234 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 405854 708358
rect 401514 706758 402134 707750
rect 401514 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 402134 706758
rect 401514 706438 402134 706522
rect 401514 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 402134 706438
rect 390954 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 391574 680614
rect 390954 680294 391574 680378
rect 390954 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 391574 680294
rect 390954 644614 391574 680058
rect 390954 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 391574 644614
rect 390954 644294 391574 644378
rect 390954 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 391574 644294
rect 390954 608614 391574 644058
rect 390954 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 391574 608614
rect 390954 608294 391574 608378
rect 390954 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 391574 608294
rect 390954 572614 391574 608058
rect 390954 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 391574 572614
rect 390954 572294 391574 572378
rect 390954 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 391574 572294
rect 390954 536614 391574 572058
rect 390954 536378 390986 536614
rect 391222 536378 391306 536614
rect 391542 536378 391574 536614
rect 390954 536294 391574 536378
rect 390954 536058 390986 536294
rect 391222 536058 391306 536294
rect 391542 536058 391574 536294
rect 390954 500614 391574 536058
rect 390954 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 391574 500614
rect 390954 500294 391574 500378
rect 390954 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 391574 500294
rect 390954 464614 391574 500058
rect 390954 464378 390986 464614
rect 391222 464378 391306 464614
rect 391542 464378 391574 464614
rect 390954 464294 391574 464378
rect 390954 464058 390986 464294
rect 391222 464058 391306 464294
rect 391542 464058 391574 464294
rect 390954 428614 391574 464058
rect 390954 428378 390986 428614
rect 391222 428378 391306 428614
rect 391542 428378 391574 428614
rect 390954 428294 391574 428378
rect 390954 428058 390986 428294
rect 391222 428058 391306 428294
rect 391542 428058 391574 428294
rect 390954 392614 391574 428058
rect 390954 392378 390986 392614
rect 391222 392378 391306 392614
rect 391542 392378 391574 392614
rect 390954 392294 391574 392378
rect 390954 392058 390986 392294
rect 391222 392058 391306 392294
rect 391542 392058 391574 392294
rect 390954 356614 391574 392058
rect 390954 356378 390986 356614
rect 391222 356378 391306 356614
rect 391542 356378 391574 356614
rect 390954 356294 391574 356378
rect 390954 356058 390986 356294
rect 391222 356058 391306 356294
rect 391542 356058 391574 356294
rect 390954 320614 391574 356058
rect 390954 320378 390986 320614
rect 391222 320378 391306 320614
rect 391542 320378 391574 320614
rect 390954 320294 391574 320378
rect 390954 320058 390986 320294
rect 391222 320058 391306 320294
rect 391542 320058 391574 320294
rect 390954 284614 391574 320058
rect 390954 284378 390986 284614
rect 391222 284378 391306 284614
rect 391542 284378 391574 284614
rect 390954 284294 391574 284378
rect 390954 284058 390986 284294
rect 391222 284058 391306 284294
rect 391542 284058 391574 284294
rect 390954 248614 391574 284058
rect 390954 248378 390986 248614
rect 391222 248378 391306 248614
rect 391542 248378 391574 248614
rect 390954 248294 391574 248378
rect 390954 248058 390986 248294
rect 391222 248058 391306 248294
rect 391542 248058 391574 248294
rect 390954 212614 391574 248058
rect 390954 212378 390986 212614
rect 391222 212378 391306 212614
rect 391542 212378 391574 212614
rect 390954 212294 391574 212378
rect 390954 212058 390986 212294
rect 391222 212058 391306 212294
rect 391542 212058 391574 212294
rect 390954 176614 391574 212058
rect 390954 176378 390986 176614
rect 391222 176378 391306 176614
rect 391542 176378 391574 176614
rect 390954 176294 391574 176378
rect 390954 176058 390986 176294
rect 391222 176058 391306 176294
rect 391542 176058 391574 176294
rect 390954 140614 391574 176058
rect 390954 140378 390986 140614
rect 391222 140378 391306 140614
rect 391542 140378 391574 140614
rect 390954 140294 391574 140378
rect 390954 140058 390986 140294
rect 391222 140058 391306 140294
rect 391542 140058 391574 140294
rect 390954 104614 391574 140058
rect 390954 104378 390986 104614
rect 391222 104378 391306 104614
rect 391542 104378 391574 104614
rect 390954 104294 391574 104378
rect 390954 104058 390986 104294
rect 391222 104058 391306 104294
rect 391542 104058 391574 104294
rect 390954 68614 391574 104058
rect 390954 68378 390986 68614
rect 391222 68378 391306 68614
rect 391542 68378 391574 68614
rect 390954 68294 391574 68378
rect 390954 68058 390986 68294
rect 391222 68058 391306 68294
rect 391542 68058 391574 68294
rect 390954 32614 391574 68058
rect 390954 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 391574 32614
rect 390954 32294 391574 32378
rect 390954 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 391574 32294
rect 372954 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 373574 -6106
rect 372954 -6426 373574 -6342
rect 372954 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 373574 -6426
rect 372954 -7654 373574 -6662
rect 390954 -7066 391574 32058
rect 397794 704838 398414 705830
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 397794 363454 398414 398898
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 219454 398414 254898
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397794 147454 398414 182898
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -1894 398414 -902
rect 401514 691174 402134 706202
rect 401514 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 402134 691174
rect 401514 690854 402134 690938
rect 401514 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 402134 690854
rect 401514 655174 402134 690618
rect 401514 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 402134 655174
rect 401514 654854 402134 654938
rect 401514 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 402134 654854
rect 401514 619174 402134 654618
rect 401514 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 402134 619174
rect 401514 618854 402134 618938
rect 401514 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 402134 618854
rect 401514 583174 402134 618618
rect 401514 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 402134 583174
rect 401514 582854 402134 582938
rect 401514 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 402134 582854
rect 401514 547174 402134 582618
rect 401514 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 402134 547174
rect 401514 546854 402134 546938
rect 401514 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 402134 546854
rect 401514 511174 402134 546618
rect 401514 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 402134 511174
rect 401514 510854 402134 510938
rect 401514 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 402134 510854
rect 401514 475174 402134 510618
rect 401514 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 402134 475174
rect 401514 474854 402134 474938
rect 401514 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 402134 474854
rect 401514 439174 402134 474618
rect 401514 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 402134 439174
rect 401514 438854 402134 438938
rect 401514 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 402134 438854
rect 401514 403174 402134 438618
rect 401514 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 402134 403174
rect 401514 402854 402134 402938
rect 401514 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 402134 402854
rect 401514 367174 402134 402618
rect 401514 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 402134 367174
rect 401514 366854 402134 366938
rect 401514 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 402134 366854
rect 401514 331174 402134 366618
rect 401514 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 402134 331174
rect 401514 330854 402134 330938
rect 401514 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 402134 330854
rect 401514 295174 402134 330618
rect 401514 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 402134 295174
rect 401514 294854 402134 294938
rect 401514 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 402134 294854
rect 401514 259174 402134 294618
rect 401514 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 402134 259174
rect 401514 258854 402134 258938
rect 401514 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 402134 258854
rect 401514 223174 402134 258618
rect 401514 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 402134 223174
rect 401514 222854 402134 222938
rect 401514 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 402134 222854
rect 401514 187174 402134 222618
rect 401514 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 402134 187174
rect 401514 186854 402134 186938
rect 401514 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 402134 186854
rect 401514 151174 402134 186618
rect 401514 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 402134 151174
rect 401514 150854 402134 150938
rect 401514 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 402134 150854
rect 401514 115174 402134 150618
rect 401514 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 402134 115174
rect 401514 114854 402134 114938
rect 401514 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 402134 114854
rect 401514 79174 402134 114618
rect 401514 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 402134 79174
rect 401514 78854 402134 78938
rect 401514 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 402134 78854
rect 401514 43174 402134 78618
rect 401514 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 402134 43174
rect 401514 42854 402134 42938
rect 401514 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 402134 42854
rect 401514 7174 402134 42618
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 401514 -2266 402134 6618
rect 401514 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 402134 -2266
rect 401514 -2586 402134 -2502
rect 401514 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 402134 -2586
rect 401514 -3814 402134 -2822
rect 405234 694894 405854 708122
rect 405234 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 405854 694894
rect 405234 694574 405854 694658
rect 405234 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 405854 694574
rect 405234 658894 405854 694338
rect 405234 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 405854 658894
rect 405234 658574 405854 658658
rect 405234 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 405854 658574
rect 405234 622894 405854 658338
rect 405234 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 405854 622894
rect 405234 622574 405854 622658
rect 405234 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 405854 622574
rect 405234 586894 405854 622338
rect 405234 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 405854 586894
rect 405234 586574 405854 586658
rect 405234 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 405854 586574
rect 405234 550894 405854 586338
rect 405234 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 405854 550894
rect 405234 550574 405854 550658
rect 405234 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 405854 550574
rect 405234 514894 405854 550338
rect 405234 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 405854 514894
rect 405234 514574 405854 514658
rect 405234 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 405854 514574
rect 405234 478894 405854 514338
rect 405234 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 405854 478894
rect 405234 478574 405854 478658
rect 405234 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 405854 478574
rect 405234 442894 405854 478338
rect 405234 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 405854 442894
rect 405234 442574 405854 442658
rect 405234 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 405854 442574
rect 405234 406894 405854 442338
rect 405234 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 405854 406894
rect 405234 406574 405854 406658
rect 405234 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 405854 406574
rect 405234 370894 405854 406338
rect 405234 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 405854 370894
rect 405234 370574 405854 370658
rect 405234 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 405854 370574
rect 405234 334894 405854 370338
rect 405234 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 405854 334894
rect 405234 334574 405854 334658
rect 405234 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 405854 334574
rect 405234 298894 405854 334338
rect 405234 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 405854 298894
rect 405234 298574 405854 298658
rect 405234 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 405854 298574
rect 405234 262894 405854 298338
rect 405234 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 405854 262894
rect 405234 262574 405854 262658
rect 405234 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 405854 262574
rect 405234 226894 405854 262338
rect 405234 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 405854 226894
rect 405234 226574 405854 226658
rect 405234 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 405854 226574
rect 405234 190894 405854 226338
rect 405234 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 405854 190894
rect 405234 190574 405854 190658
rect 405234 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 405854 190574
rect 405234 154894 405854 190338
rect 405234 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 405854 154894
rect 405234 154574 405854 154658
rect 405234 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 405854 154574
rect 405234 118894 405854 154338
rect 405234 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 405854 118894
rect 405234 118574 405854 118658
rect 405234 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 405854 118574
rect 405234 82894 405854 118338
rect 405234 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 405854 82894
rect 405234 82574 405854 82658
rect 405234 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 405854 82574
rect 405234 46894 405854 82338
rect 405234 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 405854 46894
rect 405234 46574 405854 46658
rect 405234 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 405854 46574
rect 405234 10894 405854 46338
rect 405234 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 405854 10894
rect 405234 10574 405854 10658
rect 405234 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 405854 10574
rect 405234 -4186 405854 10338
rect 405234 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 405854 -4186
rect 405234 -4506 405854 -4422
rect 405234 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 405854 -4506
rect 405234 -5734 405854 -4742
rect 408954 698614 409574 710042
rect 426954 711558 427574 711590
rect 426954 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 427574 711558
rect 426954 711238 427574 711322
rect 426954 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 427574 711238
rect 423234 709638 423854 709670
rect 423234 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 423854 709638
rect 423234 709318 423854 709402
rect 423234 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 423854 709318
rect 419514 707718 420134 707750
rect 419514 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 420134 707718
rect 419514 707398 420134 707482
rect 419514 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 420134 707398
rect 408954 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 409574 698614
rect 408954 698294 409574 698378
rect 408954 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 409574 698294
rect 408954 662614 409574 698058
rect 408954 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 409574 662614
rect 408954 662294 409574 662378
rect 408954 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 409574 662294
rect 408954 626614 409574 662058
rect 408954 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 409574 626614
rect 408954 626294 409574 626378
rect 408954 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 409574 626294
rect 408954 590614 409574 626058
rect 408954 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 409574 590614
rect 408954 590294 409574 590378
rect 408954 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 409574 590294
rect 408954 554614 409574 590058
rect 408954 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 409574 554614
rect 408954 554294 409574 554378
rect 408954 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 409574 554294
rect 408954 518614 409574 554058
rect 408954 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 409574 518614
rect 408954 518294 409574 518378
rect 408954 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 409574 518294
rect 408954 482614 409574 518058
rect 408954 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 409574 482614
rect 408954 482294 409574 482378
rect 408954 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 409574 482294
rect 408954 446614 409574 482058
rect 408954 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 409574 446614
rect 408954 446294 409574 446378
rect 408954 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 409574 446294
rect 408954 410614 409574 446058
rect 408954 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 409574 410614
rect 408954 410294 409574 410378
rect 408954 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 409574 410294
rect 408954 374614 409574 410058
rect 408954 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 409574 374614
rect 408954 374294 409574 374378
rect 408954 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 409574 374294
rect 408954 338614 409574 374058
rect 408954 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 409574 338614
rect 408954 338294 409574 338378
rect 408954 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 409574 338294
rect 408954 302614 409574 338058
rect 408954 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 409574 302614
rect 408954 302294 409574 302378
rect 408954 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 409574 302294
rect 408954 266614 409574 302058
rect 408954 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 409574 266614
rect 408954 266294 409574 266378
rect 408954 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 409574 266294
rect 408954 230614 409574 266058
rect 408954 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 409574 230614
rect 408954 230294 409574 230378
rect 408954 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 409574 230294
rect 408954 194614 409574 230058
rect 408954 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 409574 194614
rect 408954 194294 409574 194378
rect 408954 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 409574 194294
rect 408954 158614 409574 194058
rect 408954 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 409574 158614
rect 408954 158294 409574 158378
rect 408954 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 409574 158294
rect 408954 122614 409574 158058
rect 408954 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 409574 122614
rect 408954 122294 409574 122378
rect 408954 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 409574 122294
rect 408954 86614 409574 122058
rect 408954 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 409574 86614
rect 408954 86294 409574 86378
rect 408954 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 409574 86294
rect 408954 50614 409574 86058
rect 408954 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 409574 50614
rect 408954 50294 409574 50378
rect 408954 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 409574 50294
rect 408954 14614 409574 50058
rect 408954 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 409574 14614
rect 408954 14294 409574 14378
rect 408954 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 409574 14294
rect 390954 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 391574 -7066
rect 390954 -7386 391574 -7302
rect 390954 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 391574 -7386
rect 390954 -7654 391574 -7622
rect 408954 -6106 409574 14058
rect 415794 705798 416414 705830
rect 415794 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 416414 705798
rect 415794 705478 416414 705562
rect 415794 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 416414 705478
rect 415794 669454 416414 705242
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 561454 416414 596898
rect 415794 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 416414 561454
rect 415794 561134 416414 561218
rect 415794 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 416414 561134
rect 415794 525454 416414 560898
rect 415794 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 416414 525454
rect 415794 525134 416414 525218
rect 415794 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 416414 525134
rect 415794 489454 416414 524898
rect 415794 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 416414 489454
rect 415794 489134 416414 489218
rect 415794 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 416414 489134
rect 415794 453454 416414 488898
rect 415794 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 416414 453454
rect 415794 453134 416414 453218
rect 415794 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 416414 453134
rect 415794 417454 416414 452898
rect 415794 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 416414 417454
rect 415794 417134 416414 417218
rect 415794 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 416414 417134
rect 415794 381454 416414 416898
rect 415794 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 416414 381454
rect 415794 381134 416414 381218
rect 415794 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 416414 381134
rect 415794 345454 416414 380898
rect 415794 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 416414 345454
rect 415794 345134 416414 345218
rect 415794 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 416414 345134
rect 415794 309454 416414 344898
rect 415794 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 416414 309454
rect 415794 309134 416414 309218
rect 415794 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 416414 309134
rect 415794 273454 416414 308898
rect 415794 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 416414 273454
rect 415794 273134 416414 273218
rect 415794 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 416414 273134
rect 415794 237454 416414 272898
rect 415794 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 416414 237454
rect 415794 237134 416414 237218
rect 415794 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 416414 237134
rect 415794 201454 416414 236898
rect 415794 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 416414 201454
rect 415794 201134 416414 201218
rect 415794 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 416414 201134
rect 415794 165454 416414 200898
rect 415794 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 416414 165454
rect 415794 165134 416414 165218
rect 415794 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 416414 165134
rect 415794 129454 416414 164898
rect 415794 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 416414 129454
rect 415794 129134 416414 129218
rect 415794 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 416414 129134
rect 415794 93454 416414 128898
rect 415794 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 416414 93454
rect 415794 93134 416414 93218
rect 415794 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 416414 93134
rect 415794 57454 416414 92898
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -1306 416414 20898
rect 415794 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 416414 -1306
rect 415794 -1626 416414 -1542
rect 415794 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 416414 -1626
rect 415794 -1894 416414 -1862
rect 419514 673174 420134 707162
rect 419514 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 420134 673174
rect 419514 672854 420134 672938
rect 419514 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 420134 672854
rect 419514 637174 420134 672618
rect 419514 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 420134 637174
rect 419514 636854 420134 636938
rect 419514 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 420134 636854
rect 419514 601174 420134 636618
rect 419514 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 420134 601174
rect 419514 600854 420134 600938
rect 419514 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 420134 600854
rect 419514 565174 420134 600618
rect 419514 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 420134 565174
rect 419514 564854 420134 564938
rect 419514 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 420134 564854
rect 419514 529174 420134 564618
rect 419514 528938 419546 529174
rect 419782 528938 419866 529174
rect 420102 528938 420134 529174
rect 419514 528854 420134 528938
rect 419514 528618 419546 528854
rect 419782 528618 419866 528854
rect 420102 528618 420134 528854
rect 419514 493174 420134 528618
rect 419514 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 420134 493174
rect 419514 492854 420134 492938
rect 419514 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 420134 492854
rect 419514 457174 420134 492618
rect 419514 456938 419546 457174
rect 419782 456938 419866 457174
rect 420102 456938 420134 457174
rect 419514 456854 420134 456938
rect 419514 456618 419546 456854
rect 419782 456618 419866 456854
rect 420102 456618 420134 456854
rect 419514 421174 420134 456618
rect 419514 420938 419546 421174
rect 419782 420938 419866 421174
rect 420102 420938 420134 421174
rect 419514 420854 420134 420938
rect 419514 420618 419546 420854
rect 419782 420618 419866 420854
rect 420102 420618 420134 420854
rect 419514 385174 420134 420618
rect 419514 384938 419546 385174
rect 419782 384938 419866 385174
rect 420102 384938 420134 385174
rect 419514 384854 420134 384938
rect 419514 384618 419546 384854
rect 419782 384618 419866 384854
rect 420102 384618 420134 384854
rect 419514 349174 420134 384618
rect 419514 348938 419546 349174
rect 419782 348938 419866 349174
rect 420102 348938 420134 349174
rect 419514 348854 420134 348938
rect 419514 348618 419546 348854
rect 419782 348618 419866 348854
rect 420102 348618 420134 348854
rect 419514 313174 420134 348618
rect 419514 312938 419546 313174
rect 419782 312938 419866 313174
rect 420102 312938 420134 313174
rect 419514 312854 420134 312938
rect 419514 312618 419546 312854
rect 419782 312618 419866 312854
rect 420102 312618 420134 312854
rect 419514 277174 420134 312618
rect 419514 276938 419546 277174
rect 419782 276938 419866 277174
rect 420102 276938 420134 277174
rect 419514 276854 420134 276938
rect 419514 276618 419546 276854
rect 419782 276618 419866 276854
rect 420102 276618 420134 276854
rect 419514 241174 420134 276618
rect 419514 240938 419546 241174
rect 419782 240938 419866 241174
rect 420102 240938 420134 241174
rect 419514 240854 420134 240938
rect 419514 240618 419546 240854
rect 419782 240618 419866 240854
rect 420102 240618 420134 240854
rect 419514 205174 420134 240618
rect 419514 204938 419546 205174
rect 419782 204938 419866 205174
rect 420102 204938 420134 205174
rect 419514 204854 420134 204938
rect 419514 204618 419546 204854
rect 419782 204618 419866 204854
rect 420102 204618 420134 204854
rect 419514 169174 420134 204618
rect 419514 168938 419546 169174
rect 419782 168938 419866 169174
rect 420102 168938 420134 169174
rect 419514 168854 420134 168938
rect 419514 168618 419546 168854
rect 419782 168618 419866 168854
rect 420102 168618 420134 168854
rect 419514 133174 420134 168618
rect 419514 132938 419546 133174
rect 419782 132938 419866 133174
rect 420102 132938 420134 133174
rect 419514 132854 420134 132938
rect 419514 132618 419546 132854
rect 419782 132618 419866 132854
rect 420102 132618 420134 132854
rect 419514 97174 420134 132618
rect 419514 96938 419546 97174
rect 419782 96938 419866 97174
rect 420102 96938 420134 97174
rect 419514 96854 420134 96938
rect 419514 96618 419546 96854
rect 419782 96618 419866 96854
rect 420102 96618 420134 96854
rect 419514 61174 420134 96618
rect 419514 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 420134 61174
rect 419514 60854 420134 60938
rect 419514 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 420134 60854
rect 419514 25174 420134 60618
rect 419514 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 420134 25174
rect 419514 24854 420134 24938
rect 419514 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 420134 24854
rect 419514 -3226 420134 24618
rect 419514 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 420134 -3226
rect 419514 -3546 420134 -3462
rect 419514 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 420134 -3546
rect 419514 -3814 420134 -3782
rect 423234 676894 423854 709082
rect 423234 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 423854 676894
rect 423234 676574 423854 676658
rect 423234 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 423854 676574
rect 423234 640894 423854 676338
rect 423234 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 423854 640894
rect 423234 640574 423854 640658
rect 423234 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 423854 640574
rect 423234 604894 423854 640338
rect 423234 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 423854 604894
rect 423234 604574 423854 604658
rect 423234 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 423854 604574
rect 423234 568894 423854 604338
rect 423234 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 423854 568894
rect 423234 568574 423854 568658
rect 423234 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 423854 568574
rect 423234 532894 423854 568338
rect 423234 532658 423266 532894
rect 423502 532658 423586 532894
rect 423822 532658 423854 532894
rect 423234 532574 423854 532658
rect 423234 532338 423266 532574
rect 423502 532338 423586 532574
rect 423822 532338 423854 532574
rect 423234 496894 423854 532338
rect 423234 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 423854 496894
rect 423234 496574 423854 496658
rect 423234 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 423854 496574
rect 423234 460894 423854 496338
rect 423234 460658 423266 460894
rect 423502 460658 423586 460894
rect 423822 460658 423854 460894
rect 423234 460574 423854 460658
rect 423234 460338 423266 460574
rect 423502 460338 423586 460574
rect 423822 460338 423854 460574
rect 423234 424894 423854 460338
rect 423234 424658 423266 424894
rect 423502 424658 423586 424894
rect 423822 424658 423854 424894
rect 423234 424574 423854 424658
rect 423234 424338 423266 424574
rect 423502 424338 423586 424574
rect 423822 424338 423854 424574
rect 423234 388894 423854 424338
rect 423234 388658 423266 388894
rect 423502 388658 423586 388894
rect 423822 388658 423854 388894
rect 423234 388574 423854 388658
rect 423234 388338 423266 388574
rect 423502 388338 423586 388574
rect 423822 388338 423854 388574
rect 423234 352894 423854 388338
rect 423234 352658 423266 352894
rect 423502 352658 423586 352894
rect 423822 352658 423854 352894
rect 423234 352574 423854 352658
rect 423234 352338 423266 352574
rect 423502 352338 423586 352574
rect 423822 352338 423854 352574
rect 423234 316894 423854 352338
rect 423234 316658 423266 316894
rect 423502 316658 423586 316894
rect 423822 316658 423854 316894
rect 423234 316574 423854 316658
rect 423234 316338 423266 316574
rect 423502 316338 423586 316574
rect 423822 316338 423854 316574
rect 423234 280894 423854 316338
rect 423234 280658 423266 280894
rect 423502 280658 423586 280894
rect 423822 280658 423854 280894
rect 423234 280574 423854 280658
rect 423234 280338 423266 280574
rect 423502 280338 423586 280574
rect 423822 280338 423854 280574
rect 423234 244894 423854 280338
rect 423234 244658 423266 244894
rect 423502 244658 423586 244894
rect 423822 244658 423854 244894
rect 423234 244574 423854 244658
rect 423234 244338 423266 244574
rect 423502 244338 423586 244574
rect 423822 244338 423854 244574
rect 423234 208894 423854 244338
rect 423234 208658 423266 208894
rect 423502 208658 423586 208894
rect 423822 208658 423854 208894
rect 423234 208574 423854 208658
rect 423234 208338 423266 208574
rect 423502 208338 423586 208574
rect 423822 208338 423854 208574
rect 423234 172894 423854 208338
rect 423234 172658 423266 172894
rect 423502 172658 423586 172894
rect 423822 172658 423854 172894
rect 423234 172574 423854 172658
rect 423234 172338 423266 172574
rect 423502 172338 423586 172574
rect 423822 172338 423854 172574
rect 423234 136894 423854 172338
rect 423234 136658 423266 136894
rect 423502 136658 423586 136894
rect 423822 136658 423854 136894
rect 423234 136574 423854 136658
rect 423234 136338 423266 136574
rect 423502 136338 423586 136574
rect 423822 136338 423854 136574
rect 423234 100894 423854 136338
rect 423234 100658 423266 100894
rect 423502 100658 423586 100894
rect 423822 100658 423854 100894
rect 423234 100574 423854 100658
rect 423234 100338 423266 100574
rect 423502 100338 423586 100574
rect 423822 100338 423854 100574
rect 423234 64894 423854 100338
rect 423234 64658 423266 64894
rect 423502 64658 423586 64894
rect 423822 64658 423854 64894
rect 423234 64574 423854 64658
rect 423234 64338 423266 64574
rect 423502 64338 423586 64574
rect 423822 64338 423854 64574
rect 423234 28894 423854 64338
rect 423234 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 423854 28894
rect 423234 28574 423854 28658
rect 423234 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 423854 28574
rect 423234 -5146 423854 28338
rect 423234 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 423854 -5146
rect 423234 -5466 423854 -5382
rect 423234 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 423854 -5466
rect 423234 -5734 423854 -5702
rect 426954 680614 427574 711002
rect 444954 710598 445574 711590
rect 444954 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 445574 710598
rect 444954 710278 445574 710362
rect 444954 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 445574 710278
rect 441234 708678 441854 709670
rect 441234 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 441854 708678
rect 441234 708358 441854 708442
rect 441234 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 441854 708358
rect 437514 706758 438134 707750
rect 437514 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 438134 706758
rect 437514 706438 438134 706522
rect 437514 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 438134 706438
rect 426954 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 427574 680614
rect 426954 680294 427574 680378
rect 426954 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 427574 680294
rect 426954 644614 427574 680058
rect 426954 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 427574 644614
rect 426954 644294 427574 644378
rect 426954 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 427574 644294
rect 426954 608614 427574 644058
rect 426954 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 427574 608614
rect 426954 608294 427574 608378
rect 426954 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 427574 608294
rect 426954 572614 427574 608058
rect 426954 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 427574 572614
rect 426954 572294 427574 572378
rect 426954 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 427574 572294
rect 426954 536614 427574 572058
rect 426954 536378 426986 536614
rect 427222 536378 427306 536614
rect 427542 536378 427574 536614
rect 426954 536294 427574 536378
rect 426954 536058 426986 536294
rect 427222 536058 427306 536294
rect 427542 536058 427574 536294
rect 426954 500614 427574 536058
rect 426954 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 427574 500614
rect 426954 500294 427574 500378
rect 426954 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 427574 500294
rect 426954 464614 427574 500058
rect 426954 464378 426986 464614
rect 427222 464378 427306 464614
rect 427542 464378 427574 464614
rect 426954 464294 427574 464378
rect 426954 464058 426986 464294
rect 427222 464058 427306 464294
rect 427542 464058 427574 464294
rect 426954 428614 427574 464058
rect 426954 428378 426986 428614
rect 427222 428378 427306 428614
rect 427542 428378 427574 428614
rect 426954 428294 427574 428378
rect 426954 428058 426986 428294
rect 427222 428058 427306 428294
rect 427542 428058 427574 428294
rect 426954 392614 427574 428058
rect 426954 392378 426986 392614
rect 427222 392378 427306 392614
rect 427542 392378 427574 392614
rect 426954 392294 427574 392378
rect 426954 392058 426986 392294
rect 427222 392058 427306 392294
rect 427542 392058 427574 392294
rect 426954 356614 427574 392058
rect 433794 704838 434414 705830
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 435454 434414 470898
rect 433794 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 434414 435454
rect 433794 435134 434414 435218
rect 433794 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 434414 435134
rect 433794 399454 434414 434898
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 372000 434414 398898
rect 437514 691174 438134 706202
rect 437514 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 438134 691174
rect 437514 690854 438134 690938
rect 437514 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 438134 690854
rect 437514 655174 438134 690618
rect 437514 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 438134 655174
rect 437514 654854 438134 654938
rect 437514 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 438134 654854
rect 437514 619174 438134 654618
rect 437514 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 438134 619174
rect 437514 618854 438134 618938
rect 437514 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 438134 618854
rect 437514 583174 438134 618618
rect 437514 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 438134 583174
rect 437514 582854 438134 582938
rect 437514 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 438134 582854
rect 437514 547174 438134 582618
rect 437514 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 438134 547174
rect 437514 546854 438134 546938
rect 437514 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 438134 546854
rect 437514 511174 438134 546618
rect 437514 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 438134 511174
rect 437514 510854 438134 510938
rect 437514 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 438134 510854
rect 437514 475174 438134 510618
rect 437514 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 438134 475174
rect 437514 474854 438134 474938
rect 437514 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 438134 474854
rect 437514 439174 438134 474618
rect 437514 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 438134 439174
rect 437514 438854 438134 438938
rect 437514 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 438134 438854
rect 437514 403174 438134 438618
rect 437514 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 438134 403174
rect 437514 402854 438134 402938
rect 437514 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 438134 402854
rect 437514 372000 438134 402618
rect 441234 694894 441854 708122
rect 441234 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 441854 694894
rect 441234 694574 441854 694658
rect 441234 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 441854 694574
rect 441234 658894 441854 694338
rect 441234 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 441854 658894
rect 441234 658574 441854 658658
rect 441234 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 441854 658574
rect 441234 622894 441854 658338
rect 441234 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 441854 622894
rect 441234 622574 441854 622658
rect 441234 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 441854 622574
rect 441234 586894 441854 622338
rect 441234 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 441854 586894
rect 441234 586574 441854 586658
rect 441234 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 441854 586574
rect 441234 550894 441854 586338
rect 441234 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 441854 550894
rect 441234 550574 441854 550658
rect 441234 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 441854 550574
rect 441234 514894 441854 550338
rect 441234 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 441854 514894
rect 441234 514574 441854 514658
rect 441234 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 441854 514574
rect 441234 478894 441854 514338
rect 441234 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 441854 478894
rect 441234 478574 441854 478658
rect 441234 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 441854 478574
rect 441234 442894 441854 478338
rect 441234 442658 441266 442894
rect 441502 442658 441586 442894
rect 441822 442658 441854 442894
rect 441234 442574 441854 442658
rect 441234 442338 441266 442574
rect 441502 442338 441586 442574
rect 441822 442338 441854 442574
rect 441234 406894 441854 442338
rect 441234 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 441854 406894
rect 441234 406574 441854 406658
rect 441234 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 441854 406574
rect 441234 372000 441854 406338
rect 444954 698614 445574 710042
rect 462954 711558 463574 711590
rect 462954 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 463574 711558
rect 462954 711238 463574 711322
rect 462954 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 463574 711238
rect 459234 709638 459854 709670
rect 459234 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 459854 709638
rect 459234 709318 459854 709402
rect 459234 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 459854 709318
rect 455514 707718 456134 707750
rect 455514 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 456134 707718
rect 455514 707398 456134 707482
rect 455514 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 456134 707398
rect 444954 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 445574 698614
rect 444954 698294 445574 698378
rect 444954 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 445574 698294
rect 444954 662614 445574 698058
rect 444954 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 445574 662614
rect 444954 662294 445574 662378
rect 444954 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 445574 662294
rect 444954 626614 445574 662058
rect 444954 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 445574 626614
rect 444954 626294 445574 626378
rect 444954 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 445574 626294
rect 444954 590614 445574 626058
rect 444954 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 445574 590614
rect 444954 590294 445574 590378
rect 444954 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 445574 590294
rect 444954 554614 445574 590058
rect 444954 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 445574 554614
rect 444954 554294 445574 554378
rect 444954 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 445574 554294
rect 444954 518614 445574 554058
rect 444954 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 445574 518614
rect 444954 518294 445574 518378
rect 444954 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 445574 518294
rect 444954 482614 445574 518058
rect 444954 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 445574 482614
rect 444954 482294 445574 482378
rect 444954 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 445574 482294
rect 444954 446614 445574 482058
rect 444954 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 445574 446614
rect 444954 446294 445574 446378
rect 444954 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 445574 446294
rect 444954 410614 445574 446058
rect 444954 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 445574 410614
rect 444954 410294 445574 410378
rect 444954 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 445574 410294
rect 444954 374614 445574 410058
rect 444954 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 445574 374614
rect 444954 374294 445574 374378
rect 444954 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 445574 374294
rect 434243 363454 434563 363486
rect 434243 363218 434285 363454
rect 434521 363218 434563 363454
rect 434243 363134 434563 363218
rect 434243 362898 434285 363134
rect 434521 362898 434563 363134
rect 434243 362866 434563 362898
rect 436840 363454 437160 363486
rect 436840 363218 436882 363454
rect 437118 363218 437160 363454
rect 436840 363134 437160 363218
rect 436840 362898 436882 363134
rect 437118 362898 437160 363134
rect 436840 362866 437160 362898
rect 439437 363454 439757 363486
rect 439437 363218 439479 363454
rect 439715 363218 439757 363454
rect 439437 363134 439757 363218
rect 439437 362898 439479 363134
rect 439715 362898 439757 363134
rect 439437 362866 439757 362898
rect 426954 356378 426986 356614
rect 427222 356378 427306 356614
rect 427542 356378 427574 356614
rect 426954 356294 427574 356378
rect 426954 356058 426986 356294
rect 427222 356058 427306 356294
rect 427542 356058 427574 356294
rect 426954 320614 427574 356058
rect 435541 345454 435861 345486
rect 435541 345218 435583 345454
rect 435819 345218 435861 345454
rect 435541 345134 435861 345218
rect 435541 344898 435583 345134
rect 435819 344898 435861 345134
rect 435541 344866 435861 344898
rect 438138 345454 438458 345486
rect 438138 345218 438180 345454
rect 438416 345218 438458 345454
rect 438138 345134 438458 345218
rect 438138 344898 438180 345134
rect 438416 344898 438458 345134
rect 438138 344866 438458 344898
rect 444954 338614 445574 374058
rect 444954 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 445574 338614
rect 444954 338294 445574 338378
rect 444954 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 445574 338294
rect 426954 320378 426986 320614
rect 427222 320378 427306 320614
rect 427542 320378 427574 320614
rect 426954 320294 427574 320378
rect 426954 320058 426986 320294
rect 427222 320058 427306 320294
rect 427542 320058 427574 320294
rect 426954 284614 427574 320058
rect 433794 327454 434414 338000
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 300000 434414 326898
rect 437514 331174 438134 338000
rect 437514 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 438134 331174
rect 437514 330854 438134 330938
rect 437514 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 438134 330854
rect 437514 300000 438134 330618
rect 441234 334894 441854 338000
rect 441234 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 441854 334894
rect 441234 334574 441854 334658
rect 441234 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 441854 334574
rect 441234 300000 441854 334338
rect 444954 302614 445574 338058
rect 444954 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 445574 302614
rect 444954 302294 445574 302378
rect 444954 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 445574 302294
rect 434243 291454 434563 291486
rect 434243 291218 434285 291454
rect 434521 291218 434563 291454
rect 434243 291134 434563 291218
rect 434243 290898 434285 291134
rect 434521 290898 434563 291134
rect 434243 290866 434563 290898
rect 436840 291454 437160 291486
rect 436840 291218 436882 291454
rect 437118 291218 437160 291454
rect 436840 291134 437160 291218
rect 436840 290898 436882 291134
rect 437118 290898 437160 291134
rect 436840 290866 437160 290898
rect 439437 291454 439757 291486
rect 439437 291218 439479 291454
rect 439715 291218 439757 291454
rect 439437 291134 439757 291218
rect 439437 290898 439479 291134
rect 439715 290898 439757 291134
rect 439437 290866 439757 290898
rect 426954 284378 426986 284614
rect 427222 284378 427306 284614
rect 427542 284378 427574 284614
rect 426954 284294 427574 284378
rect 426954 284058 426986 284294
rect 427222 284058 427306 284294
rect 427542 284058 427574 284294
rect 426954 248614 427574 284058
rect 435541 273454 435861 273486
rect 435541 273218 435583 273454
rect 435819 273218 435861 273454
rect 435541 273134 435861 273218
rect 435541 272898 435583 273134
rect 435819 272898 435861 273134
rect 435541 272866 435861 272898
rect 438138 273454 438458 273486
rect 438138 273218 438180 273454
rect 438416 273218 438458 273454
rect 438138 273134 438458 273218
rect 438138 272898 438180 273134
rect 438416 272898 438458 273134
rect 438138 272866 438458 272898
rect 444954 266614 445574 302058
rect 444954 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 445574 266614
rect 444954 266294 445574 266378
rect 444954 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 445574 266294
rect 426954 248378 426986 248614
rect 427222 248378 427306 248614
rect 427542 248378 427574 248614
rect 426954 248294 427574 248378
rect 426954 248058 426986 248294
rect 427222 248058 427306 248294
rect 427542 248058 427574 248294
rect 426954 212614 427574 248058
rect 433794 255454 434414 266000
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 228000 434414 254898
rect 437514 259174 438134 266000
rect 437514 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 438134 259174
rect 437514 258854 438134 258938
rect 437514 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 438134 258854
rect 437514 228000 438134 258618
rect 441234 262894 441854 266000
rect 441234 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 441854 262894
rect 441234 262574 441854 262658
rect 441234 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 441854 262574
rect 441234 228000 441854 262338
rect 444954 230614 445574 266058
rect 444954 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 445574 230614
rect 444954 230294 445574 230378
rect 444954 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 445574 230294
rect 434243 219454 434563 219486
rect 434243 219218 434285 219454
rect 434521 219218 434563 219454
rect 434243 219134 434563 219218
rect 434243 218898 434285 219134
rect 434521 218898 434563 219134
rect 434243 218866 434563 218898
rect 436840 219454 437160 219486
rect 436840 219218 436882 219454
rect 437118 219218 437160 219454
rect 436840 219134 437160 219218
rect 436840 218898 436882 219134
rect 437118 218898 437160 219134
rect 436840 218866 437160 218898
rect 439437 219454 439757 219486
rect 439437 219218 439479 219454
rect 439715 219218 439757 219454
rect 439437 219134 439757 219218
rect 439437 218898 439479 219134
rect 439715 218898 439757 219134
rect 439437 218866 439757 218898
rect 426954 212378 426986 212614
rect 427222 212378 427306 212614
rect 427542 212378 427574 212614
rect 426954 212294 427574 212378
rect 426954 212058 426986 212294
rect 427222 212058 427306 212294
rect 427542 212058 427574 212294
rect 426954 176614 427574 212058
rect 435541 201454 435861 201486
rect 435541 201218 435583 201454
rect 435819 201218 435861 201454
rect 435541 201134 435861 201218
rect 435541 200898 435583 201134
rect 435819 200898 435861 201134
rect 435541 200866 435861 200898
rect 438138 201454 438458 201486
rect 438138 201218 438180 201454
rect 438416 201218 438458 201454
rect 438138 201134 438458 201218
rect 438138 200898 438180 201134
rect 438416 200898 438458 201134
rect 438138 200866 438458 200898
rect 444954 194614 445574 230058
rect 444954 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 445574 194614
rect 444954 194294 445574 194378
rect 444954 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 445574 194294
rect 426954 176378 426986 176614
rect 427222 176378 427306 176614
rect 427542 176378 427574 176614
rect 426954 176294 427574 176378
rect 426954 176058 426986 176294
rect 427222 176058 427306 176294
rect 427542 176058 427574 176294
rect 426954 140614 427574 176058
rect 433794 183454 434414 194000
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 433794 156000 434414 182898
rect 437514 187174 438134 194000
rect 437514 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 438134 187174
rect 437514 186854 438134 186938
rect 437514 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 438134 186854
rect 437514 156000 438134 186618
rect 441234 190894 441854 194000
rect 441234 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 441854 190894
rect 441234 190574 441854 190658
rect 441234 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 441854 190574
rect 441234 156000 441854 190338
rect 444954 158614 445574 194058
rect 444954 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 445574 158614
rect 444954 158294 445574 158378
rect 444954 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 445574 158294
rect 434243 147454 434563 147486
rect 434243 147218 434285 147454
rect 434521 147218 434563 147454
rect 434243 147134 434563 147218
rect 434243 146898 434285 147134
rect 434521 146898 434563 147134
rect 434243 146866 434563 146898
rect 436840 147454 437160 147486
rect 436840 147218 436882 147454
rect 437118 147218 437160 147454
rect 436840 147134 437160 147218
rect 436840 146898 436882 147134
rect 437118 146898 437160 147134
rect 436840 146866 437160 146898
rect 439437 147454 439757 147486
rect 439437 147218 439479 147454
rect 439715 147218 439757 147454
rect 439437 147134 439757 147218
rect 439437 146898 439479 147134
rect 439715 146898 439757 147134
rect 439437 146866 439757 146898
rect 426954 140378 426986 140614
rect 427222 140378 427306 140614
rect 427542 140378 427574 140614
rect 426954 140294 427574 140378
rect 426954 140058 426986 140294
rect 427222 140058 427306 140294
rect 427542 140058 427574 140294
rect 426954 104614 427574 140058
rect 435541 129454 435861 129486
rect 435541 129218 435583 129454
rect 435819 129218 435861 129454
rect 435541 129134 435861 129218
rect 435541 128898 435583 129134
rect 435819 128898 435861 129134
rect 435541 128866 435861 128898
rect 438138 129454 438458 129486
rect 438138 129218 438180 129454
rect 438416 129218 438458 129454
rect 438138 129134 438458 129218
rect 438138 128898 438180 129134
rect 438416 128898 438458 129134
rect 438138 128866 438458 128898
rect 444954 122614 445574 158058
rect 444954 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 445574 122614
rect 444954 122294 445574 122378
rect 444954 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 445574 122294
rect 426954 104378 426986 104614
rect 427222 104378 427306 104614
rect 427542 104378 427574 104614
rect 426954 104294 427574 104378
rect 426954 104058 426986 104294
rect 427222 104058 427306 104294
rect 427542 104058 427574 104294
rect 426954 68614 427574 104058
rect 426954 68378 426986 68614
rect 427222 68378 427306 68614
rect 427542 68378 427574 68614
rect 426954 68294 427574 68378
rect 426954 68058 426986 68294
rect 427222 68058 427306 68294
rect 427542 68058 427574 68294
rect 426954 32614 427574 68058
rect 426954 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 427574 32614
rect 426954 32294 427574 32378
rect 426954 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 427574 32294
rect 408954 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 409574 -6106
rect 408954 -6426 409574 -6342
rect 408954 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 409574 -6426
rect 408954 -7654 409574 -6662
rect 426954 -7066 427574 32058
rect 433794 111454 434414 122000
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -1894 434414 -902
rect 437514 115174 438134 122000
rect 437514 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 438134 115174
rect 437514 114854 438134 114938
rect 437514 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 438134 114854
rect 437514 79174 438134 114618
rect 437514 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 438134 79174
rect 437514 78854 438134 78938
rect 437514 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 438134 78854
rect 437514 43174 438134 78618
rect 437514 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 438134 43174
rect 437514 42854 438134 42938
rect 437514 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 438134 42854
rect 437514 7174 438134 42618
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -2266 438134 6618
rect 437514 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 438134 -2266
rect 437514 -2586 438134 -2502
rect 437514 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 438134 -2586
rect 437514 -3814 438134 -2822
rect 441234 118894 441854 122000
rect 441234 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 441854 118894
rect 441234 118574 441854 118658
rect 441234 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 441854 118574
rect 441234 82894 441854 118338
rect 441234 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 441854 82894
rect 441234 82574 441854 82658
rect 441234 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 441854 82574
rect 441234 46894 441854 82338
rect 441234 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 441854 46894
rect 441234 46574 441854 46658
rect 441234 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 441854 46574
rect 441234 10894 441854 46338
rect 441234 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 441854 10894
rect 441234 10574 441854 10658
rect 441234 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 441854 10574
rect 441234 -4186 441854 10338
rect 441234 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 441854 -4186
rect 441234 -4506 441854 -4422
rect 441234 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 441854 -4506
rect 441234 -5734 441854 -4742
rect 444954 86614 445574 122058
rect 444954 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 445574 86614
rect 444954 86294 445574 86378
rect 444954 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 445574 86294
rect 444954 50614 445574 86058
rect 444954 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 445574 50614
rect 444954 50294 445574 50378
rect 444954 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 445574 50294
rect 444954 14614 445574 50058
rect 444954 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 445574 14614
rect 444954 14294 445574 14378
rect 444954 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 445574 14294
rect 426954 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 427574 -7066
rect 426954 -7386 427574 -7302
rect 426954 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 427574 -7386
rect 426954 -7654 427574 -7622
rect 444954 -6106 445574 14058
rect 451794 705798 452414 705830
rect 451794 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 452414 705798
rect 451794 705478 452414 705562
rect 451794 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 452414 705478
rect 451794 669454 452414 705242
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 453454 452414 488898
rect 451794 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 452414 453454
rect 451794 453134 452414 453218
rect 451794 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 452414 453134
rect 451794 417454 452414 452898
rect 451794 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 452414 417454
rect 451794 417134 452414 417218
rect 451794 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 452414 417134
rect 451794 381454 452414 416898
rect 451794 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 452414 381454
rect 451794 381134 452414 381218
rect 451794 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 452414 381134
rect 451794 345454 452414 380898
rect 451794 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 452414 345454
rect 451794 345134 452414 345218
rect 451794 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 452414 345134
rect 451794 309454 452414 344898
rect 451794 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 452414 309454
rect 451794 309134 452414 309218
rect 451794 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 452414 309134
rect 451794 273454 452414 308898
rect 451794 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 452414 273454
rect 451794 273134 452414 273218
rect 451794 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 452414 273134
rect 451794 237454 452414 272898
rect 451794 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 452414 237454
rect 451794 237134 452414 237218
rect 451794 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 452414 237134
rect 451794 201454 452414 236898
rect 451794 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 452414 201454
rect 451794 201134 452414 201218
rect 451794 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 452414 201134
rect 451794 165454 452414 200898
rect 451794 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 452414 165454
rect 451794 165134 452414 165218
rect 451794 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 452414 165134
rect 451794 129454 452414 164898
rect 451794 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 452414 129454
rect 451794 129134 452414 129218
rect 451794 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 452414 129134
rect 451794 93454 452414 128898
rect 451794 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 452414 93454
rect 451794 93134 452414 93218
rect 451794 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 452414 93134
rect 451794 57454 452414 92898
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -1306 452414 20898
rect 451794 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 452414 -1306
rect 451794 -1626 452414 -1542
rect 451794 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 452414 -1626
rect 451794 -1894 452414 -1862
rect 455514 673174 456134 707162
rect 455514 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 456134 673174
rect 455514 672854 456134 672938
rect 455514 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 456134 672854
rect 455514 637174 456134 672618
rect 455514 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 456134 637174
rect 455514 636854 456134 636938
rect 455514 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 456134 636854
rect 455514 601174 456134 636618
rect 455514 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 456134 601174
rect 455514 600854 456134 600938
rect 455514 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 456134 600854
rect 455514 565174 456134 600618
rect 455514 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 456134 565174
rect 455514 564854 456134 564938
rect 455514 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 456134 564854
rect 455514 529174 456134 564618
rect 455514 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 456134 529174
rect 455514 528854 456134 528938
rect 455514 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 456134 528854
rect 455514 493174 456134 528618
rect 455514 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 456134 493174
rect 455514 492854 456134 492938
rect 455514 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 456134 492854
rect 455514 457174 456134 492618
rect 455514 456938 455546 457174
rect 455782 456938 455866 457174
rect 456102 456938 456134 457174
rect 455514 456854 456134 456938
rect 455514 456618 455546 456854
rect 455782 456618 455866 456854
rect 456102 456618 456134 456854
rect 455514 421174 456134 456618
rect 455514 420938 455546 421174
rect 455782 420938 455866 421174
rect 456102 420938 456134 421174
rect 455514 420854 456134 420938
rect 455514 420618 455546 420854
rect 455782 420618 455866 420854
rect 456102 420618 456134 420854
rect 455514 385174 456134 420618
rect 455514 384938 455546 385174
rect 455782 384938 455866 385174
rect 456102 384938 456134 385174
rect 455514 384854 456134 384938
rect 455514 384618 455546 384854
rect 455782 384618 455866 384854
rect 456102 384618 456134 384854
rect 455514 349174 456134 384618
rect 455514 348938 455546 349174
rect 455782 348938 455866 349174
rect 456102 348938 456134 349174
rect 455514 348854 456134 348938
rect 455514 348618 455546 348854
rect 455782 348618 455866 348854
rect 456102 348618 456134 348854
rect 455514 313174 456134 348618
rect 455514 312938 455546 313174
rect 455782 312938 455866 313174
rect 456102 312938 456134 313174
rect 455514 312854 456134 312938
rect 455514 312618 455546 312854
rect 455782 312618 455866 312854
rect 456102 312618 456134 312854
rect 455514 277174 456134 312618
rect 455514 276938 455546 277174
rect 455782 276938 455866 277174
rect 456102 276938 456134 277174
rect 455514 276854 456134 276938
rect 455514 276618 455546 276854
rect 455782 276618 455866 276854
rect 456102 276618 456134 276854
rect 455514 241174 456134 276618
rect 455514 240938 455546 241174
rect 455782 240938 455866 241174
rect 456102 240938 456134 241174
rect 455514 240854 456134 240938
rect 455514 240618 455546 240854
rect 455782 240618 455866 240854
rect 456102 240618 456134 240854
rect 455514 205174 456134 240618
rect 455514 204938 455546 205174
rect 455782 204938 455866 205174
rect 456102 204938 456134 205174
rect 455514 204854 456134 204938
rect 455514 204618 455546 204854
rect 455782 204618 455866 204854
rect 456102 204618 456134 204854
rect 455514 169174 456134 204618
rect 455514 168938 455546 169174
rect 455782 168938 455866 169174
rect 456102 168938 456134 169174
rect 455514 168854 456134 168938
rect 455514 168618 455546 168854
rect 455782 168618 455866 168854
rect 456102 168618 456134 168854
rect 455514 133174 456134 168618
rect 455514 132938 455546 133174
rect 455782 132938 455866 133174
rect 456102 132938 456134 133174
rect 455514 132854 456134 132938
rect 455514 132618 455546 132854
rect 455782 132618 455866 132854
rect 456102 132618 456134 132854
rect 455514 97174 456134 132618
rect 455514 96938 455546 97174
rect 455782 96938 455866 97174
rect 456102 96938 456134 97174
rect 455514 96854 456134 96938
rect 455514 96618 455546 96854
rect 455782 96618 455866 96854
rect 456102 96618 456134 96854
rect 455514 61174 456134 96618
rect 455514 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 456134 61174
rect 455514 60854 456134 60938
rect 455514 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 456134 60854
rect 455514 25174 456134 60618
rect 455514 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 456134 25174
rect 455514 24854 456134 24938
rect 455514 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 456134 24854
rect 455514 -3226 456134 24618
rect 455514 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 456134 -3226
rect 455514 -3546 456134 -3462
rect 455514 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 456134 -3546
rect 455514 -3814 456134 -3782
rect 459234 676894 459854 709082
rect 459234 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 459854 676894
rect 459234 676574 459854 676658
rect 459234 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 459854 676574
rect 459234 640894 459854 676338
rect 459234 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 459854 640894
rect 459234 640574 459854 640658
rect 459234 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 459854 640574
rect 459234 604894 459854 640338
rect 459234 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 459854 604894
rect 459234 604574 459854 604658
rect 459234 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 459854 604574
rect 459234 568894 459854 604338
rect 459234 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 459854 568894
rect 459234 568574 459854 568658
rect 459234 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 459854 568574
rect 459234 532894 459854 568338
rect 459234 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 459854 532894
rect 459234 532574 459854 532658
rect 459234 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 459854 532574
rect 459234 496894 459854 532338
rect 459234 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 459854 496894
rect 459234 496574 459854 496658
rect 459234 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 459854 496574
rect 459234 460894 459854 496338
rect 459234 460658 459266 460894
rect 459502 460658 459586 460894
rect 459822 460658 459854 460894
rect 459234 460574 459854 460658
rect 459234 460338 459266 460574
rect 459502 460338 459586 460574
rect 459822 460338 459854 460574
rect 459234 424894 459854 460338
rect 459234 424658 459266 424894
rect 459502 424658 459586 424894
rect 459822 424658 459854 424894
rect 459234 424574 459854 424658
rect 459234 424338 459266 424574
rect 459502 424338 459586 424574
rect 459822 424338 459854 424574
rect 459234 388894 459854 424338
rect 459234 388658 459266 388894
rect 459502 388658 459586 388894
rect 459822 388658 459854 388894
rect 459234 388574 459854 388658
rect 459234 388338 459266 388574
rect 459502 388338 459586 388574
rect 459822 388338 459854 388574
rect 459234 352894 459854 388338
rect 459234 352658 459266 352894
rect 459502 352658 459586 352894
rect 459822 352658 459854 352894
rect 459234 352574 459854 352658
rect 459234 352338 459266 352574
rect 459502 352338 459586 352574
rect 459822 352338 459854 352574
rect 459234 316894 459854 352338
rect 459234 316658 459266 316894
rect 459502 316658 459586 316894
rect 459822 316658 459854 316894
rect 459234 316574 459854 316658
rect 459234 316338 459266 316574
rect 459502 316338 459586 316574
rect 459822 316338 459854 316574
rect 459234 280894 459854 316338
rect 459234 280658 459266 280894
rect 459502 280658 459586 280894
rect 459822 280658 459854 280894
rect 459234 280574 459854 280658
rect 459234 280338 459266 280574
rect 459502 280338 459586 280574
rect 459822 280338 459854 280574
rect 459234 244894 459854 280338
rect 459234 244658 459266 244894
rect 459502 244658 459586 244894
rect 459822 244658 459854 244894
rect 459234 244574 459854 244658
rect 459234 244338 459266 244574
rect 459502 244338 459586 244574
rect 459822 244338 459854 244574
rect 459234 208894 459854 244338
rect 459234 208658 459266 208894
rect 459502 208658 459586 208894
rect 459822 208658 459854 208894
rect 459234 208574 459854 208658
rect 459234 208338 459266 208574
rect 459502 208338 459586 208574
rect 459822 208338 459854 208574
rect 459234 172894 459854 208338
rect 459234 172658 459266 172894
rect 459502 172658 459586 172894
rect 459822 172658 459854 172894
rect 459234 172574 459854 172658
rect 459234 172338 459266 172574
rect 459502 172338 459586 172574
rect 459822 172338 459854 172574
rect 459234 136894 459854 172338
rect 459234 136658 459266 136894
rect 459502 136658 459586 136894
rect 459822 136658 459854 136894
rect 459234 136574 459854 136658
rect 459234 136338 459266 136574
rect 459502 136338 459586 136574
rect 459822 136338 459854 136574
rect 459234 100894 459854 136338
rect 459234 100658 459266 100894
rect 459502 100658 459586 100894
rect 459822 100658 459854 100894
rect 459234 100574 459854 100658
rect 459234 100338 459266 100574
rect 459502 100338 459586 100574
rect 459822 100338 459854 100574
rect 459234 64894 459854 100338
rect 459234 64658 459266 64894
rect 459502 64658 459586 64894
rect 459822 64658 459854 64894
rect 459234 64574 459854 64658
rect 459234 64338 459266 64574
rect 459502 64338 459586 64574
rect 459822 64338 459854 64574
rect 459234 28894 459854 64338
rect 459234 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 459854 28894
rect 459234 28574 459854 28658
rect 459234 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 459854 28574
rect 459234 -5146 459854 28338
rect 459234 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 459854 -5146
rect 459234 -5466 459854 -5382
rect 459234 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 459854 -5466
rect 459234 -5734 459854 -5702
rect 462954 680614 463574 711002
rect 480954 710598 481574 711590
rect 480954 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 481574 710598
rect 480954 710278 481574 710362
rect 480954 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 481574 710278
rect 477234 708678 477854 709670
rect 477234 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 477854 708678
rect 477234 708358 477854 708442
rect 477234 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 477854 708358
rect 473514 706758 474134 707750
rect 473514 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 474134 706758
rect 473514 706438 474134 706522
rect 473514 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 474134 706438
rect 462954 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 463574 680614
rect 462954 680294 463574 680378
rect 462954 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 463574 680294
rect 462954 644614 463574 680058
rect 462954 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 463574 644614
rect 462954 644294 463574 644378
rect 462954 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 463574 644294
rect 462954 608614 463574 644058
rect 462954 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 463574 608614
rect 462954 608294 463574 608378
rect 462954 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 463574 608294
rect 462954 572614 463574 608058
rect 462954 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 463574 572614
rect 462954 572294 463574 572378
rect 462954 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 463574 572294
rect 462954 536614 463574 572058
rect 462954 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 463574 536614
rect 462954 536294 463574 536378
rect 462954 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 463574 536294
rect 462954 500614 463574 536058
rect 462954 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 463574 500614
rect 462954 500294 463574 500378
rect 462954 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 463574 500294
rect 462954 464614 463574 500058
rect 462954 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 463574 464614
rect 462954 464294 463574 464378
rect 462954 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 463574 464294
rect 462954 428614 463574 464058
rect 462954 428378 462986 428614
rect 463222 428378 463306 428614
rect 463542 428378 463574 428614
rect 462954 428294 463574 428378
rect 462954 428058 462986 428294
rect 463222 428058 463306 428294
rect 463542 428058 463574 428294
rect 462954 392614 463574 428058
rect 462954 392378 462986 392614
rect 463222 392378 463306 392614
rect 463542 392378 463574 392614
rect 462954 392294 463574 392378
rect 462954 392058 462986 392294
rect 463222 392058 463306 392294
rect 463542 392058 463574 392294
rect 462954 356614 463574 392058
rect 462954 356378 462986 356614
rect 463222 356378 463306 356614
rect 463542 356378 463574 356614
rect 462954 356294 463574 356378
rect 462954 356058 462986 356294
rect 463222 356058 463306 356294
rect 463542 356058 463574 356294
rect 462954 320614 463574 356058
rect 462954 320378 462986 320614
rect 463222 320378 463306 320614
rect 463542 320378 463574 320614
rect 462954 320294 463574 320378
rect 462954 320058 462986 320294
rect 463222 320058 463306 320294
rect 463542 320058 463574 320294
rect 462954 284614 463574 320058
rect 462954 284378 462986 284614
rect 463222 284378 463306 284614
rect 463542 284378 463574 284614
rect 462954 284294 463574 284378
rect 462954 284058 462986 284294
rect 463222 284058 463306 284294
rect 463542 284058 463574 284294
rect 462954 248614 463574 284058
rect 462954 248378 462986 248614
rect 463222 248378 463306 248614
rect 463542 248378 463574 248614
rect 462954 248294 463574 248378
rect 462954 248058 462986 248294
rect 463222 248058 463306 248294
rect 463542 248058 463574 248294
rect 462954 212614 463574 248058
rect 462954 212378 462986 212614
rect 463222 212378 463306 212614
rect 463542 212378 463574 212614
rect 462954 212294 463574 212378
rect 462954 212058 462986 212294
rect 463222 212058 463306 212294
rect 463542 212058 463574 212294
rect 462954 176614 463574 212058
rect 462954 176378 462986 176614
rect 463222 176378 463306 176614
rect 463542 176378 463574 176614
rect 462954 176294 463574 176378
rect 462954 176058 462986 176294
rect 463222 176058 463306 176294
rect 463542 176058 463574 176294
rect 462954 140614 463574 176058
rect 462954 140378 462986 140614
rect 463222 140378 463306 140614
rect 463542 140378 463574 140614
rect 462954 140294 463574 140378
rect 462954 140058 462986 140294
rect 463222 140058 463306 140294
rect 463542 140058 463574 140294
rect 462954 104614 463574 140058
rect 462954 104378 462986 104614
rect 463222 104378 463306 104614
rect 463542 104378 463574 104614
rect 462954 104294 463574 104378
rect 462954 104058 462986 104294
rect 463222 104058 463306 104294
rect 463542 104058 463574 104294
rect 462954 68614 463574 104058
rect 462954 68378 462986 68614
rect 463222 68378 463306 68614
rect 463542 68378 463574 68614
rect 462954 68294 463574 68378
rect 462954 68058 462986 68294
rect 463222 68058 463306 68294
rect 463542 68058 463574 68294
rect 462954 32614 463574 68058
rect 462954 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 463574 32614
rect 462954 32294 463574 32378
rect 462954 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 463574 32294
rect 444954 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 445574 -6106
rect 444954 -6426 445574 -6342
rect 444954 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 445574 -6426
rect 444954 -7654 445574 -6662
rect 462954 -7066 463574 32058
rect 469794 704838 470414 705830
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 363454 470414 398898
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 291454 470414 326898
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -1894 470414 -902
rect 473514 691174 474134 706202
rect 473514 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 474134 691174
rect 473514 690854 474134 690938
rect 473514 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 474134 690854
rect 473514 655174 474134 690618
rect 473514 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 474134 655174
rect 473514 654854 474134 654938
rect 473514 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 474134 654854
rect 473514 619174 474134 654618
rect 473514 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 474134 619174
rect 473514 618854 474134 618938
rect 473514 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 474134 618854
rect 473514 583174 474134 618618
rect 473514 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 474134 583174
rect 473514 582854 474134 582938
rect 473514 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 474134 582854
rect 473514 547174 474134 582618
rect 473514 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 474134 547174
rect 473514 546854 474134 546938
rect 473514 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 474134 546854
rect 473514 511174 474134 546618
rect 473514 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 474134 511174
rect 473514 510854 474134 510938
rect 473514 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 474134 510854
rect 473514 475174 474134 510618
rect 473514 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 474134 475174
rect 473514 474854 474134 474938
rect 473514 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 474134 474854
rect 473514 439174 474134 474618
rect 473514 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 474134 439174
rect 473514 438854 474134 438938
rect 473514 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 474134 438854
rect 473514 403174 474134 438618
rect 473514 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 474134 403174
rect 473514 402854 474134 402938
rect 473514 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 474134 402854
rect 473514 367174 474134 402618
rect 473514 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 474134 367174
rect 473514 366854 474134 366938
rect 473514 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 474134 366854
rect 473514 331174 474134 366618
rect 473514 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 474134 331174
rect 473514 330854 474134 330938
rect 473514 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 474134 330854
rect 473514 295174 474134 330618
rect 473514 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 474134 295174
rect 473514 294854 474134 294938
rect 473514 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 474134 294854
rect 473514 259174 474134 294618
rect 473514 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 474134 259174
rect 473514 258854 474134 258938
rect 473514 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 474134 258854
rect 473514 223174 474134 258618
rect 473514 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 474134 223174
rect 473514 222854 474134 222938
rect 473514 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 474134 222854
rect 473514 187174 474134 222618
rect 473514 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 474134 187174
rect 473514 186854 474134 186938
rect 473514 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 474134 186854
rect 473514 151174 474134 186618
rect 473514 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 474134 151174
rect 473514 150854 474134 150938
rect 473514 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 474134 150854
rect 473514 115174 474134 150618
rect 473514 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 474134 115174
rect 473514 114854 474134 114938
rect 473514 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 474134 114854
rect 473514 79174 474134 114618
rect 473514 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 474134 79174
rect 473514 78854 474134 78938
rect 473514 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 474134 78854
rect 473514 43174 474134 78618
rect 473514 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 474134 43174
rect 473514 42854 474134 42938
rect 473514 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 474134 42854
rect 473514 7174 474134 42618
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -2266 474134 6618
rect 473514 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 474134 -2266
rect 473514 -2586 474134 -2502
rect 473514 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 474134 -2586
rect 473514 -3814 474134 -2822
rect 477234 694894 477854 708122
rect 477234 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 477854 694894
rect 477234 694574 477854 694658
rect 477234 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 477854 694574
rect 477234 658894 477854 694338
rect 477234 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 477854 658894
rect 477234 658574 477854 658658
rect 477234 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 477854 658574
rect 477234 622894 477854 658338
rect 477234 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 477854 622894
rect 477234 622574 477854 622658
rect 477234 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 477854 622574
rect 477234 586894 477854 622338
rect 477234 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 477854 586894
rect 477234 586574 477854 586658
rect 477234 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 477854 586574
rect 477234 550894 477854 586338
rect 477234 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 477854 550894
rect 477234 550574 477854 550658
rect 477234 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 477854 550574
rect 477234 514894 477854 550338
rect 477234 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 477854 514894
rect 477234 514574 477854 514658
rect 477234 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 477854 514574
rect 477234 478894 477854 514338
rect 477234 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 477854 478894
rect 477234 478574 477854 478658
rect 477234 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 477854 478574
rect 477234 442894 477854 478338
rect 477234 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 477854 442894
rect 477234 442574 477854 442658
rect 477234 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 477854 442574
rect 477234 406894 477854 442338
rect 477234 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 477854 406894
rect 477234 406574 477854 406658
rect 477234 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 477854 406574
rect 477234 370894 477854 406338
rect 477234 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 477854 370894
rect 477234 370574 477854 370658
rect 477234 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 477854 370574
rect 477234 334894 477854 370338
rect 477234 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 477854 334894
rect 477234 334574 477854 334658
rect 477234 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 477854 334574
rect 477234 298894 477854 334338
rect 477234 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 477854 298894
rect 477234 298574 477854 298658
rect 477234 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 477854 298574
rect 477234 262894 477854 298338
rect 477234 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 477854 262894
rect 477234 262574 477854 262658
rect 477234 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 477854 262574
rect 477234 226894 477854 262338
rect 477234 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 477854 226894
rect 477234 226574 477854 226658
rect 477234 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 477854 226574
rect 477234 190894 477854 226338
rect 477234 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 477854 190894
rect 477234 190574 477854 190658
rect 477234 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 477854 190574
rect 477234 154894 477854 190338
rect 477234 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 477854 154894
rect 477234 154574 477854 154658
rect 477234 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 477854 154574
rect 477234 118894 477854 154338
rect 477234 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 477854 118894
rect 477234 118574 477854 118658
rect 477234 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 477854 118574
rect 477234 82894 477854 118338
rect 477234 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 477854 82894
rect 477234 82574 477854 82658
rect 477234 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 477854 82574
rect 477234 46894 477854 82338
rect 477234 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 477854 46894
rect 477234 46574 477854 46658
rect 477234 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 477854 46574
rect 477234 10894 477854 46338
rect 477234 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 477854 10894
rect 477234 10574 477854 10658
rect 477234 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 477854 10574
rect 477234 -4186 477854 10338
rect 477234 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 477854 -4186
rect 477234 -4506 477854 -4422
rect 477234 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 477854 -4506
rect 477234 -5734 477854 -4742
rect 480954 698614 481574 710042
rect 498954 711558 499574 711590
rect 498954 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 499574 711558
rect 498954 711238 499574 711322
rect 498954 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 499574 711238
rect 495234 709638 495854 709670
rect 495234 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 495854 709638
rect 495234 709318 495854 709402
rect 495234 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 495854 709318
rect 491514 707718 492134 707750
rect 491514 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 492134 707718
rect 491514 707398 492134 707482
rect 491514 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 492134 707398
rect 480954 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 481574 698614
rect 480954 698294 481574 698378
rect 480954 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 481574 698294
rect 480954 662614 481574 698058
rect 480954 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 481574 662614
rect 480954 662294 481574 662378
rect 480954 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 481574 662294
rect 480954 626614 481574 662058
rect 480954 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 481574 626614
rect 480954 626294 481574 626378
rect 480954 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 481574 626294
rect 480954 590614 481574 626058
rect 480954 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 481574 590614
rect 480954 590294 481574 590378
rect 480954 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 481574 590294
rect 480954 554614 481574 590058
rect 480954 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 481574 554614
rect 480954 554294 481574 554378
rect 480954 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 481574 554294
rect 480954 518614 481574 554058
rect 480954 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 481574 518614
rect 480954 518294 481574 518378
rect 480954 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 481574 518294
rect 480954 482614 481574 518058
rect 480954 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 481574 482614
rect 480954 482294 481574 482378
rect 480954 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 481574 482294
rect 480954 446614 481574 482058
rect 480954 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 481574 446614
rect 480954 446294 481574 446378
rect 480954 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 481574 446294
rect 480954 410614 481574 446058
rect 480954 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 481574 410614
rect 480954 410294 481574 410378
rect 480954 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 481574 410294
rect 480954 374614 481574 410058
rect 480954 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 481574 374614
rect 480954 374294 481574 374378
rect 480954 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 481574 374294
rect 480954 338614 481574 374058
rect 480954 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 481574 338614
rect 480954 338294 481574 338378
rect 480954 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 481574 338294
rect 480954 302614 481574 338058
rect 480954 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 481574 302614
rect 480954 302294 481574 302378
rect 480954 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 481574 302294
rect 480954 266614 481574 302058
rect 480954 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 481574 266614
rect 480954 266294 481574 266378
rect 480954 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 481574 266294
rect 480954 230614 481574 266058
rect 480954 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 481574 230614
rect 480954 230294 481574 230378
rect 480954 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 481574 230294
rect 480954 194614 481574 230058
rect 480954 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 481574 194614
rect 480954 194294 481574 194378
rect 480954 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 481574 194294
rect 480954 158614 481574 194058
rect 480954 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 481574 158614
rect 480954 158294 481574 158378
rect 480954 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 481574 158294
rect 480954 122614 481574 158058
rect 480954 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 481574 122614
rect 480954 122294 481574 122378
rect 480954 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 481574 122294
rect 480954 86614 481574 122058
rect 480954 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 481574 86614
rect 480954 86294 481574 86378
rect 480954 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 481574 86294
rect 480954 50614 481574 86058
rect 480954 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 481574 50614
rect 480954 50294 481574 50378
rect 480954 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 481574 50294
rect 480954 14614 481574 50058
rect 480954 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 481574 14614
rect 480954 14294 481574 14378
rect 480954 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 481574 14294
rect 462954 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 463574 -7066
rect 462954 -7386 463574 -7302
rect 462954 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 463574 -7386
rect 462954 -7654 463574 -7622
rect 480954 -6106 481574 14058
rect 487794 705798 488414 705830
rect 487794 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 488414 705798
rect 487794 705478 488414 705562
rect 487794 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 488414 705478
rect 487794 669454 488414 705242
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597454 488414 632898
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 561454 488414 596898
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 453454 488414 488898
rect 487794 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 488414 453454
rect 487794 453134 488414 453218
rect 487794 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 488414 453134
rect 487794 417454 488414 452898
rect 487794 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 488414 417454
rect 487794 417134 488414 417218
rect 487794 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 488414 417134
rect 487794 381454 488414 416898
rect 487794 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 488414 381454
rect 487794 381134 488414 381218
rect 487794 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 488414 381134
rect 487794 345454 488414 380898
rect 487794 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 488414 345454
rect 487794 345134 488414 345218
rect 487794 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 488414 345134
rect 487794 309454 488414 344898
rect 487794 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 488414 309454
rect 487794 309134 488414 309218
rect 487794 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 488414 309134
rect 487794 273454 488414 308898
rect 487794 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 488414 273454
rect 487794 273134 488414 273218
rect 487794 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 488414 273134
rect 487794 237454 488414 272898
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 487794 201454 488414 236898
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 165454 488414 200898
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 129454 488414 164898
rect 487794 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 488414 129454
rect 487794 129134 488414 129218
rect 487794 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 488414 129134
rect 487794 93454 488414 128898
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -1306 488414 20898
rect 487794 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 488414 -1306
rect 487794 -1626 488414 -1542
rect 487794 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 488414 -1626
rect 487794 -1894 488414 -1862
rect 491514 673174 492134 707162
rect 491514 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 492134 673174
rect 491514 672854 492134 672938
rect 491514 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 492134 672854
rect 491514 637174 492134 672618
rect 491514 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 492134 637174
rect 491514 636854 492134 636938
rect 491514 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 492134 636854
rect 491514 601174 492134 636618
rect 491514 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 492134 601174
rect 491514 600854 492134 600938
rect 491514 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 492134 600854
rect 491514 565174 492134 600618
rect 491514 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 492134 565174
rect 491514 564854 492134 564938
rect 491514 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 492134 564854
rect 491514 529174 492134 564618
rect 491514 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 492134 529174
rect 491514 528854 492134 528938
rect 491514 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 492134 528854
rect 491514 493174 492134 528618
rect 491514 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 492134 493174
rect 491514 492854 492134 492938
rect 491514 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 492134 492854
rect 491514 457174 492134 492618
rect 491514 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 492134 457174
rect 491514 456854 492134 456938
rect 491514 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 492134 456854
rect 491514 421174 492134 456618
rect 491514 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 492134 421174
rect 491514 420854 492134 420938
rect 491514 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 492134 420854
rect 491514 385174 492134 420618
rect 491514 384938 491546 385174
rect 491782 384938 491866 385174
rect 492102 384938 492134 385174
rect 491514 384854 492134 384938
rect 491514 384618 491546 384854
rect 491782 384618 491866 384854
rect 492102 384618 492134 384854
rect 491514 349174 492134 384618
rect 491514 348938 491546 349174
rect 491782 348938 491866 349174
rect 492102 348938 492134 349174
rect 491514 348854 492134 348938
rect 491514 348618 491546 348854
rect 491782 348618 491866 348854
rect 492102 348618 492134 348854
rect 491514 313174 492134 348618
rect 491514 312938 491546 313174
rect 491782 312938 491866 313174
rect 492102 312938 492134 313174
rect 491514 312854 492134 312938
rect 491514 312618 491546 312854
rect 491782 312618 491866 312854
rect 492102 312618 492134 312854
rect 491514 277174 492134 312618
rect 491514 276938 491546 277174
rect 491782 276938 491866 277174
rect 492102 276938 492134 277174
rect 491514 276854 492134 276938
rect 491514 276618 491546 276854
rect 491782 276618 491866 276854
rect 492102 276618 492134 276854
rect 491514 241174 492134 276618
rect 491514 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 492134 241174
rect 491514 240854 492134 240938
rect 491514 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 492134 240854
rect 491514 205174 492134 240618
rect 491514 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 492134 205174
rect 491514 204854 492134 204938
rect 491514 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 492134 204854
rect 491514 169174 492134 204618
rect 491514 168938 491546 169174
rect 491782 168938 491866 169174
rect 492102 168938 492134 169174
rect 491514 168854 492134 168938
rect 491514 168618 491546 168854
rect 491782 168618 491866 168854
rect 492102 168618 492134 168854
rect 491514 133174 492134 168618
rect 491514 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 492134 133174
rect 491514 132854 492134 132938
rect 491514 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 492134 132854
rect 491514 97174 492134 132618
rect 491514 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 492134 97174
rect 491514 96854 492134 96938
rect 491514 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 492134 96854
rect 491514 61174 492134 96618
rect 491514 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 492134 61174
rect 491514 60854 492134 60938
rect 491514 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 492134 60854
rect 491514 25174 492134 60618
rect 491514 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 492134 25174
rect 491514 24854 492134 24938
rect 491514 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 492134 24854
rect 491514 -3226 492134 24618
rect 491514 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 492134 -3226
rect 491514 -3546 492134 -3462
rect 491514 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 492134 -3546
rect 491514 -3814 492134 -3782
rect 495234 676894 495854 709082
rect 495234 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 495854 676894
rect 495234 676574 495854 676658
rect 495234 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 495854 676574
rect 495234 640894 495854 676338
rect 495234 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 495854 640894
rect 495234 640574 495854 640658
rect 495234 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 495854 640574
rect 495234 604894 495854 640338
rect 495234 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 495854 604894
rect 495234 604574 495854 604658
rect 495234 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 495854 604574
rect 495234 568894 495854 604338
rect 495234 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 495854 568894
rect 495234 568574 495854 568658
rect 495234 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 495854 568574
rect 495234 532894 495854 568338
rect 495234 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 495854 532894
rect 495234 532574 495854 532658
rect 495234 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 495854 532574
rect 495234 496894 495854 532338
rect 495234 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 495854 496894
rect 495234 496574 495854 496658
rect 495234 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 495854 496574
rect 495234 460894 495854 496338
rect 495234 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 495854 460894
rect 495234 460574 495854 460658
rect 495234 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 495854 460574
rect 495234 424894 495854 460338
rect 495234 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 495854 424894
rect 495234 424574 495854 424658
rect 495234 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 495854 424574
rect 495234 388894 495854 424338
rect 495234 388658 495266 388894
rect 495502 388658 495586 388894
rect 495822 388658 495854 388894
rect 495234 388574 495854 388658
rect 495234 388338 495266 388574
rect 495502 388338 495586 388574
rect 495822 388338 495854 388574
rect 495234 352894 495854 388338
rect 495234 352658 495266 352894
rect 495502 352658 495586 352894
rect 495822 352658 495854 352894
rect 495234 352574 495854 352658
rect 495234 352338 495266 352574
rect 495502 352338 495586 352574
rect 495822 352338 495854 352574
rect 495234 316894 495854 352338
rect 495234 316658 495266 316894
rect 495502 316658 495586 316894
rect 495822 316658 495854 316894
rect 495234 316574 495854 316658
rect 495234 316338 495266 316574
rect 495502 316338 495586 316574
rect 495822 316338 495854 316574
rect 495234 280894 495854 316338
rect 495234 280658 495266 280894
rect 495502 280658 495586 280894
rect 495822 280658 495854 280894
rect 495234 280574 495854 280658
rect 495234 280338 495266 280574
rect 495502 280338 495586 280574
rect 495822 280338 495854 280574
rect 495234 244894 495854 280338
rect 495234 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 495854 244894
rect 495234 244574 495854 244658
rect 495234 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 495854 244574
rect 495234 208894 495854 244338
rect 495234 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 495854 208894
rect 495234 208574 495854 208658
rect 495234 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 495854 208574
rect 495234 172894 495854 208338
rect 495234 172658 495266 172894
rect 495502 172658 495586 172894
rect 495822 172658 495854 172894
rect 495234 172574 495854 172658
rect 495234 172338 495266 172574
rect 495502 172338 495586 172574
rect 495822 172338 495854 172574
rect 495234 136894 495854 172338
rect 495234 136658 495266 136894
rect 495502 136658 495586 136894
rect 495822 136658 495854 136894
rect 495234 136574 495854 136658
rect 495234 136338 495266 136574
rect 495502 136338 495586 136574
rect 495822 136338 495854 136574
rect 495234 100894 495854 136338
rect 495234 100658 495266 100894
rect 495502 100658 495586 100894
rect 495822 100658 495854 100894
rect 495234 100574 495854 100658
rect 495234 100338 495266 100574
rect 495502 100338 495586 100574
rect 495822 100338 495854 100574
rect 495234 64894 495854 100338
rect 495234 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 495854 64894
rect 495234 64574 495854 64658
rect 495234 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 495854 64574
rect 495234 28894 495854 64338
rect 495234 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 495854 28894
rect 495234 28574 495854 28658
rect 495234 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 495854 28574
rect 495234 -5146 495854 28338
rect 495234 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 495854 -5146
rect 495234 -5466 495854 -5382
rect 495234 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 495854 -5466
rect 495234 -5734 495854 -5702
rect 498954 680614 499574 711002
rect 516954 710598 517574 711590
rect 516954 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 517574 710598
rect 516954 710278 517574 710362
rect 516954 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 517574 710278
rect 513234 708678 513854 709670
rect 513234 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 513854 708678
rect 513234 708358 513854 708442
rect 513234 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 513854 708358
rect 509514 706758 510134 707750
rect 509514 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 510134 706758
rect 509514 706438 510134 706522
rect 509514 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 510134 706438
rect 498954 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 499574 680614
rect 498954 680294 499574 680378
rect 498954 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 499574 680294
rect 498954 644614 499574 680058
rect 498954 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 499574 644614
rect 498954 644294 499574 644378
rect 498954 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 499574 644294
rect 498954 608614 499574 644058
rect 498954 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 499574 608614
rect 498954 608294 499574 608378
rect 498954 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 499574 608294
rect 498954 572614 499574 608058
rect 498954 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 499574 572614
rect 498954 572294 499574 572378
rect 498954 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 499574 572294
rect 498954 536614 499574 572058
rect 498954 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 499574 536614
rect 498954 536294 499574 536378
rect 498954 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 499574 536294
rect 498954 500614 499574 536058
rect 498954 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 499574 500614
rect 498954 500294 499574 500378
rect 498954 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 499574 500294
rect 498954 464614 499574 500058
rect 498954 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 499574 464614
rect 498954 464294 499574 464378
rect 498954 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 499574 464294
rect 498954 428614 499574 464058
rect 498954 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 499574 428614
rect 498954 428294 499574 428378
rect 498954 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 499574 428294
rect 498954 392614 499574 428058
rect 498954 392378 498986 392614
rect 499222 392378 499306 392614
rect 499542 392378 499574 392614
rect 498954 392294 499574 392378
rect 498954 392058 498986 392294
rect 499222 392058 499306 392294
rect 499542 392058 499574 392294
rect 498954 356614 499574 392058
rect 498954 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 499574 356614
rect 498954 356294 499574 356378
rect 498954 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 499574 356294
rect 498954 320614 499574 356058
rect 498954 320378 498986 320614
rect 499222 320378 499306 320614
rect 499542 320378 499574 320614
rect 498954 320294 499574 320378
rect 498954 320058 498986 320294
rect 499222 320058 499306 320294
rect 499542 320058 499574 320294
rect 498954 284614 499574 320058
rect 498954 284378 498986 284614
rect 499222 284378 499306 284614
rect 499542 284378 499574 284614
rect 498954 284294 499574 284378
rect 498954 284058 498986 284294
rect 499222 284058 499306 284294
rect 499542 284058 499574 284294
rect 498954 248614 499574 284058
rect 498954 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 499574 248614
rect 498954 248294 499574 248378
rect 498954 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 499574 248294
rect 498954 212614 499574 248058
rect 498954 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 499574 212614
rect 498954 212294 499574 212378
rect 498954 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 499574 212294
rect 498954 176614 499574 212058
rect 498954 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 499574 176614
rect 498954 176294 499574 176378
rect 498954 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 499574 176294
rect 498954 140614 499574 176058
rect 498954 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 499574 140614
rect 498954 140294 499574 140378
rect 498954 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 499574 140294
rect 498954 104614 499574 140058
rect 498954 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 499574 104614
rect 498954 104294 499574 104378
rect 498954 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 499574 104294
rect 498954 68614 499574 104058
rect 498954 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 499574 68614
rect 498954 68294 499574 68378
rect 498954 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 499574 68294
rect 498954 32614 499574 68058
rect 498954 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 499574 32614
rect 498954 32294 499574 32378
rect 498954 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 499574 32294
rect 480954 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 481574 -6106
rect 480954 -6426 481574 -6342
rect 480954 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 481574 -6426
rect 480954 -7654 481574 -6662
rect 498954 -7066 499574 32058
rect 505794 704838 506414 705830
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -1894 506414 -902
rect 509514 691174 510134 706202
rect 509514 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 510134 691174
rect 509514 690854 510134 690938
rect 509514 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 510134 690854
rect 509514 655174 510134 690618
rect 509514 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 510134 655174
rect 509514 654854 510134 654938
rect 509514 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 510134 654854
rect 509514 619174 510134 654618
rect 509514 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 510134 619174
rect 509514 618854 510134 618938
rect 509514 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 510134 618854
rect 509514 583174 510134 618618
rect 509514 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 510134 583174
rect 509514 582854 510134 582938
rect 509514 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 510134 582854
rect 509514 547174 510134 582618
rect 509514 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 510134 547174
rect 509514 546854 510134 546938
rect 509514 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 510134 546854
rect 509514 511174 510134 546618
rect 509514 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 510134 511174
rect 509514 510854 510134 510938
rect 509514 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 510134 510854
rect 509514 475174 510134 510618
rect 509514 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 510134 475174
rect 509514 474854 510134 474938
rect 509514 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 510134 474854
rect 509514 439174 510134 474618
rect 509514 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 510134 439174
rect 509514 438854 510134 438938
rect 509514 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 510134 438854
rect 509514 403174 510134 438618
rect 509514 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 510134 403174
rect 509514 402854 510134 402938
rect 509514 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 510134 402854
rect 509514 367174 510134 402618
rect 509514 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 510134 367174
rect 509514 366854 510134 366938
rect 509514 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 510134 366854
rect 509514 331174 510134 366618
rect 509514 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 510134 331174
rect 509514 330854 510134 330938
rect 509514 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 510134 330854
rect 509514 295174 510134 330618
rect 509514 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 510134 295174
rect 509514 294854 510134 294938
rect 509514 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 510134 294854
rect 509514 259174 510134 294618
rect 509514 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 510134 259174
rect 509514 258854 510134 258938
rect 509514 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 510134 258854
rect 509514 223174 510134 258618
rect 509514 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 510134 223174
rect 509514 222854 510134 222938
rect 509514 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 510134 222854
rect 509514 187174 510134 222618
rect 509514 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 510134 187174
rect 509514 186854 510134 186938
rect 509514 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 510134 186854
rect 509514 151174 510134 186618
rect 509514 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 510134 151174
rect 509514 150854 510134 150938
rect 509514 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 510134 150854
rect 509514 115174 510134 150618
rect 509514 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 510134 115174
rect 509514 114854 510134 114938
rect 509514 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 510134 114854
rect 509514 79174 510134 114618
rect 509514 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 510134 79174
rect 509514 78854 510134 78938
rect 509514 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 510134 78854
rect 509514 43174 510134 78618
rect 509514 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 510134 43174
rect 509514 42854 510134 42938
rect 509514 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 510134 42854
rect 509514 7174 510134 42618
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -2266 510134 6618
rect 509514 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 510134 -2266
rect 509514 -2586 510134 -2502
rect 509514 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 510134 -2586
rect 509514 -3814 510134 -2822
rect 513234 694894 513854 708122
rect 513234 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 513854 694894
rect 513234 694574 513854 694658
rect 513234 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 513854 694574
rect 513234 658894 513854 694338
rect 513234 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 513854 658894
rect 513234 658574 513854 658658
rect 513234 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 513854 658574
rect 513234 622894 513854 658338
rect 513234 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 513854 622894
rect 513234 622574 513854 622658
rect 513234 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 513854 622574
rect 513234 586894 513854 622338
rect 513234 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 513854 586894
rect 513234 586574 513854 586658
rect 513234 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 513854 586574
rect 513234 550894 513854 586338
rect 513234 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 513854 550894
rect 513234 550574 513854 550658
rect 513234 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 513854 550574
rect 513234 514894 513854 550338
rect 513234 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 513854 514894
rect 513234 514574 513854 514658
rect 513234 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 513854 514574
rect 513234 478894 513854 514338
rect 513234 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 513854 478894
rect 513234 478574 513854 478658
rect 513234 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 513854 478574
rect 513234 442894 513854 478338
rect 513234 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 513854 442894
rect 513234 442574 513854 442658
rect 513234 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 513854 442574
rect 513234 406894 513854 442338
rect 513234 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 513854 406894
rect 513234 406574 513854 406658
rect 513234 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 513854 406574
rect 513234 370894 513854 406338
rect 513234 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 513854 370894
rect 513234 370574 513854 370658
rect 513234 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 513854 370574
rect 513234 334894 513854 370338
rect 513234 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 513854 334894
rect 513234 334574 513854 334658
rect 513234 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 513854 334574
rect 513234 298894 513854 334338
rect 513234 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 513854 298894
rect 513234 298574 513854 298658
rect 513234 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 513854 298574
rect 513234 262894 513854 298338
rect 513234 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 513854 262894
rect 513234 262574 513854 262658
rect 513234 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 513854 262574
rect 513234 226894 513854 262338
rect 513234 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 513854 226894
rect 513234 226574 513854 226658
rect 513234 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 513854 226574
rect 513234 190894 513854 226338
rect 513234 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 513854 190894
rect 513234 190574 513854 190658
rect 513234 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 513854 190574
rect 513234 154894 513854 190338
rect 513234 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 513854 154894
rect 513234 154574 513854 154658
rect 513234 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 513854 154574
rect 513234 118894 513854 154338
rect 513234 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 513854 118894
rect 513234 118574 513854 118658
rect 513234 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 513854 118574
rect 513234 82894 513854 118338
rect 513234 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 513854 82894
rect 513234 82574 513854 82658
rect 513234 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 513854 82574
rect 513234 46894 513854 82338
rect 513234 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 513854 46894
rect 513234 46574 513854 46658
rect 513234 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 513854 46574
rect 513234 10894 513854 46338
rect 513234 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 513854 10894
rect 513234 10574 513854 10658
rect 513234 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 513854 10574
rect 513234 -4186 513854 10338
rect 513234 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 513854 -4186
rect 513234 -4506 513854 -4422
rect 513234 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 513854 -4506
rect 513234 -5734 513854 -4742
rect 516954 698614 517574 710042
rect 534954 711558 535574 711590
rect 534954 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 535574 711558
rect 534954 711238 535574 711322
rect 534954 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 535574 711238
rect 531234 709638 531854 709670
rect 531234 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 531854 709638
rect 531234 709318 531854 709402
rect 531234 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 531854 709318
rect 527514 707718 528134 707750
rect 527514 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 528134 707718
rect 527514 707398 528134 707482
rect 527514 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 528134 707398
rect 516954 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 517574 698614
rect 516954 698294 517574 698378
rect 516954 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 517574 698294
rect 516954 662614 517574 698058
rect 516954 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 517574 662614
rect 516954 662294 517574 662378
rect 516954 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 517574 662294
rect 516954 626614 517574 662058
rect 516954 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 517574 626614
rect 516954 626294 517574 626378
rect 516954 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 517574 626294
rect 516954 590614 517574 626058
rect 516954 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 517574 590614
rect 516954 590294 517574 590378
rect 516954 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 517574 590294
rect 516954 554614 517574 590058
rect 516954 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 517574 554614
rect 516954 554294 517574 554378
rect 516954 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 517574 554294
rect 516954 518614 517574 554058
rect 516954 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 517574 518614
rect 516954 518294 517574 518378
rect 516954 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 517574 518294
rect 516954 482614 517574 518058
rect 516954 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 517574 482614
rect 516954 482294 517574 482378
rect 516954 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 517574 482294
rect 516954 446614 517574 482058
rect 516954 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 517574 446614
rect 516954 446294 517574 446378
rect 516954 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 517574 446294
rect 516954 410614 517574 446058
rect 516954 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 517574 410614
rect 516954 410294 517574 410378
rect 516954 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 517574 410294
rect 516954 374614 517574 410058
rect 516954 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 517574 374614
rect 516954 374294 517574 374378
rect 516954 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 517574 374294
rect 516954 338614 517574 374058
rect 516954 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 517574 338614
rect 516954 338294 517574 338378
rect 516954 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 517574 338294
rect 516954 302614 517574 338058
rect 516954 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 517574 302614
rect 516954 302294 517574 302378
rect 516954 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 517574 302294
rect 516954 266614 517574 302058
rect 516954 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 517574 266614
rect 516954 266294 517574 266378
rect 516954 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 517574 266294
rect 516954 230614 517574 266058
rect 516954 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 517574 230614
rect 516954 230294 517574 230378
rect 516954 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 517574 230294
rect 516954 194614 517574 230058
rect 516954 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 517574 194614
rect 516954 194294 517574 194378
rect 516954 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 517574 194294
rect 516954 158614 517574 194058
rect 516954 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 517574 158614
rect 516954 158294 517574 158378
rect 516954 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 517574 158294
rect 516954 122614 517574 158058
rect 516954 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 517574 122614
rect 516954 122294 517574 122378
rect 516954 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 517574 122294
rect 516954 86614 517574 122058
rect 516954 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 517574 86614
rect 516954 86294 517574 86378
rect 516954 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 517574 86294
rect 516954 50614 517574 86058
rect 516954 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 517574 50614
rect 516954 50294 517574 50378
rect 516954 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 517574 50294
rect 516954 14614 517574 50058
rect 516954 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 517574 14614
rect 516954 14294 517574 14378
rect 516954 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 517574 14294
rect 498954 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 499574 -7066
rect 498954 -7386 499574 -7302
rect 498954 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 499574 -7386
rect 498954 -7654 499574 -7622
rect 516954 -6106 517574 14058
rect 523794 705798 524414 705830
rect 523794 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 524414 705798
rect 523794 705478 524414 705562
rect 523794 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 524414 705478
rect 523794 669454 524414 705242
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -1306 524414 20898
rect 523794 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 524414 -1306
rect 523794 -1626 524414 -1542
rect 523794 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 524414 -1626
rect 523794 -1894 524414 -1862
rect 527514 673174 528134 707162
rect 527514 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 528134 673174
rect 527514 672854 528134 672938
rect 527514 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 528134 672854
rect 527514 637174 528134 672618
rect 527514 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 528134 637174
rect 527514 636854 528134 636938
rect 527514 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 528134 636854
rect 527514 601174 528134 636618
rect 527514 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 528134 601174
rect 527514 600854 528134 600938
rect 527514 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 528134 600854
rect 527514 565174 528134 600618
rect 527514 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 528134 565174
rect 527514 564854 528134 564938
rect 527514 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 528134 564854
rect 527514 529174 528134 564618
rect 527514 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 528134 529174
rect 527514 528854 528134 528938
rect 527514 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 528134 528854
rect 527514 493174 528134 528618
rect 527514 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 528134 493174
rect 527514 492854 528134 492938
rect 527514 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 528134 492854
rect 527514 457174 528134 492618
rect 527514 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 528134 457174
rect 527514 456854 528134 456938
rect 527514 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 528134 456854
rect 527514 421174 528134 456618
rect 527514 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 528134 421174
rect 527514 420854 528134 420938
rect 527514 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 528134 420854
rect 527514 385174 528134 420618
rect 527514 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 528134 385174
rect 527514 384854 528134 384938
rect 527514 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 528134 384854
rect 527514 349174 528134 384618
rect 527514 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 528134 349174
rect 527514 348854 528134 348938
rect 527514 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 528134 348854
rect 527514 313174 528134 348618
rect 527514 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 528134 313174
rect 527514 312854 528134 312938
rect 527514 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 528134 312854
rect 527514 277174 528134 312618
rect 527514 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 528134 277174
rect 527514 276854 528134 276938
rect 527514 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 528134 276854
rect 527514 241174 528134 276618
rect 527514 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 528134 241174
rect 527514 240854 528134 240938
rect 527514 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 528134 240854
rect 527514 205174 528134 240618
rect 527514 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 528134 205174
rect 527514 204854 528134 204938
rect 527514 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 528134 204854
rect 527514 169174 528134 204618
rect 527514 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 528134 169174
rect 527514 168854 528134 168938
rect 527514 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 528134 168854
rect 527514 133174 528134 168618
rect 527514 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 528134 133174
rect 527514 132854 528134 132938
rect 527514 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 528134 132854
rect 527514 97174 528134 132618
rect 527514 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 528134 97174
rect 527514 96854 528134 96938
rect 527514 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 528134 96854
rect 527514 61174 528134 96618
rect 527514 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 528134 61174
rect 527514 60854 528134 60938
rect 527514 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 528134 60854
rect 527514 25174 528134 60618
rect 527514 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 528134 25174
rect 527514 24854 528134 24938
rect 527514 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 528134 24854
rect 527514 -3226 528134 24618
rect 527514 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 528134 -3226
rect 527514 -3546 528134 -3462
rect 527514 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 528134 -3546
rect 527514 -3814 528134 -3782
rect 531234 676894 531854 709082
rect 531234 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 531854 676894
rect 531234 676574 531854 676658
rect 531234 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 531854 676574
rect 531234 640894 531854 676338
rect 531234 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 531854 640894
rect 531234 640574 531854 640658
rect 531234 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 531854 640574
rect 531234 604894 531854 640338
rect 531234 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 531854 604894
rect 531234 604574 531854 604658
rect 531234 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 531854 604574
rect 531234 568894 531854 604338
rect 531234 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 531854 568894
rect 531234 568574 531854 568658
rect 531234 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 531854 568574
rect 531234 532894 531854 568338
rect 531234 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 531854 532894
rect 531234 532574 531854 532658
rect 531234 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 531854 532574
rect 531234 496894 531854 532338
rect 531234 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 531854 496894
rect 531234 496574 531854 496658
rect 531234 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 531854 496574
rect 531234 460894 531854 496338
rect 531234 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 531854 460894
rect 531234 460574 531854 460658
rect 531234 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 531854 460574
rect 531234 424894 531854 460338
rect 531234 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 531854 424894
rect 531234 424574 531854 424658
rect 531234 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 531854 424574
rect 531234 388894 531854 424338
rect 531234 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 531854 388894
rect 531234 388574 531854 388658
rect 531234 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 531854 388574
rect 531234 352894 531854 388338
rect 531234 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 531854 352894
rect 531234 352574 531854 352658
rect 531234 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 531854 352574
rect 531234 316894 531854 352338
rect 531234 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 531854 316894
rect 531234 316574 531854 316658
rect 531234 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 531854 316574
rect 531234 280894 531854 316338
rect 531234 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 531854 280894
rect 531234 280574 531854 280658
rect 531234 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 531854 280574
rect 531234 244894 531854 280338
rect 531234 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 531854 244894
rect 531234 244574 531854 244658
rect 531234 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 531854 244574
rect 531234 208894 531854 244338
rect 531234 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 531854 208894
rect 531234 208574 531854 208658
rect 531234 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 531854 208574
rect 531234 172894 531854 208338
rect 531234 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 531854 172894
rect 531234 172574 531854 172658
rect 531234 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 531854 172574
rect 531234 136894 531854 172338
rect 531234 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 531854 136894
rect 531234 136574 531854 136658
rect 531234 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 531854 136574
rect 531234 100894 531854 136338
rect 531234 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 531854 100894
rect 531234 100574 531854 100658
rect 531234 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 531854 100574
rect 531234 64894 531854 100338
rect 531234 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 531854 64894
rect 531234 64574 531854 64658
rect 531234 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 531854 64574
rect 531234 28894 531854 64338
rect 531234 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 531854 28894
rect 531234 28574 531854 28658
rect 531234 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 531854 28574
rect 531234 -5146 531854 28338
rect 531234 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 531854 -5146
rect 531234 -5466 531854 -5382
rect 531234 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 531854 -5466
rect 531234 -5734 531854 -5702
rect 534954 680614 535574 711002
rect 552954 710598 553574 711590
rect 552954 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 553574 710598
rect 552954 710278 553574 710362
rect 552954 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 553574 710278
rect 549234 708678 549854 709670
rect 549234 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 549854 708678
rect 549234 708358 549854 708442
rect 549234 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 549854 708358
rect 545514 706758 546134 707750
rect 545514 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 546134 706758
rect 545514 706438 546134 706522
rect 545514 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 546134 706438
rect 534954 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 535574 680614
rect 534954 680294 535574 680378
rect 534954 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 535574 680294
rect 534954 644614 535574 680058
rect 534954 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 535574 644614
rect 534954 644294 535574 644378
rect 534954 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 535574 644294
rect 534954 608614 535574 644058
rect 534954 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 535574 608614
rect 534954 608294 535574 608378
rect 534954 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 535574 608294
rect 534954 572614 535574 608058
rect 534954 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 535574 572614
rect 534954 572294 535574 572378
rect 534954 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 535574 572294
rect 534954 536614 535574 572058
rect 534954 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 535574 536614
rect 534954 536294 535574 536378
rect 534954 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 535574 536294
rect 534954 500614 535574 536058
rect 534954 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 535574 500614
rect 534954 500294 535574 500378
rect 534954 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 535574 500294
rect 534954 464614 535574 500058
rect 534954 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 535574 464614
rect 534954 464294 535574 464378
rect 534954 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 535574 464294
rect 534954 428614 535574 464058
rect 534954 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 535574 428614
rect 534954 428294 535574 428378
rect 534954 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 535574 428294
rect 534954 392614 535574 428058
rect 534954 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 535574 392614
rect 534954 392294 535574 392378
rect 534954 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 535574 392294
rect 534954 356614 535574 392058
rect 534954 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 535574 356614
rect 534954 356294 535574 356378
rect 534954 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 535574 356294
rect 534954 320614 535574 356058
rect 534954 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 535574 320614
rect 534954 320294 535574 320378
rect 534954 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 535574 320294
rect 534954 284614 535574 320058
rect 534954 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 535574 284614
rect 534954 284294 535574 284378
rect 534954 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 535574 284294
rect 534954 248614 535574 284058
rect 534954 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 535574 248614
rect 534954 248294 535574 248378
rect 534954 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 535574 248294
rect 534954 212614 535574 248058
rect 534954 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 535574 212614
rect 534954 212294 535574 212378
rect 534954 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 535574 212294
rect 534954 176614 535574 212058
rect 534954 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 535574 176614
rect 534954 176294 535574 176378
rect 534954 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 535574 176294
rect 534954 140614 535574 176058
rect 534954 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 535574 140614
rect 534954 140294 535574 140378
rect 534954 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 535574 140294
rect 534954 104614 535574 140058
rect 534954 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 535574 104614
rect 534954 104294 535574 104378
rect 534954 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 535574 104294
rect 534954 68614 535574 104058
rect 534954 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 535574 68614
rect 534954 68294 535574 68378
rect 534954 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 535574 68294
rect 534954 32614 535574 68058
rect 534954 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 535574 32614
rect 534954 32294 535574 32378
rect 534954 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 535574 32294
rect 516954 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 517574 -6106
rect 516954 -6426 517574 -6342
rect 516954 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 517574 -6426
rect 516954 -7654 517574 -6662
rect 534954 -7066 535574 32058
rect 541794 704838 542414 705830
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -1894 542414 -902
rect 545514 691174 546134 706202
rect 545514 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 546134 691174
rect 545514 690854 546134 690938
rect 545514 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 546134 690854
rect 545514 655174 546134 690618
rect 545514 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 546134 655174
rect 545514 654854 546134 654938
rect 545514 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 546134 654854
rect 545514 619174 546134 654618
rect 545514 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 546134 619174
rect 545514 618854 546134 618938
rect 545514 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 546134 618854
rect 545514 583174 546134 618618
rect 545514 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 546134 583174
rect 545514 582854 546134 582938
rect 545514 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 546134 582854
rect 545514 547174 546134 582618
rect 545514 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 546134 547174
rect 545514 546854 546134 546938
rect 545514 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 546134 546854
rect 545514 511174 546134 546618
rect 545514 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 546134 511174
rect 545514 510854 546134 510938
rect 545514 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 546134 510854
rect 545514 475174 546134 510618
rect 545514 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 546134 475174
rect 545514 474854 546134 474938
rect 545514 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 546134 474854
rect 545514 439174 546134 474618
rect 545514 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 546134 439174
rect 545514 438854 546134 438938
rect 545514 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 546134 438854
rect 545514 403174 546134 438618
rect 545514 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 546134 403174
rect 545514 402854 546134 402938
rect 545514 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 546134 402854
rect 545514 367174 546134 402618
rect 545514 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 546134 367174
rect 545514 366854 546134 366938
rect 545514 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 546134 366854
rect 545514 331174 546134 366618
rect 545514 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 546134 331174
rect 545514 330854 546134 330938
rect 545514 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 546134 330854
rect 545514 295174 546134 330618
rect 545514 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 546134 295174
rect 545514 294854 546134 294938
rect 545514 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 546134 294854
rect 545514 259174 546134 294618
rect 545514 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 546134 259174
rect 545514 258854 546134 258938
rect 545514 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 546134 258854
rect 545514 223174 546134 258618
rect 545514 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 546134 223174
rect 545514 222854 546134 222938
rect 545514 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 546134 222854
rect 545514 187174 546134 222618
rect 545514 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 546134 187174
rect 545514 186854 546134 186938
rect 545514 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 546134 186854
rect 545514 151174 546134 186618
rect 545514 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 546134 151174
rect 545514 150854 546134 150938
rect 545514 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 546134 150854
rect 545514 115174 546134 150618
rect 545514 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 546134 115174
rect 545514 114854 546134 114938
rect 545514 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 546134 114854
rect 545514 79174 546134 114618
rect 545514 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 546134 79174
rect 545514 78854 546134 78938
rect 545514 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 546134 78854
rect 545514 43174 546134 78618
rect 545514 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 546134 43174
rect 545514 42854 546134 42938
rect 545514 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 546134 42854
rect 545514 7174 546134 42618
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -2266 546134 6618
rect 545514 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 546134 -2266
rect 545514 -2586 546134 -2502
rect 545514 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 546134 -2586
rect 545514 -3814 546134 -2822
rect 549234 694894 549854 708122
rect 549234 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 549854 694894
rect 549234 694574 549854 694658
rect 549234 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 549854 694574
rect 549234 658894 549854 694338
rect 549234 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 549854 658894
rect 549234 658574 549854 658658
rect 549234 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 549854 658574
rect 549234 622894 549854 658338
rect 549234 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 549854 622894
rect 549234 622574 549854 622658
rect 549234 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 549854 622574
rect 549234 586894 549854 622338
rect 549234 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 549854 586894
rect 549234 586574 549854 586658
rect 549234 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 549854 586574
rect 549234 550894 549854 586338
rect 549234 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 549854 550894
rect 549234 550574 549854 550658
rect 549234 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 549854 550574
rect 549234 514894 549854 550338
rect 549234 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 549854 514894
rect 549234 514574 549854 514658
rect 549234 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 549854 514574
rect 549234 478894 549854 514338
rect 549234 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 549854 478894
rect 549234 478574 549854 478658
rect 549234 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 549854 478574
rect 549234 442894 549854 478338
rect 549234 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 549854 442894
rect 549234 442574 549854 442658
rect 549234 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 549854 442574
rect 549234 406894 549854 442338
rect 549234 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 549854 406894
rect 549234 406574 549854 406658
rect 549234 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 549854 406574
rect 549234 370894 549854 406338
rect 549234 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 549854 370894
rect 549234 370574 549854 370658
rect 549234 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 549854 370574
rect 549234 334894 549854 370338
rect 549234 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 549854 334894
rect 549234 334574 549854 334658
rect 549234 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 549854 334574
rect 549234 298894 549854 334338
rect 549234 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 549854 298894
rect 549234 298574 549854 298658
rect 549234 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 549854 298574
rect 549234 262894 549854 298338
rect 549234 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 549854 262894
rect 549234 262574 549854 262658
rect 549234 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 549854 262574
rect 549234 226894 549854 262338
rect 549234 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 549854 226894
rect 549234 226574 549854 226658
rect 549234 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 549854 226574
rect 549234 190894 549854 226338
rect 549234 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 549854 190894
rect 549234 190574 549854 190658
rect 549234 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 549854 190574
rect 549234 154894 549854 190338
rect 549234 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 549854 154894
rect 549234 154574 549854 154658
rect 549234 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 549854 154574
rect 549234 118894 549854 154338
rect 549234 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 549854 118894
rect 549234 118574 549854 118658
rect 549234 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 549854 118574
rect 549234 82894 549854 118338
rect 549234 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 549854 82894
rect 549234 82574 549854 82658
rect 549234 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 549854 82574
rect 549234 46894 549854 82338
rect 549234 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 549854 46894
rect 549234 46574 549854 46658
rect 549234 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 549854 46574
rect 549234 10894 549854 46338
rect 549234 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 549854 10894
rect 549234 10574 549854 10658
rect 549234 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 549854 10574
rect 549234 -4186 549854 10338
rect 549234 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 549854 -4186
rect 549234 -4506 549854 -4422
rect 549234 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 549854 -4506
rect 549234 -5734 549854 -4742
rect 552954 698614 553574 710042
rect 570954 711558 571574 711590
rect 570954 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 571574 711558
rect 570954 711238 571574 711322
rect 570954 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 571574 711238
rect 567234 709638 567854 709670
rect 567234 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 567854 709638
rect 567234 709318 567854 709402
rect 567234 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 567854 709318
rect 563514 707718 564134 707750
rect 563514 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 564134 707718
rect 563514 707398 564134 707482
rect 563514 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 564134 707398
rect 552954 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 553574 698614
rect 552954 698294 553574 698378
rect 552954 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 553574 698294
rect 552954 662614 553574 698058
rect 552954 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 553574 662614
rect 552954 662294 553574 662378
rect 552954 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 553574 662294
rect 552954 626614 553574 662058
rect 552954 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 553574 626614
rect 552954 626294 553574 626378
rect 552954 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 553574 626294
rect 552954 590614 553574 626058
rect 552954 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 553574 590614
rect 552954 590294 553574 590378
rect 552954 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 553574 590294
rect 552954 554614 553574 590058
rect 552954 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 553574 554614
rect 552954 554294 553574 554378
rect 552954 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 553574 554294
rect 552954 518614 553574 554058
rect 552954 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 553574 518614
rect 552954 518294 553574 518378
rect 552954 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 553574 518294
rect 552954 482614 553574 518058
rect 552954 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 553574 482614
rect 552954 482294 553574 482378
rect 552954 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 553574 482294
rect 552954 446614 553574 482058
rect 552954 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 553574 446614
rect 552954 446294 553574 446378
rect 552954 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 553574 446294
rect 552954 410614 553574 446058
rect 552954 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 553574 410614
rect 552954 410294 553574 410378
rect 552954 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 553574 410294
rect 552954 374614 553574 410058
rect 552954 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 553574 374614
rect 552954 374294 553574 374378
rect 552954 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 553574 374294
rect 552954 338614 553574 374058
rect 552954 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 553574 338614
rect 552954 338294 553574 338378
rect 552954 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 553574 338294
rect 552954 302614 553574 338058
rect 552954 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 553574 302614
rect 552954 302294 553574 302378
rect 552954 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 553574 302294
rect 552954 266614 553574 302058
rect 552954 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 553574 266614
rect 552954 266294 553574 266378
rect 552954 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 553574 266294
rect 552954 230614 553574 266058
rect 552954 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 553574 230614
rect 552954 230294 553574 230378
rect 552954 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 553574 230294
rect 552954 194614 553574 230058
rect 552954 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 553574 194614
rect 552954 194294 553574 194378
rect 552954 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 553574 194294
rect 552954 158614 553574 194058
rect 552954 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 553574 158614
rect 552954 158294 553574 158378
rect 552954 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 553574 158294
rect 552954 122614 553574 158058
rect 552954 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 553574 122614
rect 552954 122294 553574 122378
rect 552954 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 553574 122294
rect 552954 86614 553574 122058
rect 552954 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 553574 86614
rect 552954 86294 553574 86378
rect 552954 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 553574 86294
rect 552954 50614 553574 86058
rect 552954 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 553574 50614
rect 552954 50294 553574 50378
rect 552954 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 553574 50294
rect 552954 14614 553574 50058
rect 552954 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 553574 14614
rect 552954 14294 553574 14378
rect 552954 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 553574 14294
rect 534954 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 535574 -7066
rect 534954 -7386 535574 -7302
rect 534954 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 535574 -7386
rect 534954 -7654 535574 -7622
rect 552954 -6106 553574 14058
rect 559794 705798 560414 705830
rect 559794 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 560414 705798
rect 559794 705478 560414 705562
rect 559794 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 560414 705478
rect 559794 669454 560414 705242
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -1306 560414 20898
rect 559794 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 560414 -1306
rect 559794 -1626 560414 -1542
rect 559794 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 560414 -1626
rect 559794 -1894 560414 -1862
rect 563514 673174 564134 707162
rect 563514 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 564134 673174
rect 563514 672854 564134 672938
rect 563514 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 564134 672854
rect 563514 637174 564134 672618
rect 563514 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 564134 637174
rect 563514 636854 564134 636938
rect 563514 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 564134 636854
rect 563514 601174 564134 636618
rect 563514 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 564134 601174
rect 563514 600854 564134 600938
rect 563514 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 564134 600854
rect 563514 565174 564134 600618
rect 563514 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 564134 565174
rect 563514 564854 564134 564938
rect 563514 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 564134 564854
rect 563514 529174 564134 564618
rect 563514 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 564134 529174
rect 563514 528854 564134 528938
rect 563514 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 564134 528854
rect 563514 493174 564134 528618
rect 563514 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 564134 493174
rect 563514 492854 564134 492938
rect 563514 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 564134 492854
rect 563514 457174 564134 492618
rect 563514 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 564134 457174
rect 563514 456854 564134 456938
rect 563514 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 564134 456854
rect 563514 421174 564134 456618
rect 563514 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 564134 421174
rect 563514 420854 564134 420938
rect 563514 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 564134 420854
rect 563514 385174 564134 420618
rect 563514 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 564134 385174
rect 563514 384854 564134 384938
rect 563514 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 564134 384854
rect 563514 349174 564134 384618
rect 563514 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 564134 349174
rect 563514 348854 564134 348938
rect 563514 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 564134 348854
rect 563514 313174 564134 348618
rect 563514 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 564134 313174
rect 563514 312854 564134 312938
rect 563514 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 564134 312854
rect 563514 277174 564134 312618
rect 563514 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 564134 277174
rect 563514 276854 564134 276938
rect 563514 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 564134 276854
rect 563514 241174 564134 276618
rect 563514 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 564134 241174
rect 563514 240854 564134 240938
rect 563514 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 564134 240854
rect 563514 205174 564134 240618
rect 563514 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 564134 205174
rect 563514 204854 564134 204938
rect 563514 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 564134 204854
rect 563514 169174 564134 204618
rect 563514 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 564134 169174
rect 563514 168854 564134 168938
rect 563514 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 564134 168854
rect 563514 133174 564134 168618
rect 563514 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 564134 133174
rect 563514 132854 564134 132938
rect 563514 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 564134 132854
rect 563514 97174 564134 132618
rect 563514 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 564134 97174
rect 563514 96854 564134 96938
rect 563514 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 564134 96854
rect 563514 61174 564134 96618
rect 563514 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 564134 61174
rect 563514 60854 564134 60938
rect 563514 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 564134 60854
rect 563514 25174 564134 60618
rect 563514 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 564134 25174
rect 563514 24854 564134 24938
rect 563514 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 564134 24854
rect 563514 -3226 564134 24618
rect 563514 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 564134 -3226
rect 563514 -3546 564134 -3462
rect 563514 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 564134 -3546
rect 563514 -3814 564134 -3782
rect 567234 676894 567854 709082
rect 567234 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 567854 676894
rect 567234 676574 567854 676658
rect 567234 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 567854 676574
rect 567234 640894 567854 676338
rect 567234 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 567854 640894
rect 567234 640574 567854 640658
rect 567234 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 567854 640574
rect 567234 604894 567854 640338
rect 567234 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 567854 604894
rect 567234 604574 567854 604658
rect 567234 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 567854 604574
rect 567234 568894 567854 604338
rect 567234 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 567854 568894
rect 567234 568574 567854 568658
rect 567234 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 567854 568574
rect 567234 532894 567854 568338
rect 567234 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 567854 532894
rect 567234 532574 567854 532658
rect 567234 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 567854 532574
rect 567234 496894 567854 532338
rect 567234 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 567854 496894
rect 567234 496574 567854 496658
rect 567234 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 567854 496574
rect 567234 460894 567854 496338
rect 567234 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 567854 460894
rect 567234 460574 567854 460658
rect 567234 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 567854 460574
rect 567234 424894 567854 460338
rect 567234 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 567854 424894
rect 567234 424574 567854 424658
rect 567234 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 567854 424574
rect 567234 388894 567854 424338
rect 567234 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 567854 388894
rect 567234 388574 567854 388658
rect 567234 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 567854 388574
rect 567234 352894 567854 388338
rect 567234 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 567854 352894
rect 567234 352574 567854 352658
rect 567234 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 567854 352574
rect 567234 316894 567854 352338
rect 567234 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 567854 316894
rect 567234 316574 567854 316658
rect 567234 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 567854 316574
rect 567234 280894 567854 316338
rect 567234 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 567854 280894
rect 567234 280574 567854 280658
rect 567234 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 567854 280574
rect 567234 244894 567854 280338
rect 567234 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 567854 244894
rect 567234 244574 567854 244658
rect 567234 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 567854 244574
rect 567234 208894 567854 244338
rect 567234 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 567854 208894
rect 567234 208574 567854 208658
rect 567234 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 567854 208574
rect 567234 172894 567854 208338
rect 567234 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 567854 172894
rect 567234 172574 567854 172658
rect 567234 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 567854 172574
rect 567234 136894 567854 172338
rect 567234 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 567854 136894
rect 567234 136574 567854 136658
rect 567234 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 567854 136574
rect 567234 100894 567854 136338
rect 567234 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 567854 100894
rect 567234 100574 567854 100658
rect 567234 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 567854 100574
rect 567234 64894 567854 100338
rect 567234 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 567854 64894
rect 567234 64574 567854 64658
rect 567234 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 567854 64574
rect 567234 28894 567854 64338
rect 567234 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 567854 28894
rect 567234 28574 567854 28658
rect 567234 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 567854 28574
rect 567234 -5146 567854 28338
rect 567234 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 567854 -5146
rect 567234 -5466 567854 -5382
rect 567234 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 567854 -5466
rect 567234 -5734 567854 -5702
rect 570954 680614 571574 711002
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 581514 706758 582134 707750
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 581514 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 582134 706758
rect 581514 706438 582134 706522
rect 581514 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 582134 706438
rect 570954 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 571574 680614
rect 570954 680294 571574 680378
rect 570954 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 571574 680294
rect 570954 644614 571574 680058
rect 570954 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 571574 644614
rect 570954 644294 571574 644378
rect 570954 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 571574 644294
rect 570954 608614 571574 644058
rect 570954 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 571574 608614
rect 570954 608294 571574 608378
rect 570954 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 571574 608294
rect 570954 572614 571574 608058
rect 570954 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 571574 572614
rect 570954 572294 571574 572378
rect 570954 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 571574 572294
rect 570954 536614 571574 572058
rect 570954 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 571574 536614
rect 570954 536294 571574 536378
rect 570954 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 571574 536294
rect 570954 500614 571574 536058
rect 570954 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 571574 500614
rect 570954 500294 571574 500378
rect 570954 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 571574 500294
rect 570954 464614 571574 500058
rect 570954 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 571574 464614
rect 570954 464294 571574 464378
rect 570954 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 571574 464294
rect 570954 428614 571574 464058
rect 570954 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 571574 428614
rect 570954 428294 571574 428378
rect 570954 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 571574 428294
rect 570954 392614 571574 428058
rect 570954 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 571574 392614
rect 570954 392294 571574 392378
rect 570954 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 571574 392294
rect 570954 356614 571574 392058
rect 570954 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 571574 356614
rect 570954 356294 571574 356378
rect 570954 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 571574 356294
rect 570954 320614 571574 356058
rect 570954 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 571574 320614
rect 570954 320294 571574 320378
rect 570954 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 571574 320294
rect 570954 284614 571574 320058
rect 570954 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 571574 284614
rect 570954 284294 571574 284378
rect 570954 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 571574 284294
rect 570954 248614 571574 284058
rect 570954 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 571574 248614
rect 570954 248294 571574 248378
rect 570954 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 571574 248294
rect 570954 212614 571574 248058
rect 570954 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 571574 212614
rect 570954 212294 571574 212378
rect 570954 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 571574 212294
rect 570954 176614 571574 212058
rect 570954 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 571574 176614
rect 570954 176294 571574 176378
rect 570954 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 571574 176294
rect 570954 140614 571574 176058
rect 570954 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 571574 140614
rect 570954 140294 571574 140378
rect 570954 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 571574 140294
rect 570954 104614 571574 140058
rect 570954 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 571574 104614
rect 570954 104294 571574 104378
rect 570954 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 571574 104294
rect 570954 68614 571574 104058
rect 570954 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 571574 68614
rect 570954 68294 571574 68378
rect 570954 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 571574 68294
rect 570954 32614 571574 68058
rect 570954 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 571574 32614
rect 570954 32294 571574 32378
rect 570954 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 571574 32294
rect 552954 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 553574 -6106
rect 552954 -6426 553574 -6342
rect 552954 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 553574 -6426
rect 552954 -7654 553574 -6662
rect 570954 -7066 571574 32058
rect 577794 704838 578414 705830
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -1894 578414 -902
rect 581514 691174 582134 706202
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -2266 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 669454 586890 705242
rect 586270 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect 586270 669134 586890 669218
rect 586270 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect 586270 633454 586890 668898
rect 586270 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect 586270 633134 586890 633218
rect 586270 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect 586270 597454 586890 632898
rect 586270 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect 586270 597134 586890 597218
rect 586270 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect 586270 561454 586890 596898
rect 586270 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect 586270 561134 586890 561218
rect 586270 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect 586270 525454 586890 560898
rect 586270 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect 586270 525134 586890 525218
rect 586270 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect 586270 489454 586890 524898
rect 586270 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect 586270 489134 586890 489218
rect 586270 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect 586270 453454 586890 488898
rect 586270 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect 586270 453134 586890 453218
rect 586270 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect 586270 417454 586890 452898
rect 586270 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect 586270 417134 586890 417218
rect 586270 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect 586270 381454 586890 416898
rect 586270 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect 586270 381134 586890 381218
rect 586270 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect 586270 345454 586890 380898
rect 586270 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect 586270 345134 586890 345218
rect 586270 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect 586270 309454 586890 344898
rect 586270 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect 586270 309134 586890 309218
rect 586270 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect 586270 273454 586890 308898
rect 586270 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect 586270 273134 586890 273218
rect 586270 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect 586270 237454 586890 272898
rect 586270 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect 586270 237134 586890 237218
rect 586270 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect 586270 201454 586890 236898
rect 586270 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect 586270 201134 586890 201218
rect 586270 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect 586270 165454 586890 200898
rect 586270 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect 586270 165134 586890 165218
rect 586270 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect 586270 129454 586890 164898
rect 586270 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect 586270 129134 586890 129218
rect 586270 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect 586270 93454 586890 128898
rect 586270 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect 586270 93134 586890 93218
rect 586270 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect 586270 57454 586890 92898
rect 586270 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect 586270 57134 586890 57218
rect 586270 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect 586270 21454 586890 56898
rect 586270 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect 586270 21134 586890 21218
rect 586270 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect 586270 -1306 586890 20898
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 691174 587850 706202
rect 587230 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 587850 691174
rect 587230 690854 587850 690938
rect 587230 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 587850 690854
rect 587230 655174 587850 690618
rect 587230 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 587850 655174
rect 587230 654854 587850 654938
rect 587230 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 587850 654854
rect 587230 619174 587850 654618
rect 587230 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 587850 619174
rect 587230 618854 587850 618938
rect 587230 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 587850 618854
rect 587230 583174 587850 618618
rect 587230 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 587850 583174
rect 587230 582854 587850 582938
rect 587230 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 587850 582854
rect 587230 547174 587850 582618
rect 587230 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 587850 547174
rect 587230 546854 587850 546938
rect 587230 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 587850 546854
rect 587230 511174 587850 546618
rect 587230 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 587850 511174
rect 587230 510854 587850 510938
rect 587230 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 587850 510854
rect 587230 475174 587850 510618
rect 587230 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 587850 475174
rect 587230 474854 587850 474938
rect 587230 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 587850 474854
rect 587230 439174 587850 474618
rect 587230 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 587850 439174
rect 587230 438854 587850 438938
rect 587230 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 587850 438854
rect 587230 403174 587850 438618
rect 587230 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 587850 403174
rect 587230 402854 587850 402938
rect 587230 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 587850 402854
rect 587230 367174 587850 402618
rect 587230 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 587850 367174
rect 587230 366854 587850 366938
rect 587230 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 587850 366854
rect 587230 331174 587850 366618
rect 587230 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 587850 331174
rect 587230 330854 587850 330938
rect 587230 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 587850 330854
rect 587230 295174 587850 330618
rect 587230 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 587850 295174
rect 587230 294854 587850 294938
rect 587230 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 587850 294854
rect 587230 259174 587850 294618
rect 587230 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 587850 259174
rect 587230 258854 587850 258938
rect 587230 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 587850 258854
rect 587230 223174 587850 258618
rect 587230 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 587850 223174
rect 587230 222854 587850 222938
rect 587230 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 587850 222854
rect 587230 187174 587850 222618
rect 587230 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 587850 187174
rect 587230 186854 587850 186938
rect 587230 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 587850 186854
rect 587230 151174 587850 186618
rect 587230 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 587850 151174
rect 587230 150854 587850 150938
rect 587230 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 587850 150854
rect 587230 115174 587850 150618
rect 587230 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 587850 115174
rect 587230 114854 587850 114938
rect 587230 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 587850 114854
rect 587230 79174 587850 114618
rect 587230 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 587850 79174
rect 587230 78854 587850 78938
rect 587230 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 587850 78854
rect 587230 43174 587850 78618
rect 587230 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 587850 43174
rect 587230 42854 587850 42938
rect 587230 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 587850 42854
rect 587230 7174 587850 42618
rect 587230 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 587850 7174
rect 587230 6854 587850 6938
rect 587230 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 587850 6854
rect 581514 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 582134 -2266
rect 581514 -2586 582134 -2502
rect 581514 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 582134 -2586
rect 581514 -3814 582134 -2822
rect 587230 -2266 587850 6618
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 673174 588810 707162
rect 588190 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect 588190 672854 588810 672938
rect 588190 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect 588190 637174 588810 672618
rect 588190 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect 588190 636854 588810 636938
rect 588190 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect 588190 601174 588810 636618
rect 588190 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect 588190 600854 588810 600938
rect 588190 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect 588190 565174 588810 600618
rect 588190 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect 588190 564854 588810 564938
rect 588190 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect 588190 529174 588810 564618
rect 588190 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect 588190 528854 588810 528938
rect 588190 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect 588190 493174 588810 528618
rect 588190 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect 588190 492854 588810 492938
rect 588190 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect 588190 457174 588810 492618
rect 588190 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect 588190 456854 588810 456938
rect 588190 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect 588190 421174 588810 456618
rect 588190 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect 588190 420854 588810 420938
rect 588190 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect 588190 385174 588810 420618
rect 588190 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect 588190 384854 588810 384938
rect 588190 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect 588190 349174 588810 384618
rect 588190 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect 588190 348854 588810 348938
rect 588190 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect 588190 313174 588810 348618
rect 588190 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect 588190 312854 588810 312938
rect 588190 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect 588190 277174 588810 312618
rect 588190 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect 588190 276854 588810 276938
rect 588190 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect 588190 241174 588810 276618
rect 588190 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect 588190 240854 588810 240938
rect 588190 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect 588190 205174 588810 240618
rect 588190 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect 588190 204854 588810 204938
rect 588190 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect 588190 169174 588810 204618
rect 588190 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect 588190 168854 588810 168938
rect 588190 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect 588190 133174 588810 168618
rect 588190 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect 588190 132854 588810 132938
rect 588190 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect 588190 97174 588810 132618
rect 588190 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect 588190 96854 588810 96938
rect 588190 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect 588190 61174 588810 96618
rect 588190 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect 588190 60854 588810 60938
rect 588190 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect 588190 25174 588810 60618
rect 588190 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect 588190 24854 588810 24938
rect 588190 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect 588190 -3226 588810 24618
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 694894 589770 708122
rect 589150 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 589770 694894
rect 589150 694574 589770 694658
rect 589150 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 589770 694574
rect 589150 658894 589770 694338
rect 589150 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 589770 658894
rect 589150 658574 589770 658658
rect 589150 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 589770 658574
rect 589150 622894 589770 658338
rect 589150 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 589770 622894
rect 589150 622574 589770 622658
rect 589150 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 589770 622574
rect 589150 586894 589770 622338
rect 589150 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 589770 586894
rect 589150 586574 589770 586658
rect 589150 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 589770 586574
rect 589150 550894 589770 586338
rect 589150 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 589770 550894
rect 589150 550574 589770 550658
rect 589150 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 589770 550574
rect 589150 514894 589770 550338
rect 589150 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 589770 514894
rect 589150 514574 589770 514658
rect 589150 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 589770 514574
rect 589150 478894 589770 514338
rect 589150 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 589770 478894
rect 589150 478574 589770 478658
rect 589150 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 589770 478574
rect 589150 442894 589770 478338
rect 589150 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 589770 442894
rect 589150 442574 589770 442658
rect 589150 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 589770 442574
rect 589150 406894 589770 442338
rect 589150 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 589770 406894
rect 589150 406574 589770 406658
rect 589150 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 589770 406574
rect 589150 370894 589770 406338
rect 589150 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 589770 370894
rect 589150 370574 589770 370658
rect 589150 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 589770 370574
rect 589150 334894 589770 370338
rect 589150 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 589770 334894
rect 589150 334574 589770 334658
rect 589150 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 589770 334574
rect 589150 298894 589770 334338
rect 589150 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 589770 298894
rect 589150 298574 589770 298658
rect 589150 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 589770 298574
rect 589150 262894 589770 298338
rect 589150 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 589770 262894
rect 589150 262574 589770 262658
rect 589150 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 589770 262574
rect 589150 226894 589770 262338
rect 589150 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 589770 226894
rect 589150 226574 589770 226658
rect 589150 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 589770 226574
rect 589150 190894 589770 226338
rect 589150 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 589770 190894
rect 589150 190574 589770 190658
rect 589150 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 589770 190574
rect 589150 154894 589770 190338
rect 589150 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 589770 154894
rect 589150 154574 589770 154658
rect 589150 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 589770 154574
rect 589150 118894 589770 154338
rect 589150 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 589770 118894
rect 589150 118574 589770 118658
rect 589150 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 589770 118574
rect 589150 82894 589770 118338
rect 589150 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 589770 82894
rect 589150 82574 589770 82658
rect 589150 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 589770 82574
rect 589150 46894 589770 82338
rect 589150 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 589770 46894
rect 589150 46574 589770 46658
rect 589150 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 589770 46574
rect 589150 10894 589770 46338
rect 589150 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 589770 10894
rect 589150 10574 589770 10658
rect 589150 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 589770 10574
rect 589150 -4186 589770 10338
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 676894 590730 709082
rect 590110 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect 590110 676574 590730 676658
rect 590110 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect 590110 640894 590730 676338
rect 590110 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect 590110 640574 590730 640658
rect 590110 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect 590110 604894 590730 640338
rect 590110 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect 590110 604574 590730 604658
rect 590110 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect 590110 568894 590730 604338
rect 590110 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect 590110 568574 590730 568658
rect 590110 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect 590110 532894 590730 568338
rect 590110 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect 590110 532574 590730 532658
rect 590110 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect 590110 496894 590730 532338
rect 590110 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect 590110 496574 590730 496658
rect 590110 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect 590110 460894 590730 496338
rect 590110 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect 590110 460574 590730 460658
rect 590110 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect 590110 424894 590730 460338
rect 590110 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect 590110 424574 590730 424658
rect 590110 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect 590110 388894 590730 424338
rect 590110 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect 590110 388574 590730 388658
rect 590110 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect 590110 352894 590730 388338
rect 590110 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect 590110 352574 590730 352658
rect 590110 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect 590110 316894 590730 352338
rect 590110 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect 590110 316574 590730 316658
rect 590110 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect 590110 280894 590730 316338
rect 590110 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect 590110 280574 590730 280658
rect 590110 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect 590110 244894 590730 280338
rect 590110 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect 590110 244574 590730 244658
rect 590110 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect 590110 208894 590730 244338
rect 590110 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect 590110 208574 590730 208658
rect 590110 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect 590110 172894 590730 208338
rect 590110 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect 590110 172574 590730 172658
rect 590110 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect 590110 136894 590730 172338
rect 590110 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect 590110 136574 590730 136658
rect 590110 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect 590110 100894 590730 136338
rect 590110 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect 590110 100574 590730 100658
rect 590110 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect 590110 64894 590730 100338
rect 590110 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect 590110 64574 590730 64658
rect 590110 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect 590110 28894 590730 64338
rect 590110 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect 590110 28574 590730 28658
rect 590110 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect 590110 -5146 590730 28338
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 698614 591690 710042
rect 591070 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 591690 698614
rect 591070 698294 591690 698378
rect 591070 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 591690 698294
rect 591070 662614 591690 698058
rect 591070 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 591690 662614
rect 591070 662294 591690 662378
rect 591070 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 591690 662294
rect 591070 626614 591690 662058
rect 591070 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 591690 626614
rect 591070 626294 591690 626378
rect 591070 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 591690 626294
rect 591070 590614 591690 626058
rect 591070 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 591690 590614
rect 591070 590294 591690 590378
rect 591070 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 591690 590294
rect 591070 554614 591690 590058
rect 591070 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 591690 554614
rect 591070 554294 591690 554378
rect 591070 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 591690 554294
rect 591070 518614 591690 554058
rect 591070 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 591690 518614
rect 591070 518294 591690 518378
rect 591070 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 591690 518294
rect 591070 482614 591690 518058
rect 591070 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 591690 482614
rect 591070 482294 591690 482378
rect 591070 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 591690 482294
rect 591070 446614 591690 482058
rect 591070 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 591690 446614
rect 591070 446294 591690 446378
rect 591070 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 591690 446294
rect 591070 410614 591690 446058
rect 591070 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 591690 410614
rect 591070 410294 591690 410378
rect 591070 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 591690 410294
rect 591070 374614 591690 410058
rect 591070 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 591690 374614
rect 591070 374294 591690 374378
rect 591070 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 591690 374294
rect 591070 338614 591690 374058
rect 591070 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 591690 338614
rect 591070 338294 591690 338378
rect 591070 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 591690 338294
rect 591070 302614 591690 338058
rect 591070 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 591690 302614
rect 591070 302294 591690 302378
rect 591070 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 591690 302294
rect 591070 266614 591690 302058
rect 591070 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 591690 266614
rect 591070 266294 591690 266378
rect 591070 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 591690 266294
rect 591070 230614 591690 266058
rect 591070 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 591690 230614
rect 591070 230294 591690 230378
rect 591070 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 591690 230294
rect 591070 194614 591690 230058
rect 591070 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 591690 194614
rect 591070 194294 591690 194378
rect 591070 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 591690 194294
rect 591070 158614 591690 194058
rect 591070 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 591690 158614
rect 591070 158294 591690 158378
rect 591070 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 591690 158294
rect 591070 122614 591690 158058
rect 591070 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 591690 122614
rect 591070 122294 591690 122378
rect 591070 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 591690 122294
rect 591070 86614 591690 122058
rect 591070 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 591690 86614
rect 591070 86294 591690 86378
rect 591070 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 591690 86294
rect 591070 50614 591690 86058
rect 591070 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 591690 50614
rect 591070 50294 591690 50378
rect 591070 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 591690 50294
rect 591070 14614 591690 50058
rect 591070 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 591690 14614
rect 591070 14294 591690 14378
rect 591070 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 591690 14294
rect 591070 -6106 591690 14058
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 680614 592650 711002
rect 592030 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect 592030 680294 592650 680378
rect 592030 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect 592030 644614 592650 680058
rect 592030 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect 592030 644294 592650 644378
rect 592030 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect 592030 608614 592650 644058
rect 592030 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect 592030 608294 592650 608378
rect 592030 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect 592030 572614 592650 608058
rect 592030 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect 592030 572294 592650 572378
rect 592030 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect 592030 536614 592650 572058
rect 592030 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect 592030 536294 592650 536378
rect 592030 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect 592030 500614 592650 536058
rect 592030 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect 592030 500294 592650 500378
rect 592030 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect 592030 464614 592650 500058
rect 592030 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect 592030 464294 592650 464378
rect 592030 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect 592030 428614 592650 464058
rect 592030 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect 592030 428294 592650 428378
rect 592030 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect 592030 392614 592650 428058
rect 592030 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect 592030 392294 592650 392378
rect 592030 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect 592030 356614 592650 392058
rect 592030 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect 592030 356294 592650 356378
rect 592030 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect 592030 320614 592650 356058
rect 592030 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect 592030 320294 592650 320378
rect 592030 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect 592030 284614 592650 320058
rect 592030 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect 592030 284294 592650 284378
rect 592030 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect 592030 248614 592650 284058
rect 592030 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect 592030 248294 592650 248378
rect 592030 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect 592030 212614 592650 248058
rect 592030 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect 592030 212294 592650 212378
rect 592030 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect 592030 176614 592650 212058
rect 592030 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect 592030 176294 592650 176378
rect 592030 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect 592030 140614 592650 176058
rect 592030 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect 592030 140294 592650 140378
rect 592030 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect 592030 104614 592650 140058
rect 592030 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect 592030 104294 592650 104378
rect 592030 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect 592030 68614 592650 104058
rect 592030 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect 592030 68294 592650 68378
rect 592030 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect 592030 32614 592650 68058
rect 592030 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect 592030 32294 592650 32378
rect 592030 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect 570954 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 571574 -7066
rect 570954 -7386 571574 -7302
rect 570954 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 571574 -7386
rect 570954 -7654 571574 -7622
rect 592030 -7066 592650 32058
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 680378 -8458 680614
rect -8374 680378 -8138 680614
rect -8694 680058 -8458 680294
rect -8374 680058 -8138 680294
rect -8694 644378 -8458 644614
rect -8374 644378 -8138 644614
rect -8694 644058 -8458 644294
rect -8374 644058 -8138 644294
rect -8694 608378 -8458 608614
rect -8374 608378 -8138 608614
rect -8694 608058 -8458 608294
rect -8374 608058 -8138 608294
rect -8694 572378 -8458 572614
rect -8374 572378 -8138 572614
rect -8694 572058 -8458 572294
rect -8374 572058 -8138 572294
rect -8694 536378 -8458 536614
rect -8374 536378 -8138 536614
rect -8694 536058 -8458 536294
rect -8374 536058 -8138 536294
rect -8694 500378 -8458 500614
rect -8374 500378 -8138 500614
rect -8694 500058 -8458 500294
rect -8374 500058 -8138 500294
rect -8694 464378 -8458 464614
rect -8374 464378 -8138 464614
rect -8694 464058 -8458 464294
rect -8374 464058 -8138 464294
rect -8694 428378 -8458 428614
rect -8374 428378 -8138 428614
rect -8694 428058 -8458 428294
rect -8374 428058 -8138 428294
rect -8694 392378 -8458 392614
rect -8374 392378 -8138 392614
rect -8694 392058 -8458 392294
rect -8374 392058 -8138 392294
rect -8694 356378 -8458 356614
rect -8374 356378 -8138 356614
rect -8694 356058 -8458 356294
rect -8374 356058 -8138 356294
rect -8694 320378 -8458 320614
rect -8374 320378 -8138 320614
rect -8694 320058 -8458 320294
rect -8374 320058 -8138 320294
rect -8694 284378 -8458 284614
rect -8374 284378 -8138 284614
rect -8694 284058 -8458 284294
rect -8374 284058 -8138 284294
rect -8694 248378 -8458 248614
rect -8374 248378 -8138 248614
rect -8694 248058 -8458 248294
rect -8374 248058 -8138 248294
rect -8694 212378 -8458 212614
rect -8374 212378 -8138 212614
rect -8694 212058 -8458 212294
rect -8374 212058 -8138 212294
rect -8694 176378 -8458 176614
rect -8374 176378 -8138 176614
rect -8694 176058 -8458 176294
rect -8374 176058 -8138 176294
rect -8694 140378 -8458 140614
rect -8374 140378 -8138 140614
rect -8694 140058 -8458 140294
rect -8374 140058 -8138 140294
rect -8694 104378 -8458 104614
rect -8374 104378 -8138 104614
rect -8694 104058 -8458 104294
rect -8374 104058 -8138 104294
rect -8694 68378 -8458 68614
rect -8374 68378 -8138 68614
rect -8694 68058 -8458 68294
rect -8374 68058 -8138 68294
rect -8694 32378 -8458 32614
rect -8374 32378 -8138 32614
rect -8694 32058 -8458 32294
rect -8374 32058 -8138 32294
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect 12986 710362 13222 710598
rect 13306 710362 13542 710598
rect 12986 710042 13222 710278
rect 13306 710042 13542 710278
rect -7734 698378 -7498 698614
rect -7414 698378 -7178 698614
rect -7734 698058 -7498 698294
rect -7414 698058 -7178 698294
rect -7734 662378 -7498 662614
rect -7414 662378 -7178 662614
rect -7734 662058 -7498 662294
rect -7414 662058 -7178 662294
rect -7734 626378 -7498 626614
rect -7414 626378 -7178 626614
rect -7734 626058 -7498 626294
rect -7414 626058 -7178 626294
rect -7734 590378 -7498 590614
rect -7414 590378 -7178 590614
rect -7734 590058 -7498 590294
rect -7414 590058 -7178 590294
rect -7734 554378 -7498 554614
rect -7414 554378 -7178 554614
rect -7734 554058 -7498 554294
rect -7414 554058 -7178 554294
rect -7734 518378 -7498 518614
rect -7414 518378 -7178 518614
rect -7734 518058 -7498 518294
rect -7414 518058 -7178 518294
rect -7734 482378 -7498 482614
rect -7414 482378 -7178 482614
rect -7734 482058 -7498 482294
rect -7414 482058 -7178 482294
rect -7734 446378 -7498 446614
rect -7414 446378 -7178 446614
rect -7734 446058 -7498 446294
rect -7414 446058 -7178 446294
rect -7734 410378 -7498 410614
rect -7414 410378 -7178 410614
rect -7734 410058 -7498 410294
rect -7414 410058 -7178 410294
rect -7734 374378 -7498 374614
rect -7414 374378 -7178 374614
rect -7734 374058 -7498 374294
rect -7414 374058 -7178 374294
rect -7734 338378 -7498 338614
rect -7414 338378 -7178 338614
rect -7734 338058 -7498 338294
rect -7414 338058 -7178 338294
rect -7734 302378 -7498 302614
rect -7414 302378 -7178 302614
rect -7734 302058 -7498 302294
rect -7414 302058 -7178 302294
rect -7734 266378 -7498 266614
rect -7414 266378 -7178 266614
rect -7734 266058 -7498 266294
rect -7414 266058 -7178 266294
rect -7734 230378 -7498 230614
rect -7414 230378 -7178 230614
rect -7734 230058 -7498 230294
rect -7414 230058 -7178 230294
rect -7734 194378 -7498 194614
rect -7414 194378 -7178 194614
rect -7734 194058 -7498 194294
rect -7414 194058 -7178 194294
rect -7734 158378 -7498 158614
rect -7414 158378 -7178 158614
rect -7734 158058 -7498 158294
rect -7414 158058 -7178 158294
rect -7734 122378 -7498 122614
rect -7414 122378 -7178 122614
rect -7734 122058 -7498 122294
rect -7414 122058 -7178 122294
rect -7734 86378 -7498 86614
rect -7414 86378 -7178 86614
rect -7734 86058 -7498 86294
rect -7414 86058 -7178 86294
rect -7734 50378 -7498 50614
rect -7414 50378 -7178 50614
rect -7734 50058 -7498 50294
rect -7414 50058 -7178 50294
rect -7734 14378 -7498 14614
rect -7414 14378 -7178 14614
rect -7734 14058 -7498 14294
rect -7414 14058 -7178 14294
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 676658 -6538 676894
rect -6454 676658 -6218 676894
rect -6774 676338 -6538 676574
rect -6454 676338 -6218 676574
rect -6774 640658 -6538 640894
rect -6454 640658 -6218 640894
rect -6774 640338 -6538 640574
rect -6454 640338 -6218 640574
rect -6774 604658 -6538 604894
rect -6454 604658 -6218 604894
rect -6774 604338 -6538 604574
rect -6454 604338 -6218 604574
rect -6774 568658 -6538 568894
rect -6454 568658 -6218 568894
rect -6774 568338 -6538 568574
rect -6454 568338 -6218 568574
rect -6774 532658 -6538 532894
rect -6454 532658 -6218 532894
rect -6774 532338 -6538 532574
rect -6454 532338 -6218 532574
rect -6774 496658 -6538 496894
rect -6454 496658 -6218 496894
rect -6774 496338 -6538 496574
rect -6454 496338 -6218 496574
rect -6774 460658 -6538 460894
rect -6454 460658 -6218 460894
rect -6774 460338 -6538 460574
rect -6454 460338 -6218 460574
rect -6774 424658 -6538 424894
rect -6454 424658 -6218 424894
rect -6774 424338 -6538 424574
rect -6454 424338 -6218 424574
rect -6774 388658 -6538 388894
rect -6454 388658 -6218 388894
rect -6774 388338 -6538 388574
rect -6454 388338 -6218 388574
rect -6774 352658 -6538 352894
rect -6454 352658 -6218 352894
rect -6774 352338 -6538 352574
rect -6454 352338 -6218 352574
rect -6774 316658 -6538 316894
rect -6454 316658 -6218 316894
rect -6774 316338 -6538 316574
rect -6454 316338 -6218 316574
rect -6774 280658 -6538 280894
rect -6454 280658 -6218 280894
rect -6774 280338 -6538 280574
rect -6454 280338 -6218 280574
rect -6774 244658 -6538 244894
rect -6454 244658 -6218 244894
rect -6774 244338 -6538 244574
rect -6454 244338 -6218 244574
rect -6774 208658 -6538 208894
rect -6454 208658 -6218 208894
rect -6774 208338 -6538 208574
rect -6454 208338 -6218 208574
rect -6774 172658 -6538 172894
rect -6454 172658 -6218 172894
rect -6774 172338 -6538 172574
rect -6454 172338 -6218 172574
rect -6774 136658 -6538 136894
rect -6454 136658 -6218 136894
rect -6774 136338 -6538 136574
rect -6454 136338 -6218 136574
rect -6774 100658 -6538 100894
rect -6454 100658 -6218 100894
rect -6774 100338 -6538 100574
rect -6454 100338 -6218 100574
rect -6774 64658 -6538 64894
rect -6454 64658 -6218 64894
rect -6774 64338 -6538 64574
rect -6454 64338 -6218 64574
rect -6774 28658 -6538 28894
rect -6454 28658 -6218 28894
rect -6774 28338 -6538 28574
rect -6454 28338 -6218 28574
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect 9266 708442 9502 708678
rect 9586 708442 9822 708678
rect 9266 708122 9502 708358
rect 9586 708122 9822 708358
rect -5814 694658 -5578 694894
rect -5494 694658 -5258 694894
rect -5814 694338 -5578 694574
rect -5494 694338 -5258 694574
rect -5814 658658 -5578 658894
rect -5494 658658 -5258 658894
rect -5814 658338 -5578 658574
rect -5494 658338 -5258 658574
rect -5814 622658 -5578 622894
rect -5494 622658 -5258 622894
rect -5814 622338 -5578 622574
rect -5494 622338 -5258 622574
rect -5814 586658 -5578 586894
rect -5494 586658 -5258 586894
rect -5814 586338 -5578 586574
rect -5494 586338 -5258 586574
rect -5814 550658 -5578 550894
rect -5494 550658 -5258 550894
rect -5814 550338 -5578 550574
rect -5494 550338 -5258 550574
rect -5814 514658 -5578 514894
rect -5494 514658 -5258 514894
rect -5814 514338 -5578 514574
rect -5494 514338 -5258 514574
rect -5814 478658 -5578 478894
rect -5494 478658 -5258 478894
rect -5814 478338 -5578 478574
rect -5494 478338 -5258 478574
rect -5814 442658 -5578 442894
rect -5494 442658 -5258 442894
rect -5814 442338 -5578 442574
rect -5494 442338 -5258 442574
rect -5814 406658 -5578 406894
rect -5494 406658 -5258 406894
rect -5814 406338 -5578 406574
rect -5494 406338 -5258 406574
rect -5814 370658 -5578 370894
rect -5494 370658 -5258 370894
rect -5814 370338 -5578 370574
rect -5494 370338 -5258 370574
rect -5814 334658 -5578 334894
rect -5494 334658 -5258 334894
rect -5814 334338 -5578 334574
rect -5494 334338 -5258 334574
rect -5814 298658 -5578 298894
rect -5494 298658 -5258 298894
rect -5814 298338 -5578 298574
rect -5494 298338 -5258 298574
rect -5814 262658 -5578 262894
rect -5494 262658 -5258 262894
rect -5814 262338 -5578 262574
rect -5494 262338 -5258 262574
rect -5814 226658 -5578 226894
rect -5494 226658 -5258 226894
rect -5814 226338 -5578 226574
rect -5494 226338 -5258 226574
rect -5814 190658 -5578 190894
rect -5494 190658 -5258 190894
rect -5814 190338 -5578 190574
rect -5494 190338 -5258 190574
rect -5814 154658 -5578 154894
rect -5494 154658 -5258 154894
rect -5814 154338 -5578 154574
rect -5494 154338 -5258 154574
rect -5814 118658 -5578 118894
rect -5494 118658 -5258 118894
rect -5814 118338 -5578 118574
rect -5494 118338 -5258 118574
rect -5814 82658 -5578 82894
rect -5494 82658 -5258 82894
rect -5814 82338 -5578 82574
rect -5494 82338 -5258 82574
rect -5814 46658 -5578 46894
rect -5494 46658 -5258 46894
rect -5814 46338 -5578 46574
rect -5494 46338 -5258 46574
rect -5814 10658 -5578 10894
rect -5494 10658 -5258 10894
rect -5814 10338 -5578 10574
rect -5494 10338 -5258 10574
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 672938 -4618 673174
rect -4534 672938 -4298 673174
rect -4854 672618 -4618 672854
rect -4534 672618 -4298 672854
rect -4854 636938 -4618 637174
rect -4534 636938 -4298 637174
rect -4854 636618 -4618 636854
rect -4534 636618 -4298 636854
rect -4854 600938 -4618 601174
rect -4534 600938 -4298 601174
rect -4854 600618 -4618 600854
rect -4534 600618 -4298 600854
rect -4854 564938 -4618 565174
rect -4534 564938 -4298 565174
rect -4854 564618 -4618 564854
rect -4534 564618 -4298 564854
rect -4854 528938 -4618 529174
rect -4534 528938 -4298 529174
rect -4854 528618 -4618 528854
rect -4534 528618 -4298 528854
rect -4854 492938 -4618 493174
rect -4534 492938 -4298 493174
rect -4854 492618 -4618 492854
rect -4534 492618 -4298 492854
rect -4854 456938 -4618 457174
rect -4534 456938 -4298 457174
rect -4854 456618 -4618 456854
rect -4534 456618 -4298 456854
rect -4854 420938 -4618 421174
rect -4534 420938 -4298 421174
rect -4854 420618 -4618 420854
rect -4534 420618 -4298 420854
rect -4854 384938 -4618 385174
rect -4534 384938 -4298 385174
rect -4854 384618 -4618 384854
rect -4534 384618 -4298 384854
rect -4854 348938 -4618 349174
rect -4534 348938 -4298 349174
rect -4854 348618 -4618 348854
rect -4534 348618 -4298 348854
rect -4854 312938 -4618 313174
rect -4534 312938 -4298 313174
rect -4854 312618 -4618 312854
rect -4534 312618 -4298 312854
rect -4854 276938 -4618 277174
rect -4534 276938 -4298 277174
rect -4854 276618 -4618 276854
rect -4534 276618 -4298 276854
rect -4854 240938 -4618 241174
rect -4534 240938 -4298 241174
rect -4854 240618 -4618 240854
rect -4534 240618 -4298 240854
rect -4854 204938 -4618 205174
rect -4534 204938 -4298 205174
rect -4854 204618 -4618 204854
rect -4534 204618 -4298 204854
rect -4854 168938 -4618 169174
rect -4534 168938 -4298 169174
rect -4854 168618 -4618 168854
rect -4534 168618 -4298 168854
rect -4854 132938 -4618 133174
rect -4534 132938 -4298 133174
rect -4854 132618 -4618 132854
rect -4534 132618 -4298 132854
rect -4854 96938 -4618 97174
rect -4534 96938 -4298 97174
rect -4854 96618 -4618 96854
rect -4534 96618 -4298 96854
rect -4854 60938 -4618 61174
rect -4534 60938 -4298 61174
rect -4854 60618 -4618 60854
rect -4534 60618 -4298 60854
rect -4854 24938 -4618 25174
rect -4534 24938 -4298 25174
rect -4854 24618 -4618 24854
rect -4534 24618 -4298 24854
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect 5546 706522 5782 706758
rect 5866 706522 6102 706758
rect 5546 706202 5782 706438
rect 5866 706202 6102 706438
rect -3894 690938 -3658 691174
rect -3574 690938 -3338 691174
rect -3894 690618 -3658 690854
rect -3574 690618 -3338 690854
rect -3894 654938 -3658 655174
rect -3574 654938 -3338 655174
rect -3894 654618 -3658 654854
rect -3574 654618 -3338 654854
rect -3894 618938 -3658 619174
rect -3574 618938 -3338 619174
rect -3894 618618 -3658 618854
rect -3574 618618 -3338 618854
rect -3894 582938 -3658 583174
rect -3574 582938 -3338 583174
rect -3894 582618 -3658 582854
rect -3574 582618 -3338 582854
rect -3894 546938 -3658 547174
rect -3574 546938 -3338 547174
rect -3894 546618 -3658 546854
rect -3574 546618 -3338 546854
rect -3894 510938 -3658 511174
rect -3574 510938 -3338 511174
rect -3894 510618 -3658 510854
rect -3574 510618 -3338 510854
rect -3894 474938 -3658 475174
rect -3574 474938 -3338 475174
rect -3894 474618 -3658 474854
rect -3574 474618 -3338 474854
rect -3894 438938 -3658 439174
rect -3574 438938 -3338 439174
rect -3894 438618 -3658 438854
rect -3574 438618 -3338 438854
rect -3894 402938 -3658 403174
rect -3574 402938 -3338 403174
rect -3894 402618 -3658 402854
rect -3574 402618 -3338 402854
rect -3894 366938 -3658 367174
rect -3574 366938 -3338 367174
rect -3894 366618 -3658 366854
rect -3574 366618 -3338 366854
rect -3894 330938 -3658 331174
rect -3574 330938 -3338 331174
rect -3894 330618 -3658 330854
rect -3574 330618 -3338 330854
rect -3894 294938 -3658 295174
rect -3574 294938 -3338 295174
rect -3894 294618 -3658 294854
rect -3574 294618 -3338 294854
rect -3894 258938 -3658 259174
rect -3574 258938 -3338 259174
rect -3894 258618 -3658 258854
rect -3574 258618 -3338 258854
rect -3894 222938 -3658 223174
rect -3574 222938 -3338 223174
rect -3894 222618 -3658 222854
rect -3574 222618 -3338 222854
rect -3894 186938 -3658 187174
rect -3574 186938 -3338 187174
rect -3894 186618 -3658 186854
rect -3574 186618 -3338 186854
rect -3894 150938 -3658 151174
rect -3574 150938 -3338 151174
rect -3894 150618 -3658 150854
rect -3574 150618 -3338 150854
rect -3894 114938 -3658 115174
rect -3574 114938 -3338 115174
rect -3894 114618 -3658 114854
rect -3574 114618 -3338 114854
rect -3894 78938 -3658 79174
rect -3574 78938 -3338 79174
rect -3894 78618 -3658 78854
rect -3574 78618 -3338 78854
rect -3894 42938 -3658 43174
rect -3574 42938 -3338 43174
rect -3894 42618 -3658 42854
rect -3574 42618 -3338 42854
rect -3894 6938 -3658 7174
rect -3574 6938 -3338 7174
rect -3894 6618 -3658 6854
rect -3574 6618 -3338 6854
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 669218 -2698 669454
rect -2614 669218 -2378 669454
rect -2934 668898 -2698 669134
rect -2614 668898 -2378 669134
rect -2934 633218 -2698 633454
rect -2614 633218 -2378 633454
rect -2934 632898 -2698 633134
rect -2614 632898 -2378 633134
rect -2934 597218 -2698 597454
rect -2614 597218 -2378 597454
rect -2934 596898 -2698 597134
rect -2614 596898 -2378 597134
rect -2934 561218 -2698 561454
rect -2614 561218 -2378 561454
rect -2934 560898 -2698 561134
rect -2614 560898 -2378 561134
rect -2934 525218 -2698 525454
rect -2614 525218 -2378 525454
rect -2934 524898 -2698 525134
rect -2614 524898 -2378 525134
rect -2934 489218 -2698 489454
rect -2614 489218 -2378 489454
rect -2934 488898 -2698 489134
rect -2614 488898 -2378 489134
rect -2934 453218 -2698 453454
rect -2614 453218 -2378 453454
rect -2934 452898 -2698 453134
rect -2614 452898 -2378 453134
rect -2934 417218 -2698 417454
rect -2614 417218 -2378 417454
rect -2934 416898 -2698 417134
rect -2614 416898 -2378 417134
rect -2934 381218 -2698 381454
rect -2614 381218 -2378 381454
rect -2934 380898 -2698 381134
rect -2614 380898 -2378 381134
rect -2934 345218 -2698 345454
rect -2614 345218 -2378 345454
rect -2934 344898 -2698 345134
rect -2614 344898 -2378 345134
rect -2934 309218 -2698 309454
rect -2614 309218 -2378 309454
rect -2934 308898 -2698 309134
rect -2614 308898 -2378 309134
rect -2934 273218 -2698 273454
rect -2614 273218 -2378 273454
rect -2934 272898 -2698 273134
rect -2614 272898 -2378 273134
rect -2934 237218 -2698 237454
rect -2614 237218 -2378 237454
rect -2934 236898 -2698 237134
rect -2614 236898 -2378 237134
rect -2934 201218 -2698 201454
rect -2614 201218 -2378 201454
rect -2934 200898 -2698 201134
rect -2614 200898 -2378 201134
rect -2934 165218 -2698 165454
rect -2614 165218 -2378 165454
rect -2934 164898 -2698 165134
rect -2614 164898 -2378 165134
rect -2934 129218 -2698 129454
rect -2614 129218 -2378 129454
rect -2934 128898 -2698 129134
rect -2614 128898 -2378 129134
rect -2934 93218 -2698 93454
rect -2614 93218 -2378 93454
rect -2934 92898 -2698 93134
rect -2614 92898 -2378 93134
rect -2934 57218 -2698 57454
rect -2614 57218 -2378 57454
rect -2934 56898 -2698 57134
rect -2614 56898 -2378 57134
rect -2934 21218 -2698 21454
rect -2614 21218 -2378 21454
rect -2934 20898 -2698 21134
rect -2614 20898 -2378 21134
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect 5546 -2502 5782 -2266
rect 5866 -2502 6102 -2266
rect 5546 -2822 5782 -2586
rect 5866 -2822 6102 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect 9266 694658 9502 694894
rect 9586 694658 9822 694894
rect 9266 694338 9502 694574
rect 9586 694338 9822 694574
rect 9266 658658 9502 658894
rect 9586 658658 9822 658894
rect 9266 658338 9502 658574
rect 9586 658338 9822 658574
rect 9266 622658 9502 622894
rect 9586 622658 9822 622894
rect 9266 622338 9502 622574
rect 9586 622338 9822 622574
rect 9266 586658 9502 586894
rect 9586 586658 9822 586894
rect 9266 586338 9502 586574
rect 9586 586338 9822 586574
rect 9266 550658 9502 550894
rect 9586 550658 9822 550894
rect 9266 550338 9502 550574
rect 9586 550338 9822 550574
rect 9266 514658 9502 514894
rect 9586 514658 9822 514894
rect 9266 514338 9502 514574
rect 9586 514338 9822 514574
rect 9266 478658 9502 478894
rect 9586 478658 9822 478894
rect 9266 478338 9502 478574
rect 9586 478338 9822 478574
rect 9266 442658 9502 442894
rect 9586 442658 9822 442894
rect 9266 442338 9502 442574
rect 9586 442338 9822 442574
rect 9266 406658 9502 406894
rect 9586 406658 9822 406894
rect 9266 406338 9502 406574
rect 9586 406338 9822 406574
rect 9266 370658 9502 370894
rect 9586 370658 9822 370894
rect 9266 370338 9502 370574
rect 9586 370338 9822 370574
rect 9266 334658 9502 334894
rect 9586 334658 9822 334894
rect 9266 334338 9502 334574
rect 9586 334338 9822 334574
rect 9266 298658 9502 298894
rect 9586 298658 9822 298894
rect 9266 298338 9502 298574
rect 9586 298338 9822 298574
rect 9266 262658 9502 262894
rect 9586 262658 9822 262894
rect 9266 262338 9502 262574
rect 9586 262338 9822 262574
rect 9266 226658 9502 226894
rect 9586 226658 9822 226894
rect 9266 226338 9502 226574
rect 9586 226338 9822 226574
rect 9266 190658 9502 190894
rect 9586 190658 9822 190894
rect 9266 190338 9502 190574
rect 9586 190338 9822 190574
rect 9266 154658 9502 154894
rect 9586 154658 9822 154894
rect 9266 154338 9502 154574
rect 9586 154338 9822 154574
rect 9266 118658 9502 118894
rect 9586 118658 9822 118894
rect 9266 118338 9502 118574
rect 9586 118338 9822 118574
rect 9266 82658 9502 82894
rect 9586 82658 9822 82894
rect 9266 82338 9502 82574
rect 9586 82338 9822 82574
rect 9266 46658 9502 46894
rect 9586 46658 9822 46894
rect 9266 46338 9502 46574
rect 9586 46338 9822 46574
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect 9266 -4422 9502 -4186
rect 9586 -4422 9822 -4186
rect 9266 -4742 9502 -4506
rect 9586 -4742 9822 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect 30986 711322 31222 711558
rect 31306 711322 31542 711558
rect 30986 711002 31222 711238
rect 31306 711002 31542 711238
rect 27266 709402 27502 709638
rect 27586 709402 27822 709638
rect 27266 709082 27502 709318
rect 27586 709082 27822 709318
rect 23546 707482 23782 707718
rect 23866 707482 24102 707718
rect 23546 707162 23782 707398
rect 23866 707162 24102 707398
rect 12986 698378 13222 698614
rect 13306 698378 13542 698614
rect 12986 698058 13222 698294
rect 13306 698058 13542 698294
rect 12986 662378 13222 662614
rect 13306 662378 13542 662614
rect 12986 662058 13222 662294
rect 13306 662058 13542 662294
rect 12986 626378 13222 626614
rect 13306 626378 13542 626614
rect 12986 626058 13222 626294
rect 13306 626058 13542 626294
rect 12986 590378 13222 590614
rect 13306 590378 13542 590614
rect 12986 590058 13222 590294
rect 13306 590058 13542 590294
rect 12986 554378 13222 554614
rect 13306 554378 13542 554614
rect 12986 554058 13222 554294
rect 13306 554058 13542 554294
rect 12986 518378 13222 518614
rect 13306 518378 13542 518614
rect 12986 518058 13222 518294
rect 13306 518058 13542 518294
rect 12986 482378 13222 482614
rect 13306 482378 13542 482614
rect 12986 482058 13222 482294
rect 13306 482058 13542 482294
rect 12986 446378 13222 446614
rect 13306 446378 13542 446614
rect 12986 446058 13222 446294
rect 13306 446058 13542 446294
rect 12986 410378 13222 410614
rect 13306 410378 13542 410614
rect 12986 410058 13222 410294
rect 13306 410058 13542 410294
rect 12986 374378 13222 374614
rect 13306 374378 13542 374614
rect 12986 374058 13222 374294
rect 13306 374058 13542 374294
rect 12986 338378 13222 338614
rect 13306 338378 13542 338614
rect 12986 338058 13222 338294
rect 13306 338058 13542 338294
rect 12986 302378 13222 302614
rect 13306 302378 13542 302614
rect 12986 302058 13222 302294
rect 13306 302058 13542 302294
rect 12986 266378 13222 266614
rect 13306 266378 13542 266614
rect 12986 266058 13222 266294
rect 13306 266058 13542 266294
rect 12986 230378 13222 230614
rect 13306 230378 13542 230614
rect 12986 230058 13222 230294
rect 13306 230058 13542 230294
rect 12986 194378 13222 194614
rect 13306 194378 13542 194614
rect 12986 194058 13222 194294
rect 13306 194058 13542 194294
rect 12986 158378 13222 158614
rect 13306 158378 13542 158614
rect 12986 158058 13222 158294
rect 13306 158058 13542 158294
rect 12986 122378 13222 122614
rect 13306 122378 13542 122614
rect 12986 122058 13222 122294
rect 13306 122058 13542 122294
rect 12986 86378 13222 86614
rect 13306 86378 13542 86614
rect 12986 86058 13222 86294
rect 13306 86058 13542 86294
rect 12986 50378 13222 50614
rect 13306 50378 13542 50614
rect 12986 50058 13222 50294
rect 13306 50058 13542 50294
rect 12986 14378 13222 14614
rect 13306 14378 13542 14614
rect 12986 14058 13222 14294
rect 13306 14058 13542 14294
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect 19826 705562 20062 705798
rect 20146 705562 20382 705798
rect 19826 705242 20062 705478
rect 20146 705242 20382 705478
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -1542 20062 -1306
rect 20146 -1542 20382 -1306
rect 19826 -1862 20062 -1626
rect 20146 -1862 20382 -1626
rect 23546 672938 23782 673174
rect 23866 672938 24102 673174
rect 23546 672618 23782 672854
rect 23866 672618 24102 672854
rect 23546 636938 23782 637174
rect 23866 636938 24102 637174
rect 23546 636618 23782 636854
rect 23866 636618 24102 636854
rect 23546 600938 23782 601174
rect 23866 600938 24102 601174
rect 23546 600618 23782 600854
rect 23866 600618 24102 600854
rect 23546 564938 23782 565174
rect 23866 564938 24102 565174
rect 23546 564618 23782 564854
rect 23866 564618 24102 564854
rect 23546 528938 23782 529174
rect 23866 528938 24102 529174
rect 23546 528618 23782 528854
rect 23866 528618 24102 528854
rect 23546 492938 23782 493174
rect 23866 492938 24102 493174
rect 23546 492618 23782 492854
rect 23866 492618 24102 492854
rect 23546 456938 23782 457174
rect 23866 456938 24102 457174
rect 23546 456618 23782 456854
rect 23866 456618 24102 456854
rect 23546 420938 23782 421174
rect 23866 420938 24102 421174
rect 23546 420618 23782 420854
rect 23866 420618 24102 420854
rect 23546 384938 23782 385174
rect 23866 384938 24102 385174
rect 23546 384618 23782 384854
rect 23866 384618 24102 384854
rect 23546 348938 23782 349174
rect 23866 348938 24102 349174
rect 23546 348618 23782 348854
rect 23866 348618 24102 348854
rect 23546 312938 23782 313174
rect 23866 312938 24102 313174
rect 23546 312618 23782 312854
rect 23866 312618 24102 312854
rect 23546 276938 23782 277174
rect 23866 276938 24102 277174
rect 23546 276618 23782 276854
rect 23866 276618 24102 276854
rect 23546 240938 23782 241174
rect 23866 240938 24102 241174
rect 23546 240618 23782 240854
rect 23866 240618 24102 240854
rect 23546 204938 23782 205174
rect 23866 204938 24102 205174
rect 23546 204618 23782 204854
rect 23866 204618 24102 204854
rect 23546 168938 23782 169174
rect 23866 168938 24102 169174
rect 23546 168618 23782 168854
rect 23866 168618 24102 168854
rect 23546 132938 23782 133174
rect 23866 132938 24102 133174
rect 23546 132618 23782 132854
rect 23866 132618 24102 132854
rect 23546 96938 23782 97174
rect 23866 96938 24102 97174
rect 23546 96618 23782 96854
rect 23866 96618 24102 96854
rect 23546 60938 23782 61174
rect 23866 60938 24102 61174
rect 23546 60618 23782 60854
rect 23866 60618 24102 60854
rect 23546 24938 23782 25174
rect 23866 24938 24102 25174
rect 23546 24618 23782 24854
rect 23866 24618 24102 24854
rect 23546 -3462 23782 -3226
rect 23866 -3462 24102 -3226
rect 23546 -3782 23782 -3546
rect 23866 -3782 24102 -3546
rect 27266 676658 27502 676894
rect 27586 676658 27822 676894
rect 27266 676338 27502 676574
rect 27586 676338 27822 676574
rect 27266 640658 27502 640894
rect 27586 640658 27822 640894
rect 27266 640338 27502 640574
rect 27586 640338 27822 640574
rect 27266 604658 27502 604894
rect 27586 604658 27822 604894
rect 27266 604338 27502 604574
rect 27586 604338 27822 604574
rect 27266 568658 27502 568894
rect 27586 568658 27822 568894
rect 27266 568338 27502 568574
rect 27586 568338 27822 568574
rect 27266 532658 27502 532894
rect 27586 532658 27822 532894
rect 27266 532338 27502 532574
rect 27586 532338 27822 532574
rect 27266 496658 27502 496894
rect 27586 496658 27822 496894
rect 27266 496338 27502 496574
rect 27586 496338 27822 496574
rect 27266 460658 27502 460894
rect 27586 460658 27822 460894
rect 27266 460338 27502 460574
rect 27586 460338 27822 460574
rect 27266 424658 27502 424894
rect 27586 424658 27822 424894
rect 27266 424338 27502 424574
rect 27586 424338 27822 424574
rect 27266 388658 27502 388894
rect 27586 388658 27822 388894
rect 27266 388338 27502 388574
rect 27586 388338 27822 388574
rect 27266 352658 27502 352894
rect 27586 352658 27822 352894
rect 27266 352338 27502 352574
rect 27586 352338 27822 352574
rect 27266 316658 27502 316894
rect 27586 316658 27822 316894
rect 27266 316338 27502 316574
rect 27586 316338 27822 316574
rect 27266 280658 27502 280894
rect 27586 280658 27822 280894
rect 27266 280338 27502 280574
rect 27586 280338 27822 280574
rect 27266 244658 27502 244894
rect 27586 244658 27822 244894
rect 27266 244338 27502 244574
rect 27586 244338 27822 244574
rect 27266 208658 27502 208894
rect 27586 208658 27822 208894
rect 27266 208338 27502 208574
rect 27586 208338 27822 208574
rect 27266 172658 27502 172894
rect 27586 172658 27822 172894
rect 27266 172338 27502 172574
rect 27586 172338 27822 172574
rect 27266 136658 27502 136894
rect 27586 136658 27822 136894
rect 27266 136338 27502 136574
rect 27586 136338 27822 136574
rect 27266 100658 27502 100894
rect 27586 100658 27822 100894
rect 27266 100338 27502 100574
rect 27586 100338 27822 100574
rect 27266 64658 27502 64894
rect 27586 64658 27822 64894
rect 27266 64338 27502 64574
rect 27586 64338 27822 64574
rect 27266 28658 27502 28894
rect 27586 28658 27822 28894
rect 27266 28338 27502 28574
rect 27586 28338 27822 28574
rect 27266 -5382 27502 -5146
rect 27586 -5382 27822 -5146
rect 27266 -5702 27502 -5466
rect 27586 -5702 27822 -5466
rect 48986 710362 49222 710598
rect 49306 710362 49542 710598
rect 48986 710042 49222 710278
rect 49306 710042 49542 710278
rect 45266 708442 45502 708678
rect 45586 708442 45822 708678
rect 45266 708122 45502 708358
rect 45586 708122 45822 708358
rect 41546 706522 41782 706758
rect 41866 706522 42102 706758
rect 41546 706202 41782 706438
rect 41866 706202 42102 706438
rect 30986 680378 31222 680614
rect 31306 680378 31542 680614
rect 30986 680058 31222 680294
rect 31306 680058 31542 680294
rect 30986 644378 31222 644614
rect 31306 644378 31542 644614
rect 30986 644058 31222 644294
rect 31306 644058 31542 644294
rect 30986 608378 31222 608614
rect 31306 608378 31542 608614
rect 30986 608058 31222 608294
rect 31306 608058 31542 608294
rect 30986 572378 31222 572614
rect 31306 572378 31542 572614
rect 30986 572058 31222 572294
rect 31306 572058 31542 572294
rect 30986 536378 31222 536614
rect 31306 536378 31542 536614
rect 30986 536058 31222 536294
rect 31306 536058 31542 536294
rect 30986 500378 31222 500614
rect 31306 500378 31542 500614
rect 30986 500058 31222 500294
rect 31306 500058 31542 500294
rect 30986 464378 31222 464614
rect 31306 464378 31542 464614
rect 30986 464058 31222 464294
rect 31306 464058 31542 464294
rect 30986 428378 31222 428614
rect 31306 428378 31542 428614
rect 30986 428058 31222 428294
rect 31306 428058 31542 428294
rect 30986 392378 31222 392614
rect 31306 392378 31542 392614
rect 30986 392058 31222 392294
rect 31306 392058 31542 392294
rect 30986 356378 31222 356614
rect 31306 356378 31542 356614
rect 30986 356058 31222 356294
rect 31306 356058 31542 356294
rect 30986 320378 31222 320614
rect 31306 320378 31542 320614
rect 30986 320058 31222 320294
rect 31306 320058 31542 320294
rect 30986 284378 31222 284614
rect 31306 284378 31542 284614
rect 30986 284058 31222 284294
rect 31306 284058 31542 284294
rect 30986 248378 31222 248614
rect 31306 248378 31542 248614
rect 30986 248058 31222 248294
rect 31306 248058 31542 248294
rect 30986 212378 31222 212614
rect 31306 212378 31542 212614
rect 30986 212058 31222 212294
rect 31306 212058 31542 212294
rect 30986 176378 31222 176614
rect 31306 176378 31542 176614
rect 30986 176058 31222 176294
rect 31306 176058 31542 176294
rect 30986 140378 31222 140614
rect 31306 140378 31542 140614
rect 30986 140058 31222 140294
rect 31306 140058 31542 140294
rect 30986 104378 31222 104614
rect 31306 104378 31542 104614
rect 30986 104058 31222 104294
rect 31306 104058 31542 104294
rect 30986 68378 31222 68614
rect 31306 68378 31542 68614
rect 30986 68058 31222 68294
rect 31306 68058 31542 68294
rect 30986 32378 31222 32614
rect 31306 32378 31542 32614
rect 30986 32058 31222 32294
rect 31306 32058 31542 32294
rect 12986 -6342 13222 -6106
rect 13306 -6342 13542 -6106
rect 12986 -6662 13222 -6426
rect 13306 -6662 13542 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 41546 654938 41782 655174
rect 41866 654938 42102 655174
rect 41546 654618 41782 654854
rect 41866 654618 42102 654854
rect 41546 618938 41782 619174
rect 41866 618938 42102 619174
rect 41546 618618 41782 618854
rect 41866 618618 42102 618854
rect 41546 582938 41782 583174
rect 41866 582938 42102 583174
rect 41546 582618 41782 582854
rect 41866 582618 42102 582854
rect 41546 546938 41782 547174
rect 41866 546938 42102 547174
rect 41546 546618 41782 546854
rect 41866 546618 42102 546854
rect 41546 510938 41782 511174
rect 41866 510938 42102 511174
rect 41546 510618 41782 510854
rect 41866 510618 42102 510854
rect 41546 474938 41782 475174
rect 41866 474938 42102 475174
rect 41546 474618 41782 474854
rect 41866 474618 42102 474854
rect 41546 438938 41782 439174
rect 41866 438938 42102 439174
rect 41546 438618 41782 438854
rect 41866 438618 42102 438854
rect 41546 402938 41782 403174
rect 41866 402938 42102 403174
rect 41546 402618 41782 402854
rect 41866 402618 42102 402854
rect 41546 366938 41782 367174
rect 41866 366938 42102 367174
rect 41546 366618 41782 366854
rect 41866 366618 42102 366854
rect 41546 330938 41782 331174
rect 41866 330938 42102 331174
rect 41546 330618 41782 330854
rect 41866 330618 42102 330854
rect 41546 294938 41782 295174
rect 41866 294938 42102 295174
rect 41546 294618 41782 294854
rect 41866 294618 42102 294854
rect 41546 258938 41782 259174
rect 41866 258938 42102 259174
rect 41546 258618 41782 258854
rect 41866 258618 42102 258854
rect 41546 222938 41782 223174
rect 41866 222938 42102 223174
rect 41546 222618 41782 222854
rect 41866 222618 42102 222854
rect 41546 186938 41782 187174
rect 41866 186938 42102 187174
rect 41546 186618 41782 186854
rect 41866 186618 42102 186854
rect 41546 150938 41782 151174
rect 41866 150938 42102 151174
rect 41546 150618 41782 150854
rect 41866 150618 42102 150854
rect 41546 114938 41782 115174
rect 41866 114938 42102 115174
rect 41546 114618 41782 114854
rect 41866 114618 42102 114854
rect 41546 78938 41782 79174
rect 41866 78938 42102 79174
rect 41546 78618 41782 78854
rect 41866 78618 42102 78854
rect 41546 42938 41782 43174
rect 41866 42938 42102 43174
rect 41546 42618 41782 42854
rect 41866 42618 42102 42854
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 41546 -2502 41782 -2266
rect 41866 -2502 42102 -2266
rect 41546 -2822 41782 -2586
rect 41866 -2822 42102 -2586
rect 45266 694658 45502 694894
rect 45586 694658 45822 694894
rect 45266 694338 45502 694574
rect 45586 694338 45822 694574
rect 45266 658658 45502 658894
rect 45586 658658 45822 658894
rect 45266 658338 45502 658574
rect 45586 658338 45822 658574
rect 45266 622658 45502 622894
rect 45586 622658 45822 622894
rect 45266 622338 45502 622574
rect 45586 622338 45822 622574
rect 45266 586658 45502 586894
rect 45586 586658 45822 586894
rect 45266 586338 45502 586574
rect 45586 586338 45822 586574
rect 45266 550658 45502 550894
rect 45586 550658 45822 550894
rect 45266 550338 45502 550574
rect 45586 550338 45822 550574
rect 45266 514658 45502 514894
rect 45586 514658 45822 514894
rect 45266 514338 45502 514574
rect 45586 514338 45822 514574
rect 45266 478658 45502 478894
rect 45586 478658 45822 478894
rect 45266 478338 45502 478574
rect 45586 478338 45822 478574
rect 45266 442658 45502 442894
rect 45586 442658 45822 442894
rect 45266 442338 45502 442574
rect 45586 442338 45822 442574
rect 45266 406658 45502 406894
rect 45586 406658 45822 406894
rect 45266 406338 45502 406574
rect 45586 406338 45822 406574
rect 45266 370658 45502 370894
rect 45586 370658 45822 370894
rect 45266 370338 45502 370574
rect 45586 370338 45822 370574
rect 45266 334658 45502 334894
rect 45586 334658 45822 334894
rect 45266 334338 45502 334574
rect 45586 334338 45822 334574
rect 45266 298658 45502 298894
rect 45586 298658 45822 298894
rect 45266 298338 45502 298574
rect 45586 298338 45822 298574
rect 45266 262658 45502 262894
rect 45586 262658 45822 262894
rect 45266 262338 45502 262574
rect 45586 262338 45822 262574
rect 45266 226658 45502 226894
rect 45586 226658 45822 226894
rect 45266 226338 45502 226574
rect 45586 226338 45822 226574
rect 45266 190658 45502 190894
rect 45586 190658 45822 190894
rect 45266 190338 45502 190574
rect 45586 190338 45822 190574
rect 45266 154658 45502 154894
rect 45586 154658 45822 154894
rect 45266 154338 45502 154574
rect 45586 154338 45822 154574
rect 45266 118658 45502 118894
rect 45586 118658 45822 118894
rect 45266 118338 45502 118574
rect 45586 118338 45822 118574
rect 45266 82658 45502 82894
rect 45586 82658 45822 82894
rect 45266 82338 45502 82574
rect 45586 82338 45822 82574
rect 45266 46658 45502 46894
rect 45586 46658 45822 46894
rect 45266 46338 45502 46574
rect 45586 46338 45822 46574
rect 45266 10658 45502 10894
rect 45586 10658 45822 10894
rect 45266 10338 45502 10574
rect 45586 10338 45822 10574
rect 45266 -4422 45502 -4186
rect 45586 -4422 45822 -4186
rect 45266 -4742 45502 -4506
rect 45586 -4742 45822 -4506
rect 66986 711322 67222 711558
rect 67306 711322 67542 711558
rect 66986 711002 67222 711238
rect 67306 711002 67542 711238
rect 63266 709402 63502 709638
rect 63586 709402 63822 709638
rect 63266 709082 63502 709318
rect 63586 709082 63822 709318
rect 59546 707482 59782 707718
rect 59866 707482 60102 707718
rect 59546 707162 59782 707398
rect 59866 707162 60102 707398
rect 48986 698378 49222 698614
rect 49306 698378 49542 698614
rect 48986 698058 49222 698294
rect 49306 698058 49542 698294
rect 48986 662378 49222 662614
rect 49306 662378 49542 662614
rect 48986 662058 49222 662294
rect 49306 662058 49542 662294
rect 48986 626378 49222 626614
rect 49306 626378 49542 626614
rect 48986 626058 49222 626294
rect 49306 626058 49542 626294
rect 48986 590378 49222 590614
rect 49306 590378 49542 590614
rect 48986 590058 49222 590294
rect 49306 590058 49542 590294
rect 48986 554378 49222 554614
rect 49306 554378 49542 554614
rect 48986 554058 49222 554294
rect 49306 554058 49542 554294
rect 48986 518378 49222 518614
rect 49306 518378 49542 518614
rect 48986 518058 49222 518294
rect 49306 518058 49542 518294
rect 48986 482378 49222 482614
rect 49306 482378 49542 482614
rect 48986 482058 49222 482294
rect 49306 482058 49542 482294
rect 48986 446378 49222 446614
rect 49306 446378 49542 446614
rect 48986 446058 49222 446294
rect 49306 446058 49542 446294
rect 48986 410378 49222 410614
rect 49306 410378 49542 410614
rect 48986 410058 49222 410294
rect 49306 410058 49542 410294
rect 48986 374378 49222 374614
rect 49306 374378 49542 374614
rect 48986 374058 49222 374294
rect 49306 374058 49542 374294
rect 48986 338378 49222 338614
rect 49306 338378 49542 338614
rect 48986 338058 49222 338294
rect 49306 338058 49542 338294
rect 48986 302378 49222 302614
rect 49306 302378 49542 302614
rect 48986 302058 49222 302294
rect 49306 302058 49542 302294
rect 48986 266378 49222 266614
rect 49306 266378 49542 266614
rect 48986 266058 49222 266294
rect 49306 266058 49542 266294
rect 48986 230378 49222 230614
rect 49306 230378 49542 230614
rect 48986 230058 49222 230294
rect 49306 230058 49542 230294
rect 48986 194378 49222 194614
rect 49306 194378 49542 194614
rect 48986 194058 49222 194294
rect 49306 194058 49542 194294
rect 48986 158378 49222 158614
rect 49306 158378 49542 158614
rect 48986 158058 49222 158294
rect 49306 158058 49542 158294
rect 48986 122378 49222 122614
rect 49306 122378 49542 122614
rect 48986 122058 49222 122294
rect 49306 122058 49542 122294
rect 48986 86378 49222 86614
rect 49306 86378 49542 86614
rect 48986 86058 49222 86294
rect 49306 86058 49542 86294
rect 48986 50378 49222 50614
rect 49306 50378 49542 50614
rect 48986 50058 49222 50294
rect 49306 50058 49542 50294
rect 48986 14378 49222 14614
rect 49306 14378 49542 14614
rect 48986 14058 49222 14294
rect 49306 14058 49542 14294
rect 30986 -7302 31222 -7066
rect 31306 -7302 31542 -7066
rect 30986 -7622 31222 -7386
rect 31306 -7622 31542 -7386
rect 55826 705562 56062 705798
rect 56146 705562 56382 705798
rect 55826 705242 56062 705478
rect 56146 705242 56382 705478
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -1542 56062 -1306
rect 56146 -1542 56382 -1306
rect 55826 -1862 56062 -1626
rect 56146 -1862 56382 -1626
rect 59546 672938 59782 673174
rect 59866 672938 60102 673174
rect 59546 672618 59782 672854
rect 59866 672618 60102 672854
rect 59546 636938 59782 637174
rect 59866 636938 60102 637174
rect 59546 636618 59782 636854
rect 59866 636618 60102 636854
rect 59546 600938 59782 601174
rect 59866 600938 60102 601174
rect 59546 600618 59782 600854
rect 59866 600618 60102 600854
rect 59546 564938 59782 565174
rect 59866 564938 60102 565174
rect 59546 564618 59782 564854
rect 59866 564618 60102 564854
rect 59546 528938 59782 529174
rect 59866 528938 60102 529174
rect 59546 528618 59782 528854
rect 59866 528618 60102 528854
rect 59546 492938 59782 493174
rect 59866 492938 60102 493174
rect 59546 492618 59782 492854
rect 59866 492618 60102 492854
rect 59546 456938 59782 457174
rect 59866 456938 60102 457174
rect 59546 456618 59782 456854
rect 59866 456618 60102 456854
rect 59546 420938 59782 421174
rect 59866 420938 60102 421174
rect 59546 420618 59782 420854
rect 59866 420618 60102 420854
rect 59546 384938 59782 385174
rect 59866 384938 60102 385174
rect 59546 384618 59782 384854
rect 59866 384618 60102 384854
rect 59546 348938 59782 349174
rect 59866 348938 60102 349174
rect 59546 348618 59782 348854
rect 59866 348618 60102 348854
rect 59546 312938 59782 313174
rect 59866 312938 60102 313174
rect 59546 312618 59782 312854
rect 59866 312618 60102 312854
rect 59546 276938 59782 277174
rect 59866 276938 60102 277174
rect 59546 276618 59782 276854
rect 59866 276618 60102 276854
rect 59546 240938 59782 241174
rect 59866 240938 60102 241174
rect 59546 240618 59782 240854
rect 59866 240618 60102 240854
rect 59546 204938 59782 205174
rect 59866 204938 60102 205174
rect 59546 204618 59782 204854
rect 59866 204618 60102 204854
rect 59546 168938 59782 169174
rect 59866 168938 60102 169174
rect 59546 168618 59782 168854
rect 59866 168618 60102 168854
rect 59546 132938 59782 133174
rect 59866 132938 60102 133174
rect 59546 132618 59782 132854
rect 59866 132618 60102 132854
rect 59546 96938 59782 97174
rect 59866 96938 60102 97174
rect 59546 96618 59782 96854
rect 59866 96618 60102 96854
rect 59546 60938 59782 61174
rect 59866 60938 60102 61174
rect 59546 60618 59782 60854
rect 59866 60618 60102 60854
rect 59546 24938 59782 25174
rect 59866 24938 60102 25174
rect 59546 24618 59782 24854
rect 59866 24618 60102 24854
rect 59546 -3462 59782 -3226
rect 59866 -3462 60102 -3226
rect 59546 -3782 59782 -3546
rect 59866 -3782 60102 -3546
rect 63266 676658 63502 676894
rect 63586 676658 63822 676894
rect 63266 676338 63502 676574
rect 63586 676338 63822 676574
rect 63266 640658 63502 640894
rect 63586 640658 63822 640894
rect 63266 640338 63502 640574
rect 63586 640338 63822 640574
rect 63266 604658 63502 604894
rect 63586 604658 63822 604894
rect 63266 604338 63502 604574
rect 63586 604338 63822 604574
rect 63266 568658 63502 568894
rect 63586 568658 63822 568894
rect 63266 568338 63502 568574
rect 63586 568338 63822 568574
rect 63266 532658 63502 532894
rect 63586 532658 63822 532894
rect 63266 532338 63502 532574
rect 63586 532338 63822 532574
rect 63266 496658 63502 496894
rect 63586 496658 63822 496894
rect 63266 496338 63502 496574
rect 63586 496338 63822 496574
rect 63266 460658 63502 460894
rect 63586 460658 63822 460894
rect 63266 460338 63502 460574
rect 63586 460338 63822 460574
rect 63266 424658 63502 424894
rect 63586 424658 63822 424894
rect 63266 424338 63502 424574
rect 63586 424338 63822 424574
rect 63266 388658 63502 388894
rect 63586 388658 63822 388894
rect 63266 388338 63502 388574
rect 63586 388338 63822 388574
rect 63266 352658 63502 352894
rect 63586 352658 63822 352894
rect 63266 352338 63502 352574
rect 63586 352338 63822 352574
rect 63266 316658 63502 316894
rect 63586 316658 63822 316894
rect 63266 316338 63502 316574
rect 63586 316338 63822 316574
rect 63266 280658 63502 280894
rect 63586 280658 63822 280894
rect 63266 280338 63502 280574
rect 63586 280338 63822 280574
rect 63266 244658 63502 244894
rect 63586 244658 63822 244894
rect 63266 244338 63502 244574
rect 63586 244338 63822 244574
rect 63266 208658 63502 208894
rect 63586 208658 63822 208894
rect 63266 208338 63502 208574
rect 63586 208338 63822 208574
rect 63266 172658 63502 172894
rect 63586 172658 63822 172894
rect 63266 172338 63502 172574
rect 63586 172338 63822 172574
rect 63266 136658 63502 136894
rect 63586 136658 63822 136894
rect 63266 136338 63502 136574
rect 63586 136338 63822 136574
rect 63266 100658 63502 100894
rect 63586 100658 63822 100894
rect 63266 100338 63502 100574
rect 63586 100338 63822 100574
rect 63266 64658 63502 64894
rect 63586 64658 63822 64894
rect 63266 64338 63502 64574
rect 63586 64338 63822 64574
rect 63266 28658 63502 28894
rect 63586 28658 63822 28894
rect 63266 28338 63502 28574
rect 63586 28338 63822 28574
rect 63266 -5382 63502 -5146
rect 63586 -5382 63822 -5146
rect 63266 -5702 63502 -5466
rect 63586 -5702 63822 -5466
rect 84986 710362 85222 710598
rect 85306 710362 85542 710598
rect 84986 710042 85222 710278
rect 85306 710042 85542 710278
rect 81266 708442 81502 708678
rect 81586 708442 81822 708678
rect 81266 708122 81502 708358
rect 81586 708122 81822 708358
rect 77546 706522 77782 706758
rect 77866 706522 78102 706758
rect 77546 706202 77782 706438
rect 77866 706202 78102 706438
rect 66986 680378 67222 680614
rect 67306 680378 67542 680614
rect 66986 680058 67222 680294
rect 67306 680058 67542 680294
rect 66986 644378 67222 644614
rect 67306 644378 67542 644614
rect 66986 644058 67222 644294
rect 67306 644058 67542 644294
rect 66986 608378 67222 608614
rect 67306 608378 67542 608614
rect 66986 608058 67222 608294
rect 67306 608058 67542 608294
rect 66986 572378 67222 572614
rect 67306 572378 67542 572614
rect 66986 572058 67222 572294
rect 67306 572058 67542 572294
rect 66986 536378 67222 536614
rect 67306 536378 67542 536614
rect 66986 536058 67222 536294
rect 67306 536058 67542 536294
rect 66986 500378 67222 500614
rect 67306 500378 67542 500614
rect 66986 500058 67222 500294
rect 67306 500058 67542 500294
rect 66986 464378 67222 464614
rect 67306 464378 67542 464614
rect 66986 464058 67222 464294
rect 67306 464058 67542 464294
rect 66986 428378 67222 428614
rect 67306 428378 67542 428614
rect 66986 428058 67222 428294
rect 67306 428058 67542 428294
rect 66986 392378 67222 392614
rect 67306 392378 67542 392614
rect 66986 392058 67222 392294
rect 67306 392058 67542 392294
rect 66986 356378 67222 356614
rect 67306 356378 67542 356614
rect 66986 356058 67222 356294
rect 67306 356058 67542 356294
rect 66986 320378 67222 320614
rect 67306 320378 67542 320614
rect 66986 320058 67222 320294
rect 67306 320058 67542 320294
rect 66986 284378 67222 284614
rect 67306 284378 67542 284614
rect 66986 284058 67222 284294
rect 67306 284058 67542 284294
rect 66986 248378 67222 248614
rect 67306 248378 67542 248614
rect 66986 248058 67222 248294
rect 67306 248058 67542 248294
rect 66986 212378 67222 212614
rect 67306 212378 67542 212614
rect 66986 212058 67222 212294
rect 67306 212058 67542 212294
rect 66986 176378 67222 176614
rect 67306 176378 67542 176614
rect 66986 176058 67222 176294
rect 67306 176058 67542 176294
rect 66986 140378 67222 140614
rect 67306 140378 67542 140614
rect 66986 140058 67222 140294
rect 67306 140058 67542 140294
rect 66986 104378 67222 104614
rect 67306 104378 67542 104614
rect 66986 104058 67222 104294
rect 67306 104058 67542 104294
rect 66986 68378 67222 68614
rect 67306 68378 67542 68614
rect 66986 68058 67222 68294
rect 67306 68058 67542 68294
rect 66986 32378 67222 32614
rect 67306 32378 67542 32614
rect 66986 32058 67222 32294
rect 67306 32058 67542 32294
rect 48986 -6342 49222 -6106
rect 49306 -6342 49542 -6106
rect 48986 -6662 49222 -6426
rect 49306 -6662 49542 -6426
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 73826 579218 74062 579454
rect 74146 579218 74382 579454
rect 73826 578898 74062 579134
rect 74146 578898 74382 579134
rect 73826 543218 74062 543454
rect 74146 543218 74382 543454
rect 73826 542898 74062 543134
rect 74146 542898 74382 543134
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 73826 435218 74062 435454
rect 74146 435218 74382 435454
rect 73826 434898 74062 435134
rect 74146 434898 74382 435134
rect 73826 399218 74062 399454
rect 74146 399218 74382 399454
rect 73826 398898 74062 399134
rect 74146 398898 74382 399134
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 73826 327218 74062 327454
rect 74146 327218 74382 327454
rect 73826 326898 74062 327134
rect 74146 326898 74382 327134
rect 73826 291218 74062 291454
rect 74146 291218 74382 291454
rect 73826 290898 74062 291134
rect 74146 290898 74382 291134
rect 73826 255218 74062 255454
rect 74146 255218 74382 255454
rect 73826 254898 74062 255134
rect 74146 254898 74382 255134
rect 73826 219218 74062 219454
rect 74146 219218 74382 219454
rect 73826 218898 74062 219134
rect 74146 218898 74382 219134
rect 73826 183218 74062 183454
rect 74146 183218 74382 183454
rect 73826 182898 74062 183134
rect 74146 182898 74382 183134
rect 73826 147218 74062 147454
rect 74146 147218 74382 147454
rect 73826 146898 74062 147134
rect 74146 146898 74382 147134
rect 73826 111218 74062 111454
rect 74146 111218 74382 111454
rect 73826 110898 74062 111134
rect 74146 110898 74382 111134
rect 73826 75218 74062 75454
rect 74146 75218 74382 75454
rect 73826 74898 74062 75134
rect 74146 74898 74382 75134
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 77546 654938 77782 655174
rect 77866 654938 78102 655174
rect 77546 654618 77782 654854
rect 77866 654618 78102 654854
rect 77546 618938 77782 619174
rect 77866 618938 78102 619174
rect 77546 618618 77782 618854
rect 77866 618618 78102 618854
rect 77546 582938 77782 583174
rect 77866 582938 78102 583174
rect 77546 582618 77782 582854
rect 77866 582618 78102 582854
rect 77546 546938 77782 547174
rect 77866 546938 78102 547174
rect 77546 546618 77782 546854
rect 77866 546618 78102 546854
rect 77546 510938 77782 511174
rect 77866 510938 78102 511174
rect 77546 510618 77782 510854
rect 77866 510618 78102 510854
rect 77546 474938 77782 475174
rect 77866 474938 78102 475174
rect 77546 474618 77782 474854
rect 77866 474618 78102 474854
rect 77546 438938 77782 439174
rect 77866 438938 78102 439174
rect 77546 438618 77782 438854
rect 77866 438618 78102 438854
rect 77546 402938 77782 403174
rect 77866 402938 78102 403174
rect 77546 402618 77782 402854
rect 77866 402618 78102 402854
rect 77546 366938 77782 367174
rect 77866 366938 78102 367174
rect 77546 366618 77782 366854
rect 77866 366618 78102 366854
rect 77546 330938 77782 331174
rect 77866 330938 78102 331174
rect 77546 330618 77782 330854
rect 77866 330618 78102 330854
rect 77546 294938 77782 295174
rect 77866 294938 78102 295174
rect 77546 294618 77782 294854
rect 77866 294618 78102 294854
rect 77546 258938 77782 259174
rect 77866 258938 78102 259174
rect 77546 258618 77782 258854
rect 77866 258618 78102 258854
rect 77546 222938 77782 223174
rect 77866 222938 78102 223174
rect 77546 222618 77782 222854
rect 77866 222618 78102 222854
rect 77546 186938 77782 187174
rect 77866 186938 78102 187174
rect 77546 186618 77782 186854
rect 77866 186618 78102 186854
rect 77546 150938 77782 151174
rect 77866 150938 78102 151174
rect 77546 150618 77782 150854
rect 77866 150618 78102 150854
rect 77546 114938 77782 115174
rect 77866 114938 78102 115174
rect 77546 114618 77782 114854
rect 77866 114618 78102 114854
rect 77546 78938 77782 79174
rect 77866 78938 78102 79174
rect 77546 78618 77782 78854
rect 77866 78618 78102 78854
rect 77546 42938 77782 43174
rect 77866 42938 78102 43174
rect 77546 42618 77782 42854
rect 77866 42618 78102 42854
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 77546 -2502 77782 -2266
rect 77866 -2502 78102 -2266
rect 77546 -2822 77782 -2586
rect 77866 -2822 78102 -2586
rect 81266 694658 81502 694894
rect 81586 694658 81822 694894
rect 81266 694338 81502 694574
rect 81586 694338 81822 694574
rect 81266 658658 81502 658894
rect 81586 658658 81822 658894
rect 81266 658338 81502 658574
rect 81586 658338 81822 658574
rect 81266 622658 81502 622894
rect 81586 622658 81822 622894
rect 81266 622338 81502 622574
rect 81586 622338 81822 622574
rect 81266 586658 81502 586894
rect 81586 586658 81822 586894
rect 81266 586338 81502 586574
rect 81586 586338 81822 586574
rect 81266 550658 81502 550894
rect 81586 550658 81822 550894
rect 81266 550338 81502 550574
rect 81586 550338 81822 550574
rect 81266 514658 81502 514894
rect 81586 514658 81822 514894
rect 81266 514338 81502 514574
rect 81586 514338 81822 514574
rect 81266 478658 81502 478894
rect 81586 478658 81822 478894
rect 81266 478338 81502 478574
rect 81586 478338 81822 478574
rect 81266 442658 81502 442894
rect 81586 442658 81822 442894
rect 81266 442338 81502 442574
rect 81586 442338 81822 442574
rect 81266 406658 81502 406894
rect 81586 406658 81822 406894
rect 81266 406338 81502 406574
rect 81586 406338 81822 406574
rect 81266 370658 81502 370894
rect 81586 370658 81822 370894
rect 81266 370338 81502 370574
rect 81586 370338 81822 370574
rect 81266 334658 81502 334894
rect 81586 334658 81822 334894
rect 81266 334338 81502 334574
rect 81586 334338 81822 334574
rect 81266 298658 81502 298894
rect 81586 298658 81822 298894
rect 81266 298338 81502 298574
rect 81586 298338 81822 298574
rect 81266 262658 81502 262894
rect 81586 262658 81822 262894
rect 81266 262338 81502 262574
rect 81586 262338 81822 262574
rect 81266 226658 81502 226894
rect 81586 226658 81822 226894
rect 81266 226338 81502 226574
rect 81586 226338 81822 226574
rect 81266 190658 81502 190894
rect 81586 190658 81822 190894
rect 81266 190338 81502 190574
rect 81586 190338 81822 190574
rect 81266 154658 81502 154894
rect 81586 154658 81822 154894
rect 81266 154338 81502 154574
rect 81586 154338 81822 154574
rect 81266 118658 81502 118894
rect 81586 118658 81822 118894
rect 81266 118338 81502 118574
rect 81586 118338 81822 118574
rect 81266 82658 81502 82894
rect 81586 82658 81822 82894
rect 81266 82338 81502 82574
rect 81586 82338 81822 82574
rect 81266 46658 81502 46894
rect 81586 46658 81822 46894
rect 81266 46338 81502 46574
rect 81586 46338 81822 46574
rect 81266 10658 81502 10894
rect 81586 10658 81822 10894
rect 81266 10338 81502 10574
rect 81586 10338 81822 10574
rect 81266 -4422 81502 -4186
rect 81586 -4422 81822 -4186
rect 81266 -4742 81502 -4506
rect 81586 -4742 81822 -4506
rect 102986 711322 103222 711558
rect 103306 711322 103542 711558
rect 102986 711002 103222 711238
rect 103306 711002 103542 711238
rect 99266 709402 99502 709638
rect 99586 709402 99822 709638
rect 99266 709082 99502 709318
rect 99586 709082 99822 709318
rect 95546 707482 95782 707718
rect 95866 707482 96102 707718
rect 95546 707162 95782 707398
rect 95866 707162 96102 707398
rect 84986 698378 85222 698614
rect 85306 698378 85542 698614
rect 84986 698058 85222 698294
rect 85306 698058 85542 698294
rect 84986 662378 85222 662614
rect 85306 662378 85542 662614
rect 84986 662058 85222 662294
rect 85306 662058 85542 662294
rect 84986 626378 85222 626614
rect 85306 626378 85542 626614
rect 84986 626058 85222 626294
rect 85306 626058 85542 626294
rect 84986 590378 85222 590614
rect 85306 590378 85542 590614
rect 84986 590058 85222 590294
rect 85306 590058 85542 590294
rect 84986 554378 85222 554614
rect 85306 554378 85542 554614
rect 84986 554058 85222 554294
rect 85306 554058 85542 554294
rect 84986 518378 85222 518614
rect 85306 518378 85542 518614
rect 84986 518058 85222 518294
rect 85306 518058 85542 518294
rect 84986 482378 85222 482614
rect 85306 482378 85542 482614
rect 84986 482058 85222 482294
rect 85306 482058 85542 482294
rect 84986 446378 85222 446614
rect 85306 446378 85542 446614
rect 84986 446058 85222 446294
rect 85306 446058 85542 446294
rect 84986 410378 85222 410614
rect 85306 410378 85542 410614
rect 84986 410058 85222 410294
rect 85306 410058 85542 410294
rect 84986 374378 85222 374614
rect 85306 374378 85542 374614
rect 84986 374058 85222 374294
rect 85306 374058 85542 374294
rect 84986 338378 85222 338614
rect 85306 338378 85542 338614
rect 84986 338058 85222 338294
rect 85306 338058 85542 338294
rect 84986 302378 85222 302614
rect 85306 302378 85542 302614
rect 84986 302058 85222 302294
rect 85306 302058 85542 302294
rect 84986 266378 85222 266614
rect 85306 266378 85542 266614
rect 84986 266058 85222 266294
rect 85306 266058 85542 266294
rect 84986 230378 85222 230614
rect 85306 230378 85542 230614
rect 84986 230058 85222 230294
rect 85306 230058 85542 230294
rect 84986 194378 85222 194614
rect 85306 194378 85542 194614
rect 84986 194058 85222 194294
rect 85306 194058 85542 194294
rect 84986 158378 85222 158614
rect 85306 158378 85542 158614
rect 84986 158058 85222 158294
rect 85306 158058 85542 158294
rect 84986 122378 85222 122614
rect 85306 122378 85542 122614
rect 84986 122058 85222 122294
rect 85306 122058 85542 122294
rect 84986 86378 85222 86614
rect 85306 86378 85542 86614
rect 84986 86058 85222 86294
rect 85306 86058 85542 86294
rect 84986 50378 85222 50614
rect 85306 50378 85542 50614
rect 84986 50058 85222 50294
rect 85306 50058 85542 50294
rect 84986 14378 85222 14614
rect 85306 14378 85542 14614
rect 84986 14058 85222 14294
rect 85306 14058 85542 14294
rect 66986 -7302 67222 -7066
rect 67306 -7302 67542 -7066
rect 66986 -7622 67222 -7386
rect 67306 -7622 67542 -7386
rect 91826 705562 92062 705798
rect 92146 705562 92382 705798
rect 91826 705242 92062 705478
rect 92146 705242 92382 705478
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 91826 561218 92062 561454
rect 92146 561218 92382 561454
rect 91826 560898 92062 561134
rect 92146 560898 92382 561134
rect 91826 525218 92062 525454
rect 92146 525218 92382 525454
rect 91826 524898 92062 525134
rect 92146 524898 92382 525134
rect 91826 489218 92062 489454
rect 92146 489218 92382 489454
rect 91826 488898 92062 489134
rect 92146 488898 92382 489134
rect 91826 453218 92062 453454
rect 92146 453218 92382 453454
rect 91826 452898 92062 453134
rect 92146 452898 92382 453134
rect 91826 417218 92062 417454
rect 92146 417218 92382 417454
rect 91826 416898 92062 417134
rect 92146 416898 92382 417134
rect 91826 381218 92062 381454
rect 92146 381218 92382 381454
rect 91826 380898 92062 381134
rect 92146 380898 92382 381134
rect 91826 345218 92062 345454
rect 92146 345218 92382 345454
rect 91826 344898 92062 345134
rect 92146 344898 92382 345134
rect 91826 309218 92062 309454
rect 92146 309218 92382 309454
rect 91826 308898 92062 309134
rect 92146 308898 92382 309134
rect 91826 273218 92062 273454
rect 92146 273218 92382 273454
rect 91826 272898 92062 273134
rect 92146 272898 92382 273134
rect 91826 237218 92062 237454
rect 92146 237218 92382 237454
rect 91826 236898 92062 237134
rect 92146 236898 92382 237134
rect 91826 201218 92062 201454
rect 92146 201218 92382 201454
rect 91826 200898 92062 201134
rect 92146 200898 92382 201134
rect 91826 165218 92062 165454
rect 92146 165218 92382 165454
rect 91826 164898 92062 165134
rect 92146 164898 92382 165134
rect 91826 129218 92062 129454
rect 92146 129218 92382 129454
rect 91826 128898 92062 129134
rect 92146 128898 92382 129134
rect 91826 93218 92062 93454
rect 92146 93218 92382 93454
rect 91826 92898 92062 93134
rect 92146 92898 92382 93134
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -1542 92062 -1306
rect 92146 -1542 92382 -1306
rect 91826 -1862 92062 -1626
rect 92146 -1862 92382 -1626
rect 95546 672938 95782 673174
rect 95866 672938 96102 673174
rect 95546 672618 95782 672854
rect 95866 672618 96102 672854
rect 95546 636938 95782 637174
rect 95866 636938 96102 637174
rect 95546 636618 95782 636854
rect 95866 636618 96102 636854
rect 95546 600938 95782 601174
rect 95866 600938 96102 601174
rect 95546 600618 95782 600854
rect 95866 600618 96102 600854
rect 95546 564938 95782 565174
rect 95866 564938 96102 565174
rect 95546 564618 95782 564854
rect 95866 564618 96102 564854
rect 95546 528938 95782 529174
rect 95866 528938 96102 529174
rect 95546 528618 95782 528854
rect 95866 528618 96102 528854
rect 95546 492938 95782 493174
rect 95866 492938 96102 493174
rect 95546 492618 95782 492854
rect 95866 492618 96102 492854
rect 95546 456938 95782 457174
rect 95866 456938 96102 457174
rect 95546 456618 95782 456854
rect 95866 456618 96102 456854
rect 95546 420938 95782 421174
rect 95866 420938 96102 421174
rect 95546 420618 95782 420854
rect 95866 420618 96102 420854
rect 95546 384938 95782 385174
rect 95866 384938 96102 385174
rect 95546 384618 95782 384854
rect 95866 384618 96102 384854
rect 95546 348938 95782 349174
rect 95866 348938 96102 349174
rect 95546 348618 95782 348854
rect 95866 348618 96102 348854
rect 95546 312938 95782 313174
rect 95866 312938 96102 313174
rect 95546 312618 95782 312854
rect 95866 312618 96102 312854
rect 95546 276938 95782 277174
rect 95866 276938 96102 277174
rect 95546 276618 95782 276854
rect 95866 276618 96102 276854
rect 95546 240938 95782 241174
rect 95866 240938 96102 241174
rect 95546 240618 95782 240854
rect 95866 240618 96102 240854
rect 95546 204938 95782 205174
rect 95866 204938 96102 205174
rect 95546 204618 95782 204854
rect 95866 204618 96102 204854
rect 95546 168938 95782 169174
rect 95866 168938 96102 169174
rect 95546 168618 95782 168854
rect 95866 168618 96102 168854
rect 95546 132938 95782 133174
rect 95866 132938 96102 133174
rect 95546 132618 95782 132854
rect 95866 132618 96102 132854
rect 95546 96938 95782 97174
rect 95866 96938 96102 97174
rect 95546 96618 95782 96854
rect 95866 96618 96102 96854
rect 95546 60938 95782 61174
rect 95866 60938 96102 61174
rect 95546 60618 95782 60854
rect 95866 60618 96102 60854
rect 95546 24938 95782 25174
rect 95866 24938 96102 25174
rect 95546 24618 95782 24854
rect 95866 24618 96102 24854
rect 95546 -3462 95782 -3226
rect 95866 -3462 96102 -3226
rect 95546 -3782 95782 -3546
rect 95866 -3782 96102 -3546
rect 99266 676658 99502 676894
rect 99586 676658 99822 676894
rect 99266 676338 99502 676574
rect 99586 676338 99822 676574
rect 99266 640658 99502 640894
rect 99586 640658 99822 640894
rect 99266 640338 99502 640574
rect 99586 640338 99822 640574
rect 99266 604658 99502 604894
rect 99586 604658 99822 604894
rect 99266 604338 99502 604574
rect 99586 604338 99822 604574
rect 99266 568658 99502 568894
rect 99586 568658 99822 568894
rect 99266 568338 99502 568574
rect 99586 568338 99822 568574
rect 99266 532658 99502 532894
rect 99586 532658 99822 532894
rect 99266 532338 99502 532574
rect 99586 532338 99822 532574
rect 99266 496658 99502 496894
rect 99586 496658 99822 496894
rect 99266 496338 99502 496574
rect 99586 496338 99822 496574
rect 99266 460658 99502 460894
rect 99586 460658 99822 460894
rect 99266 460338 99502 460574
rect 99586 460338 99822 460574
rect 99266 424658 99502 424894
rect 99586 424658 99822 424894
rect 99266 424338 99502 424574
rect 99586 424338 99822 424574
rect 99266 388658 99502 388894
rect 99586 388658 99822 388894
rect 99266 388338 99502 388574
rect 99586 388338 99822 388574
rect 99266 352658 99502 352894
rect 99586 352658 99822 352894
rect 99266 352338 99502 352574
rect 99586 352338 99822 352574
rect 99266 316658 99502 316894
rect 99586 316658 99822 316894
rect 99266 316338 99502 316574
rect 99586 316338 99822 316574
rect 99266 280658 99502 280894
rect 99586 280658 99822 280894
rect 99266 280338 99502 280574
rect 99586 280338 99822 280574
rect 99266 244658 99502 244894
rect 99586 244658 99822 244894
rect 99266 244338 99502 244574
rect 99586 244338 99822 244574
rect 99266 208658 99502 208894
rect 99586 208658 99822 208894
rect 99266 208338 99502 208574
rect 99586 208338 99822 208574
rect 99266 172658 99502 172894
rect 99586 172658 99822 172894
rect 99266 172338 99502 172574
rect 99586 172338 99822 172574
rect 99266 136658 99502 136894
rect 99586 136658 99822 136894
rect 99266 136338 99502 136574
rect 99586 136338 99822 136574
rect 99266 100658 99502 100894
rect 99586 100658 99822 100894
rect 99266 100338 99502 100574
rect 99586 100338 99822 100574
rect 99266 64658 99502 64894
rect 99586 64658 99822 64894
rect 99266 64338 99502 64574
rect 99586 64338 99822 64574
rect 99266 28658 99502 28894
rect 99586 28658 99822 28894
rect 99266 28338 99502 28574
rect 99586 28338 99822 28574
rect 99266 -5382 99502 -5146
rect 99586 -5382 99822 -5146
rect 99266 -5702 99502 -5466
rect 99586 -5702 99822 -5466
rect 120986 710362 121222 710598
rect 121306 710362 121542 710598
rect 120986 710042 121222 710278
rect 121306 710042 121542 710278
rect 117266 708442 117502 708678
rect 117586 708442 117822 708678
rect 117266 708122 117502 708358
rect 117586 708122 117822 708358
rect 113546 706522 113782 706758
rect 113866 706522 114102 706758
rect 113546 706202 113782 706438
rect 113866 706202 114102 706438
rect 102986 680378 103222 680614
rect 103306 680378 103542 680614
rect 102986 680058 103222 680294
rect 103306 680058 103542 680294
rect 102986 644378 103222 644614
rect 103306 644378 103542 644614
rect 102986 644058 103222 644294
rect 103306 644058 103542 644294
rect 102986 608378 103222 608614
rect 103306 608378 103542 608614
rect 102986 608058 103222 608294
rect 103306 608058 103542 608294
rect 102986 572378 103222 572614
rect 103306 572378 103542 572614
rect 102986 572058 103222 572294
rect 103306 572058 103542 572294
rect 102986 536378 103222 536614
rect 103306 536378 103542 536614
rect 102986 536058 103222 536294
rect 103306 536058 103542 536294
rect 102986 500378 103222 500614
rect 103306 500378 103542 500614
rect 102986 500058 103222 500294
rect 103306 500058 103542 500294
rect 102986 464378 103222 464614
rect 103306 464378 103542 464614
rect 102986 464058 103222 464294
rect 103306 464058 103542 464294
rect 102986 428378 103222 428614
rect 103306 428378 103542 428614
rect 102986 428058 103222 428294
rect 103306 428058 103542 428294
rect 102986 392378 103222 392614
rect 103306 392378 103542 392614
rect 102986 392058 103222 392294
rect 103306 392058 103542 392294
rect 102986 356378 103222 356614
rect 103306 356378 103542 356614
rect 102986 356058 103222 356294
rect 103306 356058 103542 356294
rect 102986 320378 103222 320614
rect 103306 320378 103542 320614
rect 102986 320058 103222 320294
rect 103306 320058 103542 320294
rect 102986 284378 103222 284614
rect 103306 284378 103542 284614
rect 102986 284058 103222 284294
rect 103306 284058 103542 284294
rect 102986 248378 103222 248614
rect 103306 248378 103542 248614
rect 102986 248058 103222 248294
rect 103306 248058 103542 248294
rect 102986 212378 103222 212614
rect 103306 212378 103542 212614
rect 102986 212058 103222 212294
rect 103306 212058 103542 212294
rect 102986 176378 103222 176614
rect 103306 176378 103542 176614
rect 102986 176058 103222 176294
rect 103306 176058 103542 176294
rect 102986 140378 103222 140614
rect 103306 140378 103542 140614
rect 102986 140058 103222 140294
rect 103306 140058 103542 140294
rect 102986 104378 103222 104614
rect 103306 104378 103542 104614
rect 102986 104058 103222 104294
rect 103306 104058 103542 104294
rect 102986 68378 103222 68614
rect 103306 68378 103542 68614
rect 102986 68058 103222 68294
rect 103306 68058 103542 68294
rect 102986 32378 103222 32614
rect 103306 32378 103542 32614
rect 102986 32058 103222 32294
rect 103306 32058 103542 32294
rect 84986 -6342 85222 -6106
rect 85306 -6342 85542 -6106
rect 84986 -6662 85222 -6426
rect 85306 -6662 85542 -6426
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 109826 507218 110062 507454
rect 110146 507218 110382 507454
rect 109826 506898 110062 507134
rect 110146 506898 110382 507134
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 109826 435218 110062 435454
rect 110146 435218 110382 435454
rect 109826 434898 110062 435134
rect 110146 434898 110382 435134
rect 109826 399218 110062 399454
rect 110146 399218 110382 399454
rect 109826 398898 110062 399134
rect 110146 398898 110382 399134
rect 109826 363218 110062 363454
rect 110146 363218 110382 363454
rect 109826 362898 110062 363134
rect 110146 362898 110382 363134
rect 109826 327218 110062 327454
rect 110146 327218 110382 327454
rect 109826 326898 110062 327134
rect 110146 326898 110382 327134
rect 109826 291218 110062 291454
rect 110146 291218 110382 291454
rect 109826 290898 110062 291134
rect 110146 290898 110382 291134
rect 109826 255218 110062 255454
rect 110146 255218 110382 255454
rect 109826 254898 110062 255134
rect 110146 254898 110382 255134
rect 109826 219218 110062 219454
rect 110146 219218 110382 219454
rect 109826 218898 110062 219134
rect 110146 218898 110382 219134
rect 109826 183218 110062 183454
rect 110146 183218 110382 183454
rect 109826 182898 110062 183134
rect 110146 182898 110382 183134
rect 109826 147218 110062 147454
rect 110146 147218 110382 147454
rect 109826 146898 110062 147134
rect 110146 146898 110382 147134
rect 109826 111218 110062 111454
rect 110146 111218 110382 111454
rect 109826 110898 110062 111134
rect 110146 110898 110382 111134
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 690938 113782 691174
rect 113866 690938 114102 691174
rect 113546 690618 113782 690854
rect 113866 690618 114102 690854
rect 113546 654938 113782 655174
rect 113866 654938 114102 655174
rect 113546 654618 113782 654854
rect 113866 654618 114102 654854
rect 113546 618938 113782 619174
rect 113866 618938 114102 619174
rect 113546 618618 113782 618854
rect 113866 618618 114102 618854
rect 113546 582938 113782 583174
rect 113866 582938 114102 583174
rect 113546 582618 113782 582854
rect 113866 582618 114102 582854
rect 113546 546938 113782 547174
rect 113866 546938 114102 547174
rect 113546 546618 113782 546854
rect 113866 546618 114102 546854
rect 113546 510938 113782 511174
rect 113866 510938 114102 511174
rect 113546 510618 113782 510854
rect 113866 510618 114102 510854
rect 113546 474938 113782 475174
rect 113866 474938 114102 475174
rect 113546 474618 113782 474854
rect 113866 474618 114102 474854
rect 113546 438938 113782 439174
rect 113866 438938 114102 439174
rect 113546 438618 113782 438854
rect 113866 438618 114102 438854
rect 113546 402938 113782 403174
rect 113866 402938 114102 403174
rect 113546 402618 113782 402854
rect 113866 402618 114102 402854
rect 113546 366938 113782 367174
rect 113866 366938 114102 367174
rect 113546 366618 113782 366854
rect 113866 366618 114102 366854
rect 113546 330938 113782 331174
rect 113866 330938 114102 331174
rect 113546 330618 113782 330854
rect 113866 330618 114102 330854
rect 113546 294938 113782 295174
rect 113866 294938 114102 295174
rect 113546 294618 113782 294854
rect 113866 294618 114102 294854
rect 113546 258938 113782 259174
rect 113866 258938 114102 259174
rect 113546 258618 113782 258854
rect 113866 258618 114102 258854
rect 113546 222938 113782 223174
rect 113866 222938 114102 223174
rect 113546 222618 113782 222854
rect 113866 222618 114102 222854
rect 113546 186938 113782 187174
rect 113866 186938 114102 187174
rect 113546 186618 113782 186854
rect 113866 186618 114102 186854
rect 113546 150938 113782 151174
rect 113866 150938 114102 151174
rect 113546 150618 113782 150854
rect 113866 150618 114102 150854
rect 113546 114938 113782 115174
rect 113866 114938 114102 115174
rect 113546 114618 113782 114854
rect 113866 114618 114102 114854
rect 113546 78938 113782 79174
rect 113866 78938 114102 79174
rect 113546 78618 113782 78854
rect 113866 78618 114102 78854
rect 113546 42938 113782 43174
rect 113866 42938 114102 43174
rect 113546 42618 113782 42854
rect 113866 42618 114102 42854
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 113546 -2502 113782 -2266
rect 113866 -2502 114102 -2266
rect 113546 -2822 113782 -2586
rect 113866 -2822 114102 -2586
rect 117266 694658 117502 694894
rect 117586 694658 117822 694894
rect 117266 694338 117502 694574
rect 117586 694338 117822 694574
rect 117266 658658 117502 658894
rect 117586 658658 117822 658894
rect 117266 658338 117502 658574
rect 117586 658338 117822 658574
rect 117266 622658 117502 622894
rect 117586 622658 117822 622894
rect 117266 622338 117502 622574
rect 117586 622338 117822 622574
rect 117266 586658 117502 586894
rect 117586 586658 117822 586894
rect 117266 586338 117502 586574
rect 117586 586338 117822 586574
rect 117266 550658 117502 550894
rect 117586 550658 117822 550894
rect 117266 550338 117502 550574
rect 117586 550338 117822 550574
rect 117266 514658 117502 514894
rect 117586 514658 117822 514894
rect 117266 514338 117502 514574
rect 117586 514338 117822 514574
rect 117266 478658 117502 478894
rect 117586 478658 117822 478894
rect 117266 478338 117502 478574
rect 117586 478338 117822 478574
rect 117266 442658 117502 442894
rect 117586 442658 117822 442894
rect 117266 442338 117502 442574
rect 117586 442338 117822 442574
rect 117266 406658 117502 406894
rect 117586 406658 117822 406894
rect 117266 406338 117502 406574
rect 117586 406338 117822 406574
rect 117266 370658 117502 370894
rect 117586 370658 117822 370894
rect 117266 370338 117502 370574
rect 117586 370338 117822 370574
rect 117266 334658 117502 334894
rect 117586 334658 117822 334894
rect 117266 334338 117502 334574
rect 117586 334338 117822 334574
rect 117266 298658 117502 298894
rect 117586 298658 117822 298894
rect 117266 298338 117502 298574
rect 117586 298338 117822 298574
rect 117266 262658 117502 262894
rect 117586 262658 117822 262894
rect 117266 262338 117502 262574
rect 117586 262338 117822 262574
rect 117266 226658 117502 226894
rect 117586 226658 117822 226894
rect 117266 226338 117502 226574
rect 117586 226338 117822 226574
rect 117266 190658 117502 190894
rect 117586 190658 117822 190894
rect 117266 190338 117502 190574
rect 117586 190338 117822 190574
rect 117266 154658 117502 154894
rect 117586 154658 117822 154894
rect 117266 154338 117502 154574
rect 117586 154338 117822 154574
rect 117266 118658 117502 118894
rect 117586 118658 117822 118894
rect 117266 118338 117502 118574
rect 117586 118338 117822 118574
rect 117266 82658 117502 82894
rect 117586 82658 117822 82894
rect 117266 82338 117502 82574
rect 117586 82338 117822 82574
rect 117266 46658 117502 46894
rect 117586 46658 117822 46894
rect 117266 46338 117502 46574
rect 117586 46338 117822 46574
rect 117266 10658 117502 10894
rect 117586 10658 117822 10894
rect 117266 10338 117502 10574
rect 117586 10338 117822 10574
rect 117266 -4422 117502 -4186
rect 117586 -4422 117822 -4186
rect 117266 -4742 117502 -4506
rect 117586 -4742 117822 -4506
rect 138986 711322 139222 711558
rect 139306 711322 139542 711558
rect 138986 711002 139222 711238
rect 139306 711002 139542 711238
rect 135266 709402 135502 709638
rect 135586 709402 135822 709638
rect 135266 709082 135502 709318
rect 135586 709082 135822 709318
rect 131546 707482 131782 707718
rect 131866 707482 132102 707718
rect 131546 707162 131782 707398
rect 131866 707162 132102 707398
rect 120986 698378 121222 698614
rect 121306 698378 121542 698614
rect 120986 698058 121222 698294
rect 121306 698058 121542 698294
rect 120986 662378 121222 662614
rect 121306 662378 121542 662614
rect 120986 662058 121222 662294
rect 121306 662058 121542 662294
rect 120986 626378 121222 626614
rect 121306 626378 121542 626614
rect 120986 626058 121222 626294
rect 121306 626058 121542 626294
rect 120986 590378 121222 590614
rect 121306 590378 121542 590614
rect 120986 590058 121222 590294
rect 121306 590058 121542 590294
rect 120986 554378 121222 554614
rect 121306 554378 121542 554614
rect 120986 554058 121222 554294
rect 121306 554058 121542 554294
rect 120986 518378 121222 518614
rect 121306 518378 121542 518614
rect 120986 518058 121222 518294
rect 121306 518058 121542 518294
rect 120986 482378 121222 482614
rect 121306 482378 121542 482614
rect 120986 482058 121222 482294
rect 121306 482058 121542 482294
rect 120986 446378 121222 446614
rect 121306 446378 121542 446614
rect 120986 446058 121222 446294
rect 121306 446058 121542 446294
rect 120986 410378 121222 410614
rect 121306 410378 121542 410614
rect 120986 410058 121222 410294
rect 121306 410058 121542 410294
rect 120986 374378 121222 374614
rect 121306 374378 121542 374614
rect 120986 374058 121222 374294
rect 121306 374058 121542 374294
rect 120986 338378 121222 338614
rect 121306 338378 121542 338614
rect 120986 338058 121222 338294
rect 121306 338058 121542 338294
rect 120986 302378 121222 302614
rect 121306 302378 121542 302614
rect 120986 302058 121222 302294
rect 121306 302058 121542 302294
rect 120986 266378 121222 266614
rect 121306 266378 121542 266614
rect 120986 266058 121222 266294
rect 121306 266058 121542 266294
rect 120986 230378 121222 230614
rect 121306 230378 121542 230614
rect 120986 230058 121222 230294
rect 121306 230058 121542 230294
rect 120986 194378 121222 194614
rect 121306 194378 121542 194614
rect 120986 194058 121222 194294
rect 121306 194058 121542 194294
rect 120986 158378 121222 158614
rect 121306 158378 121542 158614
rect 120986 158058 121222 158294
rect 121306 158058 121542 158294
rect 120986 122378 121222 122614
rect 121306 122378 121542 122614
rect 120986 122058 121222 122294
rect 121306 122058 121542 122294
rect 120986 86378 121222 86614
rect 121306 86378 121542 86614
rect 120986 86058 121222 86294
rect 121306 86058 121542 86294
rect 120986 50378 121222 50614
rect 121306 50378 121542 50614
rect 120986 50058 121222 50294
rect 121306 50058 121542 50294
rect 120986 14378 121222 14614
rect 121306 14378 121542 14614
rect 120986 14058 121222 14294
rect 121306 14058 121542 14294
rect 102986 -7302 103222 -7066
rect 103306 -7302 103542 -7066
rect 102986 -7622 103222 -7386
rect 103306 -7622 103542 -7386
rect 127826 705562 128062 705798
rect 128146 705562 128382 705798
rect 127826 705242 128062 705478
rect 128146 705242 128382 705478
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 127826 561218 128062 561454
rect 128146 561218 128382 561454
rect 127826 560898 128062 561134
rect 128146 560898 128382 561134
rect 127826 525218 128062 525454
rect 128146 525218 128382 525454
rect 127826 524898 128062 525134
rect 128146 524898 128382 525134
rect 127826 489218 128062 489454
rect 128146 489218 128382 489454
rect 127826 488898 128062 489134
rect 128146 488898 128382 489134
rect 127826 453218 128062 453454
rect 128146 453218 128382 453454
rect 127826 452898 128062 453134
rect 128146 452898 128382 453134
rect 127826 417218 128062 417454
rect 128146 417218 128382 417454
rect 127826 416898 128062 417134
rect 128146 416898 128382 417134
rect 127826 381218 128062 381454
rect 128146 381218 128382 381454
rect 127826 380898 128062 381134
rect 128146 380898 128382 381134
rect 127826 345218 128062 345454
rect 128146 345218 128382 345454
rect 127826 344898 128062 345134
rect 128146 344898 128382 345134
rect 127826 309218 128062 309454
rect 128146 309218 128382 309454
rect 127826 308898 128062 309134
rect 128146 308898 128382 309134
rect 127826 273218 128062 273454
rect 128146 273218 128382 273454
rect 127826 272898 128062 273134
rect 128146 272898 128382 273134
rect 127826 237218 128062 237454
rect 128146 237218 128382 237454
rect 127826 236898 128062 237134
rect 128146 236898 128382 237134
rect 127826 201218 128062 201454
rect 128146 201218 128382 201454
rect 127826 200898 128062 201134
rect 128146 200898 128382 201134
rect 127826 165218 128062 165454
rect 128146 165218 128382 165454
rect 127826 164898 128062 165134
rect 128146 164898 128382 165134
rect 127826 129218 128062 129454
rect 128146 129218 128382 129454
rect 127826 128898 128062 129134
rect 128146 128898 128382 129134
rect 127826 93218 128062 93454
rect 128146 93218 128382 93454
rect 127826 92898 128062 93134
rect 128146 92898 128382 93134
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -1542 128062 -1306
rect 128146 -1542 128382 -1306
rect 127826 -1862 128062 -1626
rect 128146 -1862 128382 -1626
rect 131546 672938 131782 673174
rect 131866 672938 132102 673174
rect 131546 672618 131782 672854
rect 131866 672618 132102 672854
rect 131546 636938 131782 637174
rect 131866 636938 132102 637174
rect 131546 636618 131782 636854
rect 131866 636618 132102 636854
rect 131546 600938 131782 601174
rect 131866 600938 132102 601174
rect 131546 600618 131782 600854
rect 131866 600618 132102 600854
rect 131546 564938 131782 565174
rect 131866 564938 132102 565174
rect 131546 564618 131782 564854
rect 131866 564618 132102 564854
rect 131546 528938 131782 529174
rect 131866 528938 132102 529174
rect 131546 528618 131782 528854
rect 131866 528618 132102 528854
rect 131546 492938 131782 493174
rect 131866 492938 132102 493174
rect 131546 492618 131782 492854
rect 131866 492618 132102 492854
rect 131546 456938 131782 457174
rect 131866 456938 132102 457174
rect 131546 456618 131782 456854
rect 131866 456618 132102 456854
rect 131546 420938 131782 421174
rect 131866 420938 132102 421174
rect 131546 420618 131782 420854
rect 131866 420618 132102 420854
rect 131546 384938 131782 385174
rect 131866 384938 132102 385174
rect 131546 384618 131782 384854
rect 131866 384618 132102 384854
rect 131546 348938 131782 349174
rect 131866 348938 132102 349174
rect 131546 348618 131782 348854
rect 131866 348618 132102 348854
rect 131546 312938 131782 313174
rect 131866 312938 132102 313174
rect 131546 312618 131782 312854
rect 131866 312618 132102 312854
rect 131546 276938 131782 277174
rect 131866 276938 132102 277174
rect 131546 276618 131782 276854
rect 131866 276618 132102 276854
rect 131546 240938 131782 241174
rect 131866 240938 132102 241174
rect 131546 240618 131782 240854
rect 131866 240618 132102 240854
rect 131546 204938 131782 205174
rect 131866 204938 132102 205174
rect 131546 204618 131782 204854
rect 131866 204618 132102 204854
rect 131546 168938 131782 169174
rect 131866 168938 132102 169174
rect 131546 168618 131782 168854
rect 131866 168618 132102 168854
rect 131546 132938 131782 133174
rect 131866 132938 132102 133174
rect 131546 132618 131782 132854
rect 131866 132618 132102 132854
rect 131546 96938 131782 97174
rect 131866 96938 132102 97174
rect 131546 96618 131782 96854
rect 131866 96618 132102 96854
rect 131546 60938 131782 61174
rect 131866 60938 132102 61174
rect 131546 60618 131782 60854
rect 131866 60618 132102 60854
rect 131546 24938 131782 25174
rect 131866 24938 132102 25174
rect 131546 24618 131782 24854
rect 131866 24618 132102 24854
rect 131546 -3462 131782 -3226
rect 131866 -3462 132102 -3226
rect 131546 -3782 131782 -3546
rect 131866 -3782 132102 -3546
rect 135266 676658 135502 676894
rect 135586 676658 135822 676894
rect 135266 676338 135502 676574
rect 135586 676338 135822 676574
rect 135266 640658 135502 640894
rect 135586 640658 135822 640894
rect 135266 640338 135502 640574
rect 135586 640338 135822 640574
rect 135266 604658 135502 604894
rect 135586 604658 135822 604894
rect 135266 604338 135502 604574
rect 135586 604338 135822 604574
rect 135266 568658 135502 568894
rect 135586 568658 135822 568894
rect 135266 568338 135502 568574
rect 135586 568338 135822 568574
rect 135266 532658 135502 532894
rect 135586 532658 135822 532894
rect 135266 532338 135502 532574
rect 135586 532338 135822 532574
rect 135266 496658 135502 496894
rect 135586 496658 135822 496894
rect 135266 496338 135502 496574
rect 135586 496338 135822 496574
rect 135266 460658 135502 460894
rect 135586 460658 135822 460894
rect 135266 460338 135502 460574
rect 135586 460338 135822 460574
rect 135266 424658 135502 424894
rect 135586 424658 135822 424894
rect 135266 424338 135502 424574
rect 135586 424338 135822 424574
rect 135266 388658 135502 388894
rect 135586 388658 135822 388894
rect 135266 388338 135502 388574
rect 135586 388338 135822 388574
rect 135266 352658 135502 352894
rect 135586 352658 135822 352894
rect 135266 352338 135502 352574
rect 135586 352338 135822 352574
rect 135266 316658 135502 316894
rect 135586 316658 135822 316894
rect 135266 316338 135502 316574
rect 135586 316338 135822 316574
rect 135266 280658 135502 280894
rect 135586 280658 135822 280894
rect 135266 280338 135502 280574
rect 135586 280338 135822 280574
rect 135266 244658 135502 244894
rect 135586 244658 135822 244894
rect 135266 244338 135502 244574
rect 135586 244338 135822 244574
rect 135266 208658 135502 208894
rect 135586 208658 135822 208894
rect 135266 208338 135502 208574
rect 135586 208338 135822 208574
rect 135266 172658 135502 172894
rect 135586 172658 135822 172894
rect 135266 172338 135502 172574
rect 135586 172338 135822 172574
rect 135266 136658 135502 136894
rect 135586 136658 135822 136894
rect 135266 136338 135502 136574
rect 135586 136338 135822 136574
rect 135266 100658 135502 100894
rect 135586 100658 135822 100894
rect 135266 100338 135502 100574
rect 135586 100338 135822 100574
rect 135266 64658 135502 64894
rect 135586 64658 135822 64894
rect 135266 64338 135502 64574
rect 135586 64338 135822 64574
rect 135266 28658 135502 28894
rect 135586 28658 135822 28894
rect 135266 28338 135502 28574
rect 135586 28338 135822 28574
rect 135266 -5382 135502 -5146
rect 135586 -5382 135822 -5146
rect 135266 -5702 135502 -5466
rect 135586 -5702 135822 -5466
rect 156986 710362 157222 710598
rect 157306 710362 157542 710598
rect 156986 710042 157222 710278
rect 157306 710042 157542 710278
rect 153266 708442 153502 708678
rect 153586 708442 153822 708678
rect 153266 708122 153502 708358
rect 153586 708122 153822 708358
rect 149546 706522 149782 706758
rect 149866 706522 150102 706758
rect 149546 706202 149782 706438
rect 149866 706202 150102 706438
rect 138986 680378 139222 680614
rect 139306 680378 139542 680614
rect 138986 680058 139222 680294
rect 139306 680058 139542 680294
rect 138986 644378 139222 644614
rect 139306 644378 139542 644614
rect 138986 644058 139222 644294
rect 139306 644058 139542 644294
rect 138986 608378 139222 608614
rect 139306 608378 139542 608614
rect 138986 608058 139222 608294
rect 139306 608058 139542 608294
rect 138986 572378 139222 572614
rect 139306 572378 139542 572614
rect 138986 572058 139222 572294
rect 139306 572058 139542 572294
rect 138986 536378 139222 536614
rect 139306 536378 139542 536614
rect 138986 536058 139222 536294
rect 139306 536058 139542 536294
rect 138986 500378 139222 500614
rect 139306 500378 139542 500614
rect 138986 500058 139222 500294
rect 139306 500058 139542 500294
rect 138986 464378 139222 464614
rect 139306 464378 139542 464614
rect 138986 464058 139222 464294
rect 139306 464058 139542 464294
rect 138986 428378 139222 428614
rect 139306 428378 139542 428614
rect 138986 428058 139222 428294
rect 139306 428058 139542 428294
rect 138986 392378 139222 392614
rect 139306 392378 139542 392614
rect 138986 392058 139222 392294
rect 139306 392058 139542 392294
rect 138986 356378 139222 356614
rect 139306 356378 139542 356614
rect 138986 356058 139222 356294
rect 139306 356058 139542 356294
rect 138986 320378 139222 320614
rect 139306 320378 139542 320614
rect 138986 320058 139222 320294
rect 139306 320058 139542 320294
rect 138986 284378 139222 284614
rect 139306 284378 139542 284614
rect 138986 284058 139222 284294
rect 139306 284058 139542 284294
rect 138986 248378 139222 248614
rect 139306 248378 139542 248614
rect 138986 248058 139222 248294
rect 139306 248058 139542 248294
rect 138986 212378 139222 212614
rect 139306 212378 139542 212614
rect 138986 212058 139222 212294
rect 139306 212058 139542 212294
rect 138986 176378 139222 176614
rect 139306 176378 139542 176614
rect 138986 176058 139222 176294
rect 139306 176058 139542 176294
rect 138986 140378 139222 140614
rect 139306 140378 139542 140614
rect 138986 140058 139222 140294
rect 139306 140058 139542 140294
rect 138986 104378 139222 104614
rect 139306 104378 139542 104614
rect 138986 104058 139222 104294
rect 139306 104058 139542 104294
rect 138986 68378 139222 68614
rect 139306 68378 139542 68614
rect 138986 68058 139222 68294
rect 139306 68058 139542 68294
rect 138986 32378 139222 32614
rect 139306 32378 139542 32614
rect 138986 32058 139222 32294
rect 139306 32058 139542 32294
rect 120986 -6342 121222 -6106
rect 121306 -6342 121542 -6106
rect 120986 -6662 121222 -6426
rect 121306 -6662 121542 -6426
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 145826 507218 146062 507454
rect 146146 507218 146382 507454
rect 145826 506898 146062 507134
rect 146146 506898 146382 507134
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 145826 435218 146062 435454
rect 146146 435218 146382 435454
rect 145826 434898 146062 435134
rect 146146 434898 146382 435134
rect 145826 399218 146062 399454
rect 146146 399218 146382 399454
rect 145826 398898 146062 399134
rect 146146 398898 146382 399134
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 145826 327218 146062 327454
rect 146146 327218 146382 327454
rect 145826 326898 146062 327134
rect 146146 326898 146382 327134
rect 145826 291218 146062 291454
rect 146146 291218 146382 291454
rect 145826 290898 146062 291134
rect 146146 290898 146382 291134
rect 145826 255218 146062 255454
rect 146146 255218 146382 255454
rect 145826 254898 146062 255134
rect 146146 254898 146382 255134
rect 145826 219218 146062 219454
rect 146146 219218 146382 219454
rect 145826 218898 146062 219134
rect 146146 218898 146382 219134
rect 145826 183218 146062 183454
rect 146146 183218 146382 183454
rect 145826 182898 146062 183134
rect 146146 182898 146382 183134
rect 145826 147218 146062 147454
rect 146146 147218 146382 147454
rect 145826 146898 146062 147134
rect 146146 146898 146382 147134
rect 145826 111218 146062 111454
rect 146146 111218 146382 111454
rect 145826 110898 146062 111134
rect 146146 110898 146382 111134
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 149546 654938 149782 655174
rect 149866 654938 150102 655174
rect 149546 654618 149782 654854
rect 149866 654618 150102 654854
rect 149546 618938 149782 619174
rect 149866 618938 150102 619174
rect 149546 618618 149782 618854
rect 149866 618618 150102 618854
rect 149546 582938 149782 583174
rect 149866 582938 150102 583174
rect 149546 582618 149782 582854
rect 149866 582618 150102 582854
rect 149546 546938 149782 547174
rect 149866 546938 150102 547174
rect 149546 546618 149782 546854
rect 149866 546618 150102 546854
rect 149546 510938 149782 511174
rect 149866 510938 150102 511174
rect 149546 510618 149782 510854
rect 149866 510618 150102 510854
rect 149546 474938 149782 475174
rect 149866 474938 150102 475174
rect 149546 474618 149782 474854
rect 149866 474618 150102 474854
rect 149546 438938 149782 439174
rect 149866 438938 150102 439174
rect 149546 438618 149782 438854
rect 149866 438618 150102 438854
rect 149546 402938 149782 403174
rect 149866 402938 150102 403174
rect 149546 402618 149782 402854
rect 149866 402618 150102 402854
rect 149546 366938 149782 367174
rect 149866 366938 150102 367174
rect 149546 366618 149782 366854
rect 149866 366618 150102 366854
rect 149546 330938 149782 331174
rect 149866 330938 150102 331174
rect 149546 330618 149782 330854
rect 149866 330618 150102 330854
rect 149546 294938 149782 295174
rect 149866 294938 150102 295174
rect 149546 294618 149782 294854
rect 149866 294618 150102 294854
rect 149546 258938 149782 259174
rect 149866 258938 150102 259174
rect 149546 258618 149782 258854
rect 149866 258618 150102 258854
rect 149546 222938 149782 223174
rect 149866 222938 150102 223174
rect 149546 222618 149782 222854
rect 149866 222618 150102 222854
rect 149546 186938 149782 187174
rect 149866 186938 150102 187174
rect 149546 186618 149782 186854
rect 149866 186618 150102 186854
rect 149546 150938 149782 151174
rect 149866 150938 150102 151174
rect 149546 150618 149782 150854
rect 149866 150618 150102 150854
rect 149546 114938 149782 115174
rect 149866 114938 150102 115174
rect 149546 114618 149782 114854
rect 149866 114618 150102 114854
rect 149546 78938 149782 79174
rect 149866 78938 150102 79174
rect 149546 78618 149782 78854
rect 149866 78618 150102 78854
rect 149546 42938 149782 43174
rect 149866 42938 150102 43174
rect 149546 42618 149782 42854
rect 149866 42618 150102 42854
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 149546 -2502 149782 -2266
rect 149866 -2502 150102 -2266
rect 149546 -2822 149782 -2586
rect 149866 -2822 150102 -2586
rect 153266 694658 153502 694894
rect 153586 694658 153822 694894
rect 153266 694338 153502 694574
rect 153586 694338 153822 694574
rect 153266 658658 153502 658894
rect 153586 658658 153822 658894
rect 153266 658338 153502 658574
rect 153586 658338 153822 658574
rect 153266 622658 153502 622894
rect 153586 622658 153822 622894
rect 153266 622338 153502 622574
rect 153586 622338 153822 622574
rect 153266 586658 153502 586894
rect 153586 586658 153822 586894
rect 153266 586338 153502 586574
rect 153586 586338 153822 586574
rect 153266 550658 153502 550894
rect 153586 550658 153822 550894
rect 153266 550338 153502 550574
rect 153586 550338 153822 550574
rect 153266 514658 153502 514894
rect 153586 514658 153822 514894
rect 153266 514338 153502 514574
rect 153586 514338 153822 514574
rect 153266 478658 153502 478894
rect 153586 478658 153822 478894
rect 153266 478338 153502 478574
rect 153586 478338 153822 478574
rect 153266 442658 153502 442894
rect 153586 442658 153822 442894
rect 153266 442338 153502 442574
rect 153586 442338 153822 442574
rect 153266 406658 153502 406894
rect 153586 406658 153822 406894
rect 153266 406338 153502 406574
rect 153586 406338 153822 406574
rect 153266 370658 153502 370894
rect 153586 370658 153822 370894
rect 153266 370338 153502 370574
rect 153586 370338 153822 370574
rect 153266 334658 153502 334894
rect 153586 334658 153822 334894
rect 153266 334338 153502 334574
rect 153586 334338 153822 334574
rect 153266 298658 153502 298894
rect 153586 298658 153822 298894
rect 153266 298338 153502 298574
rect 153586 298338 153822 298574
rect 153266 262658 153502 262894
rect 153586 262658 153822 262894
rect 153266 262338 153502 262574
rect 153586 262338 153822 262574
rect 153266 226658 153502 226894
rect 153586 226658 153822 226894
rect 153266 226338 153502 226574
rect 153586 226338 153822 226574
rect 153266 190658 153502 190894
rect 153586 190658 153822 190894
rect 153266 190338 153502 190574
rect 153586 190338 153822 190574
rect 153266 154658 153502 154894
rect 153586 154658 153822 154894
rect 153266 154338 153502 154574
rect 153586 154338 153822 154574
rect 153266 118658 153502 118894
rect 153586 118658 153822 118894
rect 153266 118338 153502 118574
rect 153586 118338 153822 118574
rect 153266 82658 153502 82894
rect 153586 82658 153822 82894
rect 153266 82338 153502 82574
rect 153586 82338 153822 82574
rect 153266 46658 153502 46894
rect 153586 46658 153822 46894
rect 153266 46338 153502 46574
rect 153586 46338 153822 46574
rect 153266 10658 153502 10894
rect 153586 10658 153822 10894
rect 153266 10338 153502 10574
rect 153586 10338 153822 10574
rect 153266 -4422 153502 -4186
rect 153586 -4422 153822 -4186
rect 153266 -4742 153502 -4506
rect 153586 -4742 153822 -4506
rect 174986 711322 175222 711558
rect 175306 711322 175542 711558
rect 174986 711002 175222 711238
rect 175306 711002 175542 711238
rect 171266 709402 171502 709638
rect 171586 709402 171822 709638
rect 171266 709082 171502 709318
rect 171586 709082 171822 709318
rect 167546 707482 167782 707718
rect 167866 707482 168102 707718
rect 167546 707162 167782 707398
rect 167866 707162 168102 707398
rect 156986 698378 157222 698614
rect 157306 698378 157542 698614
rect 156986 698058 157222 698294
rect 157306 698058 157542 698294
rect 156986 662378 157222 662614
rect 157306 662378 157542 662614
rect 156986 662058 157222 662294
rect 157306 662058 157542 662294
rect 156986 626378 157222 626614
rect 157306 626378 157542 626614
rect 156986 626058 157222 626294
rect 157306 626058 157542 626294
rect 156986 590378 157222 590614
rect 157306 590378 157542 590614
rect 156986 590058 157222 590294
rect 157306 590058 157542 590294
rect 156986 554378 157222 554614
rect 157306 554378 157542 554614
rect 156986 554058 157222 554294
rect 157306 554058 157542 554294
rect 156986 518378 157222 518614
rect 157306 518378 157542 518614
rect 156986 518058 157222 518294
rect 157306 518058 157542 518294
rect 156986 482378 157222 482614
rect 157306 482378 157542 482614
rect 156986 482058 157222 482294
rect 157306 482058 157542 482294
rect 156986 446378 157222 446614
rect 157306 446378 157542 446614
rect 156986 446058 157222 446294
rect 157306 446058 157542 446294
rect 156986 410378 157222 410614
rect 157306 410378 157542 410614
rect 156986 410058 157222 410294
rect 157306 410058 157542 410294
rect 156986 374378 157222 374614
rect 157306 374378 157542 374614
rect 156986 374058 157222 374294
rect 157306 374058 157542 374294
rect 156986 338378 157222 338614
rect 157306 338378 157542 338614
rect 156986 338058 157222 338294
rect 157306 338058 157542 338294
rect 156986 302378 157222 302614
rect 157306 302378 157542 302614
rect 156986 302058 157222 302294
rect 157306 302058 157542 302294
rect 156986 266378 157222 266614
rect 157306 266378 157542 266614
rect 156986 266058 157222 266294
rect 157306 266058 157542 266294
rect 156986 230378 157222 230614
rect 157306 230378 157542 230614
rect 156986 230058 157222 230294
rect 157306 230058 157542 230294
rect 156986 194378 157222 194614
rect 157306 194378 157542 194614
rect 156986 194058 157222 194294
rect 157306 194058 157542 194294
rect 163826 705562 164062 705798
rect 164146 705562 164382 705798
rect 163826 705242 164062 705478
rect 164146 705242 164382 705478
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 163826 561218 164062 561454
rect 164146 561218 164382 561454
rect 163826 560898 164062 561134
rect 164146 560898 164382 561134
rect 163826 525218 164062 525454
rect 164146 525218 164382 525454
rect 163826 524898 164062 525134
rect 164146 524898 164382 525134
rect 163826 489218 164062 489454
rect 164146 489218 164382 489454
rect 163826 488898 164062 489134
rect 164146 488898 164382 489134
rect 163826 453218 164062 453454
rect 164146 453218 164382 453454
rect 163826 452898 164062 453134
rect 164146 452898 164382 453134
rect 163826 417218 164062 417454
rect 164146 417218 164382 417454
rect 163826 416898 164062 417134
rect 164146 416898 164382 417134
rect 163826 381218 164062 381454
rect 164146 381218 164382 381454
rect 163826 380898 164062 381134
rect 164146 380898 164382 381134
rect 163826 345218 164062 345454
rect 164146 345218 164382 345454
rect 163826 344898 164062 345134
rect 164146 344898 164382 345134
rect 163826 309218 164062 309454
rect 164146 309218 164382 309454
rect 163826 308898 164062 309134
rect 164146 308898 164382 309134
rect 163826 273218 164062 273454
rect 164146 273218 164382 273454
rect 163826 272898 164062 273134
rect 164146 272898 164382 273134
rect 163826 237218 164062 237454
rect 164146 237218 164382 237454
rect 163826 236898 164062 237134
rect 164146 236898 164382 237134
rect 163826 201218 164062 201454
rect 164146 201218 164382 201454
rect 163826 200898 164062 201134
rect 164146 200898 164382 201134
rect 167546 672938 167782 673174
rect 167866 672938 168102 673174
rect 167546 672618 167782 672854
rect 167866 672618 168102 672854
rect 167546 636938 167782 637174
rect 167866 636938 168102 637174
rect 167546 636618 167782 636854
rect 167866 636618 168102 636854
rect 167546 600938 167782 601174
rect 167866 600938 168102 601174
rect 167546 600618 167782 600854
rect 167866 600618 168102 600854
rect 167546 564938 167782 565174
rect 167866 564938 168102 565174
rect 167546 564618 167782 564854
rect 167866 564618 168102 564854
rect 167546 528938 167782 529174
rect 167866 528938 168102 529174
rect 167546 528618 167782 528854
rect 167866 528618 168102 528854
rect 167546 492938 167782 493174
rect 167866 492938 168102 493174
rect 167546 492618 167782 492854
rect 167866 492618 168102 492854
rect 167546 456938 167782 457174
rect 167866 456938 168102 457174
rect 167546 456618 167782 456854
rect 167866 456618 168102 456854
rect 167546 420938 167782 421174
rect 167866 420938 168102 421174
rect 167546 420618 167782 420854
rect 167866 420618 168102 420854
rect 167546 384938 167782 385174
rect 167866 384938 168102 385174
rect 167546 384618 167782 384854
rect 167866 384618 168102 384854
rect 167546 348938 167782 349174
rect 167866 348938 168102 349174
rect 167546 348618 167782 348854
rect 167866 348618 168102 348854
rect 167546 312938 167782 313174
rect 167866 312938 168102 313174
rect 167546 312618 167782 312854
rect 167866 312618 168102 312854
rect 167546 276938 167782 277174
rect 167866 276938 168102 277174
rect 167546 276618 167782 276854
rect 167866 276618 168102 276854
rect 167546 240938 167782 241174
rect 167866 240938 168102 241174
rect 167546 240618 167782 240854
rect 167866 240618 168102 240854
rect 167546 204938 167782 205174
rect 167866 204938 168102 205174
rect 167546 204618 167782 204854
rect 167866 204618 168102 204854
rect 171266 676658 171502 676894
rect 171586 676658 171822 676894
rect 171266 676338 171502 676574
rect 171586 676338 171822 676574
rect 171266 640658 171502 640894
rect 171586 640658 171822 640894
rect 171266 640338 171502 640574
rect 171586 640338 171822 640574
rect 171266 604658 171502 604894
rect 171586 604658 171822 604894
rect 171266 604338 171502 604574
rect 171586 604338 171822 604574
rect 171266 568658 171502 568894
rect 171586 568658 171822 568894
rect 171266 568338 171502 568574
rect 171586 568338 171822 568574
rect 171266 532658 171502 532894
rect 171586 532658 171822 532894
rect 171266 532338 171502 532574
rect 171586 532338 171822 532574
rect 171266 496658 171502 496894
rect 171586 496658 171822 496894
rect 171266 496338 171502 496574
rect 171586 496338 171822 496574
rect 171266 460658 171502 460894
rect 171586 460658 171822 460894
rect 171266 460338 171502 460574
rect 171586 460338 171822 460574
rect 171266 424658 171502 424894
rect 171586 424658 171822 424894
rect 171266 424338 171502 424574
rect 171586 424338 171822 424574
rect 171266 388658 171502 388894
rect 171586 388658 171822 388894
rect 171266 388338 171502 388574
rect 171586 388338 171822 388574
rect 171266 352658 171502 352894
rect 171586 352658 171822 352894
rect 171266 352338 171502 352574
rect 171586 352338 171822 352574
rect 171266 316658 171502 316894
rect 171586 316658 171822 316894
rect 171266 316338 171502 316574
rect 171586 316338 171822 316574
rect 171266 280658 171502 280894
rect 171586 280658 171822 280894
rect 171266 280338 171502 280574
rect 171586 280338 171822 280574
rect 171266 244658 171502 244894
rect 171586 244658 171822 244894
rect 171266 244338 171502 244574
rect 171586 244338 171822 244574
rect 171266 208658 171502 208894
rect 171586 208658 171822 208894
rect 171266 208338 171502 208574
rect 171586 208338 171822 208574
rect 192986 710362 193222 710598
rect 193306 710362 193542 710598
rect 192986 710042 193222 710278
rect 193306 710042 193542 710278
rect 189266 708442 189502 708678
rect 189586 708442 189822 708678
rect 189266 708122 189502 708358
rect 189586 708122 189822 708358
rect 185546 706522 185782 706758
rect 185866 706522 186102 706758
rect 185546 706202 185782 706438
rect 185866 706202 186102 706438
rect 174986 680378 175222 680614
rect 175306 680378 175542 680614
rect 174986 680058 175222 680294
rect 175306 680058 175542 680294
rect 174986 644378 175222 644614
rect 175306 644378 175542 644614
rect 174986 644058 175222 644294
rect 175306 644058 175542 644294
rect 174986 608378 175222 608614
rect 175306 608378 175542 608614
rect 174986 608058 175222 608294
rect 175306 608058 175542 608294
rect 174986 572378 175222 572614
rect 175306 572378 175542 572614
rect 174986 572058 175222 572294
rect 175306 572058 175542 572294
rect 174986 536378 175222 536614
rect 175306 536378 175542 536614
rect 174986 536058 175222 536294
rect 175306 536058 175542 536294
rect 174986 500378 175222 500614
rect 175306 500378 175542 500614
rect 174986 500058 175222 500294
rect 175306 500058 175542 500294
rect 174986 464378 175222 464614
rect 175306 464378 175542 464614
rect 174986 464058 175222 464294
rect 175306 464058 175542 464294
rect 174986 428378 175222 428614
rect 175306 428378 175542 428614
rect 174986 428058 175222 428294
rect 175306 428058 175542 428294
rect 174986 392378 175222 392614
rect 175306 392378 175542 392614
rect 174986 392058 175222 392294
rect 175306 392058 175542 392294
rect 174986 356378 175222 356614
rect 175306 356378 175542 356614
rect 174986 356058 175222 356294
rect 175306 356058 175542 356294
rect 174986 320378 175222 320614
rect 175306 320378 175542 320614
rect 174986 320058 175222 320294
rect 175306 320058 175542 320294
rect 174986 284378 175222 284614
rect 175306 284378 175542 284614
rect 174986 284058 175222 284294
rect 175306 284058 175542 284294
rect 174986 248378 175222 248614
rect 175306 248378 175542 248614
rect 174986 248058 175222 248294
rect 175306 248058 175542 248294
rect 174986 212378 175222 212614
rect 175306 212378 175542 212614
rect 174986 212058 175222 212294
rect 175306 212058 175542 212294
rect 162285 183218 162521 183454
rect 162285 182898 162521 183134
rect 164882 183218 165118 183454
rect 164882 182898 165118 183134
rect 167479 183218 167715 183454
rect 167479 182898 167715 183134
rect 174986 176378 175222 176614
rect 175306 176378 175542 176614
rect 174986 176058 175222 176294
rect 175306 176058 175542 176294
rect 163583 165218 163819 165454
rect 163583 164898 163819 165134
rect 166180 165218 166416 165454
rect 166180 164898 166416 165134
rect 156986 158378 157222 158614
rect 157306 158378 157542 158614
rect 156986 158058 157222 158294
rect 157306 158058 157542 158294
rect 162285 147218 162521 147454
rect 162285 146898 162521 147134
rect 164882 147218 165118 147454
rect 164882 146898 165118 147134
rect 167479 147218 167715 147454
rect 167479 146898 167715 147134
rect 174986 140378 175222 140614
rect 175306 140378 175542 140614
rect 174986 140058 175222 140294
rect 175306 140058 175542 140294
rect 163583 129218 163819 129454
rect 163583 128898 163819 129134
rect 166180 129218 166416 129454
rect 166180 128898 166416 129134
rect 156986 122378 157222 122614
rect 157306 122378 157542 122614
rect 156986 122058 157222 122294
rect 157306 122058 157542 122294
rect 156986 86378 157222 86614
rect 157306 86378 157542 86614
rect 156986 86058 157222 86294
rect 157306 86058 157542 86294
rect 156986 50378 157222 50614
rect 157306 50378 157542 50614
rect 156986 50058 157222 50294
rect 157306 50058 157542 50294
rect 156986 14378 157222 14614
rect 157306 14378 157542 14614
rect 156986 14058 157222 14294
rect 157306 14058 157542 14294
rect 138986 -7302 139222 -7066
rect 139306 -7302 139542 -7066
rect 138986 -7622 139222 -7386
rect 139306 -7622 139542 -7386
rect 163826 93218 164062 93454
rect 164146 93218 164382 93454
rect 163826 92898 164062 93134
rect 164146 92898 164382 93134
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -1542 164062 -1306
rect 164146 -1542 164382 -1306
rect 163826 -1862 164062 -1626
rect 164146 -1862 164382 -1626
rect 167546 96938 167782 97174
rect 167866 96938 168102 97174
rect 167546 96618 167782 96854
rect 167866 96618 168102 96854
rect 167546 60938 167782 61174
rect 167866 60938 168102 61174
rect 167546 60618 167782 60854
rect 167866 60618 168102 60854
rect 167546 24938 167782 25174
rect 167866 24938 168102 25174
rect 167546 24618 167782 24854
rect 167866 24618 168102 24854
rect 167546 -3462 167782 -3226
rect 167866 -3462 168102 -3226
rect 167546 -3782 167782 -3546
rect 167866 -3782 168102 -3546
rect 171266 100658 171502 100894
rect 171586 100658 171822 100894
rect 171266 100338 171502 100574
rect 171586 100338 171822 100574
rect 171266 64658 171502 64894
rect 171586 64658 171822 64894
rect 171266 64338 171502 64574
rect 171586 64338 171822 64574
rect 171266 28658 171502 28894
rect 171586 28658 171822 28894
rect 171266 28338 171502 28574
rect 171586 28338 171822 28574
rect 171266 -5382 171502 -5146
rect 171586 -5382 171822 -5146
rect 171266 -5702 171502 -5466
rect 171586 -5702 171822 -5466
rect 174986 104378 175222 104614
rect 175306 104378 175542 104614
rect 174986 104058 175222 104294
rect 175306 104058 175542 104294
rect 174986 68378 175222 68614
rect 175306 68378 175542 68614
rect 174986 68058 175222 68294
rect 175306 68058 175542 68294
rect 174986 32378 175222 32614
rect 175306 32378 175542 32614
rect 174986 32058 175222 32294
rect 175306 32058 175542 32294
rect 156986 -6342 157222 -6106
rect 157306 -6342 157542 -6106
rect 156986 -6662 157222 -6426
rect 157306 -6662 157542 -6426
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 181826 435218 182062 435454
rect 182146 435218 182382 435454
rect 181826 434898 182062 435134
rect 182146 434898 182382 435134
rect 181826 399218 182062 399454
rect 182146 399218 182382 399454
rect 181826 398898 182062 399134
rect 182146 398898 182382 399134
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 181826 327218 182062 327454
rect 182146 327218 182382 327454
rect 181826 326898 182062 327134
rect 182146 326898 182382 327134
rect 181826 291218 182062 291454
rect 182146 291218 182382 291454
rect 181826 290898 182062 291134
rect 182146 290898 182382 291134
rect 181826 255218 182062 255454
rect 182146 255218 182382 255454
rect 181826 254898 182062 255134
rect 182146 254898 182382 255134
rect 181826 219218 182062 219454
rect 182146 219218 182382 219454
rect 181826 218898 182062 219134
rect 182146 218898 182382 219134
rect 181826 183218 182062 183454
rect 182146 183218 182382 183454
rect 181826 182898 182062 183134
rect 182146 182898 182382 183134
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 181826 111218 182062 111454
rect 182146 111218 182382 111454
rect 181826 110898 182062 111134
rect 182146 110898 182382 111134
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 185546 690938 185782 691174
rect 185866 690938 186102 691174
rect 185546 690618 185782 690854
rect 185866 690618 186102 690854
rect 185546 654938 185782 655174
rect 185866 654938 186102 655174
rect 185546 654618 185782 654854
rect 185866 654618 186102 654854
rect 185546 618938 185782 619174
rect 185866 618938 186102 619174
rect 185546 618618 185782 618854
rect 185866 618618 186102 618854
rect 185546 582938 185782 583174
rect 185866 582938 186102 583174
rect 185546 582618 185782 582854
rect 185866 582618 186102 582854
rect 185546 546938 185782 547174
rect 185866 546938 186102 547174
rect 185546 546618 185782 546854
rect 185866 546618 186102 546854
rect 185546 510938 185782 511174
rect 185866 510938 186102 511174
rect 185546 510618 185782 510854
rect 185866 510618 186102 510854
rect 185546 474938 185782 475174
rect 185866 474938 186102 475174
rect 185546 474618 185782 474854
rect 185866 474618 186102 474854
rect 185546 438938 185782 439174
rect 185866 438938 186102 439174
rect 185546 438618 185782 438854
rect 185866 438618 186102 438854
rect 185546 402938 185782 403174
rect 185866 402938 186102 403174
rect 185546 402618 185782 402854
rect 185866 402618 186102 402854
rect 185546 366938 185782 367174
rect 185866 366938 186102 367174
rect 185546 366618 185782 366854
rect 185866 366618 186102 366854
rect 185546 330938 185782 331174
rect 185866 330938 186102 331174
rect 185546 330618 185782 330854
rect 185866 330618 186102 330854
rect 185546 294938 185782 295174
rect 185866 294938 186102 295174
rect 185546 294618 185782 294854
rect 185866 294618 186102 294854
rect 185546 258938 185782 259174
rect 185866 258938 186102 259174
rect 185546 258618 185782 258854
rect 185866 258618 186102 258854
rect 185546 222938 185782 223174
rect 185866 222938 186102 223174
rect 185546 222618 185782 222854
rect 185866 222618 186102 222854
rect 185546 186938 185782 187174
rect 185866 186938 186102 187174
rect 185546 186618 185782 186854
rect 185866 186618 186102 186854
rect 185546 150938 185782 151174
rect 185866 150938 186102 151174
rect 185546 150618 185782 150854
rect 185866 150618 186102 150854
rect 185546 114938 185782 115174
rect 185866 114938 186102 115174
rect 185546 114618 185782 114854
rect 185866 114618 186102 114854
rect 185546 78938 185782 79174
rect 185866 78938 186102 79174
rect 185546 78618 185782 78854
rect 185866 78618 186102 78854
rect 185546 42938 185782 43174
rect 185866 42938 186102 43174
rect 185546 42618 185782 42854
rect 185866 42618 186102 42854
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 185546 -2502 185782 -2266
rect 185866 -2502 186102 -2266
rect 185546 -2822 185782 -2586
rect 185866 -2822 186102 -2586
rect 189266 694658 189502 694894
rect 189586 694658 189822 694894
rect 189266 694338 189502 694574
rect 189586 694338 189822 694574
rect 189266 658658 189502 658894
rect 189586 658658 189822 658894
rect 189266 658338 189502 658574
rect 189586 658338 189822 658574
rect 189266 622658 189502 622894
rect 189586 622658 189822 622894
rect 189266 622338 189502 622574
rect 189586 622338 189822 622574
rect 189266 586658 189502 586894
rect 189586 586658 189822 586894
rect 189266 586338 189502 586574
rect 189586 586338 189822 586574
rect 189266 550658 189502 550894
rect 189586 550658 189822 550894
rect 189266 550338 189502 550574
rect 189586 550338 189822 550574
rect 189266 514658 189502 514894
rect 189586 514658 189822 514894
rect 189266 514338 189502 514574
rect 189586 514338 189822 514574
rect 189266 478658 189502 478894
rect 189586 478658 189822 478894
rect 189266 478338 189502 478574
rect 189586 478338 189822 478574
rect 189266 442658 189502 442894
rect 189586 442658 189822 442894
rect 189266 442338 189502 442574
rect 189586 442338 189822 442574
rect 189266 406658 189502 406894
rect 189586 406658 189822 406894
rect 189266 406338 189502 406574
rect 189586 406338 189822 406574
rect 189266 370658 189502 370894
rect 189586 370658 189822 370894
rect 189266 370338 189502 370574
rect 189586 370338 189822 370574
rect 189266 334658 189502 334894
rect 189586 334658 189822 334894
rect 189266 334338 189502 334574
rect 189586 334338 189822 334574
rect 189266 298658 189502 298894
rect 189586 298658 189822 298894
rect 189266 298338 189502 298574
rect 189586 298338 189822 298574
rect 189266 262658 189502 262894
rect 189586 262658 189822 262894
rect 189266 262338 189502 262574
rect 189586 262338 189822 262574
rect 189266 226658 189502 226894
rect 189586 226658 189822 226894
rect 189266 226338 189502 226574
rect 189586 226338 189822 226574
rect 189266 190658 189502 190894
rect 189586 190658 189822 190894
rect 189266 190338 189502 190574
rect 189586 190338 189822 190574
rect 189266 154658 189502 154894
rect 189586 154658 189822 154894
rect 189266 154338 189502 154574
rect 189586 154338 189822 154574
rect 189266 118658 189502 118894
rect 189586 118658 189822 118894
rect 189266 118338 189502 118574
rect 189586 118338 189822 118574
rect 189266 82658 189502 82894
rect 189586 82658 189822 82894
rect 189266 82338 189502 82574
rect 189586 82338 189822 82574
rect 189266 46658 189502 46894
rect 189586 46658 189822 46894
rect 189266 46338 189502 46574
rect 189586 46338 189822 46574
rect 189266 10658 189502 10894
rect 189586 10658 189822 10894
rect 189266 10338 189502 10574
rect 189586 10338 189822 10574
rect 189266 -4422 189502 -4186
rect 189586 -4422 189822 -4186
rect 189266 -4742 189502 -4506
rect 189586 -4742 189822 -4506
rect 210986 711322 211222 711558
rect 211306 711322 211542 711558
rect 210986 711002 211222 711238
rect 211306 711002 211542 711238
rect 207266 709402 207502 709638
rect 207586 709402 207822 709638
rect 207266 709082 207502 709318
rect 207586 709082 207822 709318
rect 203546 707482 203782 707718
rect 203866 707482 204102 707718
rect 203546 707162 203782 707398
rect 203866 707162 204102 707398
rect 192986 698378 193222 698614
rect 193306 698378 193542 698614
rect 192986 698058 193222 698294
rect 193306 698058 193542 698294
rect 192986 662378 193222 662614
rect 193306 662378 193542 662614
rect 192986 662058 193222 662294
rect 193306 662058 193542 662294
rect 192986 626378 193222 626614
rect 193306 626378 193542 626614
rect 192986 626058 193222 626294
rect 193306 626058 193542 626294
rect 192986 590378 193222 590614
rect 193306 590378 193542 590614
rect 192986 590058 193222 590294
rect 193306 590058 193542 590294
rect 192986 554378 193222 554614
rect 193306 554378 193542 554614
rect 192986 554058 193222 554294
rect 193306 554058 193542 554294
rect 192986 518378 193222 518614
rect 193306 518378 193542 518614
rect 192986 518058 193222 518294
rect 193306 518058 193542 518294
rect 192986 482378 193222 482614
rect 193306 482378 193542 482614
rect 192986 482058 193222 482294
rect 193306 482058 193542 482294
rect 192986 446378 193222 446614
rect 193306 446378 193542 446614
rect 192986 446058 193222 446294
rect 193306 446058 193542 446294
rect 192986 410378 193222 410614
rect 193306 410378 193542 410614
rect 192986 410058 193222 410294
rect 193306 410058 193542 410294
rect 192986 374378 193222 374614
rect 193306 374378 193542 374614
rect 192986 374058 193222 374294
rect 193306 374058 193542 374294
rect 192986 338378 193222 338614
rect 193306 338378 193542 338614
rect 192986 338058 193222 338294
rect 193306 338058 193542 338294
rect 192986 302378 193222 302614
rect 193306 302378 193542 302614
rect 192986 302058 193222 302294
rect 193306 302058 193542 302294
rect 199826 705562 200062 705798
rect 200146 705562 200382 705798
rect 199826 705242 200062 705478
rect 200146 705242 200382 705478
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 199826 561218 200062 561454
rect 200146 561218 200382 561454
rect 199826 560898 200062 561134
rect 200146 560898 200382 561134
rect 199826 525218 200062 525454
rect 200146 525218 200382 525454
rect 199826 524898 200062 525134
rect 200146 524898 200382 525134
rect 199826 489218 200062 489454
rect 200146 489218 200382 489454
rect 199826 488898 200062 489134
rect 200146 488898 200382 489134
rect 199826 453218 200062 453454
rect 200146 453218 200382 453454
rect 199826 452898 200062 453134
rect 200146 452898 200382 453134
rect 199826 417218 200062 417454
rect 200146 417218 200382 417454
rect 199826 416898 200062 417134
rect 200146 416898 200382 417134
rect 199826 381218 200062 381454
rect 200146 381218 200382 381454
rect 199826 380898 200062 381134
rect 200146 380898 200382 381134
rect 199826 345218 200062 345454
rect 200146 345218 200382 345454
rect 199826 344898 200062 345134
rect 200146 344898 200382 345134
rect 199826 309218 200062 309454
rect 200146 309218 200382 309454
rect 199826 308898 200062 309134
rect 200146 308898 200382 309134
rect 203546 672938 203782 673174
rect 203866 672938 204102 673174
rect 203546 672618 203782 672854
rect 203866 672618 204102 672854
rect 203546 636938 203782 637174
rect 203866 636938 204102 637174
rect 203546 636618 203782 636854
rect 203866 636618 204102 636854
rect 203546 600938 203782 601174
rect 203866 600938 204102 601174
rect 203546 600618 203782 600854
rect 203866 600618 204102 600854
rect 203546 564938 203782 565174
rect 203866 564938 204102 565174
rect 203546 564618 203782 564854
rect 203866 564618 204102 564854
rect 203546 528938 203782 529174
rect 203866 528938 204102 529174
rect 203546 528618 203782 528854
rect 203866 528618 204102 528854
rect 203546 492938 203782 493174
rect 203866 492938 204102 493174
rect 203546 492618 203782 492854
rect 203866 492618 204102 492854
rect 203546 456938 203782 457174
rect 203866 456938 204102 457174
rect 203546 456618 203782 456854
rect 203866 456618 204102 456854
rect 203546 420938 203782 421174
rect 203866 420938 204102 421174
rect 203546 420618 203782 420854
rect 203866 420618 204102 420854
rect 203546 384938 203782 385174
rect 203866 384938 204102 385174
rect 203546 384618 203782 384854
rect 203866 384618 204102 384854
rect 203546 348938 203782 349174
rect 203866 348938 204102 349174
rect 203546 348618 203782 348854
rect 203866 348618 204102 348854
rect 203546 312938 203782 313174
rect 203866 312938 204102 313174
rect 203546 312618 203782 312854
rect 203866 312618 204102 312854
rect 207266 676658 207502 676894
rect 207586 676658 207822 676894
rect 207266 676338 207502 676574
rect 207586 676338 207822 676574
rect 207266 640658 207502 640894
rect 207586 640658 207822 640894
rect 207266 640338 207502 640574
rect 207586 640338 207822 640574
rect 207266 604658 207502 604894
rect 207586 604658 207822 604894
rect 207266 604338 207502 604574
rect 207586 604338 207822 604574
rect 207266 568658 207502 568894
rect 207586 568658 207822 568894
rect 207266 568338 207502 568574
rect 207586 568338 207822 568574
rect 207266 532658 207502 532894
rect 207586 532658 207822 532894
rect 207266 532338 207502 532574
rect 207586 532338 207822 532574
rect 207266 496658 207502 496894
rect 207586 496658 207822 496894
rect 207266 496338 207502 496574
rect 207586 496338 207822 496574
rect 207266 460658 207502 460894
rect 207586 460658 207822 460894
rect 207266 460338 207502 460574
rect 207586 460338 207822 460574
rect 207266 424658 207502 424894
rect 207586 424658 207822 424894
rect 207266 424338 207502 424574
rect 207586 424338 207822 424574
rect 207266 388658 207502 388894
rect 207586 388658 207822 388894
rect 207266 388338 207502 388574
rect 207586 388338 207822 388574
rect 207266 352658 207502 352894
rect 207586 352658 207822 352894
rect 207266 352338 207502 352574
rect 207586 352338 207822 352574
rect 207266 316658 207502 316894
rect 207586 316658 207822 316894
rect 207266 316338 207502 316574
rect 207586 316338 207822 316574
rect 228986 710362 229222 710598
rect 229306 710362 229542 710598
rect 228986 710042 229222 710278
rect 229306 710042 229542 710278
rect 225266 708442 225502 708678
rect 225586 708442 225822 708678
rect 225266 708122 225502 708358
rect 225586 708122 225822 708358
rect 221546 706522 221782 706758
rect 221866 706522 222102 706758
rect 221546 706202 221782 706438
rect 221866 706202 222102 706438
rect 210986 680378 211222 680614
rect 211306 680378 211542 680614
rect 210986 680058 211222 680294
rect 211306 680058 211542 680294
rect 210986 644378 211222 644614
rect 211306 644378 211542 644614
rect 210986 644058 211222 644294
rect 211306 644058 211542 644294
rect 210986 608378 211222 608614
rect 211306 608378 211542 608614
rect 210986 608058 211222 608294
rect 211306 608058 211542 608294
rect 210986 572378 211222 572614
rect 211306 572378 211542 572614
rect 210986 572058 211222 572294
rect 211306 572058 211542 572294
rect 210986 536378 211222 536614
rect 211306 536378 211542 536614
rect 210986 536058 211222 536294
rect 211306 536058 211542 536294
rect 210986 500378 211222 500614
rect 211306 500378 211542 500614
rect 210986 500058 211222 500294
rect 211306 500058 211542 500294
rect 210986 464378 211222 464614
rect 211306 464378 211542 464614
rect 210986 464058 211222 464294
rect 211306 464058 211542 464294
rect 210986 428378 211222 428614
rect 211306 428378 211542 428614
rect 210986 428058 211222 428294
rect 211306 428058 211542 428294
rect 210986 392378 211222 392614
rect 211306 392378 211542 392614
rect 210986 392058 211222 392294
rect 211306 392058 211542 392294
rect 210986 356378 211222 356614
rect 211306 356378 211542 356614
rect 210986 356058 211222 356294
rect 211306 356058 211542 356294
rect 210986 320378 211222 320614
rect 211306 320378 211542 320614
rect 210986 320058 211222 320294
rect 211306 320058 211542 320294
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 217826 543218 218062 543454
rect 218146 543218 218382 543454
rect 217826 542898 218062 543134
rect 218146 542898 218382 543134
rect 217826 507218 218062 507454
rect 218146 507218 218382 507454
rect 217826 506898 218062 507134
rect 218146 506898 218382 507134
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 217826 435218 218062 435454
rect 218146 435218 218382 435454
rect 217826 434898 218062 435134
rect 218146 434898 218382 435134
rect 217826 399218 218062 399454
rect 218146 399218 218382 399454
rect 217826 398898 218062 399134
rect 218146 398898 218382 399134
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 217826 327218 218062 327454
rect 218146 327218 218382 327454
rect 217826 326898 218062 327134
rect 218146 326898 218382 327134
rect 221546 690938 221782 691174
rect 221866 690938 222102 691174
rect 221546 690618 221782 690854
rect 221866 690618 222102 690854
rect 221546 654938 221782 655174
rect 221866 654938 222102 655174
rect 221546 654618 221782 654854
rect 221866 654618 222102 654854
rect 221546 618938 221782 619174
rect 221866 618938 222102 619174
rect 221546 618618 221782 618854
rect 221866 618618 222102 618854
rect 221546 582938 221782 583174
rect 221866 582938 222102 583174
rect 221546 582618 221782 582854
rect 221866 582618 222102 582854
rect 221546 546938 221782 547174
rect 221866 546938 222102 547174
rect 221546 546618 221782 546854
rect 221866 546618 222102 546854
rect 221546 510938 221782 511174
rect 221866 510938 222102 511174
rect 221546 510618 221782 510854
rect 221866 510618 222102 510854
rect 221546 474938 221782 475174
rect 221866 474938 222102 475174
rect 221546 474618 221782 474854
rect 221866 474618 222102 474854
rect 221546 438938 221782 439174
rect 221866 438938 222102 439174
rect 221546 438618 221782 438854
rect 221866 438618 222102 438854
rect 221546 402938 221782 403174
rect 221866 402938 222102 403174
rect 221546 402618 221782 402854
rect 221866 402618 222102 402854
rect 221546 366938 221782 367174
rect 221866 366938 222102 367174
rect 221546 366618 221782 366854
rect 221866 366618 222102 366854
rect 221546 330938 221782 331174
rect 221866 330938 222102 331174
rect 221546 330618 221782 330854
rect 221866 330618 222102 330854
rect 225266 694658 225502 694894
rect 225586 694658 225822 694894
rect 225266 694338 225502 694574
rect 225586 694338 225822 694574
rect 225266 658658 225502 658894
rect 225586 658658 225822 658894
rect 225266 658338 225502 658574
rect 225586 658338 225822 658574
rect 225266 622658 225502 622894
rect 225586 622658 225822 622894
rect 225266 622338 225502 622574
rect 225586 622338 225822 622574
rect 225266 586658 225502 586894
rect 225586 586658 225822 586894
rect 225266 586338 225502 586574
rect 225586 586338 225822 586574
rect 225266 550658 225502 550894
rect 225586 550658 225822 550894
rect 225266 550338 225502 550574
rect 225586 550338 225822 550574
rect 225266 514658 225502 514894
rect 225586 514658 225822 514894
rect 225266 514338 225502 514574
rect 225586 514338 225822 514574
rect 225266 478658 225502 478894
rect 225586 478658 225822 478894
rect 225266 478338 225502 478574
rect 225586 478338 225822 478574
rect 225266 442658 225502 442894
rect 225586 442658 225822 442894
rect 225266 442338 225502 442574
rect 225586 442338 225822 442574
rect 225266 406658 225502 406894
rect 225586 406658 225822 406894
rect 225266 406338 225502 406574
rect 225586 406338 225822 406574
rect 225266 370658 225502 370894
rect 225586 370658 225822 370894
rect 225266 370338 225502 370574
rect 225586 370338 225822 370574
rect 225266 334658 225502 334894
rect 225586 334658 225822 334894
rect 225266 334338 225502 334574
rect 225586 334338 225822 334574
rect 246986 711322 247222 711558
rect 247306 711322 247542 711558
rect 246986 711002 247222 711238
rect 247306 711002 247542 711238
rect 243266 709402 243502 709638
rect 243586 709402 243822 709638
rect 243266 709082 243502 709318
rect 243586 709082 243822 709318
rect 239546 707482 239782 707718
rect 239866 707482 240102 707718
rect 239546 707162 239782 707398
rect 239866 707162 240102 707398
rect 228986 698378 229222 698614
rect 229306 698378 229542 698614
rect 228986 698058 229222 698294
rect 229306 698058 229542 698294
rect 228986 662378 229222 662614
rect 229306 662378 229542 662614
rect 228986 662058 229222 662294
rect 229306 662058 229542 662294
rect 228986 626378 229222 626614
rect 229306 626378 229542 626614
rect 228986 626058 229222 626294
rect 229306 626058 229542 626294
rect 228986 590378 229222 590614
rect 229306 590378 229542 590614
rect 228986 590058 229222 590294
rect 229306 590058 229542 590294
rect 228986 554378 229222 554614
rect 229306 554378 229542 554614
rect 228986 554058 229222 554294
rect 229306 554058 229542 554294
rect 228986 518378 229222 518614
rect 229306 518378 229542 518614
rect 228986 518058 229222 518294
rect 229306 518058 229542 518294
rect 228986 482378 229222 482614
rect 229306 482378 229542 482614
rect 228986 482058 229222 482294
rect 229306 482058 229542 482294
rect 228986 446378 229222 446614
rect 229306 446378 229542 446614
rect 228986 446058 229222 446294
rect 229306 446058 229542 446294
rect 228986 410378 229222 410614
rect 229306 410378 229542 410614
rect 228986 410058 229222 410294
rect 229306 410058 229542 410294
rect 228986 374378 229222 374614
rect 229306 374378 229542 374614
rect 228986 374058 229222 374294
rect 229306 374058 229542 374294
rect 228986 338378 229222 338614
rect 229306 338378 229542 338614
rect 228986 338058 229222 338294
rect 229306 338058 229542 338294
rect 228986 302378 229222 302614
rect 229306 302378 229542 302614
rect 228986 302058 229222 302294
rect 229306 302058 229542 302294
rect 235826 705562 236062 705798
rect 236146 705562 236382 705798
rect 235826 705242 236062 705478
rect 236146 705242 236382 705478
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 235826 561218 236062 561454
rect 236146 561218 236382 561454
rect 235826 560898 236062 561134
rect 236146 560898 236382 561134
rect 235826 525218 236062 525454
rect 236146 525218 236382 525454
rect 235826 524898 236062 525134
rect 236146 524898 236382 525134
rect 235826 489218 236062 489454
rect 236146 489218 236382 489454
rect 235826 488898 236062 489134
rect 236146 488898 236382 489134
rect 235826 453218 236062 453454
rect 236146 453218 236382 453454
rect 235826 452898 236062 453134
rect 236146 452898 236382 453134
rect 235826 417218 236062 417454
rect 236146 417218 236382 417454
rect 235826 416898 236062 417134
rect 236146 416898 236382 417134
rect 235826 381218 236062 381454
rect 236146 381218 236382 381454
rect 235826 380898 236062 381134
rect 236146 380898 236382 381134
rect 235826 345218 236062 345454
rect 236146 345218 236382 345454
rect 235826 344898 236062 345134
rect 236146 344898 236382 345134
rect 235826 309218 236062 309454
rect 236146 309218 236382 309454
rect 235826 308898 236062 309134
rect 236146 308898 236382 309134
rect 239546 672938 239782 673174
rect 239866 672938 240102 673174
rect 239546 672618 239782 672854
rect 239866 672618 240102 672854
rect 239546 636938 239782 637174
rect 239866 636938 240102 637174
rect 239546 636618 239782 636854
rect 239866 636618 240102 636854
rect 239546 600938 239782 601174
rect 239866 600938 240102 601174
rect 239546 600618 239782 600854
rect 239866 600618 240102 600854
rect 239546 564938 239782 565174
rect 239866 564938 240102 565174
rect 239546 564618 239782 564854
rect 239866 564618 240102 564854
rect 239546 528938 239782 529174
rect 239866 528938 240102 529174
rect 239546 528618 239782 528854
rect 239866 528618 240102 528854
rect 239546 492938 239782 493174
rect 239866 492938 240102 493174
rect 239546 492618 239782 492854
rect 239866 492618 240102 492854
rect 239546 456938 239782 457174
rect 239866 456938 240102 457174
rect 239546 456618 239782 456854
rect 239866 456618 240102 456854
rect 239546 420938 239782 421174
rect 239866 420938 240102 421174
rect 239546 420618 239782 420854
rect 239866 420618 240102 420854
rect 239546 384938 239782 385174
rect 239866 384938 240102 385174
rect 239546 384618 239782 384854
rect 239866 384618 240102 384854
rect 239546 348938 239782 349174
rect 239866 348938 240102 349174
rect 239546 348618 239782 348854
rect 239866 348618 240102 348854
rect 239546 312938 239782 313174
rect 239866 312938 240102 313174
rect 239546 312618 239782 312854
rect 239866 312618 240102 312854
rect 243266 676658 243502 676894
rect 243586 676658 243822 676894
rect 243266 676338 243502 676574
rect 243586 676338 243822 676574
rect 243266 640658 243502 640894
rect 243586 640658 243822 640894
rect 243266 640338 243502 640574
rect 243586 640338 243822 640574
rect 243266 604658 243502 604894
rect 243586 604658 243822 604894
rect 243266 604338 243502 604574
rect 243586 604338 243822 604574
rect 243266 568658 243502 568894
rect 243586 568658 243822 568894
rect 243266 568338 243502 568574
rect 243586 568338 243822 568574
rect 243266 532658 243502 532894
rect 243586 532658 243822 532894
rect 243266 532338 243502 532574
rect 243586 532338 243822 532574
rect 243266 496658 243502 496894
rect 243586 496658 243822 496894
rect 243266 496338 243502 496574
rect 243586 496338 243822 496574
rect 243266 460658 243502 460894
rect 243586 460658 243822 460894
rect 243266 460338 243502 460574
rect 243586 460338 243822 460574
rect 243266 424658 243502 424894
rect 243586 424658 243822 424894
rect 243266 424338 243502 424574
rect 243586 424338 243822 424574
rect 243266 388658 243502 388894
rect 243586 388658 243822 388894
rect 243266 388338 243502 388574
rect 243586 388338 243822 388574
rect 243266 352658 243502 352894
rect 243586 352658 243822 352894
rect 243266 352338 243502 352574
rect 243586 352338 243822 352574
rect 243266 316658 243502 316894
rect 243586 316658 243822 316894
rect 243266 316338 243502 316574
rect 243586 316338 243822 316574
rect 264986 710362 265222 710598
rect 265306 710362 265542 710598
rect 264986 710042 265222 710278
rect 265306 710042 265542 710278
rect 261266 708442 261502 708678
rect 261586 708442 261822 708678
rect 261266 708122 261502 708358
rect 261586 708122 261822 708358
rect 257546 706522 257782 706758
rect 257866 706522 258102 706758
rect 257546 706202 257782 706438
rect 257866 706202 258102 706438
rect 246986 680378 247222 680614
rect 247306 680378 247542 680614
rect 246986 680058 247222 680294
rect 247306 680058 247542 680294
rect 246986 644378 247222 644614
rect 247306 644378 247542 644614
rect 246986 644058 247222 644294
rect 247306 644058 247542 644294
rect 246986 608378 247222 608614
rect 247306 608378 247542 608614
rect 246986 608058 247222 608294
rect 247306 608058 247542 608294
rect 246986 572378 247222 572614
rect 247306 572378 247542 572614
rect 246986 572058 247222 572294
rect 247306 572058 247542 572294
rect 246986 536378 247222 536614
rect 247306 536378 247542 536614
rect 246986 536058 247222 536294
rect 247306 536058 247542 536294
rect 246986 500378 247222 500614
rect 247306 500378 247542 500614
rect 246986 500058 247222 500294
rect 247306 500058 247542 500294
rect 246986 464378 247222 464614
rect 247306 464378 247542 464614
rect 246986 464058 247222 464294
rect 247306 464058 247542 464294
rect 246986 428378 247222 428614
rect 247306 428378 247542 428614
rect 246986 428058 247222 428294
rect 247306 428058 247542 428294
rect 246986 392378 247222 392614
rect 247306 392378 247542 392614
rect 246986 392058 247222 392294
rect 247306 392058 247542 392294
rect 246986 356378 247222 356614
rect 247306 356378 247542 356614
rect 246986 356058 247222 356294
rect 247306 356058 247542 356294
rect 246986 320378 247222 320614
rect 247306 320378 247542 320614
rect 246986 320058 247222 320294
rect 247306 320058 247542 320294
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 253826 543218 254062 543454
rect 254146 543218 254382 543454
rect 253826 542898 254062 543134
rect 254146 542898 254382 543134
rect 253826 507218 254062 507454
rect 254146 507218 254382 507454
rect 253826 506898 254062 507134
rect 254146 506898 254382 507134
rect 253826 471218 254062 471454
rect 254146 471218 254382 471454
rect 253826 470898 254062 471134
rect 254146 470898 254382 471134
rect 253826 435218 254062 435454
rect 254146 435218 254382 435454
rect 253826 434898 254062 435134
rect 254146 434898 254382 435134
rect 253826 399218 254062 399454
rect 254146 399218 254382 399454
rect 253826 398898 254062 399134
rect 254146 398898 254382 399134
rect 253826 363218 254062 363454
rect 254146 363218 254382 363454
rect 253826 362898 254062 363134
rect 254146 362898 254382 363134
rect 253826 327218 254062 327454
rect 254146 327218 254382 327454
rect 253826 326898 254062 327134
rect 254146 326898 254382 327134
rect 257546 690938 257782 691174
rect 257866 690938 258102 691174
rect 257546 690618 257782 690854
rect 257866 690618 258102 690854
rect 257546 654938 257782 655174
rect 257866 654938 258102 655174
rect 257546 654618 257782 654854
rect 257866 654618 258102 654854
rect 257546 618938 257782 619174
rect 257866 618938 258102 619174
rect 257546 618618 257782 618854
rect 257866 618618 258102 618854
rect 257546 582938 257782 583174
rect 257866 582938 258102 583174
rect 257546 582618 257782 582854
rect 257866 582618 258102 582854
rect 257546 546938 257782 547174
rect 257866 546938 258102 547174
rect 257546 546618 257782 546854
rect 257866 546618 258102 546854
rect 257546 510938 257782 511174
rect 257866 510938 258102 511174
rect 257546 510618 257782 510854
rect 257866 510618 258102 510854
rect 257546 474938 257782 475174
rect 257866 474938 258102 475174
rect 257546 474618 257782 474854
rect 257866 474618 258102 474854
rect 257546 438938 257782 439174
rect 257866 438938 258102 439174
rect 257546 438618 257782 438854
rect 257866 438618 258102 438854
rect 257546 402938 257782 403174
rect 257866 402938 258102 403174
rect 257546 402618 257782 402854
rect 257866 402618 258102 402854
rect 257546 366938 257782 367174
rect 257866 366938 258102 367174
rect 257546 366618 257782 366854
rect 257866 366618 258102 366854
rect 257546 330938 257782 331174
rect 257866 330938 258102 331174
rect 257546 330618 257782 330854
rect 257866 330618 258102 330854
rect 261266 694658 261502 694894
rect 261586 694658 261822 694894
rect 261266 694338 261502 694574
rect 261586 694338 261822 694574
rect 261266 658658 261502 658894
rect 261586 658658 261822 658894
rect 261266 658338 261502 658574
rect 261586 658338 261822 658574
rect 261266 622658 261502 622894
rect 261586 622658 261822 622894
rect 261266 622338 261502 622574
rect 261586 622338 261822 622574
rect 261266 586658 261502 586894
rect 261586 586658 261822 586894
rect 261266 586338 261502 586574
rect 261586 586338 261822 586574
rect 261266 550658 261502 550894
rect 261586 550658 261822 550894
rect 261266 550338 261502 550574
rect 261586 550338 261822 550574
rect 261266 514658 261502 514894
rect 261586 514658 261822 514894
rect 261266 514338 261502 514574
rect 261586 514338 261822 514574
rect 261266 478658 261502 478894
rect 261586 478658 261822 478894
rect 261266 478338 261502 478574
rect 261586 478338 261822 478574
rect 261266 442658 261502 442894
rect 261586 442658 261822 442894
rect 261266 442338 261502 442574
rect 261586 442338 261822 442574
rect 261266 406658 261502 406894
rect 261586 406658 261822 406894
rect 261266 406338 261502 406574
rect 261586 406338 261822 406574
rect 261266 370658 261502 370894
rect 261586 370658 261822 370894
rect 261266 370338 261502 370574
rect 261586 370338 261822 370574
rect 261266 334658 261502 334894
rect 261586 334658 261822 334894
rect 261266 334338 261502 334574
rect 261586 334338 261822 334574
rect 282986 711322 283222 711558
rect 283306 711322 283542 711558
rect 282986 711002 283222 711238
rect 283306 711002 283542 711238
rect 279266 709402 279502 709638
rect 279586 709402 279822 709638
rect 279266 709082 279502 709318
rect 279586 709082 279822 709318
rect 275546 707482 275782 707718
rect 275866 707482 276102 707718
rect 275546 707162 275782 707398
rect 275866 707162 276102 707398
rect 264986 698378 265222 698614
rect 265306 698378 265542 698614
rect 264986 698058 265222 698294
rect 265306 698058 265542 698294
rect 264986 662378 265222 662614
rect 265306 662378 265542 662614
rect 264986 662058 265222 662294
rect 265306 662058 265542 662294
rect 264986 626378 265222 626614
rect 265306 626378 265542 626614
rect 264986 626058 265222 626294
rect 265306 626058 265542 626294
rect 264986 590378 265222 590614
rect 265306 590378 265542 590614
rect 264986 590058 265222 590294
rect 265306 590058 265542 590294
rect 264986 554378 265222 554614
rect 265306 554378 265542 554614
rect 264986 554058 265222 554294
rect 265306 554058 265542 554294
rect 264986 518378 265222 518614
rect 265306 518378 265542 518614
rect 264986 518058 265222 518294
rect 265306 518058 265542 518294
rect 264986 482378 265222 482614
rect 265306 482378 265542 482614
rect 264986 482058 265222 482294
rect 265306 482058 265542 482294
rect 264986 446378 265222 446614
rect 265306 446378 265542 446614
rect 264986 446058 265222 446294
rect 265306 446058 265542 446294
rect 264986 410378 265222 410614
rect 265306 410378 265542 410614
rect 264986 410058 265222 410294
rect 265306 410058 265542 410294
rect 264986 374378 265222 374614
rect 265306 374378 265542 374614
rect 264986 374058 265222 374294
rect 265306 374058 265542 374294
rect 264986 338378 265222 338614
rect 265306 338378 265542 338614
rect 264986 338058 265222 338294
rect 265306 338058 265542 338294
rect 264986 302378 265222 302614
rect 265306 302378 265542 302614
rect 264986 302058 265222 302294
rect 265306 302058 265542 302294
rect 271826 705562 272062 705798
rect 272146 705562 272382 705798
rect 271826 705242 272062 705478
rect 272146 705242 272382 705478
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 271826 561218 272062 561454
rect 272146 561218 272382 561454
rect 271826 560898 272062 561134
rect 272146 560898 272382 561134
rect 271826 525218 272062 525454
rect 272146 525218 272382 525454
rect 271826 524898 272062 525134
rect 272146 524898 272382 525134
rect 271826 489218 272062 489454
rect 272146 489218 272382 489454
rect 271826 488898 272062 489134
rect 272146 488898 272382 489134
rect 271826 453218 272062 453454
rect 272146 453218 272382 453454
rect 271826 452898 272062 453134
rect 272146 452898 272382 453134
rect 271826 417218 272062 417454
rect 272146 417218 272382 417454
rect 271826 416898 272062 417134
rect 272146 416898 272382 417134
rect 271826 381218 272062 381454
rect 272146 381218 272382 381454
rect 271826 380898 272062 381134
rect 272146 380898 272382 381134
rect 271826 345218 272062 345454
rect 272146 345218 272382 345454
rect 271826 344898 272062 345134
rect 272146 344898 272382 345134
rect 271826 309218 272062 309454
rect 272146 309218 272382 309454
rect 271826 308898 272062 309134
rect 272146 308898 272382 309134
rect 275546 672938 275782 673174
rect 275866 672938 276102 673174
rect 275546 672618 275782 672854
rect 275866 672618 276102 672854
rect 275546 636938 275782 637174
rect 275866 636938 276102 637174
rect 275546 636618 275782 636854
rect 275866 636618 276102 636854
rect 275546 600938 275782 601174
rect 275866 600938 276102 601174
rect 275546 600618 275782 600854
rect 275866 600618 276102 600854
rect 275546 564938 275782 565174
rect 275866 564938 276102 565174
rect 275546 564618 275782 564854
rect 275866 564618 276102 564854
rect 275546 528938 275782 529174
rect 275866 528938 276102 529174
rect 275546 528618 275782 528854
rect 275866 528618 276102 528854
rect 275546 492938 275782 493174
rect 275866 492938 276102 493174
rect 275546 492618 275782 492854
rect 275866 492618 276102 492854
rect 275546 456938 275782 457174
rect 275866 456938 276102 457174
rect 275546 456618 275782 456854
rect 275866 456618 276102 456854
rect 275546 420938 275782 421174
rect 275866 420938 276102 421174
rect 275546 420618 275782 420854
rect 275866 420618 276102 420854
rect 275546 384938 275782 385174
rect 275866 384938 276102 385174
rect 275546 384618 275782 384854
rect 275866 384618 276102 384854
rect 275546 348938 275782 349174
rect 275866 348938 276102 349174
rect 275546 348618 275782 348854
rect 275866 348618 276102 348854
rect 275546 312938 275782 313174
rect 275866 312938 276102 313174
rect 275546 312618 275782 312854
rect 275866 312618 276102 312854
rect 279266 676658 279502 676894
rect 279586 676658 279822 676894
rect 279266 676338 279502 676574
rect 279586 676338 279822 676574
rect 279266 640658 279502 640894
rect 279586 640658 279822 640894
rect 279266 640338 279502 640574
rect 279586 640338 279822 640574
rect 279266 604658 279502 604894
rect 279586 604658 279822 604894
rect 279266 604338 279502 604574
rect 279586 604338 279822 604574
rect 279266 568658 279502 568894
rect 279586 568658 279822 568894
rect 279266 568338 279502 568574
rect 279586 568338 279822 568574
rect 279266 532658 279502 532894
rect 279586 532658 279822 532894
rect 279266 532338 279502 532574
rect 279586 532338 279822 532574
rect 279266 496658 279502 496894
rect 279586 496658 279822 496894
rect 279266 496338 279502 496574
rect 279586 496338 279822 496574
rect 279266 460658 279502 460894
rect 279586 460658 279822 460894
rect 279266 460338 279502 460574
rect 279586 460338 279822 460574
rect 279266 424658 279502 424894
rect 279586 424658 279822 424894
rect 279266 424338 279502 424574
rect 279586 424338 279822 424574
rect 279266 388658 279502 388894
rect 279586 388658 279822 388894
rect 279266 388338 279502 388574
rect 279586 388338 279822 388574
rect 279266 352658 279502 352894
rect 279586 352658 279822 352894
rect 279266 352338 279502 352574
rect 279586 352338 279822 352574
rect 279266 316658 279502 316894
rect 279586 316658 279822 316894
rect 279266 316338 279502 316574
rect 279586 316338 279822 316574
rect 300986 710362 301222 710598
rect 301306 710362 301542 710598
rect 300986 710042 301222 710278
rect 301306 710042 301542 710278
rect 297266 708442 297502 708678
rect 297586 708442 297822 708678
rect 297266 708122 297502 708358
rect 297586 708122 297822 708358
rect 293546 706522 293782 706758
rect 293866 706522 294102 706758
rect 293546 706202 293782 706438
rect 293866 706202 294102 706438
rect 282986 680378 283222 680614
rect 283306 680378 283542 680614
rect 282986 680058 283222 680294
rect 283306 680058 283542 680294
rect 282986 644378 283222 644614
rect 283306 644378 283542 644614
rect 282986 644058 283222 644294
rect 283306 644058 283542 644294
rect 282986 608378 283222 608614
rect 283306 608378 283542 608614
rect 282986 608058 283222 608294
rect 283306 608058 283542 608294
rect 282986 572378 283222 572614
rect 283306 572378 283542 572614
rect 282986 572058 283222 572294
rect 283306 572058 283542 572294
rect 282986 536378 283222 536614
rect 283306 536378 283542 536614
rect 282986 536058 283222 536294
rect 283306 536058 283542 536294
rect 282986 500378 283222 500614
rect 283306 500378 283542 500614
rect 282986 500058 283222 500294
rect 283306 500058 283542 500294
rect 282986 464378 283222 464614
rect 283306 464378 283542 464614
rect 282986 464058 283222 464294
rect 283306 464058 283542 464294
rect 282986 428378 283222 428614
rect 283306 428378 283542 428614
rect 282986 428058 283222 428294
rect 283306 428058 283542 428294
rect 282986 392378 283222 392614
rect 283306 392378 283542 392614
rect 282986 392058 283222 392294
rect 283306 392058 283542 392294
rect 282986 356378 283222 356614
rect 283306 356378 283542 356614
rect 282986 356058 283222 356294
rect 283306 356058 283542 356294
rect 282986 320378 283222 320614
rect 283306 320378 283542 320614
rect 282986 320058 283222 320294
rect 283306 320058 283542 320294
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 289826 507218 290062 507454
rect 290146 507218 290382 507454
rect 289826 506898 290062 507134
rect 290146 506898 290382 507134
rect 289826 471218 290062 471454
rect 290146 471218 290382 471454
rect 289826 470898 290062 471134
rect 290146 470898 290382 471134
rect 289826 435218 290062 435454
rect 290146 435218 290382 435454
rect 289826 434898 290062 435134
rect 290146 434898 290382 435134
rect 289826 399218 290062 399454
rect 290146 399218 290382 399454
rect 289826 398898 290062 399134
rect 290146 398898 290382 399134
rect 289826 363218 290062 363454
rect 290146 363218 290382 363454
rect 289826 362898 290062 363134
rect 290146 362898 290382 363134
rect 289826 327218 290062 327454
rect 290146 327218 290382 327454
rect 289826 326898 290062 327134
rect 290146 326898 290382 327134
rect 293546 690938 293782 691174
rect 293866 690938 294102 691174
rect 293546 690618 293782 690854
rect 293866 690618 294102 690854
rect 293546 654938 293782 655174
rect 293866 654938 294102 655174
rect 293546 654618 293782 654854
rect 293866 654618 294102 654854
rect 293546 618938 293782 619174
rect 293866 618938 294102 619174
rect 293546 618618 293782 618854
rect 293866 618618 294102 618854
rect 293546 582938 293782 583174
rect 293866 582938 294102 583174
rect 293546 582618 293782 582854
rect 293866 582618 294102 582854
rect 293546 546938 293782 547174
rect 293866 546938 294102 547174
rect 293546 546618 293782 546854
rect 293866 546618 294102 546854
rect 293546 510938 293782 511174
rect 293866 510938 294102 511174
rect 293546 510618 293782 510854
rect 293866 510618 294102 510854
rect 293546 474938 293782 475174
rect 293866 474938 294102 475174
rect 293546 474618 293782 474854
rect 293866 474618 294102 474854
rect 293546 438938 293782 439174
rect 293866 438938 294102 439174
rect 293546 438618 293782 438854
rect 293866 438618 294102 438854
rect 293546 402938 293782 403174
rect 293866 402938 294102 403174
rect 293546 402618 293782 402854
rect 293866 402618 294102 402854
rect 293546 366938 293782 367174
rect 293866 366938 294102 367174
rect 293546 366618 293782 366854
rect 293866 366618 294102 366854
rect 293546 330938 293782 331174
rect 293866 330938 294102 331174
rect 293546 330618 293782 330854
rect 293866 330618 294102 330854
rect 297266 694658 297502 694894
rect 297586 694658 297822 694894
rect 297266 694338 297502 694574
rect 297586 694338 297822 694574
rect 297266 658658 297502 658894
rect 297586 658658 297822 658894
rect 297266 658338 297502 658574
rect 297586 658338 297822 658574
rect 297266 622658 297502 622894
rect 297586 622658 297822 622894
rect 297266 622338 297502 622574
rect 297586 622338 297822 622574
rect 297266 586658 297502 586894
rect 297586 586658 297822 586894
rect 297266 586338 297502 586574
rect 297586 586338 297822 586574
rect 297266 550658 297502 550894
rect 297586 550658 297822 550894
rect 297266 550338 297502 550574
rect 297586 550338 297822 550574
rect 297266 514658 297502 514894
rect 297586 514658 297822 514894
rect 297266 514338 297502 514574
rect 297586 514338 297822 514574
rect 297266 478658 297502 478894
rect 297586 478658 297822 478894
rect 297266 478338 297502 478574
rect 297586 478338 297822 478574
rect 297266 442658 297502 442894
rect 297586 442658 297822 442894
rect 297266 442338 297502 442574
rect 297586 442338 297822 442574
rect 297266 406658 297502 406894
rect 297586 406658 297822 406894
rect 297266 406338 297502 406574
rect 297586 406338 297822 406574
rect 297266 370658 297502 370894
rect 297586 370658 297822 370894
rect 297266 370338 297502 370574
rect 297586 370338 297822 370574
rect 297266 334658 297502 334894
rect 297586 334658 297822 334894
rect 297266 334338 297502 334574
rect 297586 334338 297822 334574
rect 318986 711322 319222 711558
rect 319306 711322 319542 711558
rect 318986 711002 319222 711238
rect 319306 711002 319542 711238
rect 315266 709402 315502 709638
rect 315586 709402 315822 709638
rect 315266 709082 315502 709318
rect 315586 709082 315822 709318
rect 311546 707482 311782 707718
rect 311866 707482 312102 707718
rect 311546 707162 311782 707398
rect 311866 707162 312102 707398
rect 300986 698378 301222 698614
rect 301306 698378 301542 698614
rect 300986 698058 301222 698294
rect 301306 698058 301542 698294
rect 300986 662378 301222 662614
rect 301306 662378 301542 662614
rect 300986 662058 301222 662294
rect 301306 662058 301542 662294
rect 300986 626378 301222 626614
rect 301306 626378 301542 626614
rect 300986 626058 301222 626294
rect 301306 626058 301542 626294
rect 300986 590378 301222 590614
rect 301306 590378 301542 590614
rect 300986 590058 301222 590294
rect 301306 590058 301542 590294
rect 300986 554378 301222 554614
rect 301306 554378 301542 554614
rect 300986 554058 301222 554294
rect 301306 554058 301542 554294
rect 300986 518378 301222 518614
rect 301306 518378 301542 518614
rect 300986 518058 301222 518294
rect 301306 518058 301542 518294
rect 300986 482378 301222 482614
rect 301306 482378 301542 482614
rect 300986 482058 301222 482294
rect 301306 482058 301542 482294
rect 300986 446378 301222 446614
rect 301306 446378 301542 446614
rect 300986 446058 301222 446294
rect 301306 446058 301542 446294
rect 300986 410378 301222 410614
rect 301306 410378 301542 410614
rect 300986 410058 301222 410294
rect 301306 410058 301542 410294
rect 300986 374378 301222 374614
rect 301306 374378 301542 374614
rect 300986 374058 301222 374294
rect 301306 374058 301542 374294
rect 300986 338378 301222 338614
rect 301306 338378 301542 338614
rect 300986 338058 301222 338294
rect 301306 338058 301542 338294
rect 300986 302378 301222 302614
rect 301306 302378 301542 302614
rect 300986 302058 301222 302294
rect 301306 302058 301542 302294
rect 307826 705562 308062 705798
rect 308146 705562 308382 705798
rect 307826 705242 308062 705478
rect 308146 705242 308382 705478
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 307826 561218 308062 561454
rect 308146 561218 308382 561454
rect 307826 560898 308062 561134
rect 308146 560898 308382 561134
rect 307826 525218 308062 525454
rect 308146 525218 308382 525454
rect 307826 524898 308062 525134
rect 308146 524898 308382 525134
rect 307826 489218 308062 489454
rect 308146 489218 308382 489454
rect 307826 488898 308062 489134
rect 308146 488898 308382 489134
rect 307826 453218 308062 453454
rect 308146 453218 308382 453454
rect 307826 452898 308062 453134
rect 308146 452898 308382 453134
rect 307826 417218 308062 417454
rect 308146 417218 308382 417454
rect 307826 416898 308062 417134
rect 308146 416898 308382 417134
rect 307826 381218 308062 381454
rect 308146 381218 308382 381454
rect 307826 380898 308062 381134
rect 308146 380898 308382 381134
rect 307826 345218 308062 345454
rect 308146 345218 308382 345454
rect 307826 344898 308062 345134
rect 308146 344898 308382 345134
rect 307826 309218 308062 309454
rect 308146 309218 308382 309454
rect 307826 308898 308062 309134
rect 308146 308898 308382 309134
rect 204250 291218 204486 291454
rect 204250 290898 204486 291134
rect 234970 291218 235206 291454
rect 234970 290898 235206 291134
rect 265690 291218 265926 291454
rect 265690 290898 265926 291134
rect 296410 291218 296646 291454
rect 296410 290898 296646 291134
rect 219610 273218 219846 273454
rect 219610 272898 219846 273134
rect 250330 273218 250566 273454
rect 250330 272898 250566 273134
rect 281050 273218 281286 273454
rect 281050 272898 281286 273134
rect 307826 273218 308062 273454
rect 308146 273218 308382 273454
rect 307826 272898 308062 273134
rect 308146 272898 308382 273134
rect 192986 266378 193222 266614
rect 193306 266378 193542 266614
rect 192986 266058 193222 266294
rect 193306 266058 193542 266294
rect 204250 255218 204486 255454
rect 204250 254898 204486 255134
rect 234970 255218 235206 255454
rect 234970 254898 235206 255134
rect 265690 255218 265926 255454
rect 265690 254898 265926 255134
rect 296410 255218 296646 255454
rect 296410 254898 296646 255134
rect 219610 237218 219846 237454
rect 219610 236898 219846 237134
rect 250330 237218 250566 237454
rect 250330 236898 250566 237134
rect 281050 237218 281286 237454
rect 281050 236898 281286 237134
rect 307826 237218 308062 237454
rect 308146 237218 308382 237454
rect 307826 236898 308062 237134
rect 308146 236898 308382 237134
rect 192986 230378 193222 230614
rect 193306 230378 193542 230614
rect 192986 230058 193222 230294
rect 193306 230058 193542 230294
rect 204250 219218 204486 219454
rect 204250 218898 204486 219134
rect 234970 219218 235206 219454
rect 234970 218898 235206 219134
rect 265690 219218 265926 219454
rect 265690 218898 265926 219134
rect 296410 219218 296646 219454
rect 296410 218898 296646 219134
rect 219610 201218 219846 201454
rect 219610 200898 219846 201134
rect 250330 201218 250566 201454
rect 250330 200898 250566 201134
rect 281050 201218 281286 201454
rect 281050 200898 281286 201134
rect 307826 201218 308062 201454
rect 308146 201218 308382 201454
rect 307826 200898 308062 201134
rect 308146 200898 308382 201134
rect 192986 194378 193222 194614
rect 193306 194378 193542 194614
rect 192986 194058 193222 194294
rect 193306 194058 193542 194294
rect 204250 183218 204486 183454
rect 204250 182898 204486 183134
rect 234970 183218 235206 183454
rect 234970 182898 235206 183134
rect 265690 183218 265926 183454
rect 265690 182898 265926 183134
rect 296410 183218 296646 183454
rect 296410 182898 296646 183134
rect 219610 165218 219846 165454
rect 219610 164898 219846 165134
rect 250330 165218 250566 165454
rect 250330 164898 250566 165134
rect 281050 165218 281286 165454
rect 281050 164898 281286 165134
rect 307826 165218 308062 165454
rect 308146 165218 308382 165454
rect 307826 164898 308062 165134
rect 308146 164898 308382 165134
rect 192986 158378 193222 158614
rect 193306 158378 193542 158614
rect 192986 158058 193222 158294
rect 193306 158058 193542 158294
rect 204250 147218 204486 147454
rect 204250 146898 204486 147134
rect 234970 147218 235206 147454
rect 234970 146898 235206 147134
rect 265690 147218 265926 147454
rect 265690 146898 265926 147134
rect 296410 147218 296646 147454
rect 296410 146898 296646 147134
rect 219610 129218 219846 129454
rect 219610 128898 219846 129134
rect 250330 129218 250566 129454
rect 250330 128898 250566 129134
rect 281050 129218 281286 129454
rect 281050 128898 281286 129134
rect 307826 129218 308062 129454
rect 308146 129218 308382 129454
rect 307826 128898 308062 129134
rect 308146 128898 308382 129134
rect 192986 122378 193222 122614
rect 193306 122378 193542 122614
rect 192986 122058 193222 122294
rect 193306 122058 193542 122294
rect 204250 111218 204486 111454
rect 204250 110898 204486 111134
rect 234970 111218 235206 111454
rect 234970 110898 235206 111134
rect 265690 111218 265926 111454
rect 265690 110898 265926 111134
rect 296410 111218 296646 111454
rect 296410 110898 296646 111134
rect 192986 86378 193222 86614
rect 193306 86378 193542 86614
rect 192986 86058 193222 86294
rect 193306 86058 193542 86294
rect 192986 50378 193222 50614
rect 193306 50378 193542 50614
rect 192986 50058 193222 50294
rect 193306 50058 193542 50294
rect 192986 14378 193222 14614
rect 193306 14378 193542 14614
rect 192986 14058 193222 14294
rect 193306 14058 193542 14294
rect 174986 -7302 175222 -7066
rect 175306 -7302 175542 -7066
rect 174986 -7622 175222 -7386
rect 175306 -7622 175542 -7386
rect 199826 93218 200062 93454
rect 200146 93218 200382 93454
rect 199826 92898 200062 93134
rect 200146 92898 200382 93134
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -1542 200062 -1306
rect 200146 -1542 200382 -1306
rect 199826 -1862 200062 -1626
rect 200146 -1862 200382 -1626
rect 203546 96938 203782 97174
rect 203866 96938 204102 97174
rect 203546 96618 203782 96854
rect 203866 96618 204102 96854
rect 203546 60938 203782 61174
rect 203866 60938 204102 61174
rect 203546 60618 203782 60854
rect 203866 60618 204102 60854
rect 203546 24938 203782 25174
rect 203866 24938 204102 25174
rect 203546 24618 203782 24854
rect 203866 24618 204102 24854
rect 203546 -3462 203782 -3226
rect 203866 -3462 204102 -3226
rect 203546 -3782 203782 -3546
rect 203866 -3782 204102 -3546
rect 207266 64658 207502 64894
rect 207586 64658 207822 64894
rect 207266 64338 207502 64574
rect 207586 64338 207822 64574
rect 207266 28658 207502 28894
rect 207586 28658 207822 28894
rect 207266 28338 207502 28574
rect 207586 28338 207822 28574
rect 207266 -5382 207502 -5146
rect 207586 -5382 207822 -5146
rect 207266 -5702 207502 -5466
rect 207586 -5702 207822 -5466
rect 210986 68378 211222 68614
rect 211306 68378 211542 68614
rect 210986 68058 211222 68294
rect 211306 68058 211542 68294
rect 210986 32378 211222 32614
rect 211306 32378 211542 32614
rect 210986 32058 211222 32294
rect 211306 32058 211542 32294
rect 192986 -6342 193222 -6106
rect 193306 -6342 193542 -6106
rect 192986 -6662 193222 -6426
rect 193306 -6662 193542 -6426
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 221546 78938 221782 79174
rect 221866 78938 222102 79174
rect 221546 78618 221782 78854
rect 221866 78618 222102 78854
rect 221546 42938 221782 43174
rect 221866 42938 222102 43174
rect 221546 42618 221782 42854
rect 221866 42618 222102 42854
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 221546 -2502 221782 -2266
rect 221866 -2502 222102 -2266
rect 221546 -2822 221782 -2586
rect 221866 -2822 222102 -2586
rect 225266 82658 225502 82894
rect 225586 82658 225822 82894
rect 225266 82338 225502 82574
rect 225586 82338 225822 82574
rect 225266 46658 225502 46894
rect 225586 46658 225822 46894
rect 225266 46338 225502 46574
rect 225586 46338 225822 46574
rect 225266 10658 225502 10894
rect 225586 10658 225822 10894
rect 225266 10338 225502 10574
rect 225586 10338 225822 10574
rect 225266 -4422 225502 -4186
rect 225586 -4422 225822 -4186
rect 225266 -4742 225502 -4506
rect 225586 -4742 225822 -4506
rect 228986 86378 229222 86614
rect 229306 86378 229542 86614
rect 228986 86058 229222 86294
rect 229306 86058 229542 86294
rect 228986 50378 229222 50614
rect 229306 50378 229542 50614
rect 228986 50058 229222 50294
rect 229306 50058 229542 50294
rect 228986 14378 229222 14614
rect 229306 14378 229542 14614
rect 228986 14058 229222 14294
rect 229306 14058 229542 14294
rect 210986 -7302 211222 -7066
rect 211306 -7302 211542 -7066
rect 210986 -7622 211222 -7386
rect 211306 -7622 211542 -7386
rect 235826 93218 236062 93454
rect 236146 93218 236382 93454
rect 235826 92898 236062 93134
rect 236146 92898 236382 93134
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -1542 236062 -1306
rect 236146 -1542 236382 -1306
rect 235826 -1862 236062 -1626
rect 236146 -1862 236382 -1626
rect 239546 96938 239782 97174
rect 239866 96938 240102 97174
rect 239546 96618 239782 96854
rect 239866 96618 240102 96854
rect 239546 60938 239782 61174
rect 239866 60938 240102 61174
rect 239546 60618 239782 60854
rect 239866 60618 240102 60854
rect 239546 24938 239782 25174
rect 239866 24938 240102 25174
rect 239546 24618 239782 24854
rect 239866 24618 240102 24854
rect 239546 -3462 239782 -3226
rect 239866 -3462 240102 -3226
rect 239546 -3782 239782 -3546
rect 239866 -3782 240102 -3546
rect 243266 64658 243502 64894
rect 243586 64658 243822 64894
rect 243266 64338 243502 64574
rect 243586 64338 243822 64574
rect 243266 28658 243502 28894
rect 243586 28658 243822 28894
rect 243266 28338 243502 28574
rect 243586 28338 243822 28574
rect 243266 -5382 243502 -5146
rect 243586 -5382 243822 -5146
rect 243266 -5702 243502 -5466
rect 243586 -5702 243822 -5466
rect 246986 68378 247222 68614
rect 247306 68378 247542 68614
rect 246986 68058 247222 68294
rect 247306 68058 247542 68294
rect 246986 32378 247222 32614
rect 247306 32378 247542 32614
rect 246986 32058 247222 32294
rect 247306 32058 247542 32294
rect 228986 -6342 229222 -6106
rect 229306 -6342 229542 -6106
rect 228986 -6662 229222 -6426
rect 229306 -6662 229542 -6426
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 257546 78938 257782 79174
rect 257866 78938 258102 79174
rect 257546 78618 257782 78854
rect 257866 78618 258102 78854
rect 257546 42938 257782 43174
rect 257866 42938 258102 43174
rect 257546 42618 257782 42854
rect 257866 42618 258102 42854
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 257546 -2502 257782 -2266
rect 257866 -2502 258102 -2266
rect 257546 -2822 257782 -2586
rect 257866 -2822 258102 -2586
rect 261266 82658 261502 82894
rect 261586 82658 261822 82894
rect 261266 82338 261502 82574
rect 261586 82338 261822 82574
rect 261266 46658 261502 46894
rect 261586 46658 261822 46894
rect 261266 46338 261502 46574
rect 261586 46338 261822 46574
rect 261266 10658 261502 10894
rect 261586 10658 261822 10894
rect 261266 10338 261502 10574
rect 261586 10338 261822 10574
rect 261266 -4422 261502 -4186
rect 261586 -4422 261822 -4186
rect 261266 -4742 261502 -4506
rect 261586 -4742 261822 -4506
rect 264986 86378 265222 86614
rect 265306 86378 265542 86614
rect 264986 86058 265222 86294
rect 265306 86058 265542 86294
rect 264986 50378 265222 50614
rect 265306 50378 265542 50614
rect 264986 50058 265222 50294
rect 265306 50058 265542 50294
rect 264986 14378 265222 14614
rect 265306 14378 265542 14614
rect 264986 14058 265222 14294
rect 265306 14058 265542 14294
rect 246986 -7302 247222 -7066
rect 247306 -7302 247542 -7066
rect 246986 -7622 247222 -7386
rect 247306 -7622 247542 -7386
rect 271826 93218 272062 93454
rect 272146 93218 272382 93454
rect 271826 92898 272062 93134
rect 272146 92898 272382 93134
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -1542 272062 -1306
rect 272146 -1542 272382 -1306
rect 271826 -1862 272062 -1626
rect 272146 -1862 272382 -1626
rect 275546 96938 275782 97174
rect 275866 96938 276102 97174
rect 275546 96618 275782 96854
rect 275866 96618 276102 96854
rect 275546 60938 275782 61174
rect 275866 60938 276102 61174
rect 275546 60618 275782 60854
rect 275866 60618 276102 60854
rect 275546 24938 275782 25174
rect 275866 24938 276102 25174
rect 275546 24618 275782 24854
rect 275866 24618 276102 24854
rect 275546 -3462 275782 -3226
rect 275866 -3462 276102 -3226
rect 275546 -3782 275782 -3546
rect 275866 -3782 276102 -3546
rect 279266 64658 279502 64894
rect 279586 64658 279822 64894
rect 279266 64338 279502 64574
rect 279586 64338 279822 64574
rect 279266 28658 279502 28894
rect 279586 28658 279822 28894
rect 279266 28338 279502 28574
rect 279586 28338 279822 28574
rect 279266 -5382 279502 -5146
rect 279586 -5382 279822 -5146
rect 279266 -5702 279502 -5466
rect 279586 -5702 279822 -5466
rect 282986 68378 283222 68614
rect 283306 68378 283542 68614
rect 282986 68058 283222 68294
rect 283306 68058 283542 68294
rect 282986 32378 283222 32614
rect 283306 32378 283542 32614
rect 282986 32058 283222 32294
rect 283306 32058 283542 32294
rect 264986 -6342 265222 -6106
rect 265306 -6342 265542 -6106
rect 264986 -6662 265222 -6426
rect 265306 -6662 265542 -6426
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 293546 78938 293782 79174
rect 293866 78938 294102 79174
rect 293546 78618 293782 78854
rect 293866 78618 294102 78854
rect 293546 42938 293782 43174
rect 293866 42938 294102 43174
rect 293546 42618 293782 42854
rect 293866 42618 294102 42854
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 293546 -2502 293782 -2266
rect 293866 -2502 294102 -2266
rect 293546 -2822 293782 -2586
rect 293866 -2822 294102 -2586
rect 297266 82658 297502 82894
rect 297586 82658 297822 82894
rect 297266 82338 297502 82574
rect 297586 82338 297822 82574
rect 297266 46658 297502 46894
rect 297586 46658 297822 46894
rect 297266 46338 297502 46574
rect 297586 46338 297822 46574
rect 297266 10658 297502 10894
rect 297586 10658 297822 10894
rect 297266 10338 297502 10574
rect 297586 10338 297822 10574
rect 297266 -4422 297502 -4186
rect 297586 -4422 297822 -4186
rect 297266 -4742 297502 -4506
rect 297586 -4742 297822 -4506
rect 300986 86378 301222 86614
rect 301306 86378 301542 86614
rect 300986 86058 301222 86294
rect 301306 86058 301542 86294
rect 300986 50378 301222 50614
rect 301306 50378 301542 50614
rect 300986 50058 301222 50294
rect 301306 50058 301542 50294
rect 300986 14378 301222 14614
rect 301306 14378 301542 14614
rect 300986 14058 301222 14294
rect 301306 14058 301542 14294
rect 282986 -7302 283222 -7066
rect 283306 -7302 283542 -7066
rect 282986 -7622 283222 -7386
rect 283306 -7622 283542 -7386
rect 307826 93218 308062 93454
rect 308146 93218 308382 93454
rect 307826 92898 308062 93134
rect 308146 92898 308382 93134
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -1542 308062 -1306
rect 308146 -1542 308382 -1306
rect 307826 -1862 308062 -1626
rect 308146 -1862 308382 -1626
rect 311546 672938 311782 673174
rect 311866 672938 312102 673174
rect 311546 672618 311782 672854
rect 311866 672618 312102 672854
rect 311546 636938 311782 637174
rect 311866 636938 312102 637174
rect 311546 636618 311782 636854
rect 311866 636618 312102 636854
rect 311546 600938 311782 601174
rect 311866 600938 312102 601174
rect 311546 600618 311782 600854
rect 311866 600618 312102 600854
rect 311546 564938 311782 565174
rect 311866 564938 312102 565174
rect 311546 564618 311782 564854
rect 311866 564618 312102 564854
rect 311546 528938 311782 529174
rect 311866 528938 312102 529174
rect 311546 528618 311782 528854
rect 311866 528618 312102 528854
rect 311546 492938 311782 493174
rect 311866 492938 312102 493174
rect 311546 492618 311782 492854
rect 311866 492618 312102 492854
rect 311546 456938 311782 457174
rect 311866 456938 312102 457174
rect 311546 456618 311782 456854
rect 311866 456618 312102 456854
rect 311546 420938 311782 421174
rect 311866 420938 312102 421174
rect 311546 420618 311782 420854
rect 311866 420618 312102 420854
rect 311546 384938 311782 385174
rect 311866 384938 312102 385174
rect 311546 384618 311782 384854
rect 311866 384618 312102 384854
rect 311546 348938 311782 349174
rect 311866 348938 312102 349174
rect 311546 348618 311782 348854
rect 311866 348618 312102 348854
rect 311546 312938 311782 313174
rect 311866 312938 312102 313174
rect 311546 312618 311782 312854
rect 311866 312618 312102 312854
rect 311546 276938 311782 277174
rect 311866 276938 312102 277174
rect 311546 276618 311782 276854
rect 311866 276618 312102 276854
rect 311546 240938 311782 241174
rect 311866 240938 312102 241174
rect 311546 240618 311782 240854
rect 311866 240618 312102 240854
rect 311546 204938 311782 205174
rect 311866 204938 312102 205174
rect 311546 204618 311782 204854
rect 311866 204618 312102 204854
rect 311546 168938 311782 169174
rect 311866 168938 312102 169174
rect 311546 168618 311782 168854
rect 311866 168618 312102 168854
rect 311546 132938 311782 133174
rect 311866 132938 312102 133174
rect 311546 132618 311782 132854
rect 311866 132618 312102 132854
rect 311546 96938 311782 97174
rect 311866 96938 312102 97174
rect 311546 96618 311782 96854
rect 311866 96618 312102 96854
rect 311546 60938 311782 61174
rect 311866 60938 312102 61174
rect 311546 60618 311782 60854
rect 311866 60618 312102 60854
rect 311546 24938 311782 25174
rect 311866 24938 312102 25174
rect 311546 24618 311782 24854
rect 311866 24618 312102 24854
rect 311546 -3462 311782 -3226
rect 311866 -3462 312102 -3226
rect 311546 -3782 311782 -3546
rect 311866 -3782 312102 -3546
rect 315266 676658 315502 676894
rect 315586 676658 315822 676894
rect 315266 676338 315502 676574
rect 315586 676338 315822 676574
rect 315266 640658 315502 640894
rect 315586 640658 315822 640894
rect 315266 640338 315502 640574
rect 315586 640338 315822 640574
rect 315266 604658 315502 604894
rect 315586 604658 315822 604894
rect 315266 604338 315502 604574
rect 315586 604338 315822 604574
rect 315266 568658 315502 568894
rect 315586 568658 315822 568894
rect 315266 568338 315502 568574
rect 315586 568338 315822 568574
rect 315266 532658 315502 532894
rect 315586 532658 315822 532894
rect 315266 532338 315502 532574
rect 315586 532338 315822 532574
rect 315266 496658 315502 496894
rect 315586 496658 315822 496894
rect 315266 496338 315502 496574
rect 315586 496338 315822 496574
rect 315266 460658 315502 460894
rect 315586 460658 315822 460894
rect 315266 460338 315502 460574
rect 315586 460338 315822 460574
rect 315266 424658 315502 424894
rect 315586 424658 315822 424894
rect 315266 424338 315502 424574
rect 315586 424338 315822 424574
rect 315266 388658 315502 388894
rect 315586 388658 315822 388894
rect 315266 388338 315502 388574
rect 315586 388338 315822 388574
rect 315266 352658 315502 352894
rect 315586 352658 315822 352894
rect 315266 352338 315502 352574
rect 315586 352338 315822 352574
rect 315266 316658 315502 316894
rect 315586 316658 315822 316894
rect 315266 316338 315502 316574
rect 315586 316338 315822 316574
rect 315266 280658 315502 280894
rect 315586 280658 315822 280894
rect 315266 280338 315502 280574
rect 315586 280338 315822 280574
rect 315266 244658 315502 244894
rect 315586 244658 315822 244894
rect 315266 244338 315502 244574
rect 315586 244338 315822 244574
rect 315266 208658 315502 208894
rect 315586 208658 315822 208894
rect 315266 208338 315502 208574
rect 315586 208338 315822 208574
rect 315266 172658 315502 172894
rect 315586 172658 315822 172894
rect 315266 172338 315502 172574
rect 315586 172338 315822 172574
rect 315266 136658 315502 136894
rect 315586 136658 315822 136894
rect 315266 136338 315502 136574
rect 315586 136338 315822 136574
rect 315266 100658 315502 100894
rect 315586 100658 315822 100894
rect 315266 100338 315502 100574
rect 315586 100338 315822 100574
rect 315266 64658 315502 64894
rect 315586 64658 315822 64894
rect 315266 64338 315502 64574
rect 315586 64338 315822 64574
rect 315266 28658 315502 28894
rect 315586 28658 315822 28894
rect 315266 28338 315502 28574
rect 315586 28338 315822 28574
rect 315266 -5382 315502 -5146
rect 315586 -5382 315822 -5146
rect 315266 -5702 315502 -5466
rect 315586 -5702 315822 -5466
rect 336986 710362 337222 710598
rect 337306 710362 337542 710598
rect 336986 710042 337222 710278
rect 337306 710042 337542 710278
rect 333266 708442 333502 708678
rect 333586 708442 333822 708678
rect 333266 708122 333502 708358
rect 333586 708122 333822 708358
rect 329546 706522 329782 706758
rect 329866 706522 330102 706758
rect 329546 706202 329782 706438
rect 329866 706202 330102 706438
rect 318986 680378 319222 680614
rect 319306 680378 319542 680614
rect 318986 680058 319222 680294
rect 319306 680058 319542 680294
rect 318986 644378 319222 644614
rect 319306 644378 319542 644614
rect 318986 644058 319222 644294
rect 319306 644058 319542 644294
rect 318986 608378 319222 608614
rect 319306 608378 319542 608614
rect 318986 608058 319222 608294
rect 319306 608058 319542 608294
rect 318986 572378 319222 572614
rect 319306 572378 319542 572614
rect 318986 572058 319222 572294
rect 319306 572058 319542 572294
rect 318986 536378 319222 536614
rect 319306 536378 319542 536614
rect 318986 536058 319222 536294
rect 319306 536058 319542 536294
rect 318986 500378 319222 500614
rect 319306 500378 319542 500614
rect 318986 500058 319222 500294
rect 319306 500058 319542 500294
rect 318986 464378 319222 464614
rect 319306 464378 319542 464614
rect 318986 464058 319222 464294
rect 319306 464058 319542 464294
rect 318986 428378 319222 428614
rect 319306 428378 319542 428614
rect 318986 428058 319222 428294
rect 319306 428058 319542 428294
rect 318986 392378 319222 392614
rect 319306 392378 319542 392614
rect 318986 392058 319222 392294
rect 319306 392058 319542 392294
rect 318986 356378 319222 356614
rect 319306 356378 319542 356614
rect 318986 356058 319222 356294
rect 319306 356058 319542 356294
rect 318986 320378 319222 320614
rect 319306 320378 319542 320614
rect 318986 320058 319222 320294
rect 319306 320058 319542 320294
rect 318986 284378 319222 284614
rect 319306 284378 319542 284614
rect 318986 284058 319222 284294
rect 319306 284058 319542 284294
rect 318986 248378 319222 248614
rect 319306 248378 319542 248614
rect 318986 248058 319222 248294
rect 319306 248058 319542 248294
rect 318986 212378 319222 212614
rect 319306 212378 319542 212614
rect 318986 212058 319222 212294
rect 319306 212058 319542 212294
rect 318986 176378 319222 176614
rect 319306 176378 319542 176614
rect 318986 176058 319222 176294
rect 319306 176058 319542 176294
rect 318986 140378 319222 140614
rect 319306 140378 319542 140614
rect 318986 140058 319222 140294
rect 319306 140058 319542 140294
rect 318986 104378 319222 104614
rect 319306 104378 319542 104614
rect 318986 104058 319222 104294
rect 319306 104058 319542 104294
rect 318986 68378 319222 68614
rect 319306 68378 319542 68614
rect 318986 68058 319222 68294
rect 319306 68058 319542 68294
rect 318986 32378 319222 32614
rect 319306 32378 319542 32614
rect 318986 32058 319222 32294
rect 319306 32058 319542 32294
rect 300986 -6342 301222 -6106
rect 301306 -6342 301542 -6106
rect 300986 -6662 301222 -6426
rect 301306 -6662 301542 -6426
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 325826 543218 326062 543454
rect 326146 543218 326382 543454
rect 325826 542898 326062 543134
rect 326146 542898 326382 543134
rect 325826 507218 326062 507454
rect 326146 507218 326382 507454
rect 325826 506898 326062 507134
rect 326146 506898 326382 507134
rect 325826 471218 326062 471454
rect 326146 471218 326382 471454
rect 325826 470898 326062 471134
rect 326146 470898 326382 471134
rect 325826 435218 326062 435454
rect 326146 435218 326382 435454
rect 325826 434898 326062 435134
rect 326146 434898 326382 435134
rect 325826 399218 326062 399454
rect 326146 399218 326382 399454
rect 325826 398898 326062 399134
rect 326146 398898 326382 399134
rect 325826 363218 326062 363454
rect 326146 363218 326382 363454
rect 325826 362898 326062 363134
rect 326146 362898 326382 363134
rect 325826 327218 326062 327454
rect 326146 327218 326382 327454
rect 325826 326898 326062 327134
rect 326146 326898 326382 327134
rect 325826 291218 326062 291454
rect 326146 291218 326382 291454
rect 325826 290898 326062 291134
rect 326146 290898 326382 291134
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 325826 219218 326062 219454
rect 326146 219218 326382 219454
rect 325826 218898 326062 219134
rect 326146 218898 326382 219134
rect 325826 183218 326062 183454
rect 326146 183218 326382 183454
rect 325826 182898 326062 183134
rect 326146 182898 326382 183134
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 325826 111218 326062 111454
rect 326146 111218 326382 111454
rect 325826 110898 326062 111134
rect 326146 110898 326382 111134
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 690938 329782 691174
rect 329866 690938 330102 691174
rect 329546 690618 329782 690854
rect 329866 690618 330102 690854
rect 329546 654938 329782 655174
rect 329866 654938 330102 655174
rect 329546 654618 329782 654854
rect 329866 654618 330102 654854
rect 329546 618938 329782 619174
rect 329866 618938 330102 619174
rect 329546 618618 329782 618854
rect 329866 618618 330102 618854
rect 329546 582938 329782 583174
rect 329866 582938 330102 583174
rect 329546 582618 329782 582854
rect 329866 582618 330102 582854
rect 329546 546938 329782 547174
rect 329866 546938 330102 547174
rect 329546 546618 329782 546854
rect 329866 546618 330102 546854
rect 329546 510938 329782 511174
rect 329866 510938 330102 511174
rect 329546 510618 329782 510854
rect 329866 510618 330102 510854
rect 329546 474938 329782 475174
rect 329866 474938 330102 475174
rect 329546 474618 329782 474854
rect 329866 474618 330102 474854
rect 329546 438938 329782 439174
rect 329866 438938 330102 439174
rect 329546 438618 329782 438854
rect 329866 438618 330102 438854
rect 329546 402938 329782 403174
rect 329866 402938 330102 403174
rect 329546 402618 329782 402854
rect 329866 402618 330102 402854
rect 329546 366938 329782 367174
rect 329866 366938 330102 367174
rect 329546 366618 329782 366854
rect 329866 366618 330102 366854
rect 329546 330938 329782 331174
rect 329866 330938 330102 331174
rect 329546 330618 329782 330854
rect 329866 330618 330102 330854
rect 329546 294938 329782 295174
rect 329866 294938 330102 295174
rect 329546 294618 329782 294854
rect 329866 294618 330102 294854
rect 329546 258938 329782 259174
rect 329866 258938 330102 259174
rect 329546 258618 329782 258854
rect 329866 258618 330102 258854
rect 329546 222938 329782 223174
rect 329866 222938 330102 223174
rect 329546 222618 329782 222854
rect 329866 222618 330102 222854
rect 329546 186938 329782 187174
rect 329866 186938 330102 187174
rect 329546 186618 329782 186854
rect 329866 186618 330102 186854
rect 329546 150938 329782 151174
rect 329866 150938 330102 151174
rect 329546 150618 329782 150854
rect 329866 150618 330102 150854
rect 329546 114938 329782 115174
rect 329866 114938 330102 115174
rect 329546 114618 329782 114854
rect 329866 114618 330102 114854
rect 329546 78938 329782 79174
rect 329866 78938 330102 79174
rect 329546 78618 329782 78854
rect 329866 78618 330102 78854
rect 329546 42938 329782 43174
rect 329866 42938 330102 43174
rect 329546 42618 329782 42854
rect 329866 42618 330102 42854
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 329546 -2502 329782 -2266
rect 329866 -2502 330102 -2266
rect 329546 -2822 329782 -2586
rect 329866 -2822 330102 -2586
rect 333266 694658 333502 694894
rect 333586 694658 333822 694894
rect 333266 694338 333502 694574
rect 333586 694338 333822 694574
rect 333266 658658 333502 658894
rect 333586 658658 333822 658894
rect 333266 658338 333502 658574
rect 333586 658338 333822 658574
rect 333266 622658 333502 622894
rect 333586 622658 333822 622894
rect 333266 622338 333502 622574
rect 333586 622338 333822 622574
rect 333266 586658 333502 586894
rect 333586 586658 333822 586894
rect 333266 586338 333502 586574
rect 333586 586338 333822 586574
rect 333266 550658 333502 550894
rect 333586 550658 333822 550894
rect 333266 550338 333502 550574
rect 333586 550338 333822 550574
rect 333266 514658 333502 514894
rect 333586 514658 333822 514894
rect 333266 514338 333502 514574
rect 333586 514338 333822 514574
rect 333266 478658 333502 478894
rect 333586 478658 333822 478894
rect 333266 478338 333502 478574
rect 333586 478338 333822 478574
rect 333266 442658 333502 442894
rect 333586 442658 333822 442894
rect 333266 442338 333502 442574
rect 333586 442338 333822 442574
rect 333266 406658 333502 406894
rect 333586 406658 333822 406894
rect 333266 406338 333502 406574
rect 333586 406338 333822 406574
rect 333266 370658 333502 370894
rect 333586 370658 333822 370894
rect 333266 370338 333502 370574
rect 333586 370338 333822 370574
rect 333266 334658 333502 334894
rect 333586 334658 333822 334894
rect 333266 334338 333502 334574
rect 333586 334338 333822 334574
rect 333266 298658 333502 298894
rect 333586 298658 333822 298894
rect 333266 298338 333502 298574
rect 333586 298338 333822 298574
rect 333266 262658 333502 262894
rect 333586 262658 333822 262894
rect 333266 262338 333502 262574
rect 333586 262338 333822 262574
rect 333266 226658 333502 226894
rect 333586 226658 333822 226894
rect 333266 226338 333502 226574
rect 333586 226338 333822 226574
rect 333266 190658 333502 190894
rect 333586 190658 333822 190894
rect 333266 190338 333502 190574
rect 333586 190338 333822 190574
rect 333266 154658 333502 154894
rect 333586 154658 333822 154894
rect 333266 154338 333502 154574
rect 333586 154338 333822 154574
rect 333266 118658 333502 118894
rect 333586 118658 333822 118894
rect 333266 118338 333502 118574
rect 333586 118338 333822 118574
rect 333266 82658 333502 82894
rect 333586 82658 333822 82894
rect 333266 82338 333502 82574
rect 333586 82338 333822 82574
rect 333266 46658 333502 46894
rect 333586 46658 333822 46894
rect 333266 46338 333502 46574
rect 333586 46338 333822 46574
rect 333266 10658 333502 10894
rect 333586 10658 333822 10894
rect 333266 10338 333502 10574
rect 333586 10338 333822 10574
rect 333266 -4422 333502 -4186
rect 333586 -4422 333822 -4186
rect 333266 -4742 333502 -4506
rect 333586 -4742 333822 -4506
rect 354986 711322 355222 711558
rect 355306 711322 355542 711558
rect 354986 711002 355222 711238
rect 355306 711002 355542 711238
rect 351266 709402 351502 709638
rect 351586 709402 351822 709638
rect 351266 709082 351502 709318
rect 351586 709082 351822 709318
rect 347546 707482 347782 707718
rect 347866 707482 348102 707718
rect 347546 707162 347782 707398
rect 347866 707162 348102 707398
rect 336986 698378 337222 698614
rect 337306 698378 337542 698614
rect 336986 698058 337222 698294
rect 337306 698058 337542 698294
rect 336986 662378 337222 662614
rect 337306 662378 337542 662614
rect 336986 662058 337222 662294
rect 337306 662058 337542 662294
rect 336986 626378 337222 626614
rect 337306 626378 337542 626614
rect 336986 626058 337222 626294
rect 337306 626058 337542 626294
rect 336986 590378 337222 590614
rect 337306 590378 337542 590614
rect 336986 590058 337222 590294
rect 337306 590058 337542 590294
rect 336986 554378 337222 554614
rect 337306 554378 337542 554614
rect 336986 554058 337222 554294
rect 337306 554058 337542 554294
rect 336986 518378 337222 518614
rect 337306 518378 337542 518614
rect 336986 518058 337222 518294
rect 337306 518058 337542 518294
rect 336986 482378 337222 482614
rect 337306 482378 337542 482614
rect 336986 482058 337222 482294
rect 337306 482058 337542 482294
rect 336986 446378 337222 446614
rect 337306 446378 337542 446614
rect 336986 446058 337222 446294
rect 337306 446058 337542 446294
rect 336986 410378 337222 410614
rect 337306 410378 337542 410614
rect 336986 410058 337222 410294
rect 337306 410058 337542 410294
rect 336986 374378 337222 374614
rect 337306 374378 337542 374614
rect 336986 374058 337222 374294
rect 337306 374058 337542 374294
rect 336986 338378 337222 338614
rect 337306 338378 337542 338614
rect 336986 338058 337222 338294
rect 337306 338058 337542 338294
rect 336986 302378 337222 302614
rect 337306 302378 337542 302614
rect 336986 302058 337222 302294
rect 337306 302058 337542 302294
rect 336986 266378 337222 266614
rect 337306 266378 337542 266614
rect 336986 266058 337222 266294
rect 337306 266058 337542 266294
rect 336986 230378 337222 230614
rect 337306 230378 337542 230614
rect 336986 230058 337222 230294
rect 337306 230058 337542 230294
rect 336986 194378 337222 194614
rect 337306 194378 337542 194614
rect 336986 194058 337222 194294
rect 337306 194058 337542 194294
rect 336986 158378 337222 158614
rect 337306 158378 337542 158614
rect 336986 158058 337222 158294
rect 337306 158058 337542 158294
rect 336986 122378 337222 122614
rect 337306 122378 337542 122614
rect 336986 122058 337222 122294
rect 337306 122058 337542 122294
rect 336986 86378 337222 86614
rect 337306 86378 337542 86614
rect 336986 86058 337222 86294
rect 337306 86058 337542 86294
rect 336986 50378 337222 50614
rect 337306 50378 337542 50614
rect 336986 50058 337222 50294
rect 337306 50058 337542 50294
rect 336986 14378 337222 14614
rect 337306 14378 337542 14614
rect 336986 14058 337222 14294
rect 337306 14058 337542 14294
rect 318986 -7302 319222 -7066
rect 319306 -7302 319542 -7066
rect 318986 -7622 319222 -7386
rect 319306 -7622 319542 -7386
rect 343826 705562 344062 705798
rect 344146 705562 344382 705798
rect 343826 705242 344062 705478
rect 344146 705242 344382 705478
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 343826 561218 344062 561454
rect 344146 561218 344382 561454
rect 343826 560898 344062 561134
rect 344146 560898 344382 561134
rect 343826 525218 344062 525454
rect 344146 525218 344382 525454
rect 343826 524898 344062 525134
rect 344146 524898 344382 525134
rect 343826 489218 344062 489454
rect 344146 489218 344382 489454
rect 343826 488898 344062 489134
rect 344146 488898 344382 489134
rect 343826 453218 344062 453454
rect 344146 453218 344382 453454
rect 343826 452898 344062 453134
rect 344146 452898 344382 453134
rect 343826 417218 344062 417454
rect 344146 417218 344382 417454
rect 343826 416898 344062 417134
rect 344146 416898 344382 417134
rect 343826 381218 344062 381454
rect 344146 381218 344382 381454
rect 343826 380898 344062 381134
rect 344146 380898 344382 381134
rect 343826 345218 344062 345454
rect 344146 345218 344382 345454
rect 343826 344898 344062 345134
rect 344146 344898 344382 345134
rect 343826 309218 344062 309454
rect 344146 309218 344382 309454
rect 343826 308898 344062 309134
rect 344146 308898 344382 309134
rect 343826 273218 344062 273454
rect 344146 273218 344382 273454
rect 343826 272898 344062 273134
rect 344146 272898 344382 273134
rect 343826 237218 344062 237454
rect 344146 237218 344382 237454
rect 343826 236898 344062 237134
rect 344146 236898 344382 237134
rect 343826 201218 344062 201454
rect 344146 201218 344382 201454
rect 343826 200898 344062 201134
rect 344146 200898 344382 201134
rect 343826 165218 344062 165454
rect 344146 165218 344382 165454
rect 343826 164898 344062 165134
rect 344146 164898 344382 165134
rect 343826 129218 344062 129454
rect 344146 129218 344382 129454
rect 343826 128898 344062 129134
rect 344146 128898 344382 129134
rect 343826 93218 344062 93454
rect 344146 93218 344382 93454
rect 343826 92898 344062 93134
rect 344146 92898 344382 93134
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -1542 344062 -1306
rect 344146 -1542 344382 -1306
rect 343826 -1862 344062 -1626
rect 344146 -1862 344382 -1626
rect 347546 672938 347782 673174
rect 347866 672938 348102 673174
rect 347546 672618 347782 672854
rect 347866 672618 348102 672854
rect 347546 636938 347782 637174
rect 347866 636938 348102 637174
rect 347546 636618 347782 636854
rect 347866 636618 348102 636854
rect 347546 600938 347782 601174
rect 347866 600938 348102 601174
rect 347546 600618 347782 600854
rect 347866 600618 348102 600854
rect 347546 564938 347782 565174
rect 347866 564938 348102 565174
rect 347546 564618 347782 564854
rect 347866 564618 348102 564854
rect 347546 528938 347782 529174
rect 347866 528938 348102 529174
rect 347546 528618 347782 528854
rect 347866 528618 348102 528854
rect 347546 492938 347782 493174
rect 347866 492938 348102 493174
rect 347546 492618 347782 492854
rect 347866 492618 348102 492854
rect 347546 456938 347782 457174
rect 347866 456938 348102 457174
rect 347546 456618 347782 456854
rect 347866 456618 348102 456854
rect 347546 420938 347782 421174
rect 347866 420938 348102 421174
rect 347546 420618 347782 420854
rect 347866 420618 348102 420854
rect 347546 384938 347782 385174
rect 347866 384938 348102 385174
rect 347546 384618 347782 384854
rect 347866 384618 348102 384854
rect 347546 348938 347782 349174
rect 347866 348938 348102 349174
rect 347546 348618 347782 348854
rect 347866 348618 348102 348854
rect 347546 312938 347782 313174
rect 347866 312938 348102 313174
rect 347546 312618 347782 312854
rect 347866 312618 348102 312854
rect 347546 276938 347782 277174
rect 347866 276938 348102 277174
rect 347546 276618 347782 276854
rect 347866 276618 348102 276854
rect 347546 240938 347782 241174
rect 347866 240938 348102 241174
rect 347546 240618 347782 240854
rect 347866 240618 348102 240854
rect 347546 204938 347782 205174
rect 347866 204938 348102 205174
rect 347546 204618 347782 204854
rect 347866 204618 348102 204854
rect 347546 168938 347782 169174
rect 347866 168938 348102 169174
rect 347546 168618 347782 168854
rect 347866 168618 348102 168854
rect 347546 132938 347782 133174
rect 347866 132938 348102 133174
rect 347546 132618 347782 132854
rect 347866 132618 348102 132854
rect 347546 96938 347782 97174
rect 347866 96938 348102 97174
rect 347546 96618 347782 96854
rect 347866 96618 348102 96854
rect 347546 60938 347782 61174
rect 347866 60938 348102 61174
rect 347546 60618 347782 60854
rect 347866 60618 348102 60854
rect 347546 24938 347782 25174
rect 347866 24938 348102 25174
rect 347546 24618 347782 24854
rect 347866 24618 348102 24854
rect 347546 -3462 347782 -3226
rect 347866 -3462 348102 -3226
rect 347546 -3782 347782 -3546
rect 347866 -3782 348102 -3546
rect 351266 676658 351502 676894
rect 351586 676658 351822 676894
rect 351266 676338 351502 676574
rect 351586 676338 351822 676574
rect 351266 640658 351502 640894
rect 351586 640658 351822 640894
rect 351266 640338 351502 640574
rect 351586 640338 351822 640574
rect 351266 604658 351502 604894
rect 351586 604658 351822 604894
rect 351266 604338 351502 604574
rect 351586 604338 351822 604574
rect 351266 568658 351502 568894
rect 351586 568658 351822 568894
rect 351266 568338 351502 568574
rect 351586 568338 351822 568574
rect 351266 532658 351502 532894
rect 351586 532658 351822 532894
rect 351266 532338 351502 532574
rect 351586 532338 351822 532574
rect 351266 496658 351502 496894
rect 351586 496658 351822 496894
rect 351266 496338 351502 496574
rect 351586 496338 351822 496574
rect 351266 460658 351502 460894
rect 351586 460658 351822 460894
rect 351266 460338 351502 460574
rect 351586 460338 351822 460574
rect 351266 424658 351502 424894
rect 351586 424658 351822 424894
rect 351266 424338 351502 424574
rect 351586 424338 351822 424574
rect 351266 388658 351502 388894
rect 351586 388658 351822 388894
rect 351266 388338 351502 388574
rect 351586 388338 351822 388574
rect 351266 352658 351502 352894
rect 351586 352658 351822 352894
rect 351266 352338 351502 352574
rect 351586 352338 351822 352574
rect 351266 316658 351502 316894
rect 351586 316658 351822 316894
rect 351266 316338 351502 316574
rect 351586 316338 351822 316574
rect 351266 280658 351502 280894
rect 351586 280658 351822 280894
rect 351266 280338 351502 280574
rect 351586 280338 351822 280574
rect 351266 244658 351502 244894
rect 351586 244658 351822 244894
rect 351266 244338 351502 244574
rect 351586 244338 351822 244574
rect 351266 208658 351502 208894
rect 351586 208658 351822 208894
rect 351266 208338 351502 208574
rect 351586 208338 351822 208574
rect 351266 172658 351502 172894
rect 351586 172658 351822 172894
rect 351266 172338 351502 172574
rect 351586 172338 351822 172574
rect 351266 136658 351502 136894
rect 351586 136658 351822 136894
rect 351266 136338 351502 136574
rect 351586 136338 351822 136574
rect 351266 100658 351502 100894
rect 351586 100658 351822 100894
rect 351266 100338 351502 100574
rect 351586 100338 351822 100574
rect 351266 64658 351502 64894
rect 351586 64658 351822 64894
rect 351266 64338 351502 64574
rect 351586 64338 351822 64574
rect 351266 28658 351502 28894
rect 351586 28658 351822 28894
rect 351266 28338 351502 28574
rect 351586 28338 351822 28574
rect 351266 -5382 351502 -5146
rect 351586 -5382 351822 -5146
rect 351266 -5702 351502 -5466
rect 351586 -5702 351822 -5466
rect 372986 710362 373222 710598
rect 373306 710362 373542 710598
rect 372986 710042 373222 710278
rect 373306 710042 373542 710278
rect 369266 708442 369502 708678
rect 369586 708442 369822 708678
rect 369266 708122 369502 708358
rect 369586 708122 369822 708358
rect 365546 706522 365782 706758
rect 365866 706522 366102 706758
rect 365546 706202 365782 706438
rect 365866 706202 366102 706438
rect 354986 680378 355222 680614
rect 355306 680378 355542 680614
rect 354986 680058 355222 680294
rect 355306 680058 355542 680294
rect 354986 644378 355222 644614
rect 355306 644378 355542 644614
rect 354986 644058 355222 644294
rect 355306 644058 355542 644294
rect 354986 608378 355222 608614
rect 355306 608378 355542 608614
rect 354986 608058 355222 608294
rect 355306 608058 355542 608294
rect 354986 572378 355222 572614
rect 355306 572378 355542 572614
rect 354986 572058 355222 572294
rect 355306 572058 355542 572294
rect 354986 536378 355222 536614
rect 355306 536378 355542 536614
rect 354986 536058 355222 536294
rect 355306 536058 355542 536294
rect 354986 500378 355222 500614
rect 355306 500378 355542 500614
rect 354986 500058 355222 500294
rect 355306 500058 355542 500294
rect 354986 464378 355222 464614
rect 355306 464378 355542 464614
rect 354986 464058 355222 464294
rect 355306 464058 355542 464294
rect 354986 428378 355222 428614
rect 355306 428378 355542 428614
rect 354986 428058 355222 428294
rect 355306 428058 355542 428294
rect 354986 392378 355222 392614
rect 355306 392378 355542 392614
rect 354986 392058 355222 392294
rect 355306 392058 355542 392294
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 361826 435218 362062 435454
rect 362146 435218 362382 435454
rect 361826 434898 362062 435134
rect 362146 434898 362382 435134
rect 361826 399218 362062 399454
rect 362146 399218 362382 399454
rect 361826 398898 362062 399134
rect 362146 398898 362382 399134
rect 365546 690938 365782 691174
rect 365866 690938 366102 691174
rect 365546 690618 365782 690854
rect 365866 690618 366102 690854
rect 365546 654938 365782 655174
rect 365866 654938 366102 655174
rect 365546 654618 365782 654854
rect 365866 654618 366102 654854
rect 365546 618938 365782 619174
rect 365866 618938 366102 619174
rect 365546 618618 365782 618854
rect 365866 618618 366102 618854
rect 365546 582938 365782 583174
rect 365866 582938 366102 583174
rect 365546 582618 365782 582854
rect 365866 582618 366102 582854
rect 365546 546938 365782 547174
rect 365866 546938 366102 547174
rect 365546 546618 365782 546854
rect 365866 546618 366102 546854
rect 365546 510938 365782 511174
rect 365866 510938 366102 511174
rect 365546 510618 365782 510854
rect 365866 510618 366102 510854
rect 365546 474938 365782 475174
rect 365866 474938 366102 475174
rect 365546 474618 365782 474854
rect 365866 474618 366102 474854
rect 365546 438938 365782 439174
rect 365866 438938 366102 439174
rect 365546 438618 365782 438854
rect 365866 438618 366102 438854
rect 365546 402938 365782 403174
rect 365866 402938 366102 403174
rect 365546 402618 365782 402854
rect 365866 402618 366102 402854
rect 369266 694658 369502 694894
rect 369586 694658 369822 694894
rect 369266 694338 369502 694574
rect 369586 694338 369822 694574
rect 369266 658658 369502 658894
rect 369586 658658 369822 658894
rect 369266 658338 369502 658574
rect 369586 658338 369822 658574
rect 369266 622658 369502 622894
rect 369586 622658 369822 622894
rect 369266 622338 369502 622574
rect 369586 622338 369822 622574
rect 369266 586658 369502 586894
rect 369586 586658 369822 586894
rect 369266 586338 369502 586574
rect 369586 586338 369822 586574
rect 369266 550658 369502 550894
rect 369586 550658 369822 550894
rect 369266 550338 369502 550574
rect 369586 550338 369822 550574
rect 369266 514658 369502 514894
rect 369586 514658 369822 514894
rect 369266 514338 369502 514574
rect 369586 514338 369822 514574
rect 369266 478658 369502 478894
rect 369586 478658 369822 478894
rect 369266 478338 369502 478574
rect 369586 478338 369822 478574
rect 369266 442658 369502 442894
rect 369586 442658 369822 442894
rect 369266 442338 369502 442574
rect 369586 442338 369822 442574
rect 369266 406658 369502 406894
rect 369586 406658 369822 406894
rect 369266 406338 369502 406574
rect 369586 406338 369822 406574
rect 390986 711322 391222 711558
rect 391306 711322 391542 711558
rect 390986 711002 391222 711238
rect 391306 711002 391542 711238
rect 387266 709402 387502 709638
rect 387586 709402 387822 709638
rect 387266 709082 387502 709318
rect 387586 709082 387822 709318
rect 383546 707482 383782 707718
rect 383866 707482 384102 707718
rect 383546 707162 383782 707398
rect 383866 707162 384102 707398
rect 372986 698378 373222 698614
rect 373306 698378 373542 698614
rect 372986 698058 373222 698294
rect 373306 698058 373542 698294
rect 372986 662378 373222 662614
rect 373306 662378 373542 662614
rect 372986 662058 373222 662294
rect 373306 662058 373542 662294
rect 372986 626378 373222 626614
rect 373306 626378 373542 626614
rect 372986 626058 373222 626294
rect 373306 626058 373542 626294
rect 372986 590378 373222 590614
rect 373306 590378 373542 590614
rect 372986 590058 373222 590294
rect 373306 590058 373542 590294
rect 372986 554378 373222 554614
rect 373306 554378 373542 554614
rect 372986 554058 373222 554294
rect 373306 554058 373542 554294
rect 372986 518378 373222 518614
rect 373306 518378 373542 518614
rect 372986 518058 373222 518294
rect 373306 518058 373542 518294
rect 372986 482378 373222 482614
rect 373306 482378 373542 482614
rect 372986 482058 373222 482294
rect 373306 482058 373542 482294
rect 372986 446378 373222 446614
rect 373306 446378 373542 446614
rect 372986 446058 373222 446294
rect 373306 446058 373542 446294
rect 372986 410378 373222 410614
rect 373306 410378 373542 410614
rect 372986 410058 373222 410294
rect 373306 410058 373542 410294
rect 372986 374378 373222 374614
rect 373306 374378 373542 374614
rect 372986 374058 373222 374294
rect 373306 374058 373542 374294
rect 362285 363218 362521 363454
rect 362285 362898 362521 363134
rect 364882 363218 365118 363454
rect 364882 362898 365118 363134
rect 367479 363218 367715 363454
rect 367479 362898 367715 363134
rect 354986 356378 355222 356614
rect 355306 356378 355542 356614
rect 354986 356058 355222 356294
rect 355306 356058 355542 356294
rect 363583 345218 363819 345454
rect 363583 344898 363819 345134
rect 366180 345218 366416 345454
rect 366180 344898 366416 345134
rect 354986 320378 355222 320614
rect 355306 320378 355542 320614
rect 354986 320058 355222 320294
rect 355306 320058 355542 320294
rect 354986 284378 355222 284614
rect 355306 284378 355542 284614
rect 354986 284058 355222 284294
rect 355306 284058 355542 284294
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 362285 291218 362521 291454
rect 362285 290898 362521 291134
rect 363583 273218 363819 273454
rect 363583 272898 363819 273134
rect 365546 330938 365782 331174
rect 365866 330938 366102 331174
rect 365546 330618 365782 330854
rect 365866 330618 366102 330854
rect 369266 334658 369502 334894
rect 369586 334658 369822 334894
rect 369266 334338 369502 334574
rect 369586 334338 369822 334574
rect 364882 291218 365118 291454
rect 364882 290898 365118 291134
rect 367479 291218 367715 291454
rect 367479 290898 367715 291134
rect 366180 273218 366416 273454
rect 366180 272898 366416 273134
rect 354986 248378 355222 248614
rect 355306 248378 355542 248614
rect 354986 248058 355222 248294
rect 355306 248058 355542 248294
rect 354986 212378 355222 212614
rect 355306 212378 355542 212614
rect 354986 212058 355222 212294
rect 355306 212058 355542 212294
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 362285 219218 362521 219454
rect 362285 218898 362521 219134
rect 363583 201218 363819 201454
rect 363583 200898 363819 201134
rect 365546 258938 365782 259174
rect 365866 258938 366102 259174
rect 365546 258618 365782 258854
rect 365866 258618 366102 258854
rect 369266 262658 369502 262894
rect 369586 262658 369822 262894
rect 369266 262338 369502 262574
rect 369586 262338 369822 262574
rect 364882 219218 365118 219454
rect 364882 218898 365118 219134
rect 367479 219218 367715 219454
rect 367479 218898 367715 219134
rect 372986 338378 373222 338614
rect 373306 338378 373542 338614
rect 372986 338058 373222 338294
rect 373306 338058 373542 338294
rect 372986 302378 373222 302614
rect 373306 302378 373542 302614
rect 372986 302058 373222 302294
rect 373306 302058 373542 302294
rect 372986 266378 373222 266614
rect 373306 266378 373542 266614
rect 372986 266058 373222 266294
rect 373306 266058 373542 266294
rect 372986 230378 373222 230614
rect 373306 230378 373542 230614
rect 372986 230058 373222 230294
rect 373306 230058 373542 230294
rect 366180 201218 366416 201454
rect 366180 200898 366416 201134
rect 354986 176378 355222 176614
rect 355306 176378 355542 176614
rect 354986 176058 355222 176294
rect 355306 176058 355542 176294
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 362285 147218 362521 147454
rect 362285 146898 362521 147134
rect 354986 140378 355222 140614
rect 355306 140378 355542 140614
rect 354986 140058 355222 140294
rect 355306 140058 355542 140294
rect 364882 147218 365118 147454
rect 364882 146898 365118 147134
rect 363583 129218 363819 129454
rect 363583 128898 363819 129134
rect 365546 186938 365782 187174
rect 365866 186938 366102 187174
rect 365546 186618 365782 186854
rect 365866 186618 366102 186854
rect 369266 190658 369502 190894
rect 369586 190658 369822 190894
rect 369266 190338 369502 190574
rect 369586 190338 369822 190574
rect 367479 147218 367715 147454
rect 367479 146898 367715 147134
rect 372986 194378 373222 194614
rect 373306 194378 373542 194614
rect 372986 194058 373222 194294
rect 373306 194058 373542 194294
rect 372986 158378 373222 158614
rect 373306 158378 373542 158614
rect 372986 158058 373222 158294
rect 373306 158058 373542 158294
rect 366180 129218 366416 129454
rect 366180 128898 366416 129134
rect 372986 122378 373222 122614
rect 373306 122378 373542 122614
rect 372986 122058 373222 122294
rect 373306 122058 373542 122294
rect 354986 104378 355222 104614
rect 355306 104378 355542 104614
rect 354986 104058 355222 104294
rect 355306 104058 355542 104294
rect 354986 68378 355222 68614
rect 355306 68378 355542 68614
rect 354986 68058 355222 68294
rect 355306 68058 355542 68294
rect 354986 32378 355222 32614
rect 355306 32378 355542 32614
rect 354986 32058 355222 32294
rect 355306 32058 355542 32294
rect 336986 -6342 337222 -6106
rect 337306 -6342 337542 -6106
rect 336986 -6662 337222 -6426
rect 337306 -6662 337542 -6426
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 365546 114938 365782 115174
rect 365866 114938 366102 115174
rect 365546 114618 365782 114854
rect 365866 114618 366102 114854
rect 365546 78938 365782 79174
rect 365866 78938 366102 79174
rect 365546 78618 365782 78854
rect 365866 78618 366102 78854
rect 365546 42938 365782 43174
rect 365866 42938 366102 43174
rect 365546 42618 365782 42854
rect 365866 42618 366102 42854
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 365546 -2502 365782 -2266
rect 365866 -2502 366102 -2266
rect 365546 -2822 365782 -2586
rect 365866 -2822 366102 -2586
rect 369266 118658 369502 118894
rect 369586 118658 369822 118894
rect 369266 118338 369502 118574
rect 369586 118338 369822 118574
rect 369266 82658 369502 82894
rect 369586 82658 369822 82894
rect 369266 82338 369502 82574
rect 369586 82338 369822 82574
rect 369266 46658 369502 46894
rect 369586 46658 369822 46894
rect 369266 46338 369502 46574
rect 369586 46338 369822 46574
rect 369266 10658 369502 10894
rect 369586 10658 369822 10894
rect 369266 10338 369502 10574
rect 369586 10338 369822 10574
rect 369266 -4422 369502 -4186
rect 369586 -4422 369822 -4186
rect 369266 -4742 369502 -4506
rect 369586 -4742 369822 -4506
rect 372986 86378 373222 86614
rect 373306 86378 373542 86614
rect 372986 86058 373222 86294
rect 373306 86058 373542 86294
rect 372986 50378 373222 50614
rect 373306 50378 373542 50614
rect 372986 50058 373222 50294
rect 373306 50058 373542 50294
rect 372986 14378 373222 14614
rect 373306 14378 373542 14614
rect 372986 14058 373222 14294
rect 373306 14058 373542 14294
rect 354986 -7302 355222 -7066
rect 355306 -7302 355542 -7066
rect 354986 -7622 355222 -7386
rect 355306 -7622 355542 -7386
rect 379826 705562 380062 705798
rect 380146 705562 380382 705798
rect 379826 705242 380062 705478
rect 380146 705242 380382 705478
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 379826 561218 380062 561454
rect 380146 561218 380382 561454
rect 379826 560898 380062 561134
rect 380146 560898 380382 561134
rect 379826 525218 380062 525454
rect 380146 525218 380382 525454
rect 379826 524898 380062 525134
rect 380146 524898 380382 525134
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 379826 453218 380062 453454
rect 380146 453218 380382 453454
rect 379826 452898 380062 453134
rect 380146 452898 380382 453134
rect 379826 417218 380062 417454
rect 380146 417218 380382 417454
rect 379826 416898 380062 417134
rect 380146 416898 380382 417134
rect 379826 381218 380062 381454
rect 380146 381218 380382 381454
rect 379826 380898 380062 381134
rect 380146 380898 380382 381134
rect 379826 345218 380062 345454
rect 380146 345218 380382 345454
rect 379826 344898 380062 345134
rect 380146 344898 380382 345134
rect 379826 309218 380062 309454
rect 380146 309218 380382 309454
rect 379826 308898 380062 309134
rect 380146 308898 380382 309134
rect 379826 273218 380062 273454
rect 380146 273218 380382 273454
rect 379826 272898 380062 273134
rect 380146 272898 380382 273134
rect 379826 237218 380062 237454
rect 380146 237218 380382 237454
rect 379826 236898 380062 237134
rect 380146 236898 380382 237134
rect 379826 201218 380062 201454
rect 380146 201218 380382 201454
rect 379826 200898 380062 201134
rect 380146 200898 380382 201134
rect 379826 165218 380062 165454
rect 380146 165218 380382 165454
rect 379826 164898 380062 165134
rect 380146 164898 380382 165134
rect 379826 129218 380062 129454
rect 380146 129218 380382 129454
rect 379826 128898 380062 129134
rect 380146 128898 380382 129134
rect 379826 93218 380062 93454
rect 380146 93218 380382 93454
rect 379826 92898 380062 93134
rect 380146 92898 380382 93134
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -1542 380062 -1306
rect 380146 -1542 380382 -1306
rect 379826 -1862 380062 -1626
rect 380146 -1862 380382 -1626
rect 383546 672938 383782 673174
rect 383866 672938 384102 673174
rect 383546 672618 383782 672854
rect 383866 672618 384102 672854
rect 383546 636938 383782 637174
rect 383866 636938 384102 637174
rect 383546 636618 383782 636854
rect 383866 636618 384102 636854
rect 383546 600938 383782 601174
rect 383866 600938 384102 601174
rect 383546 600618 383782 600854
rect 383866 600618 384102 600854
rect 383546 564938 383782 565174
rect 383866 564938 384102 565174
rect 383546 564618 383782 564854
rect 383866 564618 384102 564854
rect 383546 528938 383782 529174
rect 383866 528938 384102 529174
rect 383546 528618 383782 528854
rect 383866 528618 384102 528854
rect 383546 492938 383782 493174
rect 383866 492938 384102 493174
rect 383546 492618 383782 492854
rect 383866 492618 384102 492854
rect 383546 456938 383782 457174
rect 383866 456938 384102 457174
rect 383546 456618 383782 456854
rect 383866 456618 384102 456854
rect 383546 420938 383782 421174
rect 383866 420938 384102 421174
rect 383546 420618 383782 420854
rect 383866 420618 384102 420854
rect 383546 384938 383782 385174
rect 383866 384938 384102 385174
rect 383546 384618 383782 384854
rect 383866 384618 384102 384854
rect 383546 348938 383782 349174
rect 383866 348938 384102 349174
rect 383546 348618 383782 348854
rect 383866 348618 384102 348854
rect 383546 312938 383782 313174
rect 383866 312938 384102 313174
rect 383546 312618 383782 312854
rect 383866 312618 384102 312854
rect 383546 276938 383782 277174
rect 383866 276938 384102 277174
rect 383546 276618 383782 276854
rect 383866 276618 384102 276854
rect 383546 240938 383782 241174
rect 383866 240938 384102 241174
rect 383546 240618 383782 240854
rect 383866 240618 384102 240854
rect 383546 204938 383782 205174
rect 383866 204938 384102 205174
rect 383546 204618 383782 204854
rect 383866 204618 384102 204854
rect 383546 168938 383782 169174
rect 383866 168938 384102 169174
rect 383546 168618 383782 168854
rect 383866 168618 384102 168854
rect 383546 132938 383782 133174
rect 383866 132938 384102 133174
rect 383546 132618 383782 132854
rect 383866 132618 384102 132854
rect 383546 96938 383782 97174
rect 383866 96938 384102 97174
rect 383546 96618 383782 96854
rect 383866 96618 384102 96854
rect 383546 60938 383782 61174
rect 383866 60938 384102 61174
rect 383546 60618 383782 60854
rect 383866 60618 384102 60854
rect 383546 24938 383782 25174
rect 383866 24938 384102 25174
rect 383546 24618 383782 24854
rect 383866 24618 384102 24854
rect 383546 -3462 383782 -3226
rect 383866 -3462 384102 -3226
rect 383546 -3782 383782 -3546
rect 383866 -3782 384102 -3546
rect 387266 676658 387502 676894
rect 387586 676658 387822 676894
rect 387266 676338 387502 676574
rect 387586 676338 387822 676574
rect 387266 640658 387502 640894
rect 387586 640658 387822 640894
rect 387266 640338 387502 640574
rect 387586 640338 387822 640574
rect 387266 604658 387502 604894
rect 387586 604658 387822 604894
rect 387266 604338 387502 604574
rect 387586 604338 387822 604574
rect 387266 568658 387502 568894
rect 387586 568658 387822 568894
rect 387266 568338 387502 568574
rect 387586 568338 387822 568574
rect 387266 532658 387502 532894
rect 387586 532658 387822 532894
rect 387266 532338 387502 532574
rect 387586 532338 387822 532574
rect 387266 496658 387502 496894
rect 387586 496658 387822 496894
rect 387266 496338 387502 496574
rect 387586 496338 387822 496574
rect 387266 460658 387502 460894
rect 387586 460658 387822 460894
rect 387266 460338 387502 460574
rect 387586 460338 387822 460574
rect 387266 424658 387502 424894
rect 387586 424658 387822 424894
rect 387266 424338 387502 424574
rect 387586 424338 387822 424574
rect 387266 388658 387502 388894
rect 387586 388658 387822 388894
rect 387266 388338 387502 388574
rect 387586 388338 387822 388574
rect 387266 352658 387502 352894
rect 387586 352658 387822 352894
rect 387266 352338 387502 352574
rect 387586 352338 387822 352574
rect 387266 316658 387502 316894
rect 387586 316658 387822 316894
rect 387266 316338 387502 316574
rect 387586 316338 387822 316574
rect 387266 280658 387502 280894
rect 387586 280658 387822 280894
rect 387266 280338 387502 280574
rect 387586 280338 387822 280574
rect 387266 244658 387502 244894
rect 387586 244658 387822 244894
rect 387266 244338 387502 244574
rect 387586 244338 387822 244574
rect 387266 208658 387502 208894
rect 387586 208658 387822 208894
rect 387266 208338 387502 208574
rect 387586 208338 387822 208574
rect 387266 172658 387502 172894
rect 387586 172658 387822 172894
rect 387266 172338 387502 172574
rect 387586 172338 387822 172574
rect 387266 136658 387502 136894
rect 387586 136658 387822 136894
rect 387266 136338 387502 136574
rect 387586 136338 387822 136574
rect 387266 100658 387502 100894
rect 387586 100658 387822 100894
rect 387266 100338 387502 100574
rect 387586 100338 387822 100574
rect 387266 64658 387502 64894
rect 387586 64658 387822 64894
rect 387266 64338 387502 64574
rect 387586 64338 387822 64574
rect 387266 28658 387502 28894
rect 387586 28658 387822 28894
rect 387266 28338 387502 28574
rect 387586 28338 387822 28574
rect 387266 -5382 387502 -5146
rect 387586 -5382 387822 -5146
rect 387266 -5702 387502 -5466
rect 387586 -5702 387822 -5466
rect 408986 710362 409222 710598
rect 409306 710362 409542 710598
rect 408986 710042 409222 710278
rect 409306 710042 409542 710278
rect 405266 708442 405502 708678
rect 405586 708442 405822 708678
rect 405266 708122 405502 708358
rect 405586 708122 405822 708358
rect 401546 706522 401782 706758
rect 401866 706522 402102 706758
rect 401546 706202 401782 706438
rect 401866 706202 402102 706438
rect 390986 680378 391222 680614
rect 391306 680378 391542 680614
rect 390986 680058 391222 680294
rect 391306 680058 391542 680294
rect 390986 644378 391222 644614
rect 391306 644378 391542 644614
rect 390986 644058 391222 644294
rect 391306 644058 391542 644294
rect 390986 608378 391222 608614
rect 391306 608378 391542 608614
rect 390986 608058 391222 608294
rect 391306 608058 391542 608294
rect 390986 572378 391222 572614
rect 391306 572378 391542 572614
rect 390986 572058 391222 572294
rect 391306 572058 391542 572294
rect 390986 536378 391222 536614
rect 391306 536378 391542 536614
rect 390986 536058 391222 536294
rect 391306 536058 391542 536294
rect 390986 500378 391222 500614
rect 391306 500378 391542 500614
rect 390986 500058 391222 500294
rect 391306 500058 391542 500294
rect 390986 464378 391222 464614
rect 391306 464378 391542 464614
rect 390986 464058 391222 464294
rect 391306 464058 391542 464294
rect 390986 428378 391222 428614
rect 391306 428378 391542 428614
rect 390986 428058 391222 428294
rect 391306 428058 391542 428294
rect 390986 392378 391222 392614
rect 391306 392378 391542 392614
rect 390986 392058 391222 392294
rect 391306 392058 391542 392294
rect 390986 356378 391222 356614
rect 391306 356378 391542 356614
rect 390986 356058 391222 356294
rect 391306 356058 391542 356294
rect 390986 320378 391222 320614
rect 391306 320378 391542 320614
rect 390986 320058 391222 320294
rect 391306 320058 391542 320294
rect 390986 284378 391222 284614
rect 391306 284378 391542 284614
rect 390986 284058 391222 284294
rect 391306 284058 391542 284294
rect 390986 248378 391222 248614
rect 391306 248378 391542 248614
rect 390986 248058 391222 248294
rect 391306 248058 391542 248294
rect 390986 212378 391222 212614
rect 391306 212378 391542 212614
rect 390986 212058 391222 212294
rect 391306 212058 391542 212294
rect 390986 176378 391222 176614
rect 391306 176378 391542 176614
rect 390986 176058 391222 176294
rect 391306 176058 391542 176294
rect 390986 140378 391222 140614
rect 391306 140378 391542 140614
rect 390986 140058 391222 140294
rect 391306 140058 391542 140294
rect 390986 104378 391222 104614
rect 391306 104378 391542 104614
rect 390986 104058 391222 104294
rect 391306 104058 391542 104294
rect 390986 68378 391222 68614
rect 391306 68378 391542 68614
rect 390986 68058 391222 68294
rect 391306 68058 391542 68294
rect 390986 32378 391222 32614
rect 391306 32378 391542 32614
rect 390986 32058 391222 32294
rect 391306 32058 391542 32294
rect 372986 -6342 373222 -6106
rect 373306 -6342 373542 -6106
rect 372986 -6662 373222 -6426
rect 373306 -6662 373542 -6426
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 690938 401782 691174
rect 401866 690938 402102 691174
rect 401546 690618 401782 690854
rect 401866 690618 402102 690854
rect 401546 654938 401782 655174
rect 401866 654938 402102 655174
rect 401546 654618 401782 654854
rect 401866 654618 402102 654854
rect 401546 618938 401782 619174
rect 401866 618938 402102 619174
rect 401546 618618 401782 618854
rect 401866 618618 402102 618854
rect 401546 582938 401782 583174
rect 401866 582938 402102 583174
rect 401546 582618 401782 582854
rect 401866 582618 402102 582854
rect 401546 546938 401782 547174
rect 401866 546938 402102 547174
rect 401546 546618 401782 546854
rect 401866 546618 402102 546854
rect 401546 510938 401782 511174
rect 401866 510938 402102 511174
rect 401546 510618 401782 510854
rect 401866 510618 402102 510854
rect 401546 474938 401782 475174
rect 401866 474938 402102 475174
rect 401546 474618 401782 474854
rect 401866 474618 402102 474854
rect 401546 438938 401782 439174
rect 401866 438938 402102 439174
rect 401546 438618 401782 438854
rect 401866 438618 402102 438854
rect 401546 402938 401782 403174
rect 401866 402938 402102 403174
rect 401546 402618 401782 402854
rect 401866 402618 402102 402854
rect 401546 366938 401782 367174
rect 401866 366938 402102 367174
rect 401546 366618 401782 366854
rect 401866 366618 402102 366854
rect 401546 330938 401782 331174
rect 401866 330938 402102 331174
rect 401546 330618 401782 330854
rect 401866 330618 402102 330854
rect 401546 294938 401782 295174
rect 401866 294938 402102 295174
rect 401546 294618 401782 294854
rect 401866 294618 402102 294854
rect 401546 258938 401782 259174
rect 401866 258938 402102 259174
rect 401546 258618 401782 258854
rect 401866 258618 402102 258854
rect 401546 222938 401782 223174
rect 401866 222938 402102 223174
rect 401546 222618 401782 222854
rect 401866 222618 402102 222854
rect 401546 186938 401782 187174
rect 401866 186938 402102 187174
rect 401546 186618 401782 186854
rect 401866 186618 402102 186854
rect 401546 150938 401782 151174
rect 401866 150938 402102 151174
rect 401546 150618 401782 150854
rect 401866 150618 402102 150854
rect 401546 114938 401782 115174
rect 401866 114938 402102 115174
rect 401546 114618 401782 114854
rect 401866 114618 402102 114854
rect 401546 78938 401782 79174
rect 401866 78938 402102 79174
rect 401546 78618 401782 78854
rect 401866 78618 402102 78854
rect 401546 42938 401782 43174
rect 401866 42938 402102 43174
rect 401546 42618 401782 42854
rect 401866 42618 402102 42854
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 401546 -2502 401782 -2266
rect 401866 -2502 402102 -2266
rect 401546 -2822 401782 -2586
rect 401866 -2822 402102 -2586
rect 405266 694658 405502 694894
rect 405586 694658 405822 694894
rect 405266 694338 405502 694574
rect 405586 694338 405822 694574
rect 405266 658658 405502 658894
rect 405586 658658 405822 658894
rect 405266 658338 405502 658574
rect 405586 658338 405822 658574
rect 405266 622658 405502 622894
rect 405586 622658 405822 622894
rect 405266 622338 405502 622574
rect 405586 622338 405822 622574
rect 405266 586658 405502 586894
rect 405586 586658 405822 586894
rect 405266 586338 405502 586574
rect 405586 586338 405822 586574
rect 405266 550658 405502 550894
rect 405586 550658 405822 550894
rect 405266 550338 405502 550574
rect 405586 550338 405822 550574
rect 405266 514658 405502 514894
rect 405586 514658 405822 514894
rect 405266 514338 405502 514574
rect 405586 514338 405822 514574
rect 405266 478658 405502 478894
rect 405586 478658 405822 478894
rect 405266 478338 405502 478574
rect 405586 478338 405822 478574
rect 405266 442658 405502 442894
rect 405586 442658 405822 442894
rect 405266 442338 405502 442574
rect 405586 442338 405822 442574
rect 405266 406658 405502 406894
rect 405586 406658 405822 406894
rect 405266 406338 405502 406574
rect 405586 406338 405822 406574
rect 405266 370658 405502 370894
rect 405586 370658 405822 370894
rect 405266 370338 405502 370574
rect 405586 370338 405822 370574
rect 405266 334658 405502 334894
rect 405586 334658 405822 334894
rect 405266 334338 405502 334574
rect 405586 334338 405822 334574
rect 405266 298658 405502 298894
rect 405586 298658 405822 298894
rect 405266 298338 405502 298574
rect 405586 298338 405822 298574
rect 405266 262658 405502 262894
rect 405586 262658 405822 262894
rect 405266 262338 405502 262574
rect 405586 262338 405822 262574
rect 405266 226658 405502 226894
rect 405586 226658 405822 226894
rect 405266 226338 405502 226574
rect 405586 226338 405822 226574
rect 405266 190658 405502 190894
rect 405586 190658 405822 190894
rect 405266 190338 405502 190574
rect 405586 190338 405822 190574
rect 405266 154658 405502 154894
rect 405586 154658 405822 154894
rect 405266 154338 405502 154574
rect 405586 154338 405822 154574
rect 405266 118658 405502 118894
rect 405586 118658 405822 118894
rect 405266 118338 405502 118574
rect 405586 118338 405822 118574
rect 405266 82658 405502 82894
rect 405586 82658 405822 82894
rect 405266 82338 405502 82574
rect 405586 82338 405822 82574
rect 405266 46658 405502 46894
rect 405586 46658 405822 46894
rect 405266 46338 405502 46574
rect 405586 46338 405822 46574
rect 405266 10658 405502 10894
rect 405586 10658 405822 10894
rect 405266 10338 405502 10574
rect 405586 10338 405822 10574
rect 405266 -4422 405502 -4186
rect 405586 -4422 405822 -4186
rect 405266 -4742 405502 -4506
rect 405586 -4742 405822 -4506
rect 426986 711322 427222 711558
rect 427306 711322 427542 711558
rect 426986 711002 427222 711238
rect 427306 711002 427542 711238
rect 423266 709402 423502 709638
rect 423586 709402 423822 709638
rect 423266 709082 423502 709318
rect 423586 709082 423822 709318
rect 419546 707482 419782 707718
rect 419866 707482 420102 707718
rect 419546 707162 419782 707398
rect 419866 707162 420102 707398
rect 408986 698378 409222 698614
rect 409306 698378 409542 698614
rect 408986 698058 409222 698294
rect 409306 698058 409542 698294
rect 408986 662378 409222 662614
rect 409306 662378 409542 662614
rect 408986 662058 409222 662294
rect 409306 662058 409542 662294
rect 408986 626378 409222 626614
rect 409306 626378 409542 626614
rect 408986 626058 409222 626294
rect 409306 626058 409542 626294
rect 408986 590378 409222 590614
rect 409306 590378 409542 590614
rect 408986 590058 409222 590294
rect 409306 590058 409542 590294
rect 408986 554378 409222 554614
rect 409306 554378 409542 554614
rect 408986 554058 409222 554294
rect 409306 554058 409542 554294
rect 408986 518378 409222 518614
rect 409306 518378 409542 518614
rect 408986 518058 409222 518294
rect 409306 518058 409542 518294
rect 408986 482378 409222 482614
rect 409306 482378 409542 482614
rect 408986 482058 409222 482294
rect 409306 482058 409542 482294
rect 408986 446378 409222 446614
rect 409306 446378 409542 446614
rect 408986 446058 409222 446294
rect 409306 446058 409542 446294
rect 408986 410378 409222 410614
rect 409306 410378 409542 410614
rect 408986 410058 409222 410294
rect 409306 410058 409542 410294
rect 408986 374378 409222 374614
rect 409306 374378 409542 374614
rect 408986 374058 409222 374294
rect 409306 374058 409542 374294
rect 408986 338378 409222 338614
rect 409306 338378 409542 338614
rect 408986 338058 409222 338294
rect 409306 338058 409542 338294
rect 408986 302378 409222 302614
rect 409306 302378 409542 302614
rect 408986 302058 409222 302294
rect 409306 302058 409542 302294
rect 408986 266378 409222 266614
rect 409306 266378 409542 266614
rect 408986 266058 409222 266294
rect 409306 266058 409542 266294
rect 408986 230378 409222 230614
rect 409306 230378 409542 230614
rect 408986 230058 409222 230294
rect 409306 230058 409542 230294
rect 408986 194378 409222 194614
rect 409306 194378 409542 194614
rect 408986 194058 409222 194294
rect 409306 194058 409542 194294
rect 408986 158378 409222 158614
rect 409306 158378 409542 158614
rect 408986 158058 409222 158294
rect 409306 158058 409542 158294
rect 408986 122378 409222 122614
rect 409306 122378 409542 122614
rect 408986 122058 409222 122294
rect 409306 122058 409542 122294
rect 408986 86378 409222 86614
rect 409306 86378 409542 86614
rect 408986 86058 409222 86294
rect 409306 86058 409542 86294
rect 408986 50378 409222 50614
rect 409306 50378 409542 50614
rect 408986 50058 409222 50294
rect 409306 50058 409542 50294
rect 408986 14378 409222 14614
rect 409306 14378 409542 14614
rect 408986 14058 409222 14294
rect 409306 14058 409542 14294
rect 390986 -7302 391222 -7066
rect 391306 -7302 391542 -7066
rect 390986 -7622 391222 -7386
rect 391306 -7622 391542 -7386
rect 415826 705562 416062 705798
rect 416146 705562 416382 705798
rect 415826 705242 416062 705478
rect 416146 705242 416382 705478
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 415826 561218 416062 561454
rect 416146 561218 416382 561454
rect 415826 560898 416062 561134
rect 416146 560898 416382 561134
rect 415826 525218 416062 525454
rect 416146 525218 416382 525454
rect 415826 524898 416062 525134
rect 416146 524898 416382 525134
rect 415826 489218 416062 489454
rect 416146 489218 416382 489454
rect 415826 488898 416062 489134
rect 416146 488898 416382 489134
rect 415826 453218 416062 453454
rect 416146 453218 416382 453454
rect 415826 452898 416062 453134
rect 416146 452898 416382 453134
rect 415826 417218 416062 417454
rect 416146 417218 416382 417454
rect 415826 416898 416062 417134
rect 416146 416898 416382 417134
rect 415826 381218 416062 381454
rect 416146 381218 416382 381454
rect 415826 380898 416062 381134
rect 416146 380898 416382 381134
rect 415826 345218 416062 345454
rect 416146 345218 416382 345454
rect 415826 344898 416062 345134
rect 416146 344898 416382 345134
rect 415826 309218 416062 309454
rect 416146 309218 416382 309454
rect 415826 308898 416062 309134
rect 416146 308898 416382 309134
rect 415826 273218 416062 273454
rect 416146 273218 416382 273454
rect 415826 272898 416062 273134
rect 416146 272898 416382 273134
rect 415826 237218 416062 237454
rect 416146 237218 416382 237454
rect 415826 236898 416062 237134
rect 416146 236898 416382 237134
rect 415826 201218 416062 201454
rect 416146 201218 416382 201454
rect 415826 200898 416062 201134
rect 416146 200898 416382 201134
rect 415826 165218 416062 165454
rect 416146 165218 416382 165454
rect 415826 164898 416062 165134
rect 416146 164898 416382 165134
rect 415826 129218 416062 129454
rect 416146 129218 416382 129454
rect 415826 128898 416062 129134
rect 416146 128898 416382 129134
rect 415826 93218 416062 93454
rect 416146 93218 416382 93454
rect 415826 92898 416062 93134
rect 416146 92898 416382 93134
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -1542 416062 -1306
rect 416146 -1542 416382 -1306
rect 415826 -1862 416062 -1626
rect 416146 -1862 416382 -1626
rect 419546 672938 419782 673174
rect 419866 672938 420102 673174
rect 419546 672618 419782 672854
rect 419866 672618 420102 672854
rect 419546 636938 419782 637174
rect 419866 636938 420102 637174
rect 419546 636618 419782 636854
rect 419866 636618 420102 636854
rect 419546 600938 419782 601174
rect 419866 600938 420102 601174
rect 419546 600618 419782 600854
rect 419866 600618 420102 600854
rect 419546 564938 419782 565174
rect 419866 564938 420102 565174
rect 419546 564618 419782 564854
rect 419866 564618 420102 564854
rect 419546 528938 419782 529174
rect 419866 528938 420102 529174
rect 419546 528618 419782 528854
rect 419866 528618 420102 528854
rect 419546 492938 419782 493174
rect 419866 492938 420102 493174
rect 419546 492618 419782 492854
rect 419866 492618 420102 492854
rect 419546 456938 419782 457174
rect 419866 456938 420102 457174
rect 419546 456618 419782 456854
rect 419866 456618 420102 456854
rect 419546 420938 419782 421174
rect 419866 420938 420102 421174
rect 419546 420618 419782 420854
rect 419866 420618 420102 420854
rect 419546 384938 419782 385174
rect 419866 384938 420102 385174
rect 419546 384618 419782 384854
rect 419866 384618 420102 384854
rect 419546 348938 419782 349174
rect 419866 348938 420102 349174
rect 419546 348618 419782 348854
rect 419866 348618 420102 348854
rect 419546 312938 419782 313174
rect 419866 312938 420102 313174
rect 419546 312618 419782 312854
rect 419866 312618 420102 312854
rect 419546 276938 419782 277174
rect 419866 276938 420102 277174
rect 419546 276618 419782 276854
rect 419866 276618 420102 276854
rect 419546 240938 419782 241174
rect 419866 240938 420102 241174
rect 419546 240618 419782 240854
rect 419866 240618 420102 240854
rect 419546 204938 419782 205174
rect 419866 204938 420102 205174
rect 419546 204618 419782 204854
rect 419866 204618 420102 204854
rect 419546 168938 419782 169174
rect 419866 168938 420102 169174
rect 419546 168618 419782 168854
rect 419866 168618 420102 168854
rect 419546 132938 419782 133174
rect 419866 132938 420102 133174
rect 419546 132618 419782 132854
rect 419866 132618 420102 132854
rect 419546 96938 419782 97174
rect 419866 96938 420102 97174
rect 419546 96618 419782 96854
rect 419866 96618 420102 96854
rect 419546 60938 419782 61174
rect 419866 60938 420102 61174
rect 419546 60618 419782 60854
rect 419866 60618 420102 60854
rect 419546 24938 419782 25174
rect 419866 24938 420102 25174
rect 419546 24618 419782 24854
rect 419866 24618 420102 24854
rect 419546 -3462 419782 -3226
rect 419866 -3462 420102 -3226
rect 419546 -3782 419782 -3546
rect 419866 -3782 420102 -3546
rect 423266 676658 423502 676894
rect 423586 676658 423822 676894
rect 423266 676338 423502 676574
rect 423586 676338 423822 676574
rect 423266 640658 423502 640894
rect 423586 640658 423822 640894
rect 423266 640338 423502 640574
rect 423586 640338 423822 640574
rect 423266 604658 423502 604894
rect 423586 604658 423822 604894
rect 423266 604338 423502 604574
rect 423586 604338 423822 604574
rect 423266 568658 423502 568894
rect 423586 568658 423822 568894
rect 423266 568338 423502 568574
rect 423586 568338 423822 568574
rect 423266 532658 423502 532894
rect 423586 532658 423822 532894
rect 423266 532338 423502 532574
rect 423586 532338 423822 532574
rect 423266 496658 423502 496894
rect 423586 496658 423822 496894
rect 423266 496338 423502 496574
rect 423586 496338 423822 496574
rect 423266 460658 423502 460894
rect 423586 460658 423822 460894
rect 423266 460338 423502 460574
rect 423586 460338 423822 460574
rect 423266 424658 423502 424894
rect 423586 424658 423822 424894
rect 423266 424338 423502 424574
rect 423586 424338 423822 424574
rect 423266 388658 423502 388894
rect 423586 388658 423822 388894
rect 423266 388338 423502 388574
rect 423586 388338 423822 388574
rect 423266 352658 423502 352894
rect 423586 352658 423822 352894
rect 423266 352338 423502 352574
rect 423586 352338 423822 352574
rect 423266 316658 423502 316894
rect 423586 316658 423822 316894
rect 423266 316338 423502 316574
rect 423586 316338 423822 316574
rect 423266 280658 423502 280894
rect 423586 280658 423822 280894
rect 423266 280338 423502 280574
rect 423586 280338 423822 280574
rect 423266 244658 423502 244894
rect 423586 244658 423822 244894
rect 423266 244338 423502 244574
rect 423586 244338 423822 244574
rect 423266 208658 423502 208894
rect 423586 208658 423822 208894
rect 423266 208338 423502 208574
rect 423586 208338 423822 208574
rect 423266 172658 423502 172894
rect 423586 172658 423822 172894
rect 423266 172338 423502 172574
rect 423586 172338 423822 172574
rect 423266 136658 423502 136894
rect 423586 136658 423822 136894
rect 423266 136338 423502 136574
rect 423586 136338 423822 136574
rect 423266 100658 423502 100894
rect 423586 100658 423822 100894
rect 423266 100338 423502 100574
rect 423586 100338 423822 100574
rect 423266 64658 423502 64894
rect 423586 64658 423822 64894
rect 423266 64338 423502 64574
rect 423586 64338 423822 64574
rect 423266 28658 423502 28894
rect 423586 28658 423822 28894
rect 423266 28338 423502 28574
rect 423586 28338 423822 28574
rect 423266 -5382 423502 -5146
rect 423586 -5382 423822 -5146
rect 423266 -5702 423502 -5466
rect 423586 -5702 423822 -5466
rect 444986 710362 445222 710598
rect 445306 710362 445542 710598
rect 444986 710042 445222 710278
rect 445306 710042 445542 710278
rect 441266 708442 441502 708678
rect 441586 708442 441822 708678
rect 441266 708122 441502 708358
rect 441586 708122 441822 708358
rect 437546 706522 437782 706758
rect 437866 706522 438102 706758
rect 437546 706202 437782 706438
rect 437866 706202 438102 706438
rect 426986 680378 427222 680614
rect 427306 680378 427542 680614
rect 426986 680058 427222 680294
rect 427306 680058 427542 680294
rect 426986 644378 427222 644614
rect 427306 644378 427542 644614
rect 426986 644058 427222 644294
rect 427306 644058 427542 644294
rect 426986 608378 427222 608614
rect 427306 608378 427542 608614
rect 426986 608058 427222 608294
rect 427306 608058 427542 608294
rect 426986 572378 427222 572614
rect 427306 572378 427542 572614
rect 426986 572058 427222 572294
rect 427306 572058 427542 572294
rect 426986 536378 427222 536614
rect 427306 536378 427542 536614
rect 426986 536058 427222 536294
rect 427306 536058 427542 536294
rect 426986 500378 427222 500614
rect 427306 500378 427542 500614
rect 426986 500058 427222 500294
rect 427306 500058 427542 500294
rect 426986 464378 427222 464614
rect 427306 464378 427542 464614
rect 426986 464058 427222 464294
rect 427306 464058 427542 464294
rect 426986 428378 427222 428614
rect 427306 428378 427542 428614
rect 426986 428058 427222 428294
rect 427306 428058 427542 428294
rect 426986 392378 427222 392614
rect 427306 392378 427542 392614
rect 426986 392058 427222 392294
rect 427306 392058 427542 392294
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 433826 435218 434062 435454
rect 434146 435218 434382 435454
rect 433826 434898 434062 435134
rect 434146 434898 434382 435134
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 437546 690938 437782 691174
rect 437866 690938 438102 691174
rect 437546 690618 437782 690854
rect 437866 690618 438102 690854
rect 437546 654938 437782 655174
rect 437866 654938 438102 655174
rect 437546 654618 437782 654854
rect 437866 654618 438102 654854
rect 437546 618938 437782 619174
rect 437866 618938 438102 619174
rect 437546 618618 437782 618854
rect 437866 618618 438102 618854
rect 437546 582938 437782 583174
rect 437866 582938 438102 583174
rect 437546 582618 437782 582854
rect 437866 582618 438102 582854
rect 437546 546938 437782 547174
rect 437866 546938 438102 547174
rect 437546 546618 437782 546854
rect 437866 546618 438102 546854
rect 437546 510938 437782 511174
rect 437866 510938 438102 511174
rect 437546 510618 437782 510854
rect 437866 510618 438102 510854
rect 437546 474938 437782 475174
rect 437866 474938 438102 475174
rect 437546 474618 437782 474854
rect 437866 474618 438102 474854
rect 437546 438938 437782 439174
rect 437866 438938 438102 439174
rect 437546 438618 437782 438854
rect 437866 438618 438102 438854
rect 437546 402938 437782 403174
rect 437866 402938 438102 403174
rect 437546 402618 437782 402854
rect 437866 402618 438102 402854
rect 441266 694658 441502 694894
rect 441586 694658 441822 694894
rect 441266 694338 441502 694574
rect 441586 694338 441822 694574
rect 441266 658658 441502 658894
rect 441586 658658 441822 658894
rect 441266 658338 441502 658574
rect 441586 658338 441822 658574
rect 441266 622658 441502 622894
rect 441586 622658 441822 622894
rect 441266 622338 441502 622574
rect 441586 622338 441822 622574
rect 441266 586658 441502 586894
rect 441586 586658 441822 586894
rect 441266 586338 441502 586574
rect 441586 586338 441822 586574
rect 441266 550658 441502 550894
rect 441586 550658 441822 550894
rect 441266 550338 441502 550574
rect 441586 550338 441822 550574
rect 441266 514658 441502 514894
rect 441586 514658 441822 514894
rect 441266 514338 441502 514574
rect 441586 514338 441822 514574
rect 441266 478658 441502 478894
rect 441586 478658 441822 478894
rect 441266 478338 441502 478574
rect 441586 478338 441822 478574
rect 441266 442658 441502 442894
rect 441586 442658 441822 442894
rect 441266 442338 441502 442574
rect 441586 442338 441822 442574
rect 441266 406658 441502 406894
rect 441586 406658 441822 406894
rect 441266 406338 441502 406574
rect 441586 406338 441822 406574
rect 462986 711322 463222 711558
rect 463306 711322 463542 711558
rect 462986 711002 463222 711238
rect 463306 711002 463542 711238
rect 459266 709402 459502 709638
rect 459586 709402 459822 709638
rect 459266 709082 459502 709318
rect 459586 709082 459822 709318
rect 455546 707482 455782 707718
rect 455866 707482 456102 707718
rect 455546 707162 455782 707398
rect 455866 707162 456102 707398
rect 444986 698378 445222 698614
rect 445306 698378 445542 698614
rect 444986 698058 445222 698294
rect 445306 698058 445542 698294
rect 444986 662378 445222 662614
rect 445306 662378 445542 662614
rect 444986 662058 445222 662294
rect 445306 662058 445542 662294
rect 444986 626378 445222 626614
rect 445306 626378 445542 626614
rect 444986 626058 445222 626294
rect 445306 626058 445542 626294
rect 444986 590378 445222 590614
rect 445306 590378 445542 590614
rect 444986 590058 445222 590294
rect 445306 590058 445542 590294
rect 444986 554378 445222 554614
rect 445306 554378 445542 554614
rect 444986 554058 445222 554294
rect 445306 554058 445542 554294
rect 444986 518378 445222 518614
rect 445306 518378 445542 518614
rect 444986 518058 445222 518294
rect 445306 518058 445542 518294
rect 444986 482378 445222 482614
rect 445306 482378 445542 482614
rect 444986 482058 445222 482294
rect 445306 482058 445542 482294
rect 444986 446378 445222 446614
rect 445306 446378 445542 446614
rect 444986 446058 445222 446294
rect 445306 446058 445542 446294
rect 444986 410378 445222 410614
rect 445306 410378 445542 410614
rect 444986 410058 445222 410294
rect 445306 410058 445542 410294
rect 444986 374378 445222 374614
rect 445306 374378 445542 374614
rect 444986 374058 445222 374294
rect 445306 374058 445542 374294
rect 434285 363218 434521 363454
rect 434285 362898 434521 363134
rect 436882 363218 437118 363454
rect 436882 362898 437118 363134
rect 439479 363218 439715 363454
rect 439479 362898 439715 363134
rect 426986 356378 427222 356614
rect 427306 356378 427542 356614
rect 426986 356058 427222 356294
rect 427306 356058 427542 356294
rect 435583 345218 435819 345454
rect 435583 344898 435819 345134
rect 438180 345218 438416 345454
rect 438180 344898 438416 345134
rect 444986 338378 445222 338614
rect 445306 338378 445542 338614
rect 444986 338058 445222 338294
rect 445306 338058 445542 338294
rect 426986 320378 427222 320614
rect 427306 320378 427542 320614
rect 426986 320058 427222 320294
rect 427306 320058 427542 320294
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 437546 330938 437782 331174
rect 437866 330938 438102 331174
rect 437546 330618 437782 330854
rect 437866 330618 438102 330854
rect 441266 334658 441502 334894
rect 441586 334658 441822 334894
rect 441266 334338 441502 334574
rect 441586 334338 441822 334574
rect 444986 302378 445222 302614
rect 445306 302378 445542 302614
rect 444986 302058 445222 302294
rect 445306 302058 445542 302294
rect 434285 291218 434521 291454
rect 434285 290898 434521 291134
rect 436882 291218 437118 291454
rect 436882 290898 437118 291134
rect 439479 291218 439715 291454
rect 439479 290898 439715 291134
rect 426986 284378 427222 284614
rect 427306 284378 427542 284614
rect 426986 284058 427222 284294
rect 427306 284058 427542 284294
rect 435583 273218 435819 273454
rect 435583 272898 435819 273134
rect 438180 273218 438416 273454
rect 438180 272898 438416 273134
rect 444986 266378 445222 266614
rect 445306 266378 445542 266614
rect 444986 266058 445222 266294
rect 445306 266058 445542 266294
rect 426986 248378 427222 248614
rect 427306 248378 427542 248614
rect 426986 248058 427222 248294
rect 427306 248058 427542 248294
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 437546 258938 437782 259174
rect 437866 258938 438102 259174
rect 437546 258618 437782 258854
rect 437866 258618 438102 258854
rect 441266 262658 441502 262894
rect 441586 262658 441822 262894
rect 441266 262338 441502 262574
rect 441586 262338 441822 262574
rect 444986 230378 445222 230614
rect 445306 230378 445542 230614
rect 444986 230058 445222 230294
rect 445306 230058 445542 230294
rect 434285 219218 434521 219454
rect 434285 218898 434521 219134
rect 436882 219218 437118 219454
rect 436882 218898 437118 219134
rect 439479 219218 439715 219454
rect 439479 218898 439715 219134
rect 426986 212378 427222 212614
rect 427306 212378 427542 212614
rect 426986 212058 427222 212294
rect 427306 212058 427542 212294
rect 435583 201218 435819 201454
rect 435583 200898 435819 201134
rect 438180 201218 438416 201454
rect 438180 200898 438416 201134
rect 444986 194378 445222 194614
rect 445306 194378 445542 194614
rect 444986 194058 445222 194294
rect 445306 194058 445542 194294
rect 426986 176378 427222 176614
rect 427306 176378 427542 176614
rect 426986 176058 427222 176294
rect 427306 176058 427542 176294
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 437546 186938 437782 187174
rect 437866 186938 438102 187174
rect 437546 186618 437782 186854
rect 437866 186618 438102 186854
rect 441266 190658 441502 190894
rect 441586 190658 441822 190894
rect 441266 190338 441502 190574
rect 441586 190338 441822 190574
rect 444986 158378 445222 158614
rect 445306 158378 445542 158614
rect 444986 158058 445222 158294
rect 445306 158058 445542 158294
rect 434285 147218 434521 147454
rect 434285 146898 434521 147134
rect 436882 147218 437118 147454
rect 436882 146898 437118 147134
rect 439479 147218 439715 147454
rect 439479 146898 439715 147134
rect 426986 140378 427222 140614
rect 427306 140378 427542 140614
rect 426986 140058 427222 140294
rect 427306 140058 427542 140294
rect 435583 129218 435819 129454
rect 435583 128898 435819 129134
rect 438180 129218 438416 129454
rect 438180 128898 438416 129134
rect 444986 122378 445222 122614
rect 445306 122378 445542 122614
rect 444986 122058 445222 122294
rect 445306 122058 445542 122294
rect 426986 104378 427222 104614
rect 427306 104378 427542 104614
rect 426986 104058 427222 104294
rect 427306 104058 427542 104294
rect 426986 68378 427222 68614
rect 427306 68378 427542 68614
rect 426986 68058 427222 68294
rect 427306 68058 427542 68294
rect 426986 32378 427222 32614
rect 427306 32378 427542 32614
rect 426986 32058 427222 32294
rect 427306 32058 427542 32294
rect 408986 -6342 409222 -6106
rect 409306 -6342 409542 -6106
rect 408986 -6662 409222 -6426
rect 409306 -6662 409542 -6426
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 437546 114938 437782 115174
rect 437866 114938 438102 115174
rect 437546 114618 437782 114854
rect 437866 114618 438102 114854
rect 437546 78938 437782 79174
rect 437866 78938 438102 79174
rect 437546 78618 437782 78854
rect 437866 78618 438102 78854
rect 437546 42938 437782 43174
rect 437866 42938 438102 43174
rect 437546 42618 437782 42854
rect 437866 42618 438102 42854
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 437546 -2502 437782 -2266
rect 437866 -2502 438102 -2266
rect 437546 -2822 437782 -2586
rect 437866 -2822 438102 -2586
rect 441266 118658 441502 118894
rect 441586 118658 441822 118894
rect 441266 118338 441502 118574
rect 441586 118338 441822 118574
rect 441266 82658 441502 82894
rect 441586 82658 441822 82894
rect 441266 82338 441502 82574
rect 441586 82338 441822 82574
rect 441266 46658 441502 46894
rect 441586 46658 441822 46894
rect 441266 46338 441502 46574
rect 441586 46338 441822 46574
rect 441266 10658 441502 10894
rect 441586 10658 441822 10894
rect 441266 10338 441502 10574
rect 441586 10338 441822 10574
rect 441266 -4422 441502 -4186
rect 441586 -4422 441822 -4186
rect 441266 -4742 441502 -4506
rect 441586 -4742 441822 -4506
rect 444986 86378 445222 86614
rect 445306 86378 445542 86614
rect 444986 86058 445222 86294
rect 445306 86058 445542 86294
rect 444986 50378 445222 50614
rect 445306 50378 445542 50614
rect 444986 50058 445222 50294
rect 445306 50058 445542 50294
rect 444986 14378 445222 14614
rect 445306 14378 445542 14614
rect 444986 14058 445222 14294
rect 445306 14058 445542 14294
rect 426986 -7302 427222 -7066
rect 427306 -7302 427542 -7066
rect 426986 -7622 427222 -7386
rect 427306 -7622 427542 -7386
rect 451826 705562 452062 705798
rect 452146 705562 452382 705798
rect 451826 705242 452062 705478
rect 452146 705242 452382 705478
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 451826 453218 452062 453454
rect 452146 453218 452382 453454
rect 451826 452898 452062 453134
rect 452146 452898 452382 453134
rect 451826 417218 452062 417454
rect 452146 417218 452382 417454
rect 451826 416898 452062 417134
rect 452146 416898 452382 417134
rect 451826 381218 452062 381454
rect 452146 381218 452382 381454
rect 451826 380898 452062 381134
rect 452146 380898 452382 381134
rect 451826 345218 452062 345454
rect 452146 345218 452382 345454
rect 451826 344898 452062 345134
rect 452146 344898 452382 345134
rect 451826 309218 452062 309454
rect 452146 309218 452382 309454
rect 451826 308898 452062 309134
rect 452146 308898 452382 309134
rect 451826 273218 452062 273454
rect 452146 273218 452382 273454
rect 451826 272898 452062 273134
rect 452146 272898 452382 273134
rect 451826 237218 452062 237454
rect 452146 237218 452382 237454
rect 451826 236898 452062 237134
rect 452146 236898 452382 237134
rect 451826 201218 452062 201454
rect 452146 201218 452382 201454
rect 451826 200898 452062 201134
rect 452146 200898 452382 201134
rect 451826 165218 452062 165454
rect 452146 165218 452382 165454
rect 451826 164898 452062 165134
rect 452146 164898 452382 165134
rect 451826 129218 452062 129454
rect 452146 129218 452382 129454
rect 451826 128898 452062 129134
rect 452146 128898 452382 129134
rect 451826 93218 452062 93454
rect 452146 93218 452382 93454
rect 451826 92898 452062 93134
rect 452146 92898 452382 93134
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -1542 452062 -1306
rect 452146 -1542 452382 -1306
rect 451826 -1862 452062 -1626
rect 452146 -1862 452382 -1626
rect 455546 672938 455782 673174
rect 455866 672938 456102 673174
rect 455546 672618 455782 672854
rect 455866 672618 456102 672854
rect 455546 636938 455782 637174
rect 455866 636938 456102 637174
rect 455546 636618 455782 636854
rect 455866 636618 456102 636854
rect 455546 600938 455782 601174
rect 455866 600938 456102 601174
rect 455546 600618 455782 600854
rect 455866 600618 456102 600854
rect 455546 564938 455782 565174
rect 455866 564938 456102 565174
rect 455546 564618 455782 564854
rect 455866 564618 456102 564854
rect 455546 528938 455782 529174
rect 455866 528938 456102 529174
rect 455546 528618 455782 528854
rect 455866 528618 456102 528854
rect 455546 492938 455782 493174
rect 455866 492938 456102 493174
rect 455546 492618 455782 492854
rect 455866 492618 456102 492854
rect 455546 456938 455782 457174
rect 455866 456938 456102 457174
rect 455546 456618 455782 456854
rect 455866 456618 456102 456854
rect 455546 420938 455782 421174
rect 455866 420938 456102 421174
rect 455546 420618 455782 420854
rect 455866 420618 456102 420854
rect 455546 384938 455782 385174
rect 455866 384938 456102 385174
rect 455546 384618 455782 384854
rect 455866 384618 456102 384854
rect 455546 348938 455782 349174
rect 455866 348938 456102 349174
rect 455546 348618 455782 348854
rect 455866 348618 456102 348854
rect 455546 312938 455782 313174
rect 455866 312938 456102 313174
rect 455546 312618 455782 312854
rect 455866 312618 456102 312854
rect 455546 276938 455782 277174
rect 455866 276938 456102 277174
rect 455546 276618 455782 276854
rect 455866 276618 456102 276854
rect 455546 240938 455782 241174
rect 455866 240938 456102 241174
rect 455546 240618 455782 240854
rect 455866 240618 456102 240854
rect 455546 204938 455782 205174
rect 455866 204938 456102 205174
rect 455546 204618 455782 204854
rect 455866 204618 456102 204854
rect 455546 168938 455782 169174
rect 455866 168938 456102 169174
rect 455546 168618 455782 168854
rect 455866 168618 456102 168854
rect 455546 132938 455782 133174
rect 455866 132938 456102 133174
rect 455546 132618 455782 132854
rect 455866 132618 456102 132854
rect 455546 96938 455782 97174
rect 455866 96938 456102 97174
rect 455546 96618 455782 96854
rect 455866 96618 456102 96854
rect 455546 60938 455782 61174
rect 455866 60938 456102 61174
rect 455546 60618 455782 60854
rect 455866 60618 456102 60854
rect 455546 24938 455782 25174
rect 455866 24938 456102 25174
rect 455546 24618 455782 24854
rect 455866 24618 456102 24854
rect 455546 -3462 455782 -3226
rect 455866 -3462 456102 -3226
rect 455546 -3782 455782 -3546
rect 455866 -3782 456102 -3546
rect 459266 676658 459502 676894
rect 459586 676658 459822 676894
rect 459266 676338 459502 676574
rect 459586 676338 459822 676574
rect 459266 640658 459502 640894
rect 459586 640658 459822 640894
rect 459266 640338 459502 640574
rect 459586 640338 459822 640574
rect 459266 604658 459502 604894
rect 459586 604658 459822 604894
rect 459266 604338 459502 604574
rect 459586 604338 459822 604574
rect 459266 568658 459502 568894
rect 459586 568658 459822 568894
rect 459266 568338 459502 568574
rect 459586 568338 459822 568574
rect 459266 532658 459502 532894
rect 459586 532658 459822 532894
rect 459266 532338 459502 532574
rect 459586 532338 459822 532574
rect 459266 496658 459502 496894
rect 459586 496658 459822 496894
rect 459266 496338 459502 496574
rect 459586 496338 459822 496574
rect 459266 460658 459502 460894
rect 459586 460658 459822 460894
rect 459266 460338 459502 460574
rect 459586 460338 459822 460574
rect 459266 424658 459502 424894
rect 459586 424658 459822 424894
rect 459266 424338 459502 424574
rect 459586 424338 459822 424574
rect 459266 388658 459502 388894
rect 459586 388658 459822 388894
rect 459266 388338 459502 388574
rect 459586 388338 459822 388574
rect 459266 352658 459502 352894
rect 459586 352658 459822 352894
rect 459266 352338 459502 352574
rect 459586 352338 459822 352574
rect 459266 316658 459502 316894
rect 459586 316658 459822 316894
rect 459266 316338 459502 316574
rect 459586 316338 459822 316574
rect 459266 280658 459502 280894
rect 459586 280658 459822 280894
rect 459266 280338 459502 280574
rect 459586 280338 459822 280574
rect 459266 244658 459502 244894
rect 459586 244658 459822 244894
rect 459266 244338 459502 244574
rect 459586 244338 459822 244574
rect 459266 208658 459502 208894
rect 459586 208658 459822 208894
rect 459266 208338 459502 208574
rect 459586 208338 459822 208574
rect 459266 172658 459502 172894
rect 459586 172658 459822 172894
rect 459266 172338 459502 172574
rect 459586 172338 459822 172574
rect 459266 136658 459502 136894
rect 459586 136658 459822 136894
rect 459266 136338 459502 136574
rect 459586 136338 459822 136574
rect 459266 100658 459502 100894
rect 459586 100658 459822 100894
rect 459266 100338 459502 100574
rect 459586 100338 459822 100574
rect 459266 64658 459502 64894
rect 459586 64658 459822 64894
rect 459266 64338 459502 64574
rect 459586 64338 459822 64574
rect 459266 28658 459502 28894
rect 459586 28658 459822 28894
rect 459266 28338 459502 28574
rect 459586 28338 459822 28574
rect 459266 -5382 459502 -5146
rect 459586 -5382 459822 -5146
rect 459266 -5702 459502 -5466
rect 459586 -5702 459822 -5466
rect 480986 710362 481222 710598
rect 481306 710362 481542 710598
rect 480986 710042 481222 710278
rect 481306 710042 481542 710278
rect 477266 708442 477502 708678
rect 477586 708442 477822 708678
rect 477266 708122 477502 708358
rect 477586 708122 477822 708358
rect 473546 706522 473782 706758
rect 473866 706522 474102 706758
rect 473546 706202 473782 706438
rect 473866 706202 474102 706438
rect 462986 680378 463222 680614
rect 463306 680378 463542 680614
rect 462986 680058 463222 680294
rect 463306 680058 463542 680294
rect 462986 644378 463222 644614
rect 463306 644378 463542 644614
rect 462986 644058 463222 644294
rect 463306 644058 463542 644294
rect 462986 608378 463222 608614
rect 463306 608378 463542 608614
rect 462986 608058 463222 608294
rect 463306 608058 463542 608294
rect 462986 572378 463222 572614
rect 463306 572378 463542 572614
rect 462986 572058 463222 572294
rect 463306 572058 463542 572294
rect 462986 536378 463222 536614
rect 463306 536378 463542 536614
rect 462986 536058 463222 536294
rect 463306 536058 463542 536294
rect 462986 500378 463222 500614
rect 463306 500378 463542 500614
rect 462986 500058 463222 500294
rect 463306 500058 463542 500294
rect 462986 464378 463222 464614
rect 463306 464378 463542 464614
rect 462986 464058 463222 464294
rect 463306 464058 463542 464294
rect 462986 428378 463222 428614
rect 463306 428378 463542 428614
rect 462986 428058 463222 428294
rect 463306 428058 463542 428294
rect 462986 392378 463222 392614
rect 463306 392378 463542 392614
rect 462986 392058 463222 392294
rect 463306 392058 463542 392294
rect 462986 356378 463222 356614
rect 463306 356378 463542 356614
rect 462986 356058 463222 356294
rect 463306 356058 463542 356294
rect 462986 320378 463222 320614
rect 463306 320378 463542 320614
rect 462986 320058 463222 320294
rect 463306 320058 463542 320294
rect 462986 284378 463222 284614
rect 463306 284378 463542 284614
rect 462986 284058 463222 284294
rect 463306 284058 463542 284294
rect 462986 248378 463222 248614
rect 463306 248378 463542 248614
rect 462986 248058 463222 248294
rect 463306 248058 463542 248294
rect 462986 212378 463222 212614
rect 463306 212378 463542 212614
rect 462986 212058 463222 212294
rect 463306 212058 463542 212294
rect 462986 176378 463222 176614
rect 463306 176378 463542 176614
rect 462986 176058 463222 176294
rect 463306 176058 463542 176294
rect 462986 140378 463222 140614
rect 463306 140378 463542 140614
rect 462986 140058 463222 140294
rect 463306 140058 463542 140294
rect 462986 104378 463222 104614
rect 463306 104378 463542 104614
rect 462986 104058 463222 104294
rect 463306 104058 463542 104294
rect 462986 68378 463222 68614
rect 463306 68378 463542 68614
rect 462986 68058 463222 68294
rect 463306 68058 463542 68294
rect 462986 32378 463222 32614
rect 463306 32378 463542 32614
rect 462986 32058 463222 32294
rect 463306 32058 463542 32294
rect 444986 -6342 445222 -6106
rect 445306 -6342 445542 -6106
rect 444986 -6662 445222 -6426
rect 445306 -6662 445542 -6426
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 690938 473782 691174
rect 473866 690938 474102 691174
rect 473546 690618 473782 690854
rect 473866 690618 474102 690854
rect 473546 654938 473782 655174
rect 473866 654938 474102 655174
rect 473546 654618 473782 654854
rect 473866 654618 474102 654854
rect 473546 618938 473782 619174
rect 473866 618938 474102 619174
rect 473546 618618 473782 618854
rect 473866 618618 474102 618854
rect 473546 582938 473782 583174
rect 473866 582938 474102 583174
rect 473546 582618 473782 582854
rect 473866 582618 474102 582854
rect 473546 546938 473782 547174
rect 473866 546938 474102 547174
rect 473546 546618 473782 546854
rect 473866 546618 474102 546854
rect 473546 510938 473782 511174
rect 473866 510938 474102 511174
rect 473546 510618 473782 510854
rect 473866 510618 474102 510854
rect 473546 474938 473782 475174
rect 473866 474938 474102 475174
rect 473546 474618 473782 474854
rect 473866 474618 474102 474854
rect 473546 438938 473782 439174
rect 473866 438938 474102 439174
rect 473546 438618 473782 438854
rect 473866 438618 474102 438854
rect 473546 402938 473782 403174
rect 473866 402938 474102 403174
rect 473546 402618 473782 402854
rect 473866 402618 474102 402854
rect 473546 366938 473782 367174
rect 473866 366938 474102 367174
rect 473546 366618 473782 366854
rect 473866 366618 474102 366854
rect 473546 330938 473782 331174
rect 473866 330938 474102 331174
rect 473546 330618 473782 330854
rect 473866 330618 474102 330854
rect 473546 294938 473782 295174
rect 473866 294938 474102 295174
rect 473546 294618 473782 294854
rect 473866 294618 474102 294854
rect 473546 258938 473782 259174
rect 473866 258938 474102 259174
rect 473546 258618 473782 258854
rect 473866 258618 474102 258854
rect 473546 222938 473782 223174
rect 473866 222938 474102 223174
rect 473546 222618 473782 222854
rect 473866 222618 474102 222854
rect 473546 186938 473782 187174
rect 473866 186938 474102 187174
rect 473546 186618 473782 186854
rect 473866 186618 474102 186854
rect 473546 150938 473782 151174
rect 473866 150938 474102 151174
rect 473546 150618 473782 150854
rect 473866 150618 474102 150854
rect 473546 114938 473782 115174
rect 473866 114938 474102 115174
rect 473546 114618 473782 114854
rect 473866 114618 474102 114854
rect 473546 78938 473782 79174
rect 473866 78938 474102 79174
rect 473546 78618 473782 78854
rect 473866 78618 474102 78854
rect 473546 42938 473782 43174
rect 473866 42938 474102 43174
rect 473546 42618 473782 42854
rect 473866 42618 474102 42854
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -2502 473782 -2266
rect 473866 -2502 474102 -2266
rect 473546 -2822 473782 -2586
rect 473866 -2822 474102 -2586
rect 477266 694658 477502 694894
rect 477586 694658 477822 694894
rect 477266 694338 477502 694574
rect 477586 694338 477822 694574
rect 477266 658658 477502 658894
rect 477586 658658 477822 658894
rect 477266 658338 477502 658574
rect 477586 658338 477822 658574
rect 477266 622658 477502 622894
rect 477586 622658 477822 622894
rect 477266 622338 477502 622574
rect 477586 622338 477822 622574
rect 477266 586658 477502 586894
rect 477586 586658 477822 586894
rect 477266 586338 477502 586574
rect 477586 586338 477822 586574
rect 477266 550658 477502 550894
rect 477586 550658 477822 550894
rect 477266 550338 477502 550574
rect 477586 550338 477822 550574
rect 477266 514658 477502 514894
rect 477586 514658 477822 514894
rect 477266 514338 477502 514574
rect 477586 514338 477822 514574
rect 477266 478658 477502 478894
rect 477586 478658 477822 478894
rect 477266 478338 477502 478574
rect 477586 478338 477822 478574
rect 477266 442658 477502 442894
rect 477586 442658 477822 442894
rect 477266 442338 477502 442574
rect 477586 442338 477822 442574
rect 477266 406658 477502 406894
rect 477586 406658 477822 406894
rect 477266 406338 477502 406574
rect 477586 406338 477822 406574
rect 477266 370658 477502 370894
rect 477586 370658 477822 370894
rect 477266 370338 477502 370574
rect 477586 370338 477822 370574
rect 477266 334658 477502 334894
rect 477586 334658 477822 334894
rect 477266 334338 477502 334574
rect 477586 334338 477822 334574
rect 477266 298658 477502 298894
rect 477586 298658 477822 298894
rect 477266 298338 477502 298574
rect 477586 298338 477822 298574
rect 477266 262658 477502 262894
rect 477586 262658 477822 262894
rect 477266 262338 477502 262574
rect 477586 262338 477822 262574
rect 477266 226658 477502 226894
rect 477586 226658 477822 226894
rect 477266 226338 477502 226574
rect 477586 226338 477822 226574
rect 477266 190658 477502 190894
rect 477586 190658 477822 190894
rect 477266 190338 477502 190574
rect 477586 190338 477822 190574
rect 477266 154658 477502 154894
rect 477586 154658 477822 154894
rect 477266 154338 477502 154574
rect 477586 154338 477822 154574
rect 477266 118658 477502 118894
rect 477586 118658 477822 118894
rect 477266 118338 477502 118574
rect 477586 118338 477822 118574
rect 477266 82658 477502 82894
rect 477586 82658 477822 82894
rect 477266 82338 477502 82574
rect 477586 82338 477822 82574
rect 477266 46658 477502 46894
rect 477586 46658 477822 46894
rect 477266 46338 477502 46574
rect 477586 46338 477822 46574
rect 477266 10658 477502 10894
rect 477586 10658 477822 10894
rect 477266 10338 477502 10574
rect 477586 10338 477822 10574
rect 477266 -4422 477502 -4186
rect 477586 -4422 477822 -4186
rect 477266 -4742 477502 -4506
rect 477586 -4742 477822 -4506
rect 498986 711322 499222 711558
rect 499306 711322 499542 711558
rect 498986 711002 499222 711238
rect 499306 711002 499542 711238
rect 495266 709402 495502 709638
rect 495586 709402 495822 709638
rect 495266 709082 495502 709318
rect 495586 709082 495822 709318
rect 491546 707482 491782 707718
rect 491866 707482 492102 707718
rect 491546 707162 491782 707398
rect 491866 707162 492102 707398
rect 480986 698378 481222 698614
rect 481306 698378 481542 698614
rect 480986 698058 481222 698294
rect 481306 698058 481542 698294
rect 480986 662378 481222 662614
rect 481306 662378 481542 662614
rect 480986 662058 481222 662294
rect 481306 662058 481542 662294
rect 480986 626378 481222 626614
rect 481306 626378 481542 626614
rect 480986 626058 481222 626294
rect 481306 626058 481542 626294
rect 480986 590378 481222 590614
rect 481306 590378 481542 590614
rect 480986 590058 481222 590294
rect 481306 590058 481542 590294
rect 480986 554378 481222 554614
rect 481306 554378 481542 554614
rect 480986 554058 481222 554294
rect 481306 554058 481542 554294
rect 480986 518378 481222 518614
rect 481306 518378 481542 518614
rect 480986 518058 481222 518294
rect 481306 518058 481542 518294
rect 480986 482378 481222 482614
rect 481306 482378 481542 482614
rect 480986 482058 481222 482294
rect 481306 482058 481542 482294
rect 480986 446378 481222 446614
rect 481306 446378 481542 446614
rect 480986 446058 481222 446294
rect 481306 446058 481542 446294
rect 480986 410378 481222 410614
rect 481306 410378 481542 410614
rect 480986 410058 481222 410294
rect 481306 410058 481542 410294
rect 480986 374378 481222 374614
rect 481306 374378 481542 374614
rect 480986 374058 481222 374294
rect 481306 374058 481542 374294
rect 480986 338378 481222 338614
rect 481306 338378 481542 338614
rect 480986 338058 481222 338294
rect 481306 338058 481542 338294
rect 480986 302378 481222 302614
rect 481306 302378 481542 302614
rect 480986 302058 481222 302294
rect 481306 302058 481542 302294
rect 480986 266378 481222 266614
rect 481306 266378 481542 266614
rect 480986 266058 481222 266294
rect 481306 266058 481542 266294
rect 480986 230378 481222 230614
rect 481306 230378 481542 230614
rect 480986 230058 481222 230294
rect 481306 230058 481542 230294
rect 480986 194378 481222 194614
rect 481306 194378 481542 194614
rect 480986 194058 481222 194294
rect 481306 194058 481542 194294
rect 480986 158378 481222 158614
rect 481306 158378 481542 158614
rect 480986 158058 481222 158294
rect 481306 158058 481542 158294
rect 480986 122378 481222 122614
rect 481306 122378 481542 122614
rect 480986 122058 481222 122294
rect 481306 122058 481542 122294
rect 480986 86378 481222 86614
rect 481306 86378 481542 86614
rect 480986 86058 481222 86294
rect 481306 86058 481542 86294
rect 480986 50378 481222 50614
rect 481306 50378 481542 50614
rect 480986 50058 481222 50294
rect 481306 50058 481542 50294
rect 480986 14378 481222 14614
rect 481306 14378 481542 14614
rect 480986 14058 481222 14294
rect 481306 14058 481542 14294
rect 462986 -7302 463222 -7066
rect 463306 -7302 463542 -7066
rect 462986 -7622 463222 -7386
rect 463306 -7622 463542 -7386
rect 487826 705562 488062 705798
rect 488146 705562 488382 705798
rect 487826 705242 488062 705478
rect 488146 705242 488382 705478
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 487826 453218 488062 453454
rect 488146 453218 488382 453454
rect 487826 452898 488062 453134
rect 488146 452898 488382 453134
rect 487826 417218 488062 417454
rect 488146 417218 488382 417454
rect 487826 416898 488062 417134
rect 488146 416898 488382 417134
rect 487826 381218 488062 381454
rect 488146 381218 488382 381454
rect 487826 380898 488062 381134
rect 488146 380898 488382 381134
rect 487826 345218 488062 345454
rect 488146 345218 488382 345454
rect 487826 344898 488062 345134
rect 488146 344898 488382 345134
rect 487826 309218 488062 309454
rect 488146 309218 488382 309454
rect 487826 308898 488062 309134
rect 488146 308898 488382 309134
rect 487826 273218 488062 273454
rect 488146 273218 488382 273454
rect 487826 272898 488062 273134
rect 488146 272898 488382 273134
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 487826 129218 488062 129454
rect 488146 129218 488382 129454
rect 487826 128898 488062 129134
rect 488146 128898 488382 129134
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -1542 488062 -1306
rect 488146 -1542 488382 -1306
rect 487826 -1862 488062 -1626
rect 488146 -1862 488382 -1626
rect 491546 672938 491782 673174
rect 491866 672938 492102 673174
rect 491546 672618 491782 672854
rect 491866 672618 492102 672854
rect 491546 636938 491782 637174
rect 491866 636938 492102 637174
rect 491546 636618 491782 636854
rect 491866 636618 492102 636854
rect 491546 600938 491782 601174
rect 491866 600938 492102 601174
rect 491546 600618 491782 600854
rect 491866 600618 492102 600854
rect 491546 564938 491782 565174
rect 491866 564938 492102 565174
rect 491546 564618 491782 564854
rect 491866 564618 492102 564854
rect 491546 528938 491782 529174
rect 491866 528938 492102 529174
rect 491546 528618 491782 528854
rect 491866 528618 492102 528854
rect 491546 492938 491782 493174
rect 491866 492938 492102 493174
rect 491546 492618 491782 492854
rect 491866 492618 492102 492854
rect 491546 456938 491782 457174
rect 491866 456938 492102 457174
rect 491546 456618 491782 456854
rect 491866 456618 492102 456854
rect 491546 420938 491782 421174
rect 491866 420938 492102 421174
rect 491546 420618 491782 420854
rect 491866 420618 492102 420854
rect 491546 384938 491782 385174
rect 491866 384938 492102 385174
rect 491546 384618 491782 384854
rect 491866 384618 492102 384854
rect 491546 348938 491782 349174
rect 491866 348938 492102 349174
rect 491546 348618 491782 348854
rect 491866 348618 492102 348854
rect 491546 312938 491782 313174
rect 491866 312938 492102 313174
rect 491546 312618 491782 312854
rect 491866 312618 492102 312854
rect 491546 276938 491782 277174
rect 491866 276938 492102 277174
rect 491546 276618 491782 276854
rect 491866 276618 492102 276854
rect 491546 240938 491782 241174
rect 491866 240938 492102 241174
rect 491546 240618 491782 240854
rect 491866 240618 492102 240854
rect 491546 204938 491782 205174
rect 491866 204938 492102 205174
rect 491546 204618 491782 204854
rect 491866 204618 492102 204854
rect 491546 168938 491782 169174
rect 491866 168938 492102 169174
rect 491546 168618 491782 168854
rect 491866 168618 492102 168854
rect 491546 132938 491782 133174
rect 491866 132938 492102 133174
rect 491546 132618 491782 132854
rect 491866 132618 492102 132854
rect 491546 96938 491782 97174
rect 491866 96938 492102 97174
rect 491546 96618 491782 96854
rect 491866 96618 492102 96854
rect 491546 60938 491782 61174
rect 491866 60938 492102 61174
rect 491546 60618 491782 60854
rect 491866 60618 492102 60854
rect 491546 24938 491782 25174
rect 491866 24938 492102 25174
rect 491546 24618 491782 24854
rect 491866 24618 492102 24854
rect 491546 -3462 491782 -3226
rect 491866 -3462 492102 -3226
rect 491546 -3782 491782 -3546
rect 491866 -3782 492102 -3546
rect 495266 676658 495502 676894
rect 495586 676658 495822 676894
rect 495266 676338 495502 676574
rect 495586 676338 495822 676574
rect 495266 640658 495502 640894
rect 495586 640658 495822 640894
rect 495266 640338 495502 640574
rect 495586 640338 495822 640574
rect 495266 604658 495502 604894
rect 495586 604658 495822 604894
rect 495266 604338 495502 604574
rect 495586 604338 495822 604574
rect 495266 568658 495502 568894
rect 495586 568658 495822 568894
rect 495266 568338 495502 568574
rect 495586 568338 495822 568574
rect 495266 532658 495502 532894
rect 495586 532658 495822 532894
rect 495266 532338 495502 532574
rect 495586 532338 495822 532574
rect 495266 496658 495502 496894
rect 495586 496658 495822 496894
rect 495266 496338 495502 496574
rect 495586 496338 495822 496574
rect 495266 460658 495502 460894
rect 495586 460658 495822 460894
rect 495266 460338 495502 460574
rect 495586 460338 495822 460574
rect 495266 424658 495502 424894
rect 495586 424658 495822 424894
rect 495266 424338 495502 424574
rect 495586 424338 495822 424574
rect 495266 388658 495502 388894
rect 495586 388658 495822 388894
rect 495266 388338 495502 388574
rect 495586 388338 495822 388574
rect 495266 352658 495502 352894
rect 495586 352658 495822 352894
rect 495266 352338 495502 352574
rect 495586 352338 495822 352574
rect 495266 316658 495502 316894
rect 495586 316658 495822 316894
rect 495266 316338 495502 316574
rect 495586 316338 495822 316574
rect 495266 280658 495502 280894
rect 495586 280658 495822 280894
rect 495266 280338 495502 280574
rect 495586 280338 495822 280574
rect 495266 244658 495502 244894
rect 495586 244658 495822 244894
rect 495266 244338 495502 244574
rect 495586 244338 495822 244574
rect 495266 208658 495502 208894
rect 495586 208658 495822 208894
rect 495266 208338 495502 208574
rect 495586 208338 495822 208574
rect 495266 172658 495502 172894
rect 495586 172658 495822 172894
rect 495266 172338 495502 172574
rect 495586 172338 495822 172574
rect 495266 136658 495502 136894
rect 495586 136658 495822 136894
rect 495266 136338 495502 136574
rect 495586 136338 495822 136574
rect 495266 100658 495502 100894
rect 495586 100658 495822 100894
rect 495266 100338 495502 100574
rect 495586 100338 495822 100574
rect 495266 64658 495502 64894
rect 495586 64658 495822 64894
rect 495266 64338 495502 64574
rect 495586 64338 495822 64574
rect 495266 28658 495502 28894
rect 495586 28658 495822 28894
rect 495266 28338 495502 28574
rect 495586 28338 495822 28574
rect 495266 -5382 495502 -5146
rect 495586 -5382 495822 -5146
rect 495266 -5702 495502 -5466
rect 495586 -5702 495822 -5466
rect 516986 710362 517222 710598
rect 517306 710362 517542 710598
rect 516986 710042 517222 710278
rect 517306 710042 517542 710278
rect 513266 708442 513502 708678
rect 513586 708442 513822 708678
rect 513266 708122 513502 708358
rect 513586 708122 513822 708358
rect 509546 706522 509782 706758
rect 509866 706522 510102 706758
rect 509546 706202 509782 706438
rect 509866 706202 510102 706438
rect 498986 680378 499222 680614
rect 499306 680378 499542 680614
rect 498986 680058 499222 680294
rect 499306 680058 499542 680294
rect 498986 644378 499222 644614
rect 499306 644378 499542 644614
rect 498986 644058 499222 644294
rect 499306 644058 499542 644294
rect 498986 608378 499222 608614
rect 499306 608378 499542 608614
rect 498986 608058 499222 608294
rect 499306 608058 499542 608294
rect 498986 572378 499222 572614
rect 499306 572378 499542 572614
rect 498986 572058 499222 572294
rect 499306 572058 499542 572294
rect 498986 536378 499222 536614
rect 499306 536378 499542 536614
rect 498986 536058 499222 536294
rect 499306 536058 499542 536294
rect 498986 500378 499222 500614
rect 499306 500378 499542 500614
rect 498986 500058 499222 500294
rect 499306 500058 499542 500294
rect 498986 464378 499222 464614
rect 499306 464378 499542 464614
rect 498986 464058 499222 464294
rect 499306 464058 499542 464294
rect 498986 428378 499222 428614
rect 499306 428378 499542 428614
rect 498986 428058 499222 428294
rect 499306 428058 499542 428294
rect 498986 392378 499222 392614
rect 499306 392378 499542 392614
rect 498986 392058 499222 392294
rect 499306 392058 499542 392294
rect 498986 356378 499222 356614
rect 499306 356378 499542 356614
rect 498986 356058 499222 356294
rect 499306 356058 499542 356294
rect 498986 320378 499222 320614
rect 499306 320378 499542 320614
rect 498986 320058 499222 320294
rect 499306 320058 499542 320294
rect 498986 284378 499222 284614
rect 499306 284378 499542 284614
rect 498986 284058 499222 284294
rect 499306 284058 499542 284294
rect 498986 248378 499222 248614
rect 499306 248378 499542 248614
rect 498986 248058 499222 248294
rect 499306 248058 499542 248294
rect 498986 212378 499222 212614
rect 499306 212378 499542 212614
rect 498986 212058 499222 212294
rect 499306 212058 499542 212294
rect 498986 176378 499222 176614
rect 499306 176378 499542 176614
rect 498986 176058 499222 176294
rect 499306 176058 499542 176294
rect 498986 140378 499222 140614
rect 499306 140378 499542 140614
rect 498986 140058 499222 140294
rect 499306 140058 499542 140294
rect 498986 104378 499222 104614
rect 499306 104378 499542 104614
rect 498986 104058 499222 104294
rect 499306 104058 499542 104294
rect 498986 68378 499222 68614
rect 499306 68378 499542 68614
rect 498986 68058 499222 68294
rect 499306 68058 499542 68294
rect 498986 32378 499222 32614
rect 499306 32378 499542 32614
rect 498986 32058 499222 32294
rect 499306 32058 499542 32294
rect 480986 -6342 481222 -6106
rect 481306 -6342 481542 -6106
rect 480986 -6662 481222 -6426
rect 481306 -6662 481542 -6426
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 690938 509782 691174
rect 509866 690938 510102 691174
rect 509546 690618 509782 690854
rect 509866 690618 510102 690854
rect 509546 654938 509782 655174
rect 509866 654938 510102 655174
rect 509546 654618 509782 654854
rect 509866 654618 510102 654854
rect 509546 618938 509782 619174
rect 509866 618938 510102 619174
rect 509546 618618 509782 618854
rect 509866 618618 510102 618854
rect 509546 582938 509782 583174
rect 509866 582938 510102 583174
rect 509546 582618 509782 582854
rect 509866 582618 510102 582854
rect 509546 546938 509782 547174
rect 509866 546938 510102 547174
rect 509546 546618 509782 546854
rect 509866 546618 510102 546854
rect 509546 510938 509782 511174
rect 509866 510938 510102 511174
rect 509546 510618 509782 510854
rect 509866 510618 510102 510854
rect 509546 474938 509782 475174
rect 509866 474938 510102 475174
rect 509546 474618 509782 474854
rect 509866 474618 510102 474854
rect 509546 438938 509782 439174
rect 509866 438938 510102 439174
rect 509546 438618 509782 438854
rect 509866 438618 510102 438854
rect 509546 402938 509782 403174
rect 509866 402938 510102 403174
rect 509546 402618 509782 402854
rect 509866 402618 510102 402854
rect 509546 366938 509782 367174
rect 509866 366938 510102 367174
rect 509546 366618 509782 366854
rect 509866 366618 510102 366854
rect 509546 330938 509782 331174
rect 509866 330938 510102 331174
rect 509546 330618 509782 330854
rect 509866 330618 510102 330854
rect 509546 294938 509782 295174
rect 509866 294938 510102 295174
rect 509546 294618 509782 294854
rect 509866 294618 510102 294854
rect 509546 258938 509782 259174
rect 509866 258938 510102 259174
rect 509546 258618 509782 258854
rect 509866 258618 510102 258854
rect 509546 222938 509782 223174
rect 509866 222938 510102 223174
rect 509546 222618 509782 222854
rect 509866 222618 510102 222854
rect 509546 186938 509782 187174
rect 509866 186938 510102 187174
rect 509546 186618 509782 186854
rect 509866 186618 510102 186854
rect 509546 150938 509782 151174
rect 509866 150938 510102 151174
rect 509546 150618 509782 150854
rect 509866 150618 510102 150854
rect 509546 114938 509782 115174
rect 509866 114938 510102 115174
rect 509546 114618 509782 114854
rect 509866 114618 510102 114854
rect 509546 78938 509782 79174
rect 509866 78938 510102 79174
rect 509546 78618 509782 78854
rect 509866 78618 510102 78854
rect 509546 42938 509782 43174
rect 509866 42938 510102 43174
rect 509546 42618 509782 42854
rect 509866 42618 510102 42854
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -2502 509782 -2266
rect 509866 -2502 510102 -2266
rect 509546 -2822 509782 -2586
rect 509866 -2822 510102 -2586
rect 513266 694658 513502 694894
rect 513586 694658 513822 694894
rect 513266 694338 513502 694574
rect 513586 694338 513822 694574
rect 513266 658658 513502 658894
rect 513586 658658 513822 658894
rect 513266 658338 513502 658574
rect 513586 658338 513822 658574
rect 513266 622658 513502 622894
rect 513586 622658 513822 622894
rect 513266 622338 513502 622574
rect 513586 622338 513822 622574
rect 513266 586658 513502 586894
rect 513586 586658 513822 586894
rect 513266 586338 513502 586574
rect 513586 586338 513822 586574
rect 513266 550658 513502 550894
rect 513586 550658 513822 550894
rect 513266 550338 513502 550574
rect 513586 550338 513822 550574
rect 513266 514658 513502 514894
rect 513586 514658 513822 514894
rect 513266 514338 513502 514574
rect 513586 514338 513822 514574
rect 513266 478658 513502 478894
rect 513586 478658 513822 478894
rect 513266 478338 513502 478574
rect 513586 478338 513822 478574
rect 513266 442658 513502 442894
rect 513586 442658 513822 442894
rect 513266 442338 513502 442574
rect 513586 442338 513822 442574
rect 513266 406658 513502 406894
rect 513586 406658 513822 406894
rect 513266 406338 513502 406574
rect 513586 406338 513822 406574
rect 513266 370658 513502 370894
rect 513586 370658 513822 370894
rect 513266 370338 513502 370574
rect 513586 370338 513822 370574
rect 513266 334658 513502 334894
rect 513586 334658 513822 334894
rect 513266 334338 513502 334574
rect 513586 334338 513822 334574
rect 513266 298658 513502 298894
rect 513586 298658 513822 298894
rect 513266 298338 513502 298574
rect 513586 298338 513822 298574
rect 513266 262658 513502 262894
rect 513586 262658 513822 262894
rect 513266 262338 513502 262574
rect 513586 262338 513822 262574
rect 513266 226658 513502 226894
rect 513586 226658 513822 226894
rect 513266 226338 513502 226574
rect 513586 226338 513822 226574
rect 513266 190658 513502 190894
rect 513586 190658 513822 190894
rect 513266 190338 513502 190574
rect 513586 190338 513822 190574
rect 513266 154658 513502 154894
rect 513586 154658 513822 154894
rect 513266 154338 513502 154574
rect 513586 154338 513822 154574
rect 513266 118658 513502 118894
rect 513586 118658 513822 118894
rect 513266 118338 513502 118574
rect 513586 118338 513822 118574
rect 513266 82658 513502 82894
rect 513586 82658 513822 82894
rect 513266 82338 513502 82574
rect 513586 82338 513822 82574
rect 513266 46658 513502 46894
rect 513586 46658 513822 46894
rect 513266 46338 513502 46574
rect 513586 46338 513822 46574
rect 513266 10658 513502 10894
rect 513586 10658 513822 10894
rect 513266 10338 513502 10574
rect 513586 10338 513822 10574
rect 513266 -4422 513502 -4186
rect 513586 -4422 513822 -4186
rect 513266 -4742 513502 -4506
rect 513586 -4742 513822 -4506
rect 534986 711322 535222 711558
rect 535306 711322 535542 711558
rect 534986 711002 535222 711238
rect 535306 711002 535542 711238
rect 531266 709402 531502 709638
rect 531586 709402 531822 709638
rect 531266 709082 531502 709318
rect 531586 709082 531822 709318
rect 527546 707482 527782 707718
rect 527866 707482 528102 707718
rect 527546 707162 527782 707398
rect 527866 707162 528102 707398
rect 516986 698378 517222 698614
rect 517306 698378 517542 698614
rect 516986 698058 517222 698294
rect 517306 698058 517542 698294
rect 516986 662378 517222 662614
rect 517306 662378 517542 662614
rect 516986 662058 517222 662294
rect 517306 662058 517542 662294
rect 516986 626378 517222 626614
rect 517306 626378 517542 626614
rect 516986 626058 517222 626294
rect 517306 626058 517542 626294
rect 516986 590378 517222 590614
rect 517306 590378 517542 590614
rect 516986 590058 517222 590294
rect 517306 590058 517542 590294
rect 516986 554378 517222 554614
rect 517306 554378 517542 554614
rect 516986 554058 517222 554294
rect 517306 554058 517542 554294
rect 516986 518378 517222 518614
rect 517306 518378 517542 518614
rect 516986 518058 517222 518294
rect 517306 518058 517542 518294
rect 516986 482378 517222 482614
rect 517306 482378 517542 482614
rect 516986 482058 517222 482294
rect 517306 482058 517542 482294
rect 516986 446378 517222 446614
rect 517306 446378 517542 446614
rect 516986 446058 517222 446294
rect 517306 446058 517542 446294
rect 516986 410378 517222 410614
rect 517306 410378 517542 410614
rect 516986 410058 517222 410294
rect 517306 410058 517542 410294
rect 516986 374378 517222 374614
rect 517306 374378 517542 374614
rect 516986 374058 517222 374294
rect 517306 374058 517542 374294
rect 516986 338378 517222 338614
rect 517306 338378 517542 338614
rect 516986 338058 517222 338294
rect 517306 338058 517542 338294
rect 516986 302378 517222 302614
rect 517306 302378 517542 302614
rect 516986 302058 517222 302294
rect 517306 302058 517542 302294
rect 516986 266378 517222 266614
rect 517306 266378 517542 266614
rect 516986 266058 517222 266294
rect 517306 266058 517542 266294
rect 516986 230378 517222 230614
rect 517306 230378 517542 230614
rect 516986 230058 517222 230294
rect 517306 230058 517542 230294
rect 516986 194378 517222 194614
rect 517306 194378 517542 194614
rect 516986 194058 517222 194294
rect 517306 194058 517542 194294
rect 516986 158378 517222 158614
rect 517306 158378 517542 158614
rect 516986 158058 517222 158294
rect 517306 158058 517542 158294
rect 516986 122378 517222 122614
rect 517306 122378 517542 122614
rect 516986 122058 517222 122294
rect 517306 122058 517542 122294
rect 516986 86378 517222 86614
rect 517306 86378 517542 86614
rect 516986 86058 517222 86294
rect 517306 86058 517542 86294
rect 516986 50378 517222 50614
rect 517306 50378 517542 50614
rect 516986 50058 517222 50294
rect 517306 50058 517542 50294
rect 516986 14378 517222 14614
rect 517306 14378 517542 14614
rect 516986 14058 517222 14294
rect 517306 14058 517542 14294
rect 498986 -7302 499222 -7066
rect 499306 -7302 499542 -7066
rect 498986 -7622 499222 -7386
rect 499306 -7622 499542 -7386
rect 523826 705562 524062 705798
rect 524146 705562 524382 705798
rect 523826 705242 524062 705478
rect 524146 705242 524382 705478
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -1542 524062 -1306
rect 524146 -1542 524382 -1306
rect 523826 -1862 524062 -1626
rect 524146 -1862 524382 -1626
rect 527546 672938 527782 673174
rect 527866 672938 528102 673174
rect 527546 672618 527782 672854
rect 527866 672618 528102 672854
rect 527546 636938 527782 637174
rect 527866 636938 528102 637174
rect 527546 636618 527782 636854
rect 527866 636618 528102 636854
rect 527546 600938 527782 601174
rect 527866 600938 528102 601174
rect 527546 600618 527782 600854
rect 527866 600618 528102 600854
rect 527546 564938 527782 565174
rect 527866 564938 528102 565174
rect 527546 564618 527782 564854
rect 527866 564618 528102 564854
rect 527546 528938 527782 529174
rect 527866 528938 528102 529174
rect 527546 528618 527782 528854
rect 527866 528618 528102 528854
rect 527546 492938 527782 493174
rect 527866 492938 528102 493174
rect 527546 492618 527782 492854
rect 527866 492618 528102 492854
rect 527546 456938 527782 457174
rect 527866 456938 528102 457174
rect 527546 456618 527782 456854
rect 527866 456618 528102 456854
rect 527546 420938 527782 421174
rect 527866 420938 528102 421174
rect 527546 420618 527782 420854
rect 527866 420618 528102 420854
rect 527546 384938 527782 385174
rect 527866 384938 528102 385174
rect 527546 384618 527782 384854
rect 527866 384618 528102 384854
rect 527546 348938 527782 349174
rect 527866 348938 528102 349174
rect 527546 348618 527782 348854
rect 527866 348618 528102 348854
rect 527546 312938 527782 313174
rect 527866 312938 528102 313174
rect 527546 312618 527782 312854
rect 527866 312618 528102 312854
rect 527546 276938 527782 277174
rect 527866 276938 528102 277174
rect 527546 276618 527782 276854
rect 527866 276618 528102 276854
rect 527546 240938 527782 241174
rect 527866 240938 528102 241174
rect 527546 240618 527782 240854
rect 527866 240618 528102 240854
rect 527546 204938 527782 205174
rect 527866 204938 528102 205174
rect 527546 204618 527782 204854
rect 527866 204618 528102 204854
rect 527546 168938 527782 169174
rect 527866 168938 528102 169174
rect 527546 168618 527782 168854
rect 527866 168618 528102 168854
rect 527546 132938 527782 133174
rect 527866 132938 528102 133174
rect 527546 132618 527782 132854
rect 527866 132618 528102 132854
rect 527546 96938 527782 97174
rect 527866 96938 528102 97174
rect 527546 96618 527782 96854
rect 527866 96618 528102 96854
rect 527546 60938 527782 61174
rect 527866 60938 528102 61174
rect 527546 60618 527782 60854
rect 527866 60618 528102 60854
rect 527546 24938 527782 25174
rect 527866 24938 528102 25174
rect 527546 24618 527782 24854
rect 527866 24618 528102 24854
rect 527546 -3462 527782 -3226
rect 527866 -3462 528102 -3226
rect 527546 -3782 527782 -3546
rect 527866 -3782 528102 -3546
rect 531266 676658 531502 676894
rect 531586 676658 531822 676894
rect 531266 676338 531502 676574
rect 531586 676338 531822 676574
rect 531266 640658 531502 640894
rect 531586 640658 531822 640894
rect 531266 640338 531502 640574
rect 531586 640338 531822 640574
rect 531266 604658 531502 604894
rect 531586 604658 531822 604894
rect 531266 604338 531502 604574
rect 531586 604338 531822 604574
rect 531266 568658 531502 568894
rect 531586 568658 531822 568894
rect 531266 568338 531502 568574
rect 531586 568338 531822 568574
rect 531266 532658 531502 532894
rect 531586 532658 531822 532894
rect 531266 532338 531502 532574
rect 531586 532338 531822 532574
rect 531266 496658 531502 496894
rect 531586 496658 531822 496894
rect 531266 496338 531502 496574
rect 531586 496338 531822 496574
rect 531266 460658 531502 460894
rect 531586 460658 531822 460894
rect 531266 460338 531502 460574
rect 531586 460338 531822 460574
rect 531266 424658 531502 424894
rect 531586 424658 531822 424894
rect 531266 424338 531502 424574
rect 531586 424338 531822 424574
rect 531266 388658 531502 388894
rect 531586 388658 531822 388894
rect 531266 388338 531502 388574
rect 531586 388338 531822 388574
rect 531266 352658 531502 352894
rect 531586 352658 531822 352894
rect 531266 352338 531502 352574
rect 531586 352338 531822 352574
rect 531266 316658 531502 316894
rect 531586 316658 531822 316894
rect 531266 316338 531502 316574
rect 531586 316338 531822 316574
rect 531266 280658 531502 280894
rect 531586 280658 531822 280894
rect 531266 280338 531502 280574
rect 531586 280338 531822 280574
rect 531266 244658 531502 244894
rect 531586 244658 531822 244894
rect 531266 244338 531502 244574
rect 531586 244338 531822 244574
rect 531266 208658 531502 208894
rect 531586 208658 531822 208894
rect 531266 208338 531502 208574
rect 531586 208338 531822 208574
rect 531266 172658 531502 172894
rect 531586 172658 531822 172894
rect 531266 172338 531502 172574
rect 531586 172338 531822 172574
rect 531266 136658 531502 136894
rect 531586 136658 531822 136894
rect 531266 136338 531502 136574
rect 531586 136338 531822 136574
rect 531266 100658 531502 100894
rect 531586 100658 531822 100894
rect 531266 100338 531502 100574
rect 531586 100338 531822 100574
rect 531266 64658 531502 64894
rect 531586 64658 531822 64894
rect 531266 64338 531502 64574
rect 531586 64338 531822 64574
rect 531266 28658 531502 28894
rect 531586 28658 531822 28894
rect 531266 28338 531502 28574
rect 531586 28338 531822 28574
rect 531266 -5382 531502 -5146
rect 531586 -5382 531822 -5146
rect 531266 -5702 531502 -5466
rect 531586 -5702 531822 -5466
rect 552986 710362 553222 710598
rect 553306 710362 553542 710598
rect 552986 710042 553222 710278
rect 553306 710042 553542 710278
rect 549266 708442 549502 708678
rect 549586 708442 549822 708678
rect 549266 708122 549502 708358
rect 549586 708122 549822 708358
rect 545546 706522 545782 706758
rect 545866 706522 546102 706758
rect 545546 706202 545782 706438
rect 545866 706202 546102 706438
rect 534986 680378 535222 680614
rect 535306 680378 535542 680614
rect 534986 680058 535222 680294
rect 535306 680058 535542 680294
rect 534986 644378 535222 644614
rect 535306 644378 535542 644614
rect 534986 644058 535222 644294
rect 535306 644058 535542 644294
rect 534986 608378 535222 608614
rect 535306 608378 535542 608614
rect 534986 608058 535222 608294
rect 535306 608058 535542 608294
rect 534986 572378 535222 572614
rect 535306 572378 535542 572614
rect 534986 572058 535222 572294
rect 535306 572058 535542 572294
rect 534986 536378 535222 536614
rect 535306 536378 535542 536614
rect 534986 536058 535222 536294
rect 535306 536058 535542 536294
rect 534986 500378 535222 500614
rect 535306 500378 535542 500614
rect 534986 500058 535222 500294
rect 535306 500058 535542 500294
rect 534986 464378 535222 464614
rect 535306 464378 535542 464614
rect 534986 464058 535222 464294
rect 535306 464058 535542 464294
rect 534986 428378 535222 428614
rect 535306 428378 535542 428614
rect 534986 428058 535222 428294
rect 535306 428058 535542 428294
rect 534986 392378 535222 392614
rect 535306 392378 535542 392614
rect 534986 392058 535222 392294
rect 535306 392058 535542 392294
rect 534986 356378 535222 356614
rect 535306 356378 535542 356614
rect 534986 356058 535222 356294
rect 535306 356058 535542 356294
rect 534986 320378 535222 320614
rect 535306 320378 535542 320614
rect 534986 320058 535222 320294
rect 535306 320058 535542 320294
rect 534986 284378 535222 284614
rect 535306 284378 535542 284614
rect 534986 284058 535222 284294
rect 535306 284058 535542 284294
rect 534986 248378 535222 248614
rect 535306 248378 535542 248614
rect 534986 248058 535222 248294
rect 535306 248058 535542 248294
rect 534986 212378 535222 212614
rect 535306 212378 535542 212614
rect 534986 212058 535222 212294
rect 535306 212058 535542 212294
rect 534986 176378 535222 176614
rect 535306 176378 535542 176614
rect 534986 176058 535222 176294
rect 535306 176058 535542 176294
rect 534986 140378 535222 140614
rect 535306 140378 535542 140614
rect 534986 140058 535222 140294
rect 535306 140058 535542 140294
rect 534986 104378 535222 104614
rect 535306 104378 535542 104614
rect 534986 104058 535222 104294
rect 535306 104058 535542 104294
rect 534986 68378 535222 68614
rect 535306 68378 535542 68614
rect 534986 68058 535222 68294
rect 535306 68058 535542 68294
rect 534986 32378 535222 32614
rect 535306 32378 535542 32614
rect 534986 32058 535222 32294
rect 535306 32058 535542 32294
rect 516986 -6342 517222 -6106
rect 517306 -6342 517542 -6106
rect 516986 -6662 517222 -6426
rect 517306 -6662 517542 -6426
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 690938 545782 691174
rect 545866 690938 546102 691174
rect 545546 690618 545782 690854
rect 545866 690618 546102 690854
rect 545546 654938 545782 655174
rect 545866 654938 546102 655174
rect 545546 654618 545782 654854
rect 545866 654618 546102 654854
rect 545546 618938 545782 619174
rect 545866 618938 546102 619174
rect 545546 618618 545782 618854
rect 545866 618618 546102 618854
rect 545546 582938 545782 583174
rect 545866 582938 546102 583174
rect 545546 582618 545782 582854
rect 545866 582618 546102 582854
rect 545546 546938 545782 547174
rect 545866 546938 546102 547174
rect 545546 546618 545782 546854
rect 545866 546618 546102 546854
rect 545546 510938 545782 511174
rect 545866 510938 546102 511174
rect 545546 510618 545782 510854
rect 545866 510618 546102 510854
rect 545546 474938 545782 475174
rect 545866 474938 546102 475174
rect 545546 474618 545782 474854
rect 545866 474618 546102 474854
rect 545546 438938 545782 439174
rect 545866 438938 546102 439174
rect 545546 438618 545782 438854
rect 545866 438618 546102 438854
rect 545546 402938 545782 403174
rect 545866 402938 546102 403174
rect 545546 402618 545782 402854
rect 545866 402618 546102 402854
rect 545546 366938 545782 367174
rect 545866 366938 546102 367174
rect 545546 366618 545782 366854
rect 545866 366618 546102 366854
rect 545546 330938 545782 331174
rect 545866 330938 546102 331174
rect 545546 330618 545782 330854
rect 545866 330618 546102 330854
rect 545546 294938 545782 295174
rect 545866 294938 546102 295174
rect 545546 294618 545782 294854
rect 545866 294618 546102 294854
rect 545546 258938 545782 259174
rect 545866 258938 546102 259174
rect 545546 258618 545782 258854
rect 545866 258618 546102 258854
rect 545546 222938 545782 223174
rect 545866 222938 546102 223174
rect 545546 222618 545782 222854
rect 545866 222618 546102 222854
rect 545546 186938 545782 187174
rect 545866 186938 546102 187174
rect 545546 186618 545782 186854
rect 545866 186618 546102 186854
rect 545546 150938 545782 151174
rect 545866 150938 546102 151174
rect 545546 150618 545782 150854
rect 545866 150618 546102 150854
rect 545546 114938 545782 115174
rect 545866 114938 546102 115174
rect 545546 114618 545782 114854
rect 545866 114618 546102 114854
rect 545546 78938 545782 79174
rect 545866 78938 546102 79174
rect 545546 78618 545782 78854
rect 545866 78618 546102 78854
rect 545546 42938 545782 43174
rect 545866 42938 546102 43174
rect 545546 42618 545782 42854
rect 545866 42618 546102 42854
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -2502 545782 -2266
rect 545866 -2502 546102 -2266
rect 545546 -2822 545782 -2586
rect 545866 -2822 546102 -2586
rect 549266 694658 549502 694894
rect 549586 694658 549822 694894
rect 549266 694338 549502 694574
rect 549586 694338 549822 694574
rect 549266 658658 549502 658894
rect 549586 658658 549822 658894
rect 549266 658338 549502 658574
rect 549586 658338 549822 658574
rect 549266 622658 549502 622894
rect 549586 622658 549822 622894
rect 549266 622338 549502 622574
rect 549586 622338 549822 622574
rect 549266 586658 549502 586894
rect 549586 586658 549822 586894
rect 549266 586338 549502 586574
rect 549586 586338 549822 586574
rect 549266 550658 549502 550894
rect 549586 550658 549822 550894
rect 549266 550338 549502 550574
rect 549586 550338 549822 550574
rect 549266 514658 549502 514894
rect 549586 514658 549822 514894
rect 549266 514338 549502 514574
rect 549586 514338 549822 514574
rect 549266 478658 549502 478894
rect 549586 478658 549822 478894
rect 549266 478338 549502 478574
rect 549586 478338 549822 478574
rect 549266 442658 549502 442894
rect 549586 442658 549822 442894
rect 549266 442338 549502 442574
rect 549586 442338 549822 442574
rect 549266 406658 549502 406894
rect 549586 406658 549822 406894
rect 549266 406338 549502 406574
rect 549586 406338 549822 406574
rect 549266 370658 549502 370894
rect 549586 370658 549822 370894
rect 549266 370338 549502 370574
rect 549586 370338 549822 370574
rect 549266 334658 549502 334894
rect 549586 334658 549822 334894
rect 549266 334338 549502 334574
rect 549586 334338 549822 334574
rect 549266 298658 549502 298894
rect 549586 298658 549822 298894
rect 549266 298338 549502 298574
rect 549586 298338 549822 298574
rect 549266 262658 549502 262894
rect 549586 262658 549822 262894
rect 549266 262338 549502 262574
rect 549586 262338 549822 262574
rect 549266 226658 549502 226894
rect 549586 226658 549822 226894
rect 549266 226338 549502 226574
rect 549586 226338 549822 226574
rect 549266 190658 549502 190894
rect 549586 190658 549822 190894
rect 549266 190338 549502 190574
rect 549586 190338 549822 190574
rect 549266 154658 549502 154894
rect 549586 154658 549822 154894
rect 549266 154338 549502 154574
rect 549586 154338 549822 154574
rect 549266 118658 549502 118894
rect 549586 118658 549822 118894
rect 549266 118338 549502 118574
rect 549586 118338 549822 118574
rect 549266 82658 549502 82894
rect 549586 82658 549822 82894
rect 549266 82338 549502 82574
rect 549586 82338 549822 82574
rect 549266 46658 549502 46894
rect 549586 46658 549822 46894
rect 549266 46338 549502 46574
rect 549586 46338 549822 46574
rect 549266 10658 549502 10894
rect 549586 10658 549822 10894
rect 549266 10338 549502 10574
rect 549586 10338 549822 10574
rect 549266 -4422 549502 -4186
rect 549586 -4422 549822 -4186
rect 549266 -4742 549502 -4506
rect 549586 -4742 549822 -4506
rect 570986 711322 571222 711558
rect 571306 711322 571542 711558
rect 570986 711002 571222 711238
rect 571306 711002 571542 711238
rect 567266 709402 567502 709638
rect 567586 709402 567822 709638
rect 567266 709082 567502 709318
rect 567586 709082 567822 709318
rect 563546 707482 563782 707718
rect 563866 707482 564102 707718
rect 563546 707162 563782 707398
rect 563866 707162 564102 707398
rect 552986 698378 553222 698614
rect 553306 698378 553542 698614
rect 552986 698058 553222 698294
rect 553306 698058 553542 698294
rect 552986 662378 553222 662614
rect 553306 662378 553542 662614
rect 552986 662058 553222 662294
rect 553306 662058 553542 662294
rect 552986 626378 553222 626614
rect 553306 626378 553542 626614
rect 552986 626058 553222 626294
rect 553306 626058 553542 626294
rect 552986 590378 553222 590614
rect 553306 590378 553542 590614
rect 552986 590058 553222 590294
rect 553306 590058 553542 590294
rect 552986 554378 553222 554614
rect 553306 554378 553542 554614
rect 552986 554058 553222 554294
rect 553306 554058 553542 554294
rect 552986 518378 553222 518614
rect 553306 518378 553542 518614
rect 552986 518058 553222 518294
rect 553306 518058 553542 518294
rect 552986 482378 553222 482614
rect 553306 482378 553542 482614
rect 552986 482058 553222 482294
rect 553306 482058 553542 482294
rect 552986 446378 553222 446614
rect 553306 446378 553542 446614
rect 552986 446058 553222 446294
rect 553306 446058 553542 446294
rect 552986 410378 553222 410614
rect 553306 410378 553542 410614
rect 552986 410058 553222 410294
rect 553306 410058 553542 410294
rect 552986 374378 553222 374614
rect 553306 374378 553542 374614
rect 552986 374058 553222 374294
rect 553306 374058 553542 374294
rect 552986 338378 553222 338614
rect 553306 338378 553542 338614
rect 552986 338058 553222 338294
rect 553306 338058 553542 338294
rect 552986 302378 553222 302614
rect 553306 302378 553542 302614
rect 552986 302058 553222 302294
rect 553306 302058 553542 302294
rect 552986 266378 553222 266614
rect 553306 266378 553542 266614
rect 552986 266058 553222 266294
rect 553306 266058 553542 266294
rect 552986 230378 553222 230614
rect 553306 230378 553542 230614
rect 552986 230058 553222 230294
rect 553306 230058 553542 230294
rect 552986 194378 553222 194614
rect 553306 194378 553542 194614
rect 552986 194058 553222 194294
rect 553306 194058 553542 194294
rect 552986 158378 553222 158614
rect 553306 158378 553542 158614
rect 552986 158058 553222 158294
rect 553306 158058 553542 158294
rect 552986 122378 553222 122614
rect 553306 122378 553542 122614
rect 552986 122058 553222 122294
rect 553306 122058 553542 122294
rect 552986 86378 553222 86614
rect 553306 86378 553542 86614
rect 552986 86058 553222 86294
rect 553306 86058 553542 86294
rect 552986 50378 553222 50614
rect 553306 50378 553542 50614
rect 552986 50058 553222 50294
rect 553306 50058 553542 50294
rect 552986 14378 553222 14614
rect 553306 14378 553542 14614
rect 552986 14058 553222 14294
rect 553306 14058 553542 14294
rect 534986 -7302 535222 -7066
rect 535306 -7302 535542 -7066
rect 534986 -7622 535222 -7386
rect 535306 -7622 535542 -7386
rect 559826 705562 560062 705798
rect 560146 705562 560382 705798
rect 559826 705242 560062 705478
rect 560146 705242 560382 705478
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -1542 560062 -1306
rect 560146 -1542 560382 -1306
rect 559826 -1862 560062 -1626
rect 560146 -1862 560382 -1626
rect 563546 672938 563782 673174
rect 563866 672938 564102 673174
rect 563546 672618 563782 672854
rect 563866 672618 564102 672854
rect 563546 636938 563782 637174
rect 563866 636938 564102 637174
rect 563546 636618 563782 636854
rect 563866 636618 564102 636854
rect 563546 600938 563782 601174
rect 563866 600938 564102 601174
rect 563546 600618 563782 600854
rect 563866 600618 564102 600854
rect 563546 564938 563782 565174
rect 563866 564938 564102 565174
rect 563546 564618 563782 564854
rect 563866 564618 564102 564854
rect 563546 528938 563782 529174
rect 563866 528938 564102 529174
rect 563546 528618 563782 528854
rect 563866 528618 564102 528854
rect 563546 492938 563782 493174
rect 563866 492938 564102 493174
rect 563546 492618 563782 492854
rect 563866 492618 564102 492854
rect 563546 456938 563782 457174
rect 563866 456938 564102 457174
rect 563546 456618 563782 456854
rect 563866 456618 564102 456854
rect 563546 420938 563782 421174
rect 563866 420938 564102 421174
rect 563546 420618 563782 420854
rect 563866 420618 564102 420854
rect 563546 384938 563782 385174
rect 563866 384938 564102 385174
rect 563546 384618 563782 384854
rect 563866 384618 564102 384854
rect 563546 348938 563782 349174
rect 563866 348938 564102 349174
rect 563546 348618 563782 348854
rect 563866 348618 564102 348854
rect 563546 312938 563782 313174
rect 563866 312938 564102 313174
rect 563546 312618 563782 312854
rect 563866 312618 564102 312854
rect 563546 276938 563782 277174
rect 563866 276938 564102 277174
rect 563546 276618 563782 276854
rect 563866 276618 564102 276854
rect 563546 240938 563782 241174
rect 563866 240938 564102 241174
rect 563546 240618 563782 240854
rect 563866 240618 564102 240854
rect 563546 204938 563782 205174
rect 563866 204938 564102 205174
rect 563546 204618 563782 204854
rect 563866 204618 564102 204854
rect 563546 168938 563782 169174
rect 563866 168938 564102 169174
rect 563546 168618 563782 168854
rect 563866 168618 564102 168854
rect 563546 132938 563782 133174
rect 563866 132938 564102 133174
rect 563546 132618 563782 132854
rect 563866 132618 564102 132854
rect 563546 96938 563782 97174
rect 563866 96938 564102 97174
rect 563546 96618 563782 96854
rect 563866 96618 564102 96854
rect 563546 60938 563782 61174
rect 563866 60938 564102 61174
rect 563546 60618 563782 60854
rect 563866 60618 564102 60854
rect 563546 24938 563782 25174
rect 563866 24938 564102 25174
rect 563546 24618 563782 24854
rect 563866 24618 564102 24854
rect 563546 -3462 563782 -3226
rect 563866 -3462 564102 -3226
rect 563546 -3782 563782 -3546
rect 563866 -3782 564102 -3546
rect 567266 676658 567502 676894
rect 567586 676658 567822 676894
rect 567266 676338 567502 676574
rect 567586 676338 567822 676574
rect 567266 640658 567502 640894
rect 567586 640658 567822 640894
rect 567266 640338 567502 640574
rect 567586 640338 567822 640574
rect 567266 604658 567502 604894
rect 567586 604658 567822 604894
rect 567266 604338 567502 604574
rect 567586 604338 567822 604574
rect 567266 568658 567502 568894
rect 567586 568658 567822 568894
rect 567266 568338 567502 568574
rect 567586 568338 567822 568574
rect 567266 532658 567502 532894
rect 567586 532658 567822 532894
rect 567266 532338 567502 532574
rect 567586 532338 567822 532574
rect 567266 496658 567502 496894
rect 567586 496658 567822 496894
rect 567266 496338 567502 496574
rect 567586 496338 567822 496574
rect 567266 460658 567502 460894
rect 567586 460658 567822 460894
rect 567266 460338 567502 460574
rect 567586 460338 567822 460574
rect 567266 424658 567502 424894
rect 567586 424658 567822 424894
rect 567266 424338 567502 424574
rect 567586 424338 567822 424574
rect 567266 388658 567502 388894
rect 567586 388658 567822 388894
rect 567266 388338 567502 388574
rect 567586 388338 567822 388574
rect 567266 352658 567502 352894
rect 567586 352658 567822 352894
rect 567266 352338 567502 352574
rect 567586 352338 567822 352574
rect 567266 316658 567502 316894
rect 567586 316658 567822 316894
rect 567266 316338 567502 316574
rect 567586 316338 567822 316574
rect 567266 280658 567502 280894
rect 567586 280658 567822 280894
rect 567266 280338 567502 280574
rect 567586 280338 567822 280574
rect 567266 244658 567502 244894
rect 567586 244658 567822 244894
rect 567266 244338 567502 244574
rect 567586 244338 567822 244574
rect 567266 208658 567502 208894
rect 567586 208658 567822 208894
rect 567266 208338 567502 208574
rect 567586 208338 567822 208574
rect 567266 172658 567502 172894
rect 567586 172658 567822 172894
rect 567266 172338 567502 172574
rect 567586 172338 567822 172574
rect 567266 136658 567502 136894
rect 567586 136658 567822 136894
rect 567266 136338 567502 136574
rect 567586 136338 567822 136574
rect 567266 100658 567502 100894
rect 567586 100658 567822 100894
rect 567266 100338 567502 100574
rect 567586 100338 567822 100574
rect 567266 64658 567502 64894
rect 567586 64658 567822 64894
rect 567266 64338 567502 64574
rect 567586 64338 567822 64574
rect 567266 28658 567502 28894
rect 567586 28658 567822 28894
rect 567266 28338 567502 28574
rect 567586 28338 567822 28574
rect 567266 -5382 567502 -5146
rect 567586 -5382 567822 -5146
rect 567266 -5702 567502 -5466
rect 567586 -5702 567822 -5466
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 581546 706522 581782 706758
rect 581866 706522 582102 706758
rect 581546 706202 581782 706438
rect 581866 706202 582102 706438
rect 570986 680378 571222 680614
rect 571306 680378 571542 680614
rect 570986 680058 571222 680294
rect 571306 680058 571542 680294
rect 570986 644378 571222 644614
rect 571306 644378 571542 644614
rect 570986 644058 571222 644294
rect 571306 644058 571542 644294
rect 570986 608378 571222 608614
rect 571306 608378 571542 608614
rect 570986 608058 571222 608294
rect 571306 608058 571542 608294
rect 570986 572378 571222 572614
rect 571306 572378 571542 572614
rect 570986 572058 571222 572294
rect 571306 572058 571542 572294
rect 570986 536378 571222 536614
rect 571306 536378 571542 536614
rect 570986 536058 571222 536294
rect 571306 536058 571542 536294
rect 570986 500378 571222 500614
rect 571306 500378 571542 500614
rect 570986 500058 571222 500294
rect 571306 500058 571542 500294
rect 570986 464378 571222 464614
rect 571306 464378 571542 464614
rect 570986 464058 571222 464294
rect 571306 464058 571542 464294
rect 570986 428378 571222 428614
rect 571306 428378 571542 428614
rect 570986 428058 571222 428294
rect 571306 428058 571542 428294
rect 570986 392378 571222 392614
rect 571306 392378 571542 392614
rect 570986 392058 571222 392294
rect 571306 392058 571542 392294
rect 570986 356378 571222 356614
rect 571306 356378 571542 356614
rect 570986 356058 571222 356294
rect 571306 356058 571542 356294
rect 570986 320378 571222 320614
rect 571306 320378 571542 320614
rect 570986 320058 571222 320294
rect 571306 320058 571542 320294
rect 570986 284378 571222 284614
rect 571306 284378 571542 284614
rect 570986 284058 571222 284294
rect 571306 284058 571542 284294
rect 570986 248378 571222 248614
rect 571306 248378 571542 248614
rect 570986 248058 571222 248294
rect 571306 248058 571542 248294
rect 570986 212378 571222 212614
rect 571306 212378 571542 212614
rect 570986 212058 571222 212294
rect 571306 212058 571542 212294
rect 570986 176378 571222 176614
rect 571306 176378 571542 176614
rect 570986 176058 571222 176294
rect 571306 176058 571542 176294
rect 570986 140378 571222 140614
rect 571306 140378 571542 140614
rect 570986 140058 571222 140294
rect 571306 140058 571542 140294
rect 570986 104378 571222 104614
rect 571306 104378 571542 104614
rect 570986 104058 571222 104294
rect 571306 104058 571542 104294
rect 570986 68378 571222 68614
rect 571306 68378 571542 68614
rect 570986 68058 571222 68294
rect 571306 68058 571542 68294
rect 570986 32378 571222 32614
rect 571306 32378 571542 32614
rect 570986 32058 571222 32294
rect 571306 32058 571542 32294
rect 552986 -6342 553222 -6106
rect 553306 -6342 553542 -6106
rect 552986 -6662 553222 -6426
rect 553306 -6662 553542 -6426
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 669218 586538 669454
rect 586622 669218 586858 669454
rect 586302 668898 586538 669134
rect 586622 668898 586858 669134
rect 586302 633218 586538 633454
rect 586622 633218 586858 633454
rect 586302 632898 586538 633134
rect 586622 632898 586858 633134
rect 586302 597218 586538 597454
rect 586622 597218 586858 597454
rect 586302 596898 586538 597134
rect 586622 596898 586858 597134
rect 586302 561218 586538 561454
rect 586622 561218 586858 561454
rect 586302 560898 586538 561134
rect 586622 560898 586858 561134
rect 586302 525218 586538 525454
rect 586622 525218 586858 525454
rect 586302 524898 586538 525134
rect 586622 524898 586858 525134
rect 586302 489218 586538 489454
rect 586622 489218 586858 489454
rect 586302 488898 586538 489134
rect 586622 488898 586858 489134
rect 586302 453218 586538 453454
rect 586622 453218 586858 453454
rect 586302 452898 586538 453134
rect 586622 452898 586858 453134
rect 586302 417218 586538 417454
rect 586622 417218 586858 417454
rect 586302 416898 586538 417134
rect 586622 416898 586858 417134
rect 586302 381218 586538 381454
rect 586622 381218 586858 381454
rect 586302 380898 586538 381134
rect 586622 380898 586858 381134
rect 586302 345218 586538 345454
rect 586622 345218 586858 345454
rect 586302 344898 586538 345134
rect 586622 344898 586858 345134
rect 586302 309218 586538 309454
rect 586622 309218 586858 309454
rect 586302 308898 586538 309134
rect 586622 308898 586858 309134
rect 586302 273218 586538 273454
rect 586622 273218 586858 273454
rect 586302 272898 586538 273134
rect 586622 272898 586858 273134
rect 586302 237218 586538 237454
rect 586622 237218 586858 237454
rect 586302 236898 586538 237134
rect 586622 236898 586858 237134
rect 586302 201218 586538 201454
rect 586622 201218 586858 201454
rect 586302 200898 586538 201134
rect 586622 200898 586858 201134
rect 586302 165218 586538 165454
rect 586622 165218 586858 165454
rect 586302 164898 586538 165134
rect 586622 164898 586858 165134
rect 586302 129218 586538 129454
rect 586622 129218 586858 129454
rect 586302 128898 586538 129134
rect 586622 128898 586858 129134
rect 586302 93218 586538 93454
rect 586622 93218 586858 93454
rect 586302 92898 586538 93134
rect 586622 92898 586858 93134
rect 586302 57218 586538 57454
rect 586622 57218 586858 57454
rect 586302 56898 586538 57134
rect 586622 56898 586858 57134
rect 586302 21218 586538 21454
rect 586622 21218 586858 21454
rect 586302 20898 586538 21134
rect 586622 20898 586858 21134
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 690938 587498 691174
rect 587582 690938 587818 691174
rect 587262 690618 587498 690854
rect 587582 690618 587818 690854
rect 587262 654938 587498 655174
rect 587582 654938 587818 655174
rect 587262 654618 587498 654854
rect 587582 654618 587818 654854
rect 587262 618938 587498 619174
rect 587582 618938 587818 619174
rect 587262 618618 587498 618854
rect 587582 618618 587818 618854
rect 587262 582938 587498 583174
rect 587582 582938 587818 583174
rect 587262 582618 587498 582854
rect 587582 582618 587818 582854
rect 587262 546938 587498 547174
rect 587582 546938 587818 547174
rect 587262 546618 587498 546854
rect 587582 546618 587818 546854
rect 587262 510938 587498 511174
rect 587582 510938 587818 511174
rect 587262 510618 587498 510854
rect 587582 510618 587818 510854
rect 587262 474938 587498 475174
rect 587582 474938 587818 475174
rect 587262 474618 587498 474854
rect 587582 474618 587818 474854
rect 587262 438938 587498 439174
rect 587582 438938 587818 439174
rect 587262 438618 587498 438854
rect 587582 438618 587818 438854
rect 587262 402938 587498 403174
rect 587582 402938 587818 403174
rect 587262 402618 587498 402854
rect 587582 402618 587818 402854
rect 587262 366938 587498 367174
rect 587582 366938 587818 367174
rect 587262 366618 587498 366854
rect 587582 366618 587818 366854
rect 587262 330938 587498 331174
rect 587582 330938 587818 331174
rect 587262 330618 587498 330854
rect 587582 330618 587818 330854
rect 587262 294938 587498 295174
rect 587582 294938 587818 295174
rect 587262 294618 587498 294854
rect 587582 294618 587818 294854
rect 587262 258938 587498 259174
rect 587582 258938 587818 259174
rect 587262 258618 587498 258854
rect 587582 258618 587818 258854
rect 587262 222938 587498 223174
rect 587582 222938 587818 223174
rect 587262 222618 587498 222854
rect 587582 222618 587818 222854
rect 587262 186938 587498 187174
rect 587582 186938 587818 187174
rect 587262 186618 587498 186854
rect 587582 186618 587818 186854
rect 587262 150938 587498 151174
rect 587582 150938 587818 151174
rect 587262 150618 587498 150854
rect 587582 150618 587818 150854
rect 587262 114938 587498 115174
rect 587582 114938 587818 115174
rect 587262 114618 587498 114854
rect 587582 114618 587818 114854
rect 587262 78938 587498 79174
rect 587582 78938 587818 79174
rect 587262 78618 587498 78854
rect 587582 78618 587818 78854
rect 587262 42938 587498 43174
rect 587582 42938 587818 43174
rect 587262 42618 587498 42854
rect 587582 42618 587818 42854
rect 587262 6938 587498 7174
rect 587582 6938 587818 7174
rect 587262 6618 587498 6854
rect 587582 6618 587818 6854
rect 581546 -2502 581782 -2266
rect 581866 -2502 582102 -2266
rect 581546 -2822 581782 -2586
rect 581866 -2822 582102 -2586
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 672938 588458 673174
rect 588542 672938 588778 673174
rect 588222 672618 588458 672854
rect 588542 672618 588778 672854
rect 588222 636938 588458 637174
rect 588542 636938 588778 637174
rect 588222 636618 588458 636854
rect 588542 636618 588778 636854
rect 588222 600938 588458 601174
rect 588542 600938 588778 601174
rect 588222 600618 588458 600854
rect 588542 600618 588778 600854
rect 588222 564938 588458 565174
rect 588542 564938 588778 565174
rect 588222 564618 588458 564854
rect 588542 564618 588778 564854
rect 588222 528938 588458 529174
rect 588542 528938 588778 529174
rect 588222 528618 588458 528854
rect 588542 528618 588778 528854
rect 588222 492938 588458 493174
rect 588542 492938 588778 493174
rect 588222 492618 588458 492854
rect 588542 492618 588778 492854
rect 588222 456938 588458 457174
rect 588542 456938 588778 457174
rect 588222 456618 588458 456854
rect 588542 456618 588778 456854
rect 588222 420938 588458 421174
rect 588542 420938 588778 421174
rect 588222 420618 588458 420854
rect 588542 420618 588778 420854
rect 588222 384938 588458 385174
rect 588542 384938 588778 385174
rect 588222 384618 588458 384854
rect 588542 384618 588778 384854
rect 588222 348938 588458 349174
rect 588542 348938 588778 349174
rect 588222 348618 588458 348854
rect 588542 348618 588778 348854
rect 588222 312938 588458 313174
rect 588542 312938 588778 313174
rect 588222 312618 588458 312854
rect 588542 312618 588778 312854
rect 588222 276938 588458 277174
rect 588542 276938 588778 277174
rect 588222 276618 588458 276854
rect 588542 276618 588778 276854
rect 588222 240938 588458 241174
rect 588542 240938 588778 241174
rect 588222 240618 588458 240854
rect 588542 240618 588778 240854
rect 588222 204938 588458 205174
rect 588542 204938 588778 205174
rect 588222 204618 588458 204854
rect 588542 204618 588778 204854
rect 588222 168938 588458 169174
rect 588542 168938 588778 169174
rect 588222 168618 588458 168854
rect 588542 168618 588778 168854
rect 588222 132938 588458 133174
rect 588542 132938 588778 133174
rect 588222 132618 588458 132854
rect 588542 132618 588778 132854
rect 588222 96938 588458 97174
rect 588542 96938 588778 97174
rect 588222 96618 588458 96854
rect 588542 96618 588778 96854
rect 588222 60938 588458 61174
rect 588542 60938 588778 61174
rect 588222 60618 588458 60854
rect 588542 60618 588778 60854
rect 588222 24938 588458 25174
rect 588542 24938 588778 25174
rect 588222 24618 588458 24854
rect 588542 24618 588778 24854
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 694658 589418 694894
rect 589502 694658 589738 694894
rect 589182 694338 589418 694574
rect 589502 694338 589738 694574
rect 589182 658658 589418 658894
rect 589502 658658 589738 658894
rect 589182 658338 589418 658574
rect 589502 658338 589738 658574
rect 589182 622658 589418 622894
rect 589502 622658 589738 622894
rect 589182 622338 589418 622574
rect 589502 622338 589738 622574
rect 589182 586658 589418 586894
rect 589502 586658 589738 586894
rect 589182 586338 589418 586574
rect 589502 586338 589738 586574
rect 589182 550658 589418 550894
rect 589502 550658 589738 550894
rect 589182 550338 589418 550574
rect 589502 550338 589738 550574
rect 589182 514658 589418 514894
rect 589502 514658 589738 514894
rect 589182 514338 589418 514574
rect 589502 514338 589738 514574
rect 589182 478658 589418 478894
rect 589502 478658 589738 478894
rect 589182 478338 589418 478574
rect 589502 478338 589738 478574
rect 589182 442658 589418 442894
rect 589502 442658 589738 442894
rect 589182 442338 589418 442574
rect 589502 442338 589738 442574
rect 589182 406658 589418 406894
rect 589502 406658 589738 406894
rect 589182 406338 589418 406574
rect 589502 406338 589738 406574
rect 589182 370658 589418 370894
rect 589502 370658 589738 370894
rect 589182 370338 589418 370574
rect 589502 370338 589738 370574
rect 589182 334658 589418 334894
rect 589502 334658 589738 334894
rect 589182 334338 589418 334574
rect 589502 334338 589738 334574
rect 589182 298658 589418 298894
rect 589502 298658 589738 298894
rect 589182 298338 589418 298574
rect 589502 298338 589738 298574
rect 589182 262658 589418 262894
rect 589502 262658 589738 262894
rect 589182 262338 589418 262574
rect 589502 262338 589738 262574
rect 589182 226658 589418 226894
rect 589502 226658 589738 226894
rect 589182 226338 589418 226574
rect 589502 226338 589738 226574
rect 589182 190658 589418 190894
rect 589502 190658 589738 190894
rect 589182 190338 589418 190574
rect 589502 190338 589738 190574
rect 589182 154658 589418 154894
rect 589502 154658 589738 154894
rect 589182 154338 589418 154574
rect 589502 154338 589738 154574
rect 589182 118658 589418 118894
rect 589502 118658 589738 118894
rect 589182 118338 589418 118574
rect 589502 118338 589738 118574
rect 589182 82658 589418 82894
rect 589502 82658 589738 82894
rect 589182 82338 589418 82574
rect 589502 82338 589738 82574
rect 589182 46658 589418 46894
rect 589502 46658 589738 46894
rect 589182 46338 589418 46574
rect 589502 46338 589738 46574
rect 589182 10658 589418 10894
rect 589502 10658 589738 10894
rect 589182 10338 589418 10574
rect 589502 10338 589738 10574
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 676658 590378 676894
rect 590462 676658 590698 676894
rect 590142 676338 590378 676574
rect 590462 676338 590698 676574
rect 590142 640658 590378 640894
rect 590462 640658 590698 640894
rect 590142 640338 590378 640574
rect 590462 640338 590698 640574
rect 590142 604658 590378 604894
rect 590462 604658 590698 604894
rect 590142 604338 590378 604574
rect 590462 604338 590698 604574
rect 590142 568658 590378 568894
rect 590462 568658 590698 568894
rect 590142 568338 590378 568574
rect 590462 568338 590698 568574
rect 590142 532658 590378 532894
rect 590462 532658 590698 532894
rect 590142 532338 590378 532574
rect 590462 532338 590698 532574
rect 590142 496658 590378 496894
rect 590462 496658 590698 496894
rect 590142 496338 590378 496574
rect 590462 496338 590698 496574
rect 590142 460658 590378 460894
rect 590462 460658 590698 460894
rect 590142 460338 590378 460574
rect 590462 460338 590698 460574
rect 590142 424658 590378 424894
rect 590462 424658 590698 424894
rect 590142 424338 590378 424574
rect 590462 424338 590698 424574
rect 590142 388658 590378 388894
rect 590462 388658 590698 388894
rect 590142 388338 590378 388574
rect 590462 388338 590698 388574
rect 590142 352658 590378 352894
rect 590462 352658 590698 352894
rect 590142 352338 590378 352574
rect 590462 352338 590698 352574
rect 590142 316658 590378 316894
rect 590462 316658 590698 316894
rect 590142 316338 590378 316574
rect 590462 316338 590698 316574
rect 590142 280658 590378 280894
rect 590462 280658 590698 280894
rect 590142 280338 590378 280574
rect 590462 280338 590698 280574
rect 590142 244658 590378 244894
rect 590462 244658 590698 244894
rect 590142 244338 590378 244574
rect 590462 244338 590698 244574
rect 590142 208658 590378 208894
rect 590462 208658 590698 208894
rect 590142 208338 590378 208574
rect 590462 208338 590698 208574
rect 590142 172658 590378 172894
rect 590462 172658 590698 172894
rect 590142 172338 590378 172574
rect 590462 172338 590698 172574
rect 590142 136658 590378 136894
rect 590462 136658 590698 136894
rect 590142 136338 590378 136574
rect 590462 136338 590698 136574
rect 590142 100658 590378 100894
rect 590462 100658 590698 100894
rect 590142 100338 590378 100574
rect 590462 100338 590698 100574
rect 590142 64658 590378 64894
rect 590462 64658 590698 64894
rect 590142 64338 590378 64574
rect 590462 64338 590698 64574
rect 590142 28658 590378 28894
rect 590462 28658 590698 28894
rect 590142 28338 590378 28574
rect 590462 28338 590698 28574
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 698378 591338 698614
rect 591422 698378 591658 698614
rect 591102 698058 591338 698294
rect 591422 698058 591658 698294
rect 591102 662378 591338 662614
rect 591422 662378 591658 662614
rect 591102 662058 591338 662294
rect 591422 662058 591658 662294
rect 591102 626378 591338 626614
rect 591422 626378 591658 626614
rect 591102 626058 591338 626294
rect 591422 626058 591658 626294
rect 591102 590378 591338 590614
rect 591422 590378 591658 590614
rect 591102 590058 591338 590294
rect 591422 590058 591658 590294
rect 591102 554378 591338 554614
rect 591422 554378 591658 554614
rect 591102 554058 591338 554294
rect 591422 554058 591658 554294
rect 591102 518378 591338 518614
rect 591422 518378 591658 518614
rect 591102 518058 591338 518294
rect 591422 518058 591658 518294
rect 591102 482378 591338 482614
rect 591422 482378 591658 482614
rect 591102 482058 591338 482294
rect 591422 482058 591658 482294
rect 591102 446378 591338 446614
rect 591422 446378 591658 446614
rect 591102 446058 591338 446294
rect 591422 446058 591658 446294
rect 591102 410378 591338 410614
rect 591422 410378 591658 410614
rect 591102 410058 591338 410294
rect 591422 410058 591658 410294
rect 591102 374378 591338 374614
rect 591422 374378 591658 374614
rect 591102 374058 591338 374294
rect 591422 374058 591658 374294
rect 591102 338378 591338 338614
rect 591422 338378 591658 338614
rect 591102 338058 591338 338294
rect 591422 338058 591658 338294
rect 591102 302378 591338 302614
rect 591422 302378 591658 302614
rect 591102 302058 591338 302294
rect 591422 302058 591658 302294
rect 591102 266378 591338 266614
rect 591422 266378 591658 266614
rect 591102 266058 591338 266294
rect 591422 266058 591658 266294
rect 591102 230378 591338 230614
rect 591422 230378 591658 230614
rect 591102 230058 591338 230294
rect 591422 230058 591658 230294
rect 591102 194378 591338 194614
rect 591422 194378 591658 194614
rect 591102 194058 591338 194294
rect 591422 194058 591658 194294
rect 591102 158378 591338 158614
rect 591422 158378 591658 158614
rect 591102 158058 591338 158294
rect 591422 158058 591658 158294
rect 591102 122378 591338 122614
rect 591422 122378 591658 122614
rect 591102 122058 591338 122294
rect 591422 122058 591658 122294
rect 591102 86378 591338 86614
rect 591422 86378 591658 86614
rect 591102 86058 591338 86294
rect 591422 86058 591658 86294
rect 591102 50378 591338 50614
rect 591422 50378 591658 50614
rect 591102 50058 591338 50294
rect 591422 50058 591658 50294
rect 591102 14378 591338 14614
rect 591422 14378 591658 14614
rect 591102 14058 591338 14294
rect 591422 14058 591658 14294
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 680378 592298 680614
rect 592382 680378 592618 680614
rect 592062 680058 592298 680294
rect 592382 680058 592618 680294
rect 592062 644378 592298 644614
rect 592382 644378 592618 644614
rect 592062 644058 592298 644294
rect 592382 644058 592618 644294
rect 592062 608378 592298 608614
rect 592382 608378 592618 608614
rect 592062 608058 592298 608294
rect 592382 608058 592618 608294
rect 592062 572378 592298 572614
rect 592382 572378 592618 572614
rect 592062 572058 592298 572294
rect 592382 572058 592618 572294
rect 592062 536378 592298 536614
rect 592382 536378 592618 536614
rect 592062 536058 592298 536294
rect 592382 536058 592618 536294
rect 592062 500378 592298 500614
rect 592382 500378 592618 500614
rect 592062 500058 592298 500294
rect 592382 500058 592618 500294
rect 592062 464378 592298 464614
rect 592382 464378 592618 464614
rect 592062 464058 592298 464294
rect 592382 464058 592618 464294
rect 592062 428378 592298 428614
rect 592382 428378 592618 428614
rect 592062 428058 592298 428294
rect 592382 428058 592618 428294
rect 592062 392378 592298 392614
rect 592382 392378 592618 392614
rect 592062 392058 592298 392294
rect 592382 392058 592618 392294
rect 592062 356378 592298 356614
rect 592382 356378 592618 356614
rect 592062 356058 592298 356294
rect 592382 356058 592618 356294
rect 592062 320378 592298 320614
rect 592382 320378 592618 320614
rect 592062 320058 592298 320294
rect 592382 320058 592618 320294
rect 592062 284378 592298 284614
rect 592382 284378 592618 284614
rect 592062 284058 592298 284294
rect 592382 284058 592618 284294
rect 592062 248378 592298 248614
rect 592382 248378 592618 248614
rect 592062 248058 592298 248294
rect 592382 248058 592618 248294
rect 592062 212378 592298 212614
rect 592382 212378 592618 212614
rect 592062 212058 592298 212294
rect 592382 212058 592618 212294
rect 592062 176378 592298 176614
rect 592382 176378 592618 176614
rect 592062 176058 592298 176294
rect 592382 176058 592618 176294
rect 592062 140378 592298 140614
rect 592382 140378 592618 140614
rect 592062 140058 592298 140294
rect 592382 140058 592618 140294
rect 592062 104378 592298 104614
rect 592382 104378 592618 104614
rect 592062 104058 592298 104294
rect 592382 104058 592618 104294
rect 592062 68378 592298 68614
rect 592382 68378 592618 68614
rect 592062 68058 592298 68294
rect 592382 68058 592618 68294
rect 592062 32378 592298 32614
rect 592382 32378 592618 32614
rect 592062 32058 592298 32294
rect 592382 32058 592618 32294
rect 570986 -7302 571222 -7066
rect 571306 -7302 571542 -7066
rect 570986 -7622 571222 -7386
rect 571306 -7622 571542 -7386
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 592650 698294
rect -8726 698026 592650 698058
rect -6806 694894 590730 694926
rect -6806 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 590730 694894
rect -6806 694574 590730 694658
rect -6806 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 590730 694574
rect -6806 694306 590730 694338
rect -4886 691174 588810 691206
rect -4886 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 588810 691174
rect -4886 690854 588810 690938
rect -4886 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 588810 690854
rect -4886 690586 588810 690618
rect -2966 687454 586890 687486
rect -2966 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 586890 687454
rect -2966 687134 586890 687218
rect -2966 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 586890 687134
rect -2966 686866 586890 686898
rect -8726 680614 592650 680646
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect -8726 680294 592650 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect -8726 680026 592650 680058
rect -6806 676894 590730 676926
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect -6806 676574 590730 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect -6806 676306 590730 676338
rect -4886 673174 588810 673206
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect -4886 672854 588810 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect -4886 672586 588810 672618
rect -2966 669454 586890 669486
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect -2966 669134 586890 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect -2966 668866 586890 668898
rect -8726 662614 592650 662646
rect -8726 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 592650 662294
rect -8726 662026 592650 662058
rect -6806 658894 590730 658926
rect -6806 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 590730 658894
rect -6806 658574 590730 658658
rect -6806 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 590730 658574
rect -6806 658306 590730 658338
rect -4886 655174 588810 655206
rect -4886 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 588810 655174
rect -4886 654854 588810 654938
rect -4886 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 588810 654854
rect -4886 654586 588810 654618
rect -2966 651454 586890 651486
rect -2966 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 586890 651454
rect -2966 651134 586890 651218
rect -2966 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 586890 651134
rect -2966 650866 586890 650898
rect -8726 644614 592650 644646
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect -8726 644294 592650 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect -8726 644026 592650 644058
rect -6806 640894 590730 640926
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect -6806 640574 590730 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect -6806 640306 590730 640338
rect -4886 637174 588810 637206
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect -4886 636854 588810 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect -4886 636586 588810 636618
rect -2966 633454 586890 633486
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect -2966 633134 586890 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect -2966 632866 586890 632898
rect -8726 626614 592650 626646
rect -8726 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 592650 626294
rect -8726 626026 592650 626058
rect -6806 622894 590730 622926
rect -6806 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 590730 622894
rect -6806 622574 590730 622658
rect -6806 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 590730 622574
rect -6806 622306 590730 622338
rect -4886 619174 588810 619206
rect -4886 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 588810 619174
rect -4886 618854 588810 618938
rect -4886 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 588810 618854
rect -4886 618586 588810 618618
rect -2966 615454 586890 615486
rect -2966 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 586890 615454
rect -2966 615134 586890 615218
rect -2966 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 586890 615134
rect -2966 614866 586890 614898
rect -8726 608614 592650 608646
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect -8726 608294 592650 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect -8726 608026 592650 608058
rect -6806 604894 590730 604926
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect -6806 604574 590730 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect -6806 604306 590730 604338
rect -4886 601174 588810 601206
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect -4886 600854 588810 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect -4886 600586 588810 600618
rect -2966 597454 586890 597486
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect -2966 597134 586890 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect -2966 596866 586890 596898
rect -8726 590614 592650 590646
rect -8726 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 592650 590294
rect -8726 590026 592650 590058
rect -6806 586894 590730 586926
rect -6806 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 590730 586894
rect -6806 586574 590730 586658
rect -6806 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 590730 586574
rect -6806 586306 590730 586338
rect -4886 583174 588810 583206
rect -4886 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 77546 583174
rect 77782 582938 77866 583174
rect 78102 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 588810 583174
rect -4886 582854 588810 582938
rect -4886 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 77546 582854
rect 77782 582618 77866 582854
rect 78102 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 588810 582854
rect -4886 582586 588810 582618
rect -2966 579454 586890 579486
rect -2966 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 586890 579454
rect -2966 579134 586890 579218
rect -2966 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 586890 579134
rect -2966 578866 586890 578898
rect -8726 572614 592650 572646
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect -8726 572294 592650 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect -8726 572026 592650 572058
rect -6806 568894 590730 568926
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect -6806 568574 590730 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect -6806 568306 590730 568338
rect -4886 565174 588810 565206
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 95546 565174
rect 95782 564938 95866 565174
rect 96102 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect -4886 564854 588810 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 95546 564854
rect 95782 564618 95866 564854
rect 96102 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect -4886 564586 588810 564618
rect -2966 561454 586890 561486
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect -2966 561134 586890 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect -2966 560866 586890 560898
rect -8726 554614 592650 554646
rect -8726 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 84986 554614
rect 85222 554378 85306 554614
rect 85542 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 84986 554294
rect 85222 554058 85306 554294
rect 85542 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 592650 554294
rect -8726 554026 592650 554058
rect -6806 550894 590730 550926
rect -6806 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 81266 550894
rect 81502 550658 81586 550894
rect 81822 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 590730 550894
rect -6806 550574 590730 550658
rect -6806 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 81266 550574
rect 81502 550338 81586 550574
rect 81822 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 590730 550574
rect -6806 550306 590730 550338
rect -4886 547174 588810 547206
rect -4886 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 77546 547174
rect 77782 546938 77866 547174
rect 78102 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 588810 547174
rect -4886 546854 588810 546938
rect -4886 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 77546 546854
rect 77782 546618 77866 546854
rect 78102 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 588810 546854
rect -4886 546586 588810 546618
rect -2966 543454 586890 543486
rect -2966 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 586890 543454
rect -2966 543134 586890 543218
rect -2966 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 586890 543134
rect -2966 542866 586890 542898
rect -8726 536614 592650 536646
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 174986 536614
rect 175222 536378 175306 536614
rect 175542 536378 210986 536614
rect 211222 536378 211306 536614
rect 211542 536378 246986 536614
rect 247222 536378 247306 536614
rect 247542 536378 282986 536614
rect 283222 536378 283306 536614
rect 283542 536378 318986 536614
rect 319222 536378 319306 536614
rect 319542 536378 354986 536614
rect 355222 536378 355306 536614
rect 355542 536378 390986 536614
rect 391222 536378 391306 536614
rect 391542 536378 426986 536614
rect 427222 536378 427306 536614
rect 427542 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect -8726 536294 592650 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 174986 536294
rect 175222 536058 175306 536294
rect 175542 536058 210986 536294
rect 211222 536058 211306 536294
rect 211542 536058 246986 536294
rect 247222 536058 247306 536294
rect 247542 536058 282986 536294
rect 283222 536058 283306 536294
rect 283542 536058 318986 536294
rect 319222 536058 319306 536294
rect 319542 536058 354986 536294
rect 355222 536058 355306 536294
rect 355542 536058 390986 536294
rect 391222 536058 391306 536294
rect 391542 536058 426986 536294
rect 427222 536058 427306 536294
rect 427542 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect -8726 536026 592650 536058
rect -6806 532894 590730 532926
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 171266 532894
rect 171502 532658 171586 532894
rect 171822 532658 207266 532894
rect 207502 532658 207586 532894
rect 207822 532658 243266 532894
rect 243502 532658 243586 532894
rect 243822 532658 279266 532894
rect 279502 532658 279586 532894
rect 279822 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 351266 532894
rect 351502 532658 351586 532894
rect 351822 532658 387266 532894
rect 387502 532658 387586 532894
rect 387822 532658 423266 532894
rect 423502 532658 423586 532894
rect 423822 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect -6806 532574 590730 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 171266 532574
rect 171502 532338 171586 532574
rect 171822 532338 207266 532574
rect 207502 532338 207586 532574
rect 207822 532338 243266 532574
rect 243502 532338 243586 532574
rect 243822 532338 279266 532574
rect 279502 532338 279586 532574
rect 279822 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 351266 532574
rect 351502 532338 351586 532574
rect 351822 532338 387266 532574
rect 387502 532338 387586 532574
rect 387822 532338 423266 532574
rect 423502 532338 423586 532574
rect 423822 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect -6806 532306 590730 532338
rect -4886 529174 588810 529206
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 167546 529174
rect 167782 528938 167866 529174
rect 168102 528938 203546 529174
rect 203782 528938 203866 529174
rect 204102 528938 239546 529174
rect 239782 528938 239866 529174
rect 240102 528938 275546 529174
rect 275782 528938 275866 529174
rect 276102 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 347546 529174
rect 347782 528938 347866 529174
rect 348102 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 419546 529174
rect 419782 528938 419866 529174
rect 420102 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect -4886 528854 588810 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 167546 528854
rect 167782 528618 167866 528854
rect 168102 528618 203546 528854
rect 203782 528618 203866 528854
rect 204102 528618 239546 528854
rect 239782 528618 239866 528854
rect 240102 528618 275546 528854
rect 275782 528618 275866 528854
rect 276102 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 347546 528854
rect 347782 528618 347866 528854
rect 348102 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 419546 528854
rect 419782 528618 419866 528854
rect 420102 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect -4886 528586 588810 528618
rect -2966 525454 586890 525486
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect -2966 525134 586890 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect -2966 524866 586890 524898
rect -8726 518614 592650 518646
rect -8726 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 592650 518294
rect -8726 518026 592650 518058
rect -6806 514894 590730 514926
rect -6806 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 590730 514894
rect -6806 514574 590730 514658
rect -6806 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 590730 514574
rect -6806 514306 590730 514338
rect -4886 511174 588810 511206
rect -4886 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 588810 511174
rect -4886 510854 588810 510938
rect -4886 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 588810 510854
rect -4886 510586 588810 510618
rect -2966 507454 586890 507486
rect -2966 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 586890 507454
rect -2966 507134 586890 507218
rect -2966 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 586890 507134
rect -2966 506866 586890 506898
rect -8726 500614 592650 500646
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 138986 500614
rect 139222 500378 139306 500614
rect 139542 500378 174986 500614
rect 175222 500378 175306 500614
rect 175542 500378 210986 500614
rect 211222 500378 211306 500614
rect 211542 500378 246986 500614
rect 247222 500378 247306 500614
rect 247542 500378 282986 500614
rect 283222 500378 283306 500614
rect 283542 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect -8726 500294 592650 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 138986 500294
rect 139222 500058 139306 500294
rect 139542 500058 174986 500294
rect 175222 500058 175306 500294
rect 175542 500058 210986 500294
rect 211222 500058 211306 500294
rect 211542 500058 246986 500294
rect 247222 500058 247306 500294
rect 247542 500058 282986 500294
rect 283222 500058 283306 500294
rect 283542 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect -8726 500026 592650 500058
rect -6806 496894 590730 496926
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 171266 496894
rect 171502 496658 171586 496894
rect 171822 496658 207266 496894
rect 207502 496658 207586 496894
rect 207822 496658 243266 496894
rect 243502 496658 243586 496894
rect 243822 496658 279266 496894
rect 279502 496658 279586 496894
rect 279822 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect -6806 496574 590730 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 171266 496574
rect 171502 496338 171586 496574
rect 171822 496338 207266 496574
rect 207502 496338 207586 496574
rect 207822 496338 243266 496574
rect 243502 496338 243586 496574
rect 243822 496338 279266 496574
rect 279502 496338 279586 496574
rect 279822 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect -6806 496306 590730 496338
rect -4886 493174 588810 493206
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 167546 493174
rect 167782 492938 167866 493174
rect 168102 492938 203546 493174
rect 203782 492938 203866 493174
rect 204102 492938 239546 493174
rect 239782 492938 239866 493174
rect 240102 492938 275546 493174
rect 275782 492938 275866 493174
rect 276102 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect -4886 492854 588810 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 167546 492854
rect 167782 492618 167866 492854
rect 168102 492618 203546 492854
rect 203782 492618 203866 492854
rect 204102 492618 239546 492854
rect 239782 492618 239866 492854
rect 240102 492618 275546 492854
rect 275782 492618 275866 492854
rect 276102 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect -4886 492586 588810 492618
rect -2966 489454 586890 489486
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect -2966 489134 586890 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect -2966 488866 586890 488898
rect -8726 482614 592650 482646
rect -8726 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 592650 482294
rect -8726 482026 592650 482058
rect -6806 478894 590730 478926
rect -6806 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 590730 478894
rect -6806 478574 590730 478658
rect -6806 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 590730 478574
rect -6806 478306 590730 478338
rect -4886 475174 588810 475206
rect -4886 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 588810 475174
rect -4886 474854 588810 474938
rect -4886 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 588810 474854
rect -4886 474586 588810 474618
rect -2966 471454 586890 471486
rect -2966 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 586890 471454
rect -2966 471134 586890 471218
rect -2966 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 586890 471134
rect -2966 470866 586890 470898
rect -8726 464614 592650 464646
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 102986 464614
rect 103222 464378 103306 464614
rect 103542 464378 138986 464614
rect 139222 464378 139306 464614
rect 139542 464378 174986 464614
rect 175222 464378 175306 464614
rect 175542 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 246986 464614
rect 247222 464378 247306 464614
rect 247542 464378 282986 464614
rect 283222 464378 283306 464614
rect 283542 464378 318986 464614
rect 319222 464378 319306 464614
rect 319542 464378 354986 464614
rect 355222 464378 355306 464614
rect 355542 464378 390986 464614
rect 391222 464378 391306 464614
rect 391542 464378 426986 464614
rect 427222 464378 427306 464614
rect 427542 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect -8726 464294 592650 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 102986 464294
rect 103222 464058 103306 464294
rect 103542 464058 138986 464294
rect 139222 464058 139306 464294
rect 139542 464058 174986 464294
rect 175222 464058 175306 464294
rect 175542 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 246986 464294
rect 247222 464058 247306 464294
rect 247542 464058 282986 464294
rect 283222 464058 283306 464294
rect 283542 464058 318986 464294
rect 319222 464058 319306 464294
rect 319542 464058 354986 464294
rect 355222 464058 355306 464294
rect 355542 464058 390986 464294
rect 391222 464058 391306 464294
rect 391542 464058 426986 464294
rect 427222 464058 427306 464294
rect 427542 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect -8726 464026 592650 464058
rect -6806 460894 590730 460926
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 99266 460894
rect 99502 460658 99586 460894
rect 99822 460658 135266 460894
rect 135502 460658 135586 460894
rect 135822 460658 171266 460894
rect 171502 460658 171586 460894
rect 171822 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 243266 460894
rect 243502 460658 243586 460894
rect 243822 460658 279266 460894
rect 279502 460658 279586 460894
rect 279822 460658 315266 460894
rect 315502 460658 315586 460894
rect 315822 460658 351266 460894
rect 351502 460658 351586 460894
rect 351822 460658 387266 460894
rect 387502 460658 387586 460894
rect 387822 460658 423266 460894
rect 423502 460658 423586 460894
rect 423822 460658 459266 460894
rect 459502 460658 459586 460894
rect 459822 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect -6806 460574 590730 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 99266 460574
rect 99502 460338 99586 460574
rect 99822 460338 135266 460574
rect 135502 460338 135586 460574
rect 135822 460338 171266 460574
rect 171502 460338 171586 460574
rect 171822 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 243266 460574
rect 243502 460338 243586 460574
rect 243822 460338 279266 460574
rect 279502 460338 279586 460574
rect 279822 460338 315266 460574
rect 315502 460338 315586 460574
rect 315822 460338 351266 460574
rect 351502 460338 351586 460574
rect 351822 460338 387266 460574
rect 387502 460338 387586 460574
rect 387822 460338 423266 460574
rect 423502 460338 423586 460574
rect 423822 460338 459266 460574
rect 459502 460338 459586 460574
rect 459822 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect -6806 460306 590730 460338
rect -4886 457174 588810 457206
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 95546 457174
rect 95782 456938 95866 457174
rect 96102 456938 131546 457174
rect 131782 456938 131866 457174
rect 132102 456938 167546 457174
rect 167782 456938 167866 457174
rect 168102 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 239546 457174
rect 239782 456938 239866 457174
rect 240102 456938 275546 457174
rect 275782 456938 275866 457174
rect 276102 456938 311546 457174
rect 311782 456938 311866 457174
rect 312102 456938 347546 457174
rect 347782 456938 347866 457174
rect 348102 456938 383546 457174
rect 383782 456938 383866 457174
rect 384102 456938 419546 457174
rect 419782 456938 419866 457174
rect 420102 456938 455546 457174
rect 455782 456938 455866 457174
rect 456102 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect -4886 456854 588810 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 95546 456854
rect 95782 456618 95866 456854
rect 96102 456618 131546 456854
rect 131782 456618 131866 456854
rect 132102 456618 167546 456854
rect 167782 456618 167866 456854
rect 168102 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 239546 456854
rect 239782 456618 239866 456854
rect 240102 456618 275546 456854
rect 275782 456618 275866 456854
rect 276102 456618 311546 456854
rect 311782 456618 311866 456854
rect 312102 456618 347546 456854
rect 347782 456618 347866 456854
rect 348102 456618 383546 456854
rect 383782 456618 383866 456854
rect 384102 456618 419546 456854
rect 419782 456618 419866 456854
rect 420102 456618 455546 456854
rect 455782 456618 455866 456854
rect 456102 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect -4886 456586 588810 456618
rect -2966 453454 586890 453486
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect -2966 453134 586890 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect -2966 452866 586890 452898
rect -8726 446614 592650 446646
rect -8726 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 84986 446614
rect 85222 446378 85306 446614
rect 85542 446378 120986 446614
rect 121222 446378 121306 446614
rect 121542 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 192986 446614
rect 193222 446378 193306 446614
rect 193542 446378 228986 446614
rect 229222 446378 229306 446614
rect 229542 446378 264986 446614
rect 265222 446378 265306 446614
rect 265542 446378 300986 446614
rect 301222 446378 301306 446614
rect 301542 446378 336986 446614
rect 337222 446378 337306 446614
rect 337542 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 84986 446294
rect 85222 446058 85306 446294
rect 85542 446058 120986 446294
rect 121222 446058 121306 446294
rect 121542 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 192986 446294
rect 193222 446058 193306 446294
rect 193542 446058 228986 446294
rect 229222 446058 229306 446294
rect 229542 446058 264986 446294
rect 265222 446058 265306 446294
rect 265542 446058 300986 446294
rect 301222 446058 301306 446294
rect 301542 446058 336986 446294
rect 337222 446058 337306 446294
rect 337542 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 592650 446294
rect -8726 446026 592650 446058
rect -6806 442894 590730 442926
rect -6806 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 81266 442894
rect 81502 442658 81586 442894
rect 81822 442658 117266 442894
rect 117502 442658 117586 442894
rect 117822 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 225266 442894
rect 225502 442658 225586 442894
rect 225822 442658 261266 442894
rect 261502 442658 261586 442894
rect 261822 442658 297266 442894
rect 297502 442658 297586 442894
rect 297822 442658 333266 442894
rect 333502 442658 333586 442894
rect 333822 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 441266 442894
rect 441502 442658 441586 442894
rect 441822 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 590730 442894
rect -6806 442574 590730 442658
rect -6806 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 81266 442574
rect 81502 442338 81586 442574
rect 81822 442338 117266 442574
rect 117502 442338 117586 442574
rect 117822 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 225266 442574
rect 225502 442338 225586 442574
rect 225822 442338 261266 442574
rect 261502 442338 261586 442574
rect 261822 442338 297266 442574
rect 297502 442338 297586 442574
rect 297822 442338 333266 442574
rect 333502 442338 333586 442574
rect 333822 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 441266 442574
rect 441502 442338 441586 442574
rect 441822 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 590730 442574
rect -6806 442306 590730 442338
rect -4886 439174 588810 439206
rect -4886 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 77546 439174
rect 77782 438938 77866 439174
rect 78102 438938 113546 439174
rect 113782 438938 113866 439174
rect 114102 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 221546 439174
rect 221782 438938 221866 439174
rect 222102 438938 257546 439174
rect 257782 438938 257866 439174
rect 258102 438938 293546 439174
rect 293782 438938 293866 439174
rect 294102 438938 329546 439174
rect 329782 438938 329866 439174
rect 330102 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 588810 439174
rect -4886 438854 588810 438938
rect -4886 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 77546 438854
rect 77782 438618 77866 438854
rect 78102 438618 113546 438854
rect 113782 438618 113866 438854
rect 114102 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 221546 438854
rect 221782 438618 221866 438854
rect 222102 438618 257546 438854
rect 257782 438618 257866 438854
rect 258102 438618 293546 438854
rect 293782 438618 293866 438854
rect 294102 438618 329546 438854
rect 329782 438618 329866 438854
rect 330102 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 588810 438854
rect -4886 438586 588810 438618
rect -2966 435454 586890 435486
rect -2966 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 586890 435454
rect -2966 435134 586890 435218
rect -2966 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 586890 435134
rect -2966 434866 586890 434898
rect -8726 428614 592650 428646
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 66986 428614
rect 67222 428378 67306 428614
rect 67542 428378 102986 428614
rect 103222 428378 103306 428614
rect 103542 428378 138986 428614
rect 139222 428378 139306 428614
rect 139542 428378 174986 428614
rect 175222 428378 175306 428614
rect 175542 428378 210986 428614
rect 211222 428378 211306 428614
rect 211542 428378 246986 428614
rect 247222 428378 247306 428614
rect 247542 428378 282986 428614
rect 283222 428378 283306 428614
rect 283542 428378 318986 428614
rect 319222 428378 319306 428614
rect 319542 428378 354986 428614
rect 355222 428378 355306 428614
rect 355542 428378 390986 428614
rect 391222 428378 391306 428614
rect 391542 428378 426986 428614
rect 427222 428378 427306 428614
rect 427542 428378 462986 428614
rect 463222 428378 463306 428614
rect 463542 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect -8726 428294 592650 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 66986 428294
rect 67222 428058 67306 428294
rect 67542 428058 102986 428294
rect 103222 428058 103306 428294
rect 103542 428058 138986 428294
rect 139222 428058 139306 428294
rect 139542 428058 174986 428294
rect 175222 428058 175306 428294
rect 175542 428058 210986 428294
rect 211222 428058 211306 428294
rect 211542 428058 246986 428294
rect 247222 428058 247306 428294
rect 247542 428058 282986 428294
rect 283222 428058 283306 428294
rect 283542 428058 318986 428294
rect 319222 428058 319306 428294
rect 319542 428058 354986 428294
rect 355222 428058 355306 428294
rect 355542 428058 390986 428294
rect 391222 428058 391306 428294
rect 391542 428058 426986 428294
rect 427222 428058 427306 428294
rect 427542 428058 462986 428294
rect 463222 428058 463306 428294
rect 463542 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect -8726 428026 592650 428058
rect -6806 424894 590730 424926
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 99266 424894
rect 99502 424658 99586 424894
rect 99822 424658 135266 424894
rect 135502 424658 135586 424894
rect 135822 424658 171266 424894
rect 171502 424658 171586 424894
rect 171822 424658 207266 424894
rect 207502 424658 207586 424894
rect 207822 424658 243266 424894
rect 243502 424658 243586 424894
rect 243822 424658 279266 424894
rect 279502 424658 279586 424894
rect 279822 424658 315266 424894
rect 315502 424658 315586 424894
rect 315822 424658 351266 424894
rect 351502 424658 351586 424894
rect 351822 424658 387266 424894
rect 387502 424658 387586 424894
rect 387822 424658 423266 424894
rect 423502 424658 423586 424894
rect 423822 424658 459266 424894
rect 459502 424658 459586 424894
rect 459822 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect -6806 424574 590730 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 99266 424574
rect 99502 424338 99586 424574
rect 99822 424338 135266 424574
rect 135502 424338 135586 424574
rect 135822 424338 171266 424574
rect 171502 424338 171586 424574
rect 171822 424338 207266 424574
rect 207502 424338 207586 424574
rect 207822 424338 243266 424574
rect 243502 424338 243586 424574
rect 243822 424338 279266 424574
rect 279502 424338 279586 424574
rect 279822 424338 315266 424574
rect 315502 424338 315586 424574
rect 315822 424338 351266 424574
rect 351502 424338 351586 424574
rect 351822 424338 387266 424574
rect 387502 424338 387586 424574
rect 387822 424338 423266 424574
rect 423502 424338 423586 424574
rect 423822 424338 459266 424574
rect 459502 424338 459586 424574
rect 459822 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect -6806 424306 590730 424338
rect -4886 421174 588810 421206
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 95546 421174
rect 95782 420938 95866 421174
rect 96102 420938 131546 421174
rect 131782 420938 131866 421174
rect 132102 420938 167546 421174
rect 167782 420938 167866 421174
rect 168102 420938 203546 421174
rect 203782 420938 203866 421174
rect 204102 420938 239546 421174
rect 239782 420938 239866 421174
rect 240102 420938 275546 421174
rect 275782 420938 275866 421174
rect 276102 420938 311546 421174
rect 311782 420938 311866 421174
rect 312102 420938 347546 421174
rect 347782 420938 347866 421174
rect 348102 420938 383546 421174
rect 383782 420938 383866 421174
rect 384102 420938 419546 421174
rect 419782 420938 419866 421174
rect 420102 420938 455546 421174
rect 455782 420938 455866 421174
rect 456102 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect -4886 420854 588810 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 95546 420854
rect 95782 420618 95866 420854
rect 96102 420618 131546 420854
rect 131782 420618 131866 420854
rect 132102 420618 167546 420854
rect 167782 420618 167866 420854
rect 168102 420618 203546 420854
rect 203782 420618 203866 420854
rect 204102 420618 239546 420854
rect 239782 420618 239866 420854
rect 240102 420618 275546 420854
rect 275782 420618 275866 420854
rect 276102 420618 311546 420854
rect 311782 420618 311866 420854
rect 312102 420618 347546 420854
rect 347782 420618 347866 420854
rect 348102 420618 383546 420854
rect 383782 420618 383866 420854
rect 384102 420618 419546 420854
rect 419782 420618 419866 420854
rect 420102 420618 455546 420854
rect 455782 420618 455866 420854
rect 456102 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect -4886 420586 588810 420618
rect -2966 417454 586890 417486
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect -2966 417134 586890 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect -2966 416866 586890 416898
rect -8726 410614 592650 410646
rect -8726 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 84986 410614
rect 85222 410378 85306 410614
rect 85542 410378 120986 410614
rect 121222 410378 121306 410614
rect 121542 410378 156986 410614
rect 157222 410378 157306 410614
rect 157542 410378 192986 410614
rect 193222 410378 193306 410614
rect 193542 410378 228986 410614
rect 229222 410378 229306 410614
rect 229542 410378 264986 410614
rect 265222 410378 265306 410614
rect 265542 410378 300986 410614
rect 301222 410378 301306 410614
rect 301542 410378 336986 410614
rect 337222 410378 337306 410614
rect 337542 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 84986 410294
rect 85222 410058 85306 410294
rect 85542 410058 120986 410294
rect 121222 410058 121306 410294
rect 121542 410058 156986 410294
rect 157222 410058 157306 410294
rect 157542 410058 192986 410294
rect 193222 410058 193306 410294
rect 193542 410058 228986 410294
rect 229222 410058 229306 410294
rect 229542 410058 264986 410294
rect 265222 410058 265306 410294
rect 265542 410058 300986 410294
rect 301222 410058 301306 410294
rect 301542 410058 336986 410294
rect 337222 410058 337306 410294
rect 337542 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 592650 410294
rect -8726 410026 592650 410058
rect -6806 406894 590730 406926
rect -6806 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 81266 406894
rect 81502 406658 81586 406894
rect 81822 406658 117266 406894
rect 117502 406658 117586 406894
rect 117822 406658 153266 406894
rect 153502 406658 153586 406894
rect 153822 406658 189266 406894
rect 189502 406658 189586 406894
rect 189822 406658 225266 406894
rect 225502 406658 225586 406894
rect 225822 406658 261266 406894
rect 261502 406658 261586 406894
rect 261822 406658 297266 406894
rect 297502 406658 297586 406894
rect 297822 406658 333266 406894
rect 333502 406658 333586 406894
rect 333822 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 590730 406894
rect -6806 406574 590730 406658
rect -6806 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 81266 406574
rect 81502 406338 81586 406574
rect 81822 406338 117266 406574
rect 117502 406338 117586 406574
rect 117822 406338 153266 406574
rect 153502 406338 153586 406574
rect 153822 406338 189266 406574
rect 189502 406338 189586 406574
rect 189822 406338 225266 406574
rect 225502 406338 225586 406574
rect 225822 406338 261266 406574
rect 261502 406338 261586 406574
rect 261822 406338 297266 406574
rect 297502 406338 297586 406574
rect 297822 406338 333266 406574
rect 333502 406338 333586 406574
rect 333822 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 590730 406574
rect -6806 406306 590730 406338
rect -4886 403174 588810 403206
rect -4886 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 77546 403174
rect 77782 402938 77866 403174
rect 78102 402938 113546 403174
rect 113782 402938 113866 403174
rect 114102 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 185546 403174
rect 185782 402938 185866 403174
rect 186102 402938 221546 403174
rect 221782 402938 221866 403174
rect 222102 402938 257546 403174
rect 257782 402938 257866 403174
rect 258102 402938 293546 403174
rect 293782 402938 293866 403174
rect 294102 402938 329546 403174
rect 329782 402938 329866 403174
rect 330102 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 588810 403174
rect -4886 402854 588810 402938
rect -4886 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 77546 402854
rect 77782 402618 77866 402854
rect 78102 402618 113546 402854
rect 113782 402618 113866 402854
rect 114102 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 185546 402854
rect 185782 402618 185866 402854
rect 186102 402618 221546 402854
rect 221782 402618 221866 402854
rect 222102 402618 257546 402854
rect 257782 402618 257866 402854
rect 258102 402618 293546 402854
rect 293782 402618 293866 402854
rect 294102 402618 329546 402854
rect 329782 402618 329866 402854
rect 330102 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 588810 402854
rect -4886 402586 588810 402618
rect -2966 399454 586890 399486
rect -2966 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 586890 399454
rect -2966 399134 586890 399218
rect -2966 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 586890 399134
rect -2966 398866 586890 398898
rect -8726 392614 592650 392646
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 66986 392614
rect 67222 392378 67306 392614
rect 67542 392378 102986 392614
rect 103222 392378 103306 392614
rect 103542 392378 138986 392614
rect 139222 392378 139306 392614
rect 139542 392378 174986 392614
rect 175222 392378 175306 392614
rect 175542 392378 210986 392614
rect 211222 392378 211306 392614
rect 211542 392378 246986 392614
rect 247222 392378 247306 392614
rect 247542 392378 282986 392614
rect 283222 392378 283306 392614
rect 283542 392378 318986 392614
rect 319222 392378 319306 392614
rect 319542 392378 354986 392614
rect 355222 392378 355306 392614
rect 355542 392378 390986 392614
rect 391222 392378 391306 392614
rect 391542 392378 426986 392614
rect 427222 392378 427306 392614
rect 427542 392378 462986 392614
rect 463222 392378 463306 392614
rect 463542 392378 498986 392614
rect 499222 392378 499306 392614
rect 499542 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect -8726 392294 592650 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 66986 392294
rect 67222 392058 67306 392294
rect 67542 392058 102986 392294
rect 103222 392058 103306 392294
rect 103542 392058 138986 392294
rect 139222 392058 139306 392294
rect 139542 392058 174986 392294
rect 175222 392058 175306 392294
rect 175542 392058 210986 392294
rect 211222 392058 211306 392294
rect 211542 392058 246986 392294
rect 247222 392058 247306 392294
rect 247542 392058 282986 392294
rect 283222 392058 283306 392294
rect 283542 392058 318986 392294
rect 319222 392058 319306 392294
rect 319542 392058 354986 392294
rect 355222 392058 355306 392294
rect 355542 392058 390986 392294
rect 391222 392058 391306 392294
rect 391542 392058 426986 392294
rect 427222 392058 427306 392294
rect 427542 392058 462986 392294
rect 463222 392058 463306 392294
rect 463542 392058 498986 392294
rect 499222 392058 499306 392294
rect 499542 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect -8726 392026 592650 392058
rect -6806 388894 590730 388926
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 99266 388894
rect 99502 388658 99586 388894
rect 99822 388658 135266 388894
rect 135502 388658 135586 388894
rect 135822 388658 171266 388894
rect 171502 388658 171586 388894
rect 171822 388658 207266 388894
rect 207502 388658 207586 388894
rect 207822 388658 243266 388894
rect 243502 388658 243586 388894
rect 243822 388658 279266 388894
rect 279502 388658 279586 388894
rect 279822 388658 315266 388894
rect 315502 388658 315586 388894
rect 315822 388658 351266 388894
rect 351502 388658 351586 388894
rect 351822 388658 387266 388894
rect 387502 388658 387586 388894
rect 387822 388658 423266 388894
rect 423502 388658 423586 388894
rect 423822 388658 459266 388894
rect 459502 388658 459586 388894
rect 459822 388658 495266 388894
rect 495502 388658 495586 388894
rect 495822 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect -6806 388574 590730 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 99266 388574
rect 99502 388338 99586 388574
rect 99822 388338 135266 388574
rect 135502 388338 135586 388574
rect 135822 388338 171266 388574
rect 171502 388338 171586 388574
rect 171822 388338 207266 388574
rect 207502 388338 207586 388574
rect 207822 388338 243266 388574
rect 243502 388338 243586 388574
rect 243822 388338 279266 388574
rect 279502 388338 279586 388574
rect 279822 388338 315266 388574
rect 315502 388338 315586 388574
rect 315822 388338 351266 388574
rect 351502 388338 351586 388574
rect 351822 388338 387266 388574
rect 387502 388338 387586 388574
rect 387822 388338 423266 388574
rect 423502 388338 423586 388574
rect 423822 388338 459266 388574
rect 459502 388338 459586 388574
rect 459822 388338 495266 388574
rect 495502 388338 495586 388574
rect 495822 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect -6806 388306 590730 388338
rect -4886 385174 588810 385206
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 59546 385174
rect 59782 384938 59866 385174
rect 60102 384938 95546 385174
rect 95782 384938 95866 385174
rect 96102 384938 131546 385174
rect 131782 384938 131866 385174
rect 132102 384938 167546 385174
rect 167782 384938 167866 385174
rect 168102 384938 203546 385174
rect 203782 384938 203866 385174
rect 204102 384938 239546 385174
rect 239782 384938 239866 385174
rect 240102 384938 275546 385174
rect 275782 384938 275866 385174
rect 276102 384938 311546 385174
rect 311782 384938 311866 385174
rect 312102 384938 347546 385174
rect 347782 384938 347866 385174
rect 348102 384938 383546 385174
rect 383782 384938 383866 385174
rect 384102 384938 419546 385174
rect 419782 384938 419866 385174
rect 420102 384938 455546 385174
rect 455782 384938 455866 385174
rect 456102 384938 491546 385174
rect 491782 384938 491866 385174
rect 492102 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect -4886 384854 588810 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 59546 384854
rect 59782 384618 59866 384854
rect 60102 384618 95546 384854
rect 95782 384618 95866 384854
rect 96102 384618 131546 384854
rect 131782 384618 131866 384854
rect 132102 384618 167546 384854
rect 167782 384618 167866 384854
rect 168102 384618 203546 384854
rect 203782 384618 203866 384854
rect 204102 384618 239546 384854
rect 239782 384618 239866 384854
rect 240102 384618 275546 384854
rect 275782 384618 275866 384854
rect 276102 384618 311546 384854
rect 311782 384618 311866 384854
rect 312102 384618 347546 384854
rect 347782 384618 347866 384854
rect 348102 384618 383546 384854
rect 383782 384618 383866 384854
rect 384102 384618 419546 384854
rect 419782 384618 419866 384854
rect 420102 384618 455546 384854
rect 455782 384618 455866 384854
rect 456102 384618 491546 384854
rect 491782 384618 491866 384854
rect 492102 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect -4886 384586 588810 384618
rect -2966 381454 586890 381486
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect -2966 381134 586890 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect -2966 380866 586890 380898
rect -8726 374614 592650 374646
rect -8726 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 264986 374614
rect 265222 374378 265306 374614
rect 265542 374378 300986 374614
rect 301222 374378 301306 374614
rect 301542 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 264986 374294
rect 265222 374058 265306 374294
rect 265542 374058 300986 374294
rect 301222 374058 301306 374294
rect 301542 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 592650 374294
rect -8726 374026 592650 374058
rect -6806 370894 590730 370926
rect -6806 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 261266 370894
rect 261502 370658 261586 370894
rect 261822 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 590730 370894
rect -6806 370574 590730 370658
rect -6806 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 261266 370574
rect 261502 370338 261586 370574
rect 261822 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 590730 370574
rect -6806 370306 590730 370338
rect -4886 367174 588810 367206
rect -4886 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 257546 367174
rect 257782 366938 257866 367174
rect 258102 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 588810 367174
rect -4886 366854 588810 366938
rect -4886 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 257546 366854
rect 257782 366618 257866 366854
rect 258102 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 588810 366854
rect -4886 366586 588810 366618
rect -2966 363454 586890 363486
rect -2966 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 362285 363454
rect 362521 363218 364882 363454
rect 365118 363218 367479 363454
rect 367715 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 434285 363454
rect 434521 363218 436882 363454
rect 437118 363218 439479 363454
rect 439715 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 586890 363454
rect -2966 363134 586890 363218
rect -2966 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 362285 363134
rect 362521 362898 364882 363134
rect 365118 362898 367479 363134
rect 367715 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 434285 363134
rect 434521 362898 436882 363134
rect 437118 362898 439479 363134
rect 439715 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 586890 363134
rect -2966 362866 586890 362898
rect -8726 356614 592650 356646
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 102986 356614
rect 103222 356378 103306 356614
rect 103542 356378 138986 356614
rect 139222 356378 139306 356614
rect 139542 356378 174986 356614
rect 175222 356378 175306 356614
rect 175542 356378 210986 356614
rect 211222 356378 211306 356614
rect 211542 356378 246986 356614
rect 247222 356378 247306 356614
rect 247542 356378 282986 356614
rect 283222 356378 283306 356614
rect 283542 356378 318986 356614
rect 319222 356378 319306 356614
rect 319542 356378 354986 356614
rect 355222 356378 355306 356614
rect 355542 356378 390986 356614
rect 391222 356378 391306 356614
rect 391542 356378 426986 356614
rect 427222 356378 427306 356614
rect 427542 356378 462986 356614
rect 463222 356378 463306 356614
rect 463542 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect -8726 356294 592650 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 102986 356294
rect 103222 356058 103306 356294
rect 103542 356058 138986 356294
rect 139222 356058 139306 356294
rect 139542 356058 174986 356294
rect 175222 356058 175306 356294
rect 175542 356058 210986 356294
rect 211222 356058 211306 356294
rect 211542 356058 246986 356294
rect 247222 356058 247306 356294
rect 247542 356058 282986 356294
rect 283222 356058 283306 356294
rect 283542 356058 318986 356294
rect 319222 356058 319306 356294
rect 319542 356058 354986 356294
rect 355222 356058 355306 356294
rect 355542 356058 390986 356294
rect 391222 356058 391306 356294
rect 391542 356058 426986 356294
rect 427222 356058 427306 356294
rect 427542 356058 462986 356294
rect 463222 356058 463306 356294
rect 463542 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect -8726 356026 592650 356058
rect -6806 352894 590730 352926
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 63266 352894
rect 63502 352658 63586 352894
rect 63822 352658 99266 352894
rect 99502 352658 99586 352894
rect 99822 352658 135266 352894
rect 135502 352658 135586 352894
rect 135822 352658 171266 352894
rect 171502 352658 171586 352894
rect 171822 352658 207266 352894
rect 207502 352658 207586 352894
rect 207822 352658 243266 352894
rect 243502 352658 243586 352894
rect 243822 352658 279266 352894
rect 279502 352658 279586 352894
rect 279822 352658 315266 352894
rect 315502 352658 315586 352894
rect 315822 352658 351266 352894
rect 351502 352658 351586 352894
rect 351822 352658 387266 352894
rect 387502 352658 387586 352894
rect 387822 352658 423266 352894
rect 423502 352658 423586 352894
rect 423822 352658 459266 352894
rect 459502 352658 459586 352894
rect 459822 352658 495266 352894
rect 495502 352658 495586 352894
rect 495822 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect -6806 352574 590730 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 63266 352574
rect 63502 352338 63586 352574
rect 63822 352338 99266 352574
rect 99502 352338 99586 352574
rect 99822 352338 135266 352574
rect 135502 352338 135586 352574
rect 135822 352338 171266 352574
rect 171502 352338 171586 352574
rect 171822 352338 207266 352574
rect 207502 352338 207586 352574
rect 207822 352338 243266 352574
rect 243502 352338 243586 352574
rect 243822 352338 279266 352574
rect 279502 352338 279586 352574
rect 279822 352338 315266 352574
rect 315502 352338 315586 352574
rect 315822 352338 351266 352574
rect 351502 352338 351586 352574
rect 351822 352338 387266 352574
rect 387502 352338 387586 352574
rect 387822 352338 423266 352574
rect 423502 352338 423586 352574
rect 423822 352338 459266 352574
rect 459502 352338 459586 352574
rect 459822 352338 495266 352574
rect 495502 352338 495586 352574
rect 495822 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect -6806 352306 590730 352338
rect -4886 349174 588810 349206
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 59546 349174
rect 59782 348938 59866 349174
rect 60102 348938 95546 349174
rect 95782 348938 95866 349174
rect 96102 348938 131546 349174
rect 131782 348938 131866 349174
rect 132102 348938 167546 349174
rect 167782 348938 167866 349174
rect 168102 348938 203546 349174
rect 203782 348938 203866 349174
rect 204102 348938 239546 349174
rect 239782 348938 239866 349174
rect 240102 348938 275546 349174
rect 275782 348938 275866 349174
rect 276102 348938 311546 349174
rect 311782 348938 311866 349174
rect 312102 348938 347546 349174
rect 347782 348938 347866 349174
rect 348102 348938 383546 349174
rect 383782 348938 383866 349174
rect 384102 348938 419546 349174
rect 419782 348938 419866 349174
rect 420102 348938 455546 349174
rect 455782 348938 455866 349174
rect 456102 348938 491546 349174
rect 491782 348938 491866 349174
rect 492102 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect -4886 348854 588810 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 59546 348854
rect 59782 348618 59866 348854
rect 60102 348618 95546 348854
rect 95782 348618 95866 348854
rect 96102 348618 131546 348854
rect 131782 348618 131866 348854
rect 132102 348618 167546 348854
rect 167782 348618 167866 348854
rect 168102 348618 203546 348854
rect 203782 348618 203866 348854
rect 204102 348618 239546 348854
rect 239782 348618 239866 348854
rect 240102 348618 275546 348854
rect 275782 348618 275866 348854
rect 276102 348618 311546 348854
rect 311782 348618 311866 348854
rect 312102 348618 347546 348854
rect 347782 348618 347866 348854
rect 348102 348618 383546 348854
rect 383782 348618 383866 348854
rect 384102 348618 419546 348854
rect 419782 348618 419866 348854
rect 420102 348618 455546 348854
rect 455782 348618 455866 348854
rect 456102 348618 491546 348854
rect 491782 348618 491866 348854
rect 492102 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect -4886 348586 588810 348618
rect -2966 345454 586890 345486
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 363583 345454
rect 363819 345218 366180 345454
rect 366416 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 435583 345454
rect 435819 345218 438180 345454
rect 438416 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect -2966 345134 586890 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 363583 345134
rect 363819 344898 366180 345134
rect 366416 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 435583 345134
rect 435819 344898 438180 345134
rect 438416 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect -2966 344866 586890 344898
rect -8726 338614 592650 338646
rect -8726 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 84986 338614
rect 85222 338378 85306 338614
rect 85542 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 192986 338614
rect 193222 338378 193306 338614
rect 193542 338378 228986 338614
rect 229222 338378 229306 338614
rect 229542 338378 264986 338614
rect 265222 338378 265306 338614
rect 265542 338378 300986 338614
rect 301222 338378 301306 338614
rect 301542 338378 336986 338614
rect 337222 338378 337306 338614
rect 337542 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 84986 338294
rect 85222 338058 85306 338294
rect 85542 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 192986 338294
rect 193222 338058 193306 338294
rect 193542 338058 228986 338294
rect 229222 338058 229306 338294
rect 229542 338058 264986 338294
rect 265222 338058 265306 338294
rect 265542 338058 300986 338294
rect 301222 338058 301306 338294
rect 301542 338058 336986 338294
rect 337222 338058 337306 338294
rect 337542 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 592650 338294
rect -8726 338026 592650 338058
rect -6806 334894 590730 334926
rect -6806 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 189266 334894
rect 189502 334658 189586 334894
rect 189822 334658 225266 334894
rect 225502 334658 225586 334894
rect 225822 334658 261266 334894
rect 261502 334658 261586 334894
rect 261822 334658 297266 334894
rect 297502 334658 297586 334894
rect 297822 334658 333266 334894
rect 333502 334658 333586 334894
rect 333822 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 590730 334894
rect -6806 334574 590730 334658
rect -6806 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 189266 334574
rect 189502 334338 189586 334574
rect 189822 334338 225266 334574
rect 225502 334338 225586 334574
rect 225822 334338 261266 334574
rect 261502 334338 261586 334574
rect 261822 334338 297266 334574
rect 297502 334338 297586 334574
rect 297822 334338 333266 334574
rect 333502 334338 333586 334574
rect 333822 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 590730 334574
rect -6806 334306 590730 334338
rect -4886 331174 588810 331206
rect -4886 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 113546 331174
rect 113782 330938 113866 331174
rect 114102 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 221546 331174
rect 221782 330938 221866 331174
rect 222102 330938 257546 331174
rect 257782 330938 257866 331174
rect 258102 330938 293546 331174
rect 293782 330938 293866 331174
rect 294102 330938 329546 331174
rect 329782 330938 329866 331174
rect 330102 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 588810 331174
rect -4886 330854 588810 330938
rect -4886 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 113546 330854
rect 113782 330618 113866 330854
rect 114102 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 221546 330854
rect 221782 330618 221866 330854
rect 222102 330618 257546 330854
rect 257782 330618 257866 330854
rect 258102 330618 293546 330854
rect 293782 330618 293866 330854
rect 294102 330618 329546 330854
rect 329782 330618 329866 330854
rect 330102 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 588810 330854
rect -4886 330586 588810 330618
rect -2966 327454 586890 327486
rect -2966 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 586890 327454
rect -2966 327134 586890 327218
rect -2966 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 586890 327134
rect -2966 326866 586890 326898
rect -8726 320614 592650 320646
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 66986 320614
rect 67222 320378 67306 320614
rect 67542 320378 102986 320614
rect 103222 320378 103306 320614
rect 103542 320378 138986 320614
rect 139222 320378 139306 320614
rect 139542 320378 174986 320614
rect 175222 320378 175306 320614
rect 175542 320378 210986 320614
rect 211222 320378 211306 320614
rect 211542 320378 246986 320614
rect 247222 320378 247306 320614
rect 247542 320378 282986 320614
rect 283222 320378 283306 320614
rect 283542 320378 318986 320614
rect 319222 320378 319306 320614
rect 319542 320378 354986 320614
rect 355222 320378 355306 320614
rect 355542 320378 390986 320614
rect 391222 320378 391306 320614
rect 391542 320378 426986 320614
rect 427222 320378 427306 320614
rect 427542 320378 462986 320614
rect 463222 320378 463306 320614
rect 463542 320378 498986 320614
rect 499222 320378 499306 320614
rect 499542 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect -8726 320294 592650 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 66986 320294
rect 67222 320058 67306 320294
rect 67542 320058 102986 320294
rect 103222 320058 103306 320294
rect 103542 320058 138986 320294
rect 139222 320058 139306 320294
rect 139542 320058 174986 320294
rect 175222 320058 175306 320294
rect 175542 320058 210986 320294
rect 211222 320058 211306 320294
rect 211542 320058 246986 320294
rect 247222 320058 247306 320294
rect 247542 320058 282986 320294
rect 283222 320058 283306 320294
rect 283542 320058 318986 320294
rect 319222 320058 319306 320294
rect 319542 320058 354986 320294
rect 355222 320058 355306 320294
rect 355542 320058 390986 320294
rect 391222 320058 391306 320294
rect 391542 320058 426986 320294
rect 427222 320058 427306 320294
rect 427542 320058 462986 320294
rect 463222 320058 463306 320294
rect 463542 320058 498986 320294
rect 499222 320058 499306 320294
rect 499542 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect -8726 320026 592650 320058
rect -6806 316894 590730 316926
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 63266 316894
rect 63502 316658 63586 316894
rect 63822 316658 99266 316894
rect 99502 316658 99586 316894
rect 99822 316658 135266 316894
rect 135502 316658 135586 316894
rect 135822 316658 171266 316894
rect 171502 316658 171586 316894
rect 171822 316658 207266 316894
rect 207502 316658 207586 316894
rect 207822 316658 243266 316894
rect 243502 316658 243586 316894
rect 243822 316658 279266 316894
rect 279502 316658 279586 316894
rect 279822 316658 315266 316894
rect 315502 316658 315586 316894
rect 315822 316658 351266 316894
rect 351502 316658 351586 316894
rect 351822 316658 387266 316894
rect 387502 316658 387586 316894
rect 387822 316658 423266 316894
rect 423502 316658 423586 316894
rect 423822 316658 459266 316894
rect 459502 316658 459586 316894
rect 459822 316658 495266 316894
rect 495502 316658 495586 316894
rect 495822 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect -6806 316574 590730 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 63266 316574
rect 63502 316338 63586 316574
rect 63822 316338 99266 316574
rect 99502 316338 99586 316574
rect 99822 316338 135266 316574
rect 135502 316338 135586 316574
rect 135822 316338 171266 316574
rect 171502 316338 171586 316574
rect 171822 316338 207266 316574
rect 207502 316338 207586 316574
rect 207822 316338 243266 316574
rect 243502 316338 243586 316574
rect 243822 316338 279266 316574
rect 279502 316338 279586 316574
rect 279822 316338 315266 316574
rect 315502 316338 315586 316574
rect 315822 316338 351266 316574
rect 351502 316338 351586 316574
rect 351822 316338 387266 316574
rect 387502 316338 387586 316574
rect 387822 316338 423266 316574
rect 423502 316338 423586 316574
rect 423822 316338 459266 316574
rect 459502 316338 459586 316574
rect 459822 316338 495266 316574
rect 495502 316338 495586 316574
rect 495822 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect -6806 316306 590730 316338
rect -4886 313174 588810 313206
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 59546 313174
rect 59782 312938 59866 313174
rect 60102 312938 95546 313174
rect 95782 312938 95866 313174
rect 96102 312938 131546 313174
rect 131782 312938 131866 313174
rect 132102 312938 167546 313174
rect 167782 312938 167866 313174
rect 168102 312938 203546 313174
rect 203782 312938 203866 313174
rect 204102 312938 239546 313174
rect 239782 312938 239866 313174
rect 240102 312938 275546 313174
rect 275782 312938 275866 313174
rect 276102 312938 311546 313174
rect 311782 312938 311866 313174
rect 312102 312938 347546 313174
rect 347782 312938 347866 313174
rect 348102 312938 383546 313174
rect 383782 312938 383866 313174
rect 384102 312938 419546 313174
rect 419782 312938 419866 313174
rect 420102 312938 455546 313174
rect 455782 312938 455866 313174
rect 456102 312938 491546 313174
rect 491782 312938 491866 313174
rect 492102 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect -4886 312854 588810 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 59546 312854
rect 59782 312618 59866 312854
rect 60102 312618 95546 312854
rect 95782 312618 95866 312854
rect 96102 312618 131546 312854
rect 131782 312618 131866 312854
rect 132102 312618 167546 312854
rect 167782 312618 167866 312854
rect 168102 312618 203546 312854
rect 203782 312618 203866 312854
rect 204102 312618 239546 312854
rect 239782 312618 239866 312854
rect 240102 312618 275546 312854
rect 275782 312618 275866 312854
rect 276102 312618 311546 312854
rect 311782 312618 311866 312854
rect 312102 312618 347546 312854
rect 347782 312618 347866 312854
rect 348102 312618 383546 312854
rect 383782 312618 383866 312854
rect 384102 312618 419546 312854
rect 419782 312618 419866 312854
rect 420102 312618 455546 312854
rect 455782 312618 455866 312854
rect 456102 312618 491546 312854
rect 491782 312618 491866 312854
rect 492102 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect -4886 312586 588810 312618
rect -2966 309454 586890 309486
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect -2966 309134 586890 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect -2966 308866 586890 308898
rect -8726 302614 592650 302646
rect -8726 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 84986 302614
rect 85222 302378 85306 302614
rect 85542 302378 120986 302614
rect 121222 302378 121306 302614
rect 121542 302378 156986 302614
rect 157222 302378 157306 302614
rect 157542 302378 192986 302614
rect 193222 302378 193306 302614
rect 193542 302378 228986 302614
rect 229222 302378 229306 302614
rect 229542 302378 264986 302614
rect 265222 302378 265306 302614
rect 265542 302378 300986 302614
rect 301222 302378 301306 302614
rect 301542 302378 336986 302614
rect 337222 302378 337306 302614
rect 337542 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 84986 302294
rect 85222 302058 85306 302294
rect 85542 302058 120986 302294
rect 121222 302058 121306 302294
rect 121542 302058 156986 302294
rect 157222 302058 157306 302294
rect 157542 302058 192986 302294
rect 193222 302058 193306 302294
rect 193542 302058 228986 302294
rect 229222 302058 229306 302294
rect 229542 302058 264986 302294
rect 265222 302058 265306 302294
rect 265542 302058 300986 302294
rect 301222 302058 301306 302294
rect 301542 302058 336986 302294
rect 337222 302058 337306 302294
rect 337542 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 592650 302294
rect -8726 302026 592650 302058
rect -6806 298894 590730 298926
rect -6806 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 81266 298894
rect 81502 298658 81586 298894
rect 81822 298658 117266 298894
rect 117502 298658 117586 298894
rect 117822 298658 153266 298894
rect 153502 298658 153586 298894
rect 153822 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 333266 298894
rect 333502 298658 333586 298894
rect 333822 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 590730 298894
rect -6806 298574 590730 298658
rect -6806 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 81266 298574
rect 81502 298338 81586 298574
rect 81822 298338 117266 298574
rect 117502 298338 117586 298574
rect 117822 298338 153266 298574
rect 153502 298338 153586 298574
rect 153822 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 333266 298574
rect 333502 298338 333586 298574
rect 333822 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 590730 298574
rect -6806 298306 590730 298338
rect -4886 295174 588810 295206
rect -4886 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 77546 295174
rect 77782 294938 77866 295174
rect 78102 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 149546 295174
rect 149782 294938 149866 295174
rect 150102 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 329546 295174
rect 329782 294938 329866 295174
rect 330102 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 588810 295174
rect -4886 294854 588810 294938
rect -4886 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 77546 294854
rect 77782 294618 77866 294854
rect 78102 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 149546 294854
rect 149782 294618 149866 294854
rect 150102 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 329546 294854
rect 329782 294618 329866 294854
rect 330102 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 588810 294854
rect -4886 294586 588810 294618
rect -2966 291454 586890 291486
rect -2966 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 204250 291454
rect 204486 291218 234970 291454
rect 235206 291218 265690 291454
rect 265926 291218 296410 291454
rect 296646 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 362285 291454
rect 362521 291218 364882 291454
rect 365118 291218 367479 291454
rect 367715 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 434285 291454
rect 434521 291218 436882 291454
rect 437118 291218 439479 291454
rect 439715 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 586890 291454
rect -2966 291134 586890 291218
rect -2966 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 204250 291134
rect 204486 290898 234970 291134
rect 235206 290898 265690 291134
rect 265926 290898 296410 291134
rect 296646 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 362285 291134
rect 362521 290898 364882 291134
rect 365118 290898 367479 291134
rect 367715 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 434285 291134
rect 434521 290898 436882 291134
rect 437118 290898 439479 291134
rect 439715 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 586890 291134
rect -2966 290866 586890 290898
rect -8726 284614 592650 284646
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 66986 284614
rect 67222 284378 67306 284614
rect 67542 284378 102986 284614
rect 103222 284378 103306 284614
rect 103542 284378 138986 284614
rect 139222 284378 139306 284614
rect 139542 284378 174986 284614
rect 175222 284378 175306 284614
rect 175542 284378 318986 284614
rect 319222 284378 319306 284614
rect 319542 284378 354986 284614
rect 355222 284378 355306 284614
rect 355542 284378 390986 284614
rect 391222 284378 391306 284614
rect 391542 284378 426986 284614
rect 427222 284378 427306 284614
rect 427542 284378 462986 284614
rect 463222 284378 463306 284614
rect 463542 284378 498986 284614
rect 499222 284378 499306 284614
rect 499542 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect -8726 284294 592650 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 66986 284294
rect 67222 284058 67306 284294
rect 67542 284058 102986 284294
rect 103222 284058 103306 284294
rect 103542 284058 138986 284294
rect 139222 284058 139306 284294
rect 139542 284058 174986 284294
rect 175222 284058 175306 284294
rect 175542 284058 318986 284294
rect 319222 284058 319306 284294
rect 319542 284058 354986 284294
rect 355222 284058 355306 284294
rect 355542 284058 390986 284294
rect 391222 284058 391306 284294
rect 391542 284058 426986 284294
rect 427222 284058 427306 284294
rect 427542 284058 462986 284294
rect 463222 284058 463306 284294
rect 463542 284058 498986 284294
rect 499222 284058 499306 284294
rect 499542 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect -8726 284026 592650 284058
rect -6806 280894 590730 280926
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 63266 280894
rect 63502 280658 63586 280894
rect 63822 280658 99266 280894
rect 99502 280658 99586 280894
rect 99822 280658 135266 280894
rect 135502 280658 135586 280894
rect 135822 280658 171266 280894
rect 171502 280658 171586 280894
rect 171822 280658 315266 280894
rect 315502 280658 315586 280894
rect 315822 280658 351266 280894
rect 351502 280658 351586 280894
rect 351822 280658 387266 280894
rect 387502 280658 387586 280894
rect 387822 280658 423266 280894
rect 423502 280658 423586 280894
rect 423822 280658 459266 280894
rect 459502 280658 459586 280894
rect 459822 280658 495266 280894
rect 495502 280658 495586 280894
rect 495822 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect -6806 280574 590730 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 63266 280574
rect 63502 280338 63586 280574
rect 63822 280338 99266 280574
rect 99502 280338 99586 280574
rect 99822 280338 135266 280574
rect 135502 280338 135586 280574
rect 135822 280338 171266 280574
rect 171502 280338 171586 280574
rect 171822 280338 315266 280574
rect 315502 280338 315586 280574
rect 315822 280338 351266 280574
rect 351502 280338 351586 280574
rect 351822 280338 387266 280574
rect 387502 280338 387586 280574
rect 387822 280338 423266 280574
rect 423502 280338 423586 280574
rect 423822 280338 459266 280574
rect 459502 280338 459586 280574
rect 459822 280338 495266 280574
rect 495502 280338 495586 280574
rect 495822 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect -6806 280306 590730 280338
rect -4886 277174 588810 277206
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 59546 277174
rect 59782 276938 59866 277174
rect 60102 276938 95546 277174
rect 95782 276938 95866 277174
rect 96102 276938 131546 277174
rect 131782 276938 131866 277174
rect 132102 276938 167546 277174
rect 167782 276938 167866 277174
rect 168102 276938 311546 277174
rect 311782 276938 311866 277174
rect 312102 276938 347546 277174
rect 347782 276938 347866 277174
rect 348102 276938 383546 277174
rect 383782 276938 383866 277174
rect 384102 276938 419546 277174
rect 419782 276938 419866 277174
rect 420102 276938 455546 277174
rect 455782 276938 455866 277174
rect 456102 276938 491546 277174
rect 491782 276938 491866 277174
rect 492102 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect -4886 276854 588810 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 59546 276854
rect 59782 276618 59866 276854
rect 60102 276618 95546 276854
rect 95782 276618 95866 276854
rect 96102 276618 131546 276854
rect 131782 276618 131866 276854
rect 132102 276618 167546 276854
rect 167782 276618 167866 276854
rect 168102 276618 311546 276854
rect 311782 276618 311866 276854
rect 312102 276618 347546 276854
rect 347782 276618 347866 276854
rect 348102 276618 383546 276854
rect 383782 276618 383866 276854
rect 384102 276618 419546 276854
rect 419782 276618 419866 276854
rect 420102 276618 455546 276854
rect 455782 276618 455866 276854
rect 456102 276618 491546 276854
rect 491782 276618 491866 276854
rect 492102 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect -4886 276586 588810 276618
rect -2966 273454 586890 273486
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 219610 273454
rect 219846 273218 250330 273454
rect 250566 273218 281050 273454
rect 281286 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 363583 273454
rect 363819 273218 366180 273454
rect 366416 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 435583 273454
rect 435819 273218 438180 273454
rect 438416 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect -2966 273134 586890 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 219610 273134
rect 219846 272898 250330 273134
rect 250566 272898 281050 273134
rect 281286 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 363583 273134
rect 363819 272898 366180 273134
rect 366416 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 435583 273134
rect 435819 272898 438180 273134
rect 438416 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect -2966 272866 586890 272898
rect -8726 266614 592650 266646
rect -8726 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 84986 266614
rect 85222 266378 85306 266614
rect 85542 266378 120986 266614
rect 121222 266378 121306 266614
rect 121542 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 192986 266614
rect 193222 266378 193306 266614
rect 193542 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 84986 266294
rect 85222 266058 85306 266294
rect 85542 266058 120986 266294
rect 121222 266058 121306 266294
rect 121542 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 192986 266294
rect 193222 266058 193306 266294
rect 193542 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 592650 266294
rect -8726 266026 592650 266058
rect -6806 262894 590730 262926
rect -6806 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 81266 262894
rect 81502 262658 81586 262894
rect 81822 262658 117266 262894
rect 117502 262658 117586 262894
rect 117822 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 590730 262894
rect -6806 262574 590730 262658
rect -6806 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 81266 262574
rect 81502 262338 81586 262574
rect 81822 262338 117266 262574
rect 117502 262338 117586 262574
rect 117822 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 590730 262574
rect -6806 262306 590730 262338
rect -4886 259174 588810 259206
rect -4886 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 77546 259174
rect 77782 258938 77866 259174
rect 78102 258938 113546 259174
rect 113782 258938 113866 259174
rect 114102 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 588810 259174
rect -4886 258854 588810 258938
rect -4886 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 77546 258854
rect 77782 258618 77866 258854
rect 78102 258618 113546 258854
rect 113782 258618 113866 258854
rect 114102 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 588810 258854
rect -4886 258586 588810 258618
rect -2966 255454 586890 255486
rect -2966 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 204250 255454
rect 204486 255218 234970 255454
rect 235206 255218 265690 255454
rect 265926 255218 296410 255454
rect 296646 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 586890 255454
rect -2966 255134 586890 255218
rect -2966 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 204250 255134
rect 204486 254898 234970 255134
rect 235206 254898 265690 255134
rect 265926 254898 296410 255134
rect 296646 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 586890 255134
rect -2966 254866 586890 254898
rect -8726 248614 592650 248646
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 66986 248614
rect 67222 248378 67306 248614
rect 67542 248378 102986 248614
rect 103222 248378 103306 248614
rect 103542 248378 138986 248614
rect 139222 248378 139306 248614
rect 139542 248378 174986 248614
rect 175222 248378 175306 248614
rect 175542 248378 318986 248614
rect 319222 248378 319306 248614
rect 319542 248378 354986 248614
rect 355222 248378 355306 248614
rect 355542 248378 390986 248614
rect 391222 248378 391306 248614
rect 391542 248378 426986 248614
rect 427222 248378 427306 248614
rect 427542 248378 462986 248614
rect 463222 248378 463306 248614
rect 463542 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect -8726 248294 592650 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 66986 248294
rect 67222 248058 67306 248294
rect 67542 248058 102986 248294
rect 103222 248058 103306 248294
rect 103542 248058 138986 248294
rect 139222 248058 139306 248294
rect 139542 248058 174986 248294
rect 175222 248058 175306 248294
rect 175542 248058 318986 248294
rect 319222 248058 319306 248294
rect 319542 248058 354986 248294
rect 355222 248058 355306 248294
rect 355542 248058 390986 248294
rect 391222 248058 391306 248294
rect 391542 248058 426986 248294
rect 427222 248058 427306 248294
rect 427542 248058 462986 248294
rect 463222 248058 463306 248294
rect 463542 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect -8726 248026 592650 248058
rect -6806 244894 590730 244926
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 99266 244894
rect 99502 244658 99586 244894
rect 99822 244658 135266 244894
rect 135502 244658 135586 244894
rect 135822 244658 171266 244894
rect 171502 244658 171586 244894
rect 171822 244658 315266 244894
rect 315502 244658 315586 244894
rect 315822 244658 351266 244894
rect 351502 244658 351586 244894
rect 351822 244658 387266 244894
rect 387502 244658 387586 244894
rect 387822 244658 423266 244894
rect 423502 244658 423586 244894
rect 423822 244658 459266 244894
rect 459502 244658 459586 244894
rect 459822 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect -6806 244574 590730 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 99266 244574
rect 99502 244338 99586 244574
rect 99822 244338 135266 244574
rect 135502 244338 135586 244574
rect 135822 244338 171266 244574
rect 171502 244338 171586 244574
rect 171822 244338 315266 244574
rect 315502 244338 315586 244574
rect 315822 244338 351266 244574
rect 351502 244338 351586 244574
rect 351822 244338 387266 244574
rect 387502 244338 387586 244574
rect 387822 244338 423266 244574
rect 423502 244338 423586 244574
rect 423822 244338 459266 244574
rect 459502 244338 459586 244574
rect 459822 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect -6806 244306 590730 244338
rect -4886 241174 588810 241206
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 95546 241174
rect 95782 240938 95866 241174
rect 96102 240938 131546 241174
rect 131782 240938 131866 241174
rect 132102 240938 167546 241174
rect 167782 240938 167866 241174
rect 168102 240938 311546 241174
rect 311782 240938 311866 241174
rect 312102 240938 347546 241174
rect 347782 240938 347866 241174
rect 348102 240938 383546 241174
rect 383782 240938 383866 241174
rect 384102 240938 419546 241174
rect 419782 240938 419866 241174
rect 420102 240938 455546 241174
rect 455782 240938 455866 241174
rect 456102 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect -4886 240854 588810 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 95546 240854
rect 95782 240618 95866 240854
rect 96102 240618 131546 240854
rect 131782 240618 131866 240854
rect 132102 240618 167546 240854
rect 167782 240618 167866 240854
rect 168102 240618 311546 240854
rect 311782 240618 311866 240854
rect 312102 240618 347546 240854
rect 347782 240618 347866 240854
rect 348102 240618 383546 240854
rect 383782 240618 383866 240854
rect 384102 240618 419546 240854
rect 419782 240618 419866 240854
rect 420102 240618 455546 240854
rect 455782 240618 455866 240854
rect 456102 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect -4886 240586 588810 240618
rect -2966 237454 586890 237486
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 219610 237454
rect 219846 237218 250330 237454
rect 250566 237218 281050 237454
rect 281286 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect -2966 237134 586890 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 219610 237134
rect 219846 236898 250330 237134
rect 250566 236898 281050 237134
rect 281286 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect -2966 236866 586890 236898
rect -8726 230614 592650 230646
rect -8726 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 156986 230614
rect 157222 230378 157306 230614
rect 157542 230378 192986 230614
rect 193222 230378 193306 230614
rect 193542 230378 336986 230614
rect 337222 230378 337306 230614
rect 337542 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 156986 230294
rect 157222 230058 157306 230294
rect 157542 230058 192986 230294
rect 193222 230058 193306 230294
rect 193542 230058 336986 230294
rect 337222 230058 337306 230294
rect 337542 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 592650 230294
rect -8726 230026 592650 230058
rect -6806 226894 590730 226926
rect -6806 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 81266 226894
rect 81502 226658 81586 226894
rect 81822 226658 117266 226894
rect 117502 226658 117586 226894
rect 117822 226658 153266 226894
rect 153502 226658 153586 226894
rect 153822 226658 189266 226894
rect 189502 226658 189586 226894
rect 189822 226658 333266 226894
rect 333502 226658 333586 226894
rect 333822 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 590730 226894
rect -6806 226574 590730 226658
rect -6806 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 81266 226574
rect 81502 226338 81586 226574
rect 81822 226338 117266 226574
rect 117502 226338 117586 226574
rect 117822 226338 153266 226574
rect 153502 226338 153586 226574
rect 153822 226338 189266 226574
rect 189502 226338 189586 226574
rect 189822 226338 333266 226574
rect 333502 226338 333586 226574
rect 333822 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 590730 226574
rect -6806 226306 590730 226338
rect -4886 223174 588810 223206
rect -4886 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 113546 223174
rect 113782 222938 113866 223174
rect 114102 222938 149546 223174
rect 149782 222938 149866 223174
rect 150102 222938 185546 223174
rect 185782 222938 185866 223174
rect 186102 222938 329546 223174
rect 329782 222938 329866 223174
rect 330102 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 588810 223174
rect -4886 222854 588810 222938
rect -4886 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 113546 222854
rect 113782 222618 113866 222854
rect 114102 222618 149546 222854
rect 149782 222618 149866 222854
rect 150102 222618 185546 222854
rect 185782 222618 185866 222854
rect 186102 222618 329546 222854
rect 329782 222618 329866 222854
rect 330102 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 588810 222854
rect -4886 222586 588810 222618
rect -2966 219454 586890 219486
rect -2966 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 204250 219454
rect 204486 219218 234970 219454
rect 235206 219218 265690 219454
rect 265926 219218 296410 219454
rect 296646 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 362285 219454
rect 362521 219218 364882 219454
rect 365118 219218 367479 219454
rect 367715 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 434285 219454
rect 434521 219218 436882 219454
rect 437118 219218 439479 219454
rect 439715 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 586890 219454
rect -2966 219134 586890 219218
rect -2966 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 204250 219134
rect 204486 218898 234970 219134
rect 235206 218898 265690 219134
rect 265926 218898 296410 219134
rect 296646 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 362285 219134
rect 362521 218898 364882 219134
rect 365118 218898 367479 219134
rect 367715 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 434285 219134
rect 434521 218898 436882 219134
rect 437118 218898 439479 219134
rect 439715 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 586890 219134
rect -2966 218866 586890 218898
rect -8726 212614 592650 212646
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 66986 212614
rect 67222 212378 67306 212614
rect 67542 212378 102986 212614
rect 103222 212378 103306 212614
rect 103542 212378 138986 212614
rect 139222 212378 139306 212614
rect 139542 212378 174986 212614
rect 175222 212378 175306 212614
rect 175542 212378 318986 212614
rect 319222 212378 319306 212614
rect 319542 212378 354986 212614
rect 355222 212378 355306 212614
rect 355542 212378 390986 212614
rect 391222 212378 391306 212614
rect 391542 212378 426986 212614
rect 427222 212378 427306 212614
rect 427542 212378 462986 212614
rect 463222 212378 463306 212614
rect 463542 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect -8726 212294 592650 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 66986 212294
rect 67222 212058 67306 212294
rect 67542 212058 102986 212294
rect 103222 212058 103306 212294
rect 103542 212058 138986 212294
rect 139222 212058 139306 212294
rect 139542 212058 174986 212294
rect 175222 212058 175306 212294
rect 175542 212058 318986 212294
rect 319222 212058 319306 212294
rect 319542 212058 354986 212294
rect 355222 212058 355306 212294
rect 355542 212058 390986 212294
rect 391222 212058 391306 212294
rect 391542 212058 426986 212294
rect 427222 212058 427306 212294
rect 427542 212058 462986 212294
rect 463222 212058 463306 212294
rect 463542 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect -8726 212026 592650 212058
rect -6806 208894 590730 208926
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 63266 208894
rect 63502 208658 63586 208894
rect 63822 208658 99266 208894
rect 99502 208658 99586 208894
rect 99822 208658 135266 208894
rect 135502 208658 135586 208894
rect 135822 208658 171266 208894
rect 171502 208658 171586 208894
rect 171822 208658 315266 208894
rect 315502 208658 315586 208894
rect 315822 208658 351266 208894
rect 351502 208658 351586 208894
rect 351822 208658 387266 208894
rect 387502 208658 387586 208894
rect 387822 208658 423266 208894
rect 423502 208658 423586 208894
rect 423822 208658 459266 208894
rect 459502 208658 459586 208894
rect 459822 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect -6806 208574 590730 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 63266 208574
rect 63502 208338 63586 208574
rect 63822 208338 99266 208574
rect 99502 208338 99586 208574
rect 99822 208338 135266 208574
rect 135502 208338 135586 208574
rect 135822 208338 171266 208574
rect 171502 208338 171586 208574
rect 171822 208338 315266 208574
rect 315502 208338 315586 208574
rect 315822 208338 351266 208574
rect 351502 208338 351586 208574
rect 351822 208338 387266 208574
rect 387502 208338 387586 208574
rect 387822 208338 423266 208574
rect 423502 208338 423586 208574
rect 423822 208338 459266 208574
rect 459502 208338 459586 208574
rect 459822 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect -6806 208306 590730 208338
rect -4886 205174 588810 205206
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 59546 205174
rect 59782 204938 59866 205174
rect 60102 204938 95546 205174
rect 95782 204938 95866 205174
rect 96102 204938 131546 205174
rect 131782 204938 131866 205174
rect 132102 204938 167546 205174
rect 167782 204938 167866 205174
rect 168102 204938 311546 205174
rect 311782 204938 311866 205174
rect 312102 204938 347546 205174
rect 347782 204938 347866 205174
rect 348102 204938 383546 205174
rect 383782 204938 383866 205174
rect 384102 204938 419546 205174
rect 419782 204938 419866 205174
rect 420102 204938 455546 205174
rect 455782 204938 455866 205174
rect 456102 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect -4886 204854 588810 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 59546 204854
rect 59782 204618 59866 204854
rect 60102 204618 95546 204854
rect 95782 204618 95866 204854
rect 96102 204618 131546 204854
rect 131782 204618 131866 204854
rect 132102 204618 167546 204854
rect 167782 204618 167866 204854
rect 168102 204618 311546 204854
rect 311782 204618 311866 204854
rect 312102 204618 347546 204854
rect 347782 204618 347866 204854
rect 348102 204618 383546 204854
rect 383782 204618 383866 204854
rect 384102 204618 419546 204854
rect 419782 204618 419866 204854
rect 420102 204618 455546 204854
rect 455782 204618 455866 204854
rect 456102 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect -4886 204586 588810 204618
rect -2966 201454 586890 201486
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 219610 201454
rect 219846 201218 250330 201454
rect 250566 201218 281050 201454
rect 281286 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 363583 201454
rect 363819 201218 366180 201454
rect 366416 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 435583 201454
rect 435819 201218 438180 201454
rect 438416 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect -2966 201134 586890 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 219610 201134
rect 219846 200898 250330 201134
rect 250566 200898 281050 201134
rect 281286 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 363583 201134
rect 363819 200898 366180 201134
rect 366416 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 435583 201134
rect 435819 200898 438180 201134
rect 438416 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect -2966 200866 586890 200898
rect -8726 194614 592650 194646
rect -8726 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 120986 194614
rect 121222 194378 121306 194614
rect 121542 194378 156986 194614
rect 157222 194378 157306 194614
rect 157542 194378 192986 194614
rect 193222 194378 193306 194614
rect 193542 194378 336986 194614
rect 337222 194378 337306 194614
rect 337542 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 120986 194294
rect 121222 194058 121306 194294
rect 121542 194058 156986 194294
rect 157222 194058 157306 194294
rect 157542 194058 192986 194294
rect 193222 194058 193306 194294
rect 193542 194058 336986 194294
rect 337222 194058 337306 194294
rect 337542 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 592650 194294
rect -8726 194026 592650 194058
rect -6806 190894 590730 190926
rect -6806 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 117266 190894
rect 117502 190658 117586 190894
rect 117822 190658 153266 190894
rect 153502 190658 153586 190894
rect 153822 190658 189266 190894
rect 189502 190658 189586 190894
rect 189822 190658 333266 190894
rect 333502 190658 333586 190894
rect 333822 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 590730 190894
rect -6806 190574 590730 190658
rect -6806 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 117266 190574
rect 117502 190338 117586 190574
rect 117822 190338 153266 190574
rect 153502 190338 153586 190574
rect 153822 190338 189266 190574
rect 189502 190338 189586 190574
rect 189822 190338 333266 190574
rect 333502 190338 333586 190574
rect 333822 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 590730 190574
rect -6806 190306 590730 190338
rect -4886 187174 588810 187206
rect -4886 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 149546 187174
rect 149782 186938 149866 187174
rect 150102 186938 185546 187174
rect 185782 186938 185866 187174
rect 186102 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 588810 187174
rect -4886 186854 588810 186938
rect -4886 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 149546 186854
rect 149782 186618 149866 186854
rect 150102 186618 185546 186854
rect 185782 186618 185866 186854
rect 186102 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 588810 186854
rect -4886 186586 588810 186618
rect -2966 183454 586890 183486
rect -2966 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 162285 183454
rect 162521 183218 164882 183454
rect 165118 183218 167479 183454
rect 167715 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 204250 183454
rect 204486 183218 234970 183454
rect 235206 183218 265690 183454
rect 265926 183218 296410 183454
rect 296646 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 586890 183454
rect -2966 183134 586890 183218
rect -2966 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 162285 183134
rect 162521 182898 164882 183134
rect 165118 182898 167479 183134
rect 167715 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 204250 183134
rect 204486 182898 234970 183134
rect 235206 182898 265690 183134
rect 265926 182898 296410 183134
rect 296646 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 586890 183134
rect -2966 182866 586890 182898
rect -8726 176614 592650 176646
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 66986 176614
rect 67222 176378 67306 176614
rect 67542 176378 102986 176614
rect 103222 176378 103306 176614
rect 103542 176378 138986 176614
rect 139222 176378 139306 176614
rect 139542 176378 174986 176614
rect 175222 176378 175306 176614
rect 175542 176378 318986 176614
rect 319222 176378 319306 176614
rect 319542 176378 354986 176614
rect 355222 176378 355306 176614
rect 355542 176378 390986 176614
rect 391222 176378 391306 176614
rect 391542 176378 426986 176614
rect 427222 176378 427306 176614
rect 427542 176378 462986 176614
rect 463222 176378 463306 176614
rect 463542 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect -8726 176294 592650 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 66986 176294
rect 67222 176058 67306 176294
rect 67542 176058 102986 176294
rect 103222 176058 103306 176294
rect 103542 176058 138986 176294
rect 139222 176058 139306 176294
rect 139542 176058 174986 176294
rect 175222 176058 175306 176294
rect 175542 176058 318986 176294
rect 319222 176058 319306 176294
rect 319542 176058 354986 176294
rect 355222 176058 355306 176294
rect 355542 176058 390986 176294
rect 391222 176058 391306 176294
rect 391542 176058 426986 176294
rect 427222 176058 427306 176294
rect 427542 176058 462986 176294
rect 463222 176058 463306 176294
rect 463542 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect -8726 176026 592650 176058
rect -6806 172894 590730 172926
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 63266 172894
rect 63502 172658 63586 172894
rect 63822 172658 99266 172894
rect 99502 172658 99586 172894
rect 99822 172658 135266 172894
rect 135502 172658 135586 172894
rect 135822 172658 315266 172894
rect 315502 172658 315586 172894
rect 315822 172658 351266 172894
rect 351502 172658 351586 172894
rect 351822 172658 387266 172894
rect 387502 172658 387586 172894
rect 387822 172658 423266 172894
rect 423502 172658 423586 172894
rect 423822 172658 459266 172894
rect 459502 172658 459586 172894
rect 459822 172658 495266 172894
rect 495502 172658 495586 172894
rect 495822 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect -6806 172574 590730 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 63266 172574
rect 63502 172338 63586 172574
rect 63822 172338 99266 172574
rect 99502 172338 99586 172574
rect 99822 172338 135266 172574
rect 135502 172338 135586 172574
rect 135822 172338 315266 172574
rect 315502 172338 315586 172574
rect 315822 172338 351266 172574
rect 351502 172338 351586 172574
rect 351822 172338 387266 172574
rect 387502 172338 387586 172574
rect 387822 172338 423266 172574
rect 423502 172338 423586 172574
rect 423822 172338 459266 172574
rect 459502 172338 459586 172574
rect 459822 172338 495266 172574
rect 495502 172338 495586 172574
rect 495822 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect -6806 172306 590730 172338
rect -4886 169174 588810 169206
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 59546 169174
rect 59782 168938 59866 169174
rect 60102 168938 95546 169174
rect 95782 168938 95866 169174
rect 96102 168938 131546 169174
rect 131782 168938 131866 169174
rect 132102 168938 311546 169174
rect 311782 168938 311866 169174
rect 312102 168938 347546 169174
rect 347782 168938 347866 169174
rect 348102 168938 383546 169174
rect 383782 168938 383866 169174
rect 384102 168938 419546 169174
rect 419782 168938 419866 169174
rect 420102 168938 455546 169174
rect 455782 168938 455866 169174
rect 456102 168938 491546 169174
rect 491782 168938 491866 169174
rect 492102 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect -4886 168854 588810 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 59546 168854
rect 59782 168618 59866 168854
rect 60102 168618 95546 168854
rect 95782 168618 95866 168854
rect 96102 168618 131546 168854
rect 131782 168618 131866 168854
rect 132102 168618 311546 168854
rect 311782 168618 311866 168854
rect 312102 168618 347546 168854
rect 347782 168618 347866 168854
rect 348102 168618 383546 168854
rect 383782 168618 383866 168854
rect 384102 168618 419546 168854
rect 419782 168618 419866 168854
rect 420102 168618 455546 168854
rect 455782 168618 455866 168854
rect 456102 168618 491546 168854
rect 491782 168618 491866 168854
rect 492102 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect -4886 168586 588810 168618
rect -2966 165454 586890 165486
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 163583 165454
rect 163819 165218 166180 165454
rect 166416 165218 219610 165454
rect 219846 165218 250330 165454
rect 250566 165218 281050 165454
rect 281286 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect -2966 165134 586890 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 163583 165134
rect 163819 164898 166180 165134
rect 166416 164898 219610 165134
rect 219846 164898 250330 165134
rect 250566 164898 281050 165134
rect 281286 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect -2966 164866 586890 164898
rect -8726 158614 592650 158646
rect -8726 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 84986 158614
rect 85222 158378 85306 158614
rect 85542 158378 120986 158614
rect 121222 158378 121306 158614
rect 121542 158378 156986 158614
rect 157222 158378 157306 158614
rect 157542 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 84986 158294
rect 85222 158058 85306 158294
rect 85542 158058 120986 158294
rect 121222 158058 121306 158294
rect 121542 158058 156986 158294
rect 157222 158058 157306 158294
rect 157542 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 592650 158294
rect -8726 158026 592650 158058
rect -6806 154894 590730 154926
rect -6806 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 81266 154894
rect 81502 154658 81586 154894
rect 81822 154658 117266 154894
rect 117502 154658 117586 154894
rect 117822 154658 153266 154894
rect 153502 154658 153586 154894
rect 153822 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 590730 154894
rect -6806 154574 590730 154658
rect -6806 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 81266 154574
rect 81502 154338 81586 154574
rect 81822 154338 117266 154574
rect 117502 154338 117586 154574
rect 117822 154338 153266 154574
rect 153502 154338 153586 154574
rect 153822 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 590730 154574
rect -6806 154306 590730 154338
rect -4886 151174 588810 151206
rect -4886 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 77546 151174
rect 77782 150938 77866 151174
rect 78102 150938 113546 151174
rect 113782 150938 113866 151174
rect 114102 150938 149546 151174
rect 149782 150938 149866 151174
rect 150102 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 588810 151174
rect -4886 150854 588810 150938
rect -4886 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 77546 150854
rect 77782 150618 77866 150854
rect 78102 150618 113546 150854
rect 113782 150618 113866 150854
rect 114102 150618 149546 150854
rect 149782 150618 149866 150854
rect 150102 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 588810 150854
rect -4886 150586 588810 150618
rect -2966 147454 586890 147486
rect -2966 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 162285 147454
rect 162521 147218 164882 147454
rect 165118 147218 167479 147454
rect 167715 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 204250 147454
rect 204486 147218 234970 147454
rect 235206 147218 265690 147454
rect 265926 147218 296410 147454
rect 296646 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 362285 147454
rect 362521 147218 364882 147454
rect 365118 147218 367479 147454
rect 367715 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 434285 147454
rect 434521 147218 436882 147454
rect 437118 147218 439479 147454
rect 439715 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 586890 147454
rect -2966 147134 586890 147218
rect -2966 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 162285 147134
rect 162521 146898 164882 147134
rect 165118 146898 167479 147134
rect 167715 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 204250 147134
rect 204486 146898 234970 147134
rect 235206 146898 265690 147134
rect 265926 146898 296410 147134
rect 296646 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 362285 147134
rect 362521 146898 364882 147134
rect 365118 146898 367479 147134
rect 367715 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 434285 147134
rect 434521 146898 436882 147134
rect 437118 146898 439479 147134
rect 439715 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 586890 147134
rect -2966 146866 586890 146898
rect -8726 140614 592650 140646
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 66986 140614
rect 67222 140378 67306 140614
rect 67542 140378 102986 140614
rect 103222 140378 103306 140614
rect 103542 140378 138986 140614
rect 139222 140378 139306 140614
rect 139542 140378 174986 140614
rect 175222 140378 175306 140614
rect 175542 140378 318986 140614
rect 319222 140378 319306 140614
rect 319542 140378 354986 140614
rect 355222 140378 355306 140614
rect 355542 140378 390986 140614
rect 391222 140378 391306 140614
rect 391542 140378 426986 140614
rect 427222 140378 427306 140614
rect 427542 140378 462986 140614
rect 463222 140378 463306 140614
rect 463542 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect -8726 140294 592650 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 66986 140294
rect 67222 140058 67306 140294
rect 67542 140058 102986 140294
rect 103222 140058 103306 140294
rect 103542 140058 138986 140294
rect 139222 140058 139306 140294
rect 139542 140058 174986 140294
rect 175222 140058 175306 140294
rect 175542 140058 318986 140294
rect 319222 140058 319306 140294
rect 319542 140058 354986 140294
rect 355222 140058 355306 140294
rect 355542 140058 390986 140294
rect 391222 140058 391306 140294
rect 391542 140058 426986 140294
rect 427222 140058 427306 140294
rect 427542 140058 462986 140294
rect 463222 140058 463306 140294
rect 463542 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect -8726 140026 592650 140058
rect -6806 136894 590730 136926
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 63266 136894
rect 63502 136658 63586 136894
rect 63822 136658 99266 136894
rect 99502 136658 99586 136894
rect 99822 136658 135266 136894
rect 135502 136658 135586 136894
rect 135822 136658 315266 136894
rect 315502 136658 315586 136894
rect 315822 136658 351266 136894
rect 351502 136658 351586 136894
rect 351822 136658 387266 136894
rect 387502 136658 387586 136894
rect 387822 136658 423266 136894
rect 423502 136658 423586 136894
rect 423822 136658 459266 136894
rect 459502 136658 459586 136894
rect 459822 136658 495266 136894
rect 495502 136658 495586 136894
rect 495822 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect -6806 136574 590730 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 63266 136574
rect 63502 136338 63586 136574
rect 63822 136338 99266 136574
rect 99502 136338 99586 136574
rect 99822 136338 135266 136574
rect 135502 136338 135586 136574
rect 135822 136338 315266 136574
rect 315502 136338 315586 136574
rect 315822 136338 351266 136574
rect 351502 136338 351586 136574
rect 351822 136338 387266 136574
rect 387502 136338 387586 136574
rect 387822 136338 423266 136574
rect 423502 136338 423586 136574
rect 423822 136338 459266 136574
rect 459502 136338 459586 136574
rect 459822 136338 495266 136574
rect 495502 136338 495586 136574
rect 495822 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect -6806 136306 590730 136338
rect -4886 133174 588810 133206
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 59546 133174
rect 59782 132938 59866 133174
rect 60102 132938 95546 133174
rect 95782 132938 95866 133174
rect 96102 132938 131546 133174
rect 131782 132938 131866 133174
rect 132102 132938 311546 133174
rect 311782 132938 311866 133174
rect 312102 132938 347546 133174
rect 347782 132938 347866 133174
rect 348102 132938 383546 133174
rect 383782 132938 383866 133174
rect 384102 132938 419546 133174
rect 419782 132938 419866 133174
rect 420102 132938 455546 133174
rect 455782 132938 455866 133174
rect 456102 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect -4886 132854 588810 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 59546 132854
rect 59782 132618 59866 132854
rect 60102 132618 95546 132854
rect 95782 132618 95866 132854
rect 96102 132618 131546 132854
rect 131782 132618 131866 132854
rect 132102 132618 311546 132854
rect 311782 132618 311866 132854
rect 312102 132618 347546 132854
rect 347782 132618 347866 132854
rect 348102 132618 383546 132854
rect 383782 132618 383866 132854
rect 384102 132618 419546 132854
rect 419782 132618 419866 132854
rect 420102 132618 455546 132854
rect 455782 132618 455866 132854
rect 456102 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect -4886 132586 588810 132618
rect -2966 129454 586890 129486
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 127826 129454
rect 128062 129218 128146 129454
rect 128382 129218 163583 129454
rect 163819 129218 166180 129454
rect 166416 129218 219610 129454
rect 219846 129218 250330 129454
rect 250566 129218 281050 129454
rect 281286 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 363583 129454
rect 363819 129218 366180 129454
rect 366416 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 435583 129454
rect 435819 129218 438180 129454
rect 438416 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect -2966 129134 586890 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 127826 129134
rect 128062 128898 128146 129134
rect 128382 128898 163583 129134
rect 163819 128898 166180 129134
rect 166416 128898 219610 129134
rect 219846 128898 250330 129134
rect 250566 128898 281050 129134
rect 281286 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 363583 129134
rect 363819 128898 366180 129134
rect 366416 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 435583 129134
rect 435819 128898 438180 129134
rect 438416 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect -2966 128866 586890 128898
rect -8726 122614 592650 122646
rect -8726 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 84986 122614
rect 85222 122378 85306 122614
rect 85542 122378 120986 122614
rect 121222 122378 121306 122614
rect 121542 122378 156986 122614
rect 157222 122378 157306 122614
rect 157542 122378 192986 122614
rect 193222 122378 193306 122614
rect 193542 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 84986 122294
rect 85222 122058 85306 122294
rect 85542 122058 120986 122294
rect 121222 122058 121306 122294
rect 121542 122058 156986 122294
rect 157222 122058 157306 122294
rect 157542 122058 192986 122294
rect 193222 122058 193306 122294
rect 193542 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 592650 122294
rect -8726 122026 592650 122058
rect -6806 118894 590730 118926
rect -6806 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 81266 118894
rect 81502 118658 81586 118894
rect 81822 118658 117266 118894
rect 117502 118658 117586 118894
rect 117822 118658 153266 118894
rect 153502 118658 153586 118894
rect 153822 118658 189266 118894
rect 189502 118658 189586 118894
rect 189822 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 590730 118894
rect -6806 118574 590730 118658
rect -6806 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 81266 118574
rect 81502 118338 81586 118574
rect 81822 118338 117266 118574
rect 117502 118338 117586 118574
rect 117822 118338 153266 118574
rect 153502 118338 153586 118574
rect 153822 118338 189266 118574
rect 189502 118338 189586 118574
rect 189822 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 590730 118574
rect -6806 118306 590730 118338
rect -4886 115174 588810 115206
rect -4886 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 77546 115174
rect 77782 114938 77866 115174
rect 78102 114938 113546 115174
rect 113782 114938 113866 115174
rect 114102 114938 149546 115174
rect 149782 114938 149866 115174
rect 150102 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 588810 115174
rect -4886 114854 588810 114938
rect -4886 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 77546 114854
rect 77782 114618 77866 114854
rect 78102 114618 113546 114854
rect 113782 114618 113866 114854
rect 114102 114618 149546 114854
rect 149782 114618 149866 114854
rect 150102 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 588810 114854
rect -4886 114586 588810 114618
rect -2966 111454 586890 111486
rect -2966 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 204250 111454
rect 204486 111218 234970 111454
rect 235206 111218 265690 111454
rect 265926 111218 296410 111454
rect 296646 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 586890 111454
rect -2966 111134 586890 111218
rect -2966 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 204250 111134
rect 204486 110898 234970 111134
rect 235206 110898 265690 111134
rect 265926 110898 296410 111134
rect 296646 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 586890 111134
rect -2966 110866 586890 110898
rect -8726 104614 592650 104646
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 66986 104614
rect 67222 104378 67306 104614
rect 67542 104378 102986 104614
rect 103222 104378 103306 104614
rect 103542 104378 138986 104614
rect 139222 104378 139306 104614
rect 139542 104378 174986 104614
rect 175222 104378 175306 104614
rect 175542 104378 318986 104614
rect 319222 104378 319306 104614
rect 319542 104378 354986 104614
rect 355222 104378 355306 104614
rect 355542 104378 390986 104614
rect 391222 104378 391306 104614
rect 391542 104378 426986 104614
rect 427222 104378 427306 104614
rect 427542 104378 462986 104614
rect 463222 104378 463306 104614
rect 463542 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect -8726 104294 592650 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 66986 104294
rect 67222 104058 67306 104294
rect 67542 104058 102986 104294
rect 103222 104058 103306 104294
rect 103542 104058 138986 104294
rect 139222 104058 139306 104294
rect 139542 104058 174986 104294
rect 175222 104058 175306 104294
rect 175542 104058 318986 104294
rect 319222 104058 319306 104294
rect 319542 104058 354986 104294
rect 355222 104058 355306 104294
rect 355542 104058 390986 104294
rect 391222 104058 391306 104294
rect 391542 104058 426986 104294
rect 427222 104058 427306 104294
rect 427542 104058 462986 104294
rect 463222 104058 463306 104294
rect 463542 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect -8726 104026 592650 104058
rect -6806 100894 590730 100926
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 63266 100894
rect 63502 100658 63586 100894
rect 63822 100658 99266 100894
rect 99502 100658 99586 100894
rect 99822 100658 135266 100894
rect 135502 100658 135586 100894
rect 135822 100658 171266 100894
rect 171502 100658 171586 100894
rect 171822 100658 315266 100894
rect 315502 100658 315586 100894
rect 315822 100658 351266 100894
rect 351502 100658 351586 100894
rect 351822 100658 387266 100894
rect 387502 100658 387586 100894
rect 387822 100658 423266 100894
rect 423502 100658 423586 100894
rect 423822 100658 459266 100894
rect 459502 100658 459586 100894
rect 459822 100658 495266 100894
rect 495502 100658 495586 100894
rect 495822 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect -6806 100574 590730 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 63266 100574
rect 63502 100338 63586 100574
rect 63822 100338 99266 100574
rect 99502 100338 99586 100574
rect 99822 100338 135266 100574
rect 135502 100338 135586 100574
rect 135822 100338 171266 100574
rect 171502 100338 171586 100574
rect 171822 100338 315266 100574
rect 315502 100338 315586 100574
rect 315822 100338 351266 100574
rect 351502 100338 351586 100574
rect 351822 100338 387266 100574
rect 387502 100338 387586 100574
rect 387822 100338 423266 100574
rect 423502 100338 423586 100574
rect 423822 100338 459266 100574
rect 459502 100338 459586 100574
rect 459822 100338 495266 100574
rect 495502 100338 495586 100574
rect 495822 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect -6806 100306 590730 100338
rect -4886 97174 588810 97206
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 59546 97174
rect 59782 96938 59866 97174
rect 60102 96938 95546 97174
rect 95782 96938 95866 97174
rect 96102 96938 131546 97174
rect 131782 96938 131866 97174
rect 132102 96938 167546 97174
rect 167782 96938 167866 97174
rect 168102 96938 203546 97174
rect 203782 96938 203866 97174
rect 204102 96938 239546 97174
rect 239782 96938 239866 97174
rect 240102 96938 275546 97174
rect 275782 96938 275866 97174
rect 276102 96938 311546 97174
rect 311782 96938 311866 97174
rect 312102 96938 347546 97174
rect 347782 96938 347866 97174
rect 348102 96938 383546 97174
rect 383782 96938 383866 97174
rect 384102 96938 419546 97174
rect 419782 96938 419866 97174
rect 420102 96938 455546 97174
rect 455782 96938 455866 97174
rect 456102 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect -4886 96854 588810 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 59546 96854
rect 59782 96618 59866 96854
rect 60102 96618 95546 96854
rect 95782 96618 95866 96854
rect 96102 96618 131546 96854
rect 131782 96618 131866 96854
rect 132102 96618 167546 96854
rect 167782 96618 167866 96854
rect 168102 96618 203546 96854
rect 203782 96618 203866 96854
rect 204102 96618 239546 96854
rect 239782 96618 239866 96854
rect 240102 96618 275546 96854
rect 275782 96618 275866 96854
rect 276102 96618 311546 96854
rect 311782 96618 311866 96854
rect 312102 96618 347546 96854
rect 347782 96618 347866 96854
rect 348102 96618 383546 96854
rect 383782 96618 383866 96854
rect 384102 96618 419546 96854
rect 419782 96618 419866 96854
rect 420102 96618 455546 96854
rect 455782 96618 455866 96854
rect 456102 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect -4886 96586 588810 96618
rect -2966 93454 586890 93486
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 127826 93454
rect 128062 93218 128146 93454
rect 128382 93218 163826 93454
rect 164062 93218 164146 93454
rect 164382 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect -2966 93134 586890 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 127826 93134
rect 128062 92898 128146 93134
rect 128382 92898 163826 93134
rect 164062 92898 164146 93134
rect 164382 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect -2966 92866 586890 92898
rect -8726 86614 592650 86646
rect -8726 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 120986 86614
rect 121222 86378 121306 86614
rect 121542 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 192986 86614
rect 193222 86378 193306 86614
rect 193542 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 120986 86294
rect 121222 86058 121306 86294
rect 121542 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 192986 86294
rect 193222 86058 193306 86294
rect 193542 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 592650 86294
rect -8726 86026 592650 86058
rect -6806 82894 590730 82926
rect -6806 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 117266 82894
rect 117502 82658 117586 82894
rect 117822 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 189266 82894
rect 189502 82658 189586 82894
rect 189822 82658 225266 82894
rect 225502 82658 225586 82894
rect 225822 82658 261266 82894
rect 261502 82658 261586 82894
rect 261822 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 590730 82894
rect -6806 82574 590730 82658
rect -6806 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 117266 82574
rect 117502 82338 117586 82574
rect 117822 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 189266 82574
rect 189502 82338 189586 82574
rect 189822 82338 225266 82574
rect 225502 82338 225586 82574
rect 225822 82338 261266 82574
rect 261502 82338 261586 82574
rect 261822 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 590730 82574
rect -6806 82306 590730 82338
rect -4886 79174 588810 79206
rect -4886 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 588810 79174
rect -4886 78854 588810 78938
rect -4886 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 588810 78854
rect -4886 78586 588810 78618
rect -2966 75454 586890 75486
rect -2966 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 586890 75454
rect -2966 75134 586890 75218
rect -2966 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 586890 75134
rect -2966 74866 586890 74898
rect -8726 68614 592650 68646
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 66986 68614
rect 67222 68378 67306 68614
rect 67542 68378 102986 68614
rect 103222 68378 103306 68614
rect 103542 68378 138986 68614
rect 139222 68378 139306 68614
rect 139542 68378 174986 68614
rect 175222 68378 175306 68614
rect 175542 68378 210986 68614
rect 211222 68378 211306 68614
rect 211542 68378 246986 68614
rect 247222 68378 247306 68614
rect 247542 68378 282986 68614
rect 283222 68378 283306 68614
rect 283542 68378 318986 68614
rect 319222 68378 319306 68614
rect 319542 68378 354986 68614
rect 355222 68378 355306 68614
rect 355542 68378 390986 68614
rect 391222 68378 391306 68614
rect 391542 68378 426986 68614
rect 427222 68378 427306 68614
rect 427542 68378 462986 68614
rect 463222 68378 463306 68614
rect 463542 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect -8726 68294 592650 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 66986 68294
rect 67222 68058 67306 68294
rect 67542 68058 102986 68294
rect 103222 68058 103306 68294
rect 103542 68058 138986 68294
rect 139222 68058 139306 68294
rect 139542 68058 174986 68294
rect 175222 68058 175306 68294
rect 175542 68058 210986 68294
rect 211222 68058 211306 68294
rect 211542 68058 246986 68294
rect 247222 68058 247306 68294
rect 247542 68058 282986 68294
rect 283222 68058 283306 68294
rect 283542 68058 318986 68294
rect 319222 68058 319306 68294
rect 319542 68058 354986 68294
rect 355222 68058 355306 68294
rect 355542 68058 390986 68294
rect 391222 68058 391306 68294
rect 391542 68058 426986 68294
rect 427222 68058 427306 68294
rect 427542 68058 462986 68294
rect 463222 68058 463306 68294
rect 463542 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect -8726 68026 592650 68058
rect -6806 64894 590730 64926
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 63266 64894
rect 63502 64658 63586 64894
rect 63822 64658 99266 64894
rect 99502 64658 99586 64894
rect 99822 64658 135266 64894
rect 135502 64658 135586 64894
rect 135822 64658 171266 64894
rect 171502 64658 171586 64894
rect 171822 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 243266 64894
rect 243502 64658 243586 64894
rect 243822 64658 279266 64894
rect 279502 64658 279586 64894
rect 279822 64658 315266 64894
rect 315502 64658 315586 64894
rect 315822 64658 351266 64894
rect 351502 64658 351586 64894
rect 351822 64658 387266 64894
rect 387502 64658 387586 64894
rect 387822 64658 423266 64894
rect 423502 64658 423586 64894
rect 423822 64658 459266 64894
rect 459502 64658 459586 64894
rect 459822 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect -6806 64574 590730 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 63266 64574
rect 63502 64338 63586 64574
rect 63822 64338 99266 64574
rect 99502 64338 99586 64574
rect 99822 64338 135266 64574
rect 135502 64338 135586 64574
rect 135822 64338 171266 64574
rect 171502 64338 171586 64574
rect 171822 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 243266 64574
rect 243502 64338 243586 64574
rect 243822 64338 279266 64574
rect 279502 64338 279586 64574
rect 279822 64338 315266 64574
rect 315502 64338 315586 64574
rect 315822 64338 351266 64574
rect 351502 64338 351586 64574
rect 351822 64338 387266 64574
rect 387502 64338 387586 64574
rect 387822 64338 423266 64574
rect 423502 64338 423586 64574
rect 423822 64338 459266 64574
rect 459502 64338 459586 64574
rect 459822 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect -6806 64306 590730 64338
rect -4886 61174 588810 61206
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 59546 61174
rect 59782 60938 59866 61174
rect 60102 60938 95546 61174
rect 95782 60938 95866 61174
rect 96102 60938 131546 61174
rect 131782 60938 131866 61174
rect 132102 60938 167546 61174
rect 167782 60938 167866 61174
rect 168102 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 239546 61174
rect 239782 60938 239866 61174
rect 240102 60938 275546 61174
rect 275782 60938 275866 61174
rect 276102 60938 311546 61174
rect 311782 60938 311866 61174
rect 312102 60938 347546 61174
rect 347782 60938 347866 61174
rect 348102 60938 383546 61174
rect 383782 60938 383866 61174
rect 384102 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect -4886 60854 588810 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 59546 60854
rect 59782 60618 59866 60854
rect 60102 60618 95546 60854
rect 95782 60618 95866 60854
rect 96102 60618 131546 60854
rect 131782 60618 131866 60854
rect 132102 60618 167546 60854
rect 167782 60618 167866 60854
rect 168102 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 239546 60854
rect 239782 60618 239866 60854
rect 240102 60618 275546 60854
rect 275782 60618 275866 60854
rect 276102 60618 311546 60854
rect 311782 60618 311866 60854
rect 312102 60618 347546 60854
rect 347782 60618 347866 60854
rect 348102 60618 383546 60854
rect 383782 60618 383866 60854
rect 384102 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect -4886 60586 588810 60618
rect -2966 57454 586890 57486
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect -2966 57134 586890 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect -2966 56866 586890 56898
rect -8726 50614 592650 50646
rect -8726 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 592650 50294
rect -8726 50026 592650 50058
rect -6806 46894 590730 46926
rect -6806 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 590730 46894
rect -6806 46574 590730 46658
rect -6806 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 590730 46574
rect -6806 46306 590730 46338
rect -4886 43174 588810 43206
rect -4886 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 588810 43174
rect -4886 42854 588810 42938
rect -4886 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 588810 42854
rect -4886 42586 588810 42618
rect -2966 39454 586890 39486
rect -2966 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 586890 39454
rect -2966 39134 586890 39218
rect -2966 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 586890 39134
rect -2966 38866 586890 38898
rect -8726 32614 592650 32646
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect -8726 32294 592650 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect -8726 32026 592650 32058
rect -6806 28894 590730 28926
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect -6806 28574 590730 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect -6806 28306 590730 28338
rect -4886 25174 588810 25206
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect -4886 24854 588810 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect -4886 24586 588810 24618
rect -2966 21454 586890 21486
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect -2966 21134 586890 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect -2966 20866 586890 20898
rect -8726 14614 592650 14646
rect -8726 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 592650 14294
rect -8726 14026 592650 14058
rect -6806 10894 590730 10926
rect -6806 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 590730 10894
rect -6806 10574 590730 10658
rect -6806 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 590730 10574
rect -6806 10306 590730 10338
rect -4886 7174 588810 7206
rect -4886 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 588810 7174
rect -4886 6854 588810 6938
rect -4886 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 588810 6854
rect -4886 6586 588810 6618
rect -2966 3454 586890 3486
rect -2966 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 586890 3454
rect -2966 3134 586890 3218
rect -2966 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 586890 3134
rect -2966 2866 586890 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use digitalcore_macro  digitalcore
timestamp 1641031085
transform 1 0 200000 0 1 100000
box 0 0 100000 200000
use collapsering_macro  ring0
timestamp 1641031085
transform 1 0 160000 0 1 124000
box 934 0 10000 29776
use ringosc_macro  ring1
timestamp 1641031085
transform 1 0 160000 0 1 160000
box 934 0 10000 29504
use collapsering_macro  ring2
timestamp 1641031085
transform 1 0 360000 0 1 124000
box 934 0 10000 29776
use collapsering_macro  ring3
timestamp 1641031085
transform 1 0 360000 0 1 196000
box 934 0 10000 29776
use collapsering_macro  ring4
timestamp 1641031085
transform 1 0 360000 0 1 268000
box 934 0 10000 29776
use collapsering_macro  ring5
timestamp 1641031085
transform 1 0 360000 0 1 340000
box 934 0 10000 29776
use ringosc_macro  ring6
timestamp 1641031085
transform 1 0 432000 0 1 124000
box 934 0 10000 29504
use ringosc_macro  ring7
timestamp 1641031085
transform 1 0 432000 0 1 196000
box 934 0 10000 29504
use ringosc_macro  ring8
timestamp 1641031085
transform 1 0 432000 0 1 268000
box 934 0 10000 29504
use ringosc_macro  ring9
timestamp 1641031085
transform 1 0 432000 0 1 340000
box 934 0 10000 29504
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 38866 586890 39486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 74866 586890 75486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 110866 586890 111486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 146866 586890 147486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 182866 586890 183486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 218866 586890 219486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 254866 586890 255486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 290866 586890 291486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 326866 586890 327486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 362866 586890 363486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 398866 586890 399486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 434866 586890 435486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 470866 586890 471486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 506866 586890 507486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 542866 586890 543486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 578866 586890 579486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 614866 586890 615486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 650866 586890 651486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 686866 586890 687486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 -1894 218414 98000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 -1894 254414 98000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 -1894 290414 98000 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 -1894 362414 122000 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 -1894 434414 122000 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 156000 362414 194000 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 156000 434414 194000 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 228000 362414 266000 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 228000 434414 266000 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 300000 362414 338000 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 300000 434414 338000 6 vccd1
port 531 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 1794 -1894 2414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 -1894 38414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 -1894 74414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 -1894 110414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 -1894 146414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 -1894 182414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 302000 218414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 302000 254414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 302000 290414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 -1894 326414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 372000 362414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 -1894 398414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 372000 434414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 -1894 470414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 -1894 506414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 -1894 542414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 577794 -1894 578414 705830 6 vccd1
port 531 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 532 nsew power input
rlabel metal5 s -4886 6586 588810 7206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 42586 588810 43206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 78586 588810 79206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 114586 588810 115206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 150586 588810 151206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 186586 588810 187206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 222586 588810 223206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 258586 588810 259206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 294586 588810 295206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 330586 588810 331206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 366586 588810 367206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 402586 588810 403206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 438586 588810 439206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 474586 588810 475206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 510586 588810 511206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 546586 588810 547206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 582586 588810 583206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 618586 588810 619206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 654586 588810 655206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 690586 588810 691206 6 vccd2
port 532 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 -3814 222134 98000 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 -3814 258134 98000 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 -3814 294134 98000 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 -3814 366134 122000 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 -3814 438134 122000 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 156000 366134 194000 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 156000 438134 194000 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 228000 366134 266000 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 228000 438134 266000 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 300000 366134 338000 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 300000 438134 338000 6 vccd2
port 532 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 532 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 5514 -3814 6134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 41514 -3814 42134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 -3814 78134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 -3814 114134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 -3814 150134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 -3814 186134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 302000 222134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 302000 258134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 302000 294134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 -3814 330134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 372000 366134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 -3814 402134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 372000 438134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 -3814 474134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 -3814 510134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 545514 -3814 546134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 581514 -3814 582134 707750 6 vccd2
port 532 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 533 nsew power input
rlabel metal5 s -6806 10306 590730 10926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 46306 590730 46926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 82306 590730 82926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 118306 590730 118926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 154306 590730 154926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 190306 590730 190926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 226306 590730 226926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 262306 590730 262926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 298306 590730 298926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 334306 590730 334926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 370306 590730 370926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 406306 590730 406926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 442306 590730 442926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 478306 590730 478926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 514306 590730 514926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 550306 590730 550926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 586306 590730 586926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 622306 590730 622926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 658306 590730 658926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 694306 590730 694926 6 vdda1
port 533 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 -5734 225854 98000 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 -5734 261854 98000 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 -5734 297854 98000 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 -5734 369854 122000 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 -5734 441854 122000 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 156000 369854 194000 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 156000 441854 194000 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 228000 369854 266000 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 228000 441854 266000 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 300000 369854 338000 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 300000 441854 338000 6 vdda1
port 533 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 533 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 9234 -5734 9854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 45234 -5734 45854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 -5734 81854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 -5734 117854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 -5734 153854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 -5734 189854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 302000 225854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 302000 261854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 302000 297854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 -5734 333854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 372000 369854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 -5734 405854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 372000 441854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 -5734 477854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 -5734 513854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 549234 -5734 549854 709670 6 vdda1
port 533 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 534 nsew power input
rlabel metal5 s -8726 14026 592650 14646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 50026 592650 50646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 86026 592650 86646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 122026 592650 122646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 158026 592650 158646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 194026 592650 194646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 230026 592650 230646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 266026 592650 266646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 302026 592650 302646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 338026 592650 338646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 374026 592650 374646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 410026 592650 410646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 446026 592650 446646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 482026 592650 482646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 518026 592650 518646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 554026 592650 554646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 590026 592650 590646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 626026 592650 626646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 662026 592650 662646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 698026 592650 698646 6 vdda2
port 534 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 -7654 229574 98000 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 -7654 265574 98000 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 -7654 301574 98000 6 vdda2
port 534 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 534 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 12954 -7654 13574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 -7654 49574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 -7654 85574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 -7654 121574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 -7654 157574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 -7654 193574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 302000 229574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 302000 265574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 302000 301574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 -7654 337574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 -7654 373574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 -7654 409574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 -7654 445574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 -7654 481574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 -7654 517574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 552954 -7654 553574 711590 6 vdda2
port 534 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 28306 590730 28926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 64306 590730 64926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 100306 590730 100926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 136306 590730 136926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 172306 590730 172926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 208306 590730 208926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 244306 590730 244926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 280306 590730 280926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 316306 590730 316926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 352306 590730 352926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 388306 590730 388926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 424306 590730 424926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 460306 590730 460926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 496306 590730 496926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 532306 590730 532926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 568306 590730 568926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 604306 590730 604926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 640306 590730 640926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 676306 590730 676926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 -5734 207854 98000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 -5734 243854 98000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 -5734 279854 98000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 -5734 171854 122000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 156000 171854 158000 6 vssa1
port 535 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 535 nsew ground input
rlabel metal4 s 27234 -5734 27854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 -5734 63854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 -5734 99854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 -5734 135854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 192000 171854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 302000 207854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 302000 243854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 302000 279854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 -5734 315854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 -5734 351854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 -5734 387854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 -5734 423854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 -5734 459854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 -5734 495854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 -5734 531854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 567234 -5734 567854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 32026 592650 32646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 68026 592650 68646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 104026 592650 104646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 140026 592650 140646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 176026 592650 176646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 212026 592650 212646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 248026 592650 248646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 284026 592650 284646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 320026 592650 320646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 356026 592650 356646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 392026 592650 392646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 428026 592650 428646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 464026 592650 464646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 500026 592650 500646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 536026 592650 536646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 572026 592650 572646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 608026 592650 608646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 644026 592650 644646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 680026 592650 680646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 -7654 211574 98000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 -7654 247574 98000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 -7654 283574 98000 6 vssa2
port 536 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 536 nsew ground input
rlabel metal4 s 30954 -7654 31574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 -7654 67574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 -7654 103574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 -7654 139574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 -7654 175574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 302000 211574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 302000 247574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 302000 283574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 -7654 319574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 -7654 355574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 -7654 391574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 -7654 427574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 -7654 463574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 -7654 499574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 -7654 535574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 570954 -7654 571574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 20866 586890 21486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 56866 586890 57486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 92866 586890 93486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 128866 586890 129486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 164866 586890 165486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 200866 586890 201486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 236866 586890 237486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 272866 586890 273486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 308866 586890 309486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 344866 586890 345486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 380866 586890 381486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 416866 586890 417486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 452866 586890 453486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 488866 586890 489486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 524866 586890 525486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 560866 586890 561486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 596866 586890 597486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 632866 586890 633486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 668866 586890 669486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 -1894 200414 98000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 -1894 236414 98000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 -1894 272414 98000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 -1894 164414 122000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 156000 164414 158000 6 vssd1
port 537 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 537 nsew ground input
rlabel metal4 s 19794 -1894 20414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 -1894 56414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 -1894 92414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 -1894 128414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 192000 164414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 302000 200414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 302000 236414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 302000 272414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 -1894 308414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 -1894 344414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 -1894 380414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 -1894 416414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 -1894 452414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 -1894 488414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 -1894 524414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 559794 -1894 560414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 24586 588810 25206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 60586 588810 61206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 96586 588810 97206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 132586 588810 133206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 168586 588810 169206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 204586 588810 205206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 240586 588810 241206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 276586 588810 277206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 312586 588810 313206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 348586 588810 349206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 384586 588810 385206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 420586 588810 421206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 456586 588810 457206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 492586 588810 493206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 528586 588810 529206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 564586 588810 565206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 600586 588810 601206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 636586 588810 637206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 672586 588810 673206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 -3814 204134 98000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 -3814 240134 98000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 -3814 276134 98000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 -3814 168134 122000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 156000 168134 158000 6 vssd2
port 538 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 538 nsew ground input
rlabel metal4 s 23514 -3814 24134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 -3814 60134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 -3814 96134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 -3814 132134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 192000 168134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 302000 204134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 302000 240134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 302000 276134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 -3814 312134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 -3814 348134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 -3814 384134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 -3814 420134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 -3814 456134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 -3814 492134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 -3814 528134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 563514 -3814 564134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 539 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 540 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 541 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 542 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 543 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 544 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 545 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 546 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 547 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 548 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 549 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 550 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 551 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 552 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 553 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 554 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 555 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 556 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 557 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 558 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 559 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 560 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 561 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 562 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 563 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 564 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 565 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 566 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 567 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 568 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 569 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 570 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 571 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 572 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 573 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 574 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 575 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 576 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 577 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 578 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 579 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 580 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 581 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 582 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 583 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 584 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 585 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 586 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 587 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 588 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 589 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 590 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 591 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 592 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 593 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 594 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 595 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 596 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 597 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 598 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 599 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 600 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 601 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 602 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 603 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 604 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 605 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 606 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 607 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 608 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 609 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 610 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 611 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 612 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 613 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 614 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 615 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 616 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 617 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 618 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 619 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 620 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 621 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 622 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 623 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 624 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 625 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 626 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 627 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 628 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 629 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 630 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 631 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 632 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 633 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 634 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 635 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 636 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 637 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 638 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 639 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 640 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 641 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 642 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 643 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
