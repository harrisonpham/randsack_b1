magic
tech sky130A
magscale 1 2
timestamp 1635131530
<< metal1 >>
rect 331214 702992 331220 703044
rect 331272 703032 331278 703044
rect 332502 703032 332508 703044
rect 331272 703004 332508 703032
rect 331272 702992 331278 703004
rect 332502 702992 332508 703004
rect 332560 702992 332566 703044
rect 294598 700544 294604 700596
rect 294656 700584 294662 700596
rect 364978 700584 364984 700596
rect 294656 700556 364984 700584
rect 294656 700544 294662 700556
rect 364978 700544 364984 700556
rect 365036 700544 365042 700596
rect 298738 700476 298744 700528
rect 298796 700516 298802 700528
rect 397454 700516 397460 700528
rect 298796 700488 397460 700516
rect 298796 700476 298802 700488
rect 397454 700476 397460 700488
rect 397512 700476 397518 700528
rect 40494 700408 40500 700460
rect 40552 700448 40558 700460
rect 41322 700448 41328 700460
rect 40552 700420 41328 700448
rect 40552 700408 40558 700420
rect 41322 700408 41328 700420
rect 41380 700408 41386 700460
rect 305638 700408 305644 700460
rect 305696 700448 305702 700460
rect 494790 700448 494796 700460
rect 305696 700420 494796 700448
rect 305696 700408 305702 700420
rect 494790 700408 494796 700420
rect 494848 700408 494854 700460
rect 137830 700340 137836 700392
rect 137888 700380 137894 700392
rect 195238 700380 195244 700392
rect 137888 700352 195244 700380
rect 137888 700340 137894 700352
rect 195238 700340 195244 700352
rect 195296 700340 195302 700392
rect 244918 700340 244924 700392
rect 244976 700380 244982 700392
rect 462314 700380 462320 700392
rect 244976 700352 462320 700380
rect 244976 700340 244982 700352
rect 462314 700340 462320 700352
rect 462372 700340 462378 700392
rect 24302 700272 24308 700324
rect 24360 700312 24366 700324
rect 137278 700312 137284 700324
rect 24360 700284 137284 700312
rect 24360 700272 24366 700284
rect 137278 700272 137284 700284
rect 137336 700272 137342 700324
rect 218974 700272 218980 700324
rect 219032 700312 219038 700324
rect 240778 700312 240784 700324
rect 219032 700284 240784 700312
rect 219032 700272 219038 700284
rect 240778 700272 240784 700284
rect 240836 700272 240842 700324
rect 242158 700272 242164 700324
rect 242216 700312 242222 700324
rect 527174 700312 527180 700324
rect 242216 700284 527180 700312
rect 242216 700272 242222 700284
rect 527174 700272 527180 700284
rect 527232 700272 527238 700324
rect 559650 700272 559656 700324
rect 559708 700312 559714 700324
rect 582926 700312 582932 700324
rect 559708 700284 582932 700312
rect 559708 700272 559714 700284
rect 582926 700272 582932 700284
rect 582984 700272 582990 700324
rect 154114 699728 154120 699780
rect 154172 699768 154178 699780
rect 157978 699768 157984 699780
rect 154172 699740 157984 699768
rect 154172 699728 154178 699740
rect 157978 699728 157984 699740
rect 158036 699728 158042 699780
rect 105446 699660 105452 699712
rect 105504 699700 105510 699712
rect 106182 699700 106188 699712
rect 105504 699672 106188 699700
rect 105504 699660 105510 699672
rect 106182 699660 106188 699672
rect 106240 699660 106246 699712
rect 170306 699660 170312 699712
rect 170364 699700 170370 699712
rect 171042 699700 171048 699712
rect 170364 699672 171048 699700
rect 170364 699660 170370 699672
rect 171042 699660 171048 699672
rect 171100 699660 171106 699712
rect 235166 699660 235172 699712
rect 235224 699700 235230 699712
rect 235902 699700 235908 699712
rect 235224 699672 235908 699700
rect 235224 699660 235230 699672
rect 235902 699660 235908 699672
rect 235960 699660 235966 699712
rect 282178 699660 282184 699712
rect 282236 699700 282242 699712
rect 283834 699700 283840 699712
rect 282236 699672 283840 699700
rect 282236 699660 282242 699672
rect 283834 699660 283840 699672
rect 283892 699660 283898 699712
rect 347038 699660 347044 699712
rect 347096 699700 347102 699712
rect 348786 699700 348792 699712
rect 347096 699672 348792 699700
rect 347096 699660 347102 699672
rect 348786 699660 348792 699672
rect 348844 699660 348850 699712
rect 476758 699660 476764 699712
rect 476816 699700 476822 699712
rect 478506 699700 478512 699712
rect 476816 699672 478512 699700
rect 476816 699660 476822 699672
rect 478506 699660 478512 699672
rect 478564 699660 478570 699712
rect 266354 697552 266360 697604
rect 266412 697592 266418 697604
rect 267642 697592 267648 697604
rect 266412 697564 267648 697592
rect 266412 697552 266418 697564
rect 267642 697552 267648 697564
rect 267700 697552 267706 697604
rect 3418 683136 3424 683188
rect 3476 683176 3482 683188
rect 199378 683176 199384 683188
rect 3476 683148 199384 683176
rect 3476 683136 3482 683148
rect 199378 683136 199384 683148
rect 199436 683136 199442 683188
rect 3510 670692 3516 670744
rect 3568 670732 3574 670744
rect 260098 670732 260104 670744
rect 3568 670704 260104 670732
rect 3568 670692 3574 670704
rect 260098 670692 260104 670704
rect 260156 670692 260162 670744
rect 3418 656888 3424 656940
rect 3476 656928 3482 656940
rect 262858 656928 262864 656940
rect 3476 656900 262864 656928
rect 3476 656888 3482 656900
rect 262858 656888 262864 656900
rect 262916 656888 262922 656940
rect 251082 649272 251088 649324
rect 251140 649312 251146 649324
rect 266354 649312 266360 649324
rect 251140 649284 266360 649312
rect 251140 649272 251146 649284
rect 266354 649272 266360 649284
rect 266412 649272 266418 649324
rect 3418 632068 3424 632120
rect 3476 632108 3482 632120
rect 258718 632108 258724 632120
rect 3476 632080 258724 632108
rect 3476 632068 3482 632080
rect 258718 632068 258724 632080
rect 258776 632068 258782 632120
rect 3142 618264 3148 618316
rect 3200 618304 3206 618316
rect 231118 618304 231124 618316
rect 3200 618276 231124 618304
rect 3200 618264 3206 618276
rect 231118 618264 231124 618276
rect 231176 618264 231182 618316
rect 235902 606432 235908 606484
rect 235960 606472 235966 606484
rect 252554 606472 252560 606484
rect 235960 606444 252560 606472
rect 235960 606432 235966 606444
rect 252554 606432 252560 606444
rect 252612 606432 252618 606484
rect 3234 605820 3240 605872
rect 3292 605860 3298 605872
rect 192478 605860 192484 605872
rect 3292 605832 192484 605860
rect 3292 605820 3298 605832
rect 192478 605820 192484 605832
rect 192536 605820 192542 605872
rect 3326 579640 3332 579692
rect 3384 579680 3390 579692
rect 255958 579680 255964 579692
rect 3384 579652 255964 579680
rect 3384 579640 3390 579652
rect 255958 579640 255964 579652
rect 256016 579640 256022 579692
rect 3418 565836 3424 565888
rect 3476 565876 3482 565888
rect 39298 565876 39304 565888
rect 3476 565848 39304 565876
rect 3476 565836 3482 565848
rect 39298 565836 39304 565848
rect 39356 565836 39362 565888
rect 3418 553392 3424 553444
rect 3476 553432 3482 553444
rect 173158 553432 173164 553444
rect 3476 553404 173164 553432
rect 3476 553392 3482 553404
rect 173158 553392 173164 553404
rect 173216 553392 173222 553444
rect 3418 527144 3424 527196
rect 3476 527184 3482 527196
rect 210418 527184 210424 527196
rect 3476 527156 210424 527184
rect 3476 527144 3482 527156
rect 210418 527144 210424 527156
rect 210476 527144 210482 527196
rect 3418 514768 3424 514820
rect 3476 514808 3482 514820
rect 206278 514808 206284 514820
rect 3476 514780 206284 514808
rect 3476 514768 3482 514780
rect 206278 514768 206284 514780
rect 206336 514768 206342 514820
rect 3050 474716 3056 474768
rect 3108 474756 3114 474768
rect 197998 474756 198004 474768
rect 3108 474728 198004 474756
rect 3108 474716 3114 474728
rect 197998 474716 198004 474728
rect 198056 474716 198062 474768
rect 3510 462340 3516 462392
rect 3568 462380 3574 462392
rect 191098 462380 191104 462392
rect 3568 462352 191104 462380
rect 3568 462340 3574 462352
rect 191098 462340 191104 462352
rect 191156 462340 191162 462392
rect 238662 458804 238668 458856
rect 238720 458844 238726 458856
rect 583386 458844 583392 458856
rect 238720 458816 583392 458844
rect 238720 458804 238726 458816
rect 583386 458804 583392 458816
rect 583444 458804 583450 458856
rect 291838 456764 291844 456816
rect 291896 456804 291902 456816
rect 580166 456804 580172 456816
rect 291896 456776 580172 456804
rect 291896 456764 291902 456776
rect 580166 456764 580172 456776
rect 580224 456764 580230 456816
rect 3142 448536 3148 448588
rect 3200 448576 3206 448588
rect 166258 448576 166264 448588
rect 3200 448548 166264 448576
rect 3200 448536 3206 448548
rect 166258 448536 166264 448548
rect 166316 448536 166322 448588
rect 224862 430584 224868 430636
rect 224920 430624 224926 430636
rect 580166 430624 580172 430636
rect 224920 430596 580172 430624
rect 224920 430584 224926 430596
rect 580166 430584 580172 430596
rect 580224 430584 580230 430636
rect 3510 422288 3516 422340
rect 3568 422328 3574 422340
rect 196618 422328 196624 422340
rect 3568 422300 196624 422328
rect 3568 422288 3574 422300
rect 196618 422288 196624 422300
rect 196676 422288 196682 422340
rect 289078 418140 289084 418192
rect 289136 418180 289142 418192
rect 580166 418180 580172 418192
rect 289136 418152 580172 418180
rect 289136 418140 289142 418152
rect 580166 418140 580172 418152
rect 580224 418140 580230 418192
rect 2866 409844 2872 409896
rect 2924 409884 2930 409896
rect 249058 409884 249064 409896
rect 2924 409856 249064 409884
rect 2924 409844 2930 409856
rect 249058 409844 249064 409856
rect 249116 409844 249122 409896
rect 234522 403588 234528 403640
rect 234580 403628 234586 403640
rect 583478 403628 583484 403640
rect 234580 403600 583484 403628
rect 234580 403588 234586 403600
rect 583478 403588 583484 403600
rect 583536 403588 583542 403640
rect 3510 397468 3516 397520
rect 3568 397508 3574 397520
rect 177298 397508 177304 397520
rect 3568 397480 177304 397508
rect 3568 397468 3574 397480
rect 177298 397468 177304 397480
rect 177356 397468 177362 397520
rect 3510 371220 3516 371272
rect 3568 371260 3574 371272
rect 213178 371260 213184 371272
rect 3568 371232 213184 371260
rect 3568 371220 3574 371232
rect 213178 371220 213184 371232
rect 213236 371220 213242 371272
rect 246298 364352 246304 364404
rect 246356 364392 246362 364404
rect 580166 364392 580172 364404
rect 246356 364364 580172 364392
rect 246356 364352 246362 364364
rect 580166 364352 580172 364364
rect 580224 364352 580230 364404
rect 3142 357416 3148 357468
rect 3200 357456 3206 357468
rect 280338 357456 280344 357468
rect 3200 357428 280344 357456
rect 3200 357416 3206 357428
rect 280338 357416 280344 357428
rect 280396 357416 280402 357468
rect 231118 355308 231124 355360
rect 231176 355348 231182 355360
rect 267274 355348 267280 355360
rect 231176 355320 267280 355348
rect 231176 355308 231182 355320
rect 267274 355308 267280 355320
rect 267332 355308 267338 355360
rect 231762 353948 231768 354000
rect 231820 353988 231826 354000
rect 583662 353988 583668 354000
rect 231820 353960 583668 353988
rect 231820 353948 231826 353960
rect 583662 353948 583668 353960
rect 583720 353948 583726 354000
rect 295978 351908 295984 351960
rect 296036 351948 296042 351960
rect 579890 351948 579896 351960
rect 296036 351920 579896 351948
rect 296036 351908 296042 351920
rect 579890 351908 579896 351920
rect 579948 351908 579954 351960
rect 3326 345040 3332 345092
rect 3384 345080 3390 345092
rect 226978 345080 226984 345092
rect 3384 345052 226984 345080
rect 3384 345040 3390 345052
rect 226978 345040 226984 345052
rect 227036 345040 227042 345092
rect 39298 344292 39304 344344
rect 39356 344332 39362 344344
rect 269942 344332 269948 344344
rect 39356 344304 269948 344332
rect 39356 344292 39362 344304
rect 269942 344292 269948 344304
rect 270000 344292 270006 344344
rect 580902 343204 580908 343256
rect 580960 343244 580966 343256
rect 583478 343244 583484 343256
rect 580960 343216 583484 343244
rect 580960 343204 580966 343216
rect 583478 343204 583484 343216
rect 583536 343204 583542 343256
rect 235258 324300 235264 324352
rect 235316 324340 235322 324352
rect 580166 324340 580172 324352
rect 235316 324312 580172 324340
rect 235316 324300 235322 324312
rect 580166 324300 580172 324312
rect 580224 324300 580230 324352
rect 3326 318792 3332 318844
rect 3384 318832 3390 318844
rect 209038 318832 209044 318844
rect 3384 318804 209044 318832
rect 3384 318792 3390 318804
rect 209038 318792 209044 318804
rect 209096 318792 209102 318844
rect 249058 318044 249064 318096
rect 249116 318084 249122 318096
rect 277762 318084 277768 318096
rect 249116 318056 277768 318084
rect 249116 318044 249122 318056
rect 277762 318044 277768 318056
rect 277820 318044 277826 318096
rect 220722 311856 220728 311908
rect 220780 311896 220786 311908
rect 580166 311896 580172 311908
rect 220780 311868 580172 311896
rect 220780 311856 220786 311868
rect 580166 311856 580172 311868
rect 580224 311856 580230 311908
rect 3510 304988 3516 305040
rect 3568 305028 3574 305040
rect 200758 305028 200764 305040
rect 3568 305000 200764 305028
rect 3568 304988 3574 305000
rect 200758 304988 200764 305000
rect 200816 304988 200822 305040
rect 229002 300092 229008 300144
rect 229060 300132 229066 300144
rect 583570 300132 583576 300144
rect 229060 300104 583576 300132
rect 229060 300092 229066 300104
rect 583570 300092 583576 300104
rect 583628 300092 583634 300144
rect 252462 294584 252468 294636
rect 252520 294624 252526 294636
rect 282178 294624 282184 294636
rect 252520 294596 282184 294624
rect 252520 294584 252526 294596
rect 282178 294584 282184 294596
rect 282236 294584 282242 294636
rect 3510 292544 3516 292596
rect 3568 292584 3574 292596
rect 282086 292584 282092 292596
rect 3568 292556 282092 292584
rect 3568 292544 3574 292556
rect 282086 292544 282092 292556
rect 282144 292544 282150 292596
rect 177298 286288 177304 286340
rect 177356 286328 177362 286340
rect 276842 286328 276848 286340
rect 177356 286300 276848 286328
rect 177356 286288 177362 286300
rect 276842 286288 276848 286300
rect 276900 286288 276906 286340
rect 232498 271872 232504 271924
rect 232556 271912 232562 271924
rect 580166 271912 580172 271924
rect 232556 271884 580172 271912
rect 232556 271872 232562 271884
rect 580166 271872 580172 271884
rect 580224 271872 580230 271924
rect 3050 266364 3056 266416
rect 3108 266404 3114 266416
rect 285674 266404 285680 266416
rect 3108 266376 285680 266404
rect 3108 266364 3114 266376
rect 285674 266364 285680 266376
rect 285732 266364 285738 266416
rect 217962 258068 217968 258120
rect 218020 258108 218026 258120
rect 580166 258108 580172 258120
rect 218020 258080 580172 258108
rect 218020 258068 218026 258080
rect 580166 258068 580172 258080
rect 580224 258068 580230 258120
rect 3510 253920 3516 253972
rect 3568 253960 3574 253972
rect 285582 253960 285588 253972
rect 3568 253932 285588 253960
rect 3568 253920 3574 253932
rect 285582 253920 285588 253932
rect 285640 253920 285646 253972
rect 240042 246304 240048 246356
rect 240100 246344 240106 246356
rect 582926 246344 582932 246356
rect 240100 246316 582932 246344
rect 240100 246304 240106 246316
rect 582926 246304 582932 246316
rect 582984 246304 582990 246356
rect 3050 240116 3056 240168
rect 3108 240156 3114 240168
rect 204898 240156 204904 240168
rect 3108 240128 204904 240156
rect 3108 240116 3114 240128
rect 204898 240116 204904 240128
rect 204956 240116 204962 240168
rect 215938 231820 215944 231872
rect 215996 231860 216002 231872
rect 580166 231860 580172 231872
rect 215996 231832 580172 231860
rect 215996 231820 216002 231832
rect 580166 231820 580172 231832
rect 580224 231820 580230 231872
rect 166258 228352 166264 228404
rect 166316 228392 166322 228404
rect 274266 228392 274272 228404
rect 166316 228364 274272 228392
rect 166316 228352 166322 228364
rect 274266 228352 274272 228364
rect 274324 228352 274330 228404
rect 3418 226992 3424 227044
rect 3476 227032 3482 227044
rect 271690 227032 271696 227044
rect 3476 227004 271696 227032
rect 3476 226992 3482 227004
rect 271690 226992 271696 227004
rect 271748 226992 271754 227044
rect 89622 224204 89628 224256
rect 89680 224244 89686 224256
rect 259454 224244 259460 224256
rect 89680 224216 259460 224244
rect 89680 224204 89686 224216
rect 259454 224204 259460 224216
rect 259512 224204 259518 224256
rect 260098 224204 260104 224256
rect 260156 224244 260162 224256
rect 264698 224244 264704 224256
rect 260156 224216 264704 224244
rect 260156 224204 260162 224216
rect 264698 224204 264704 224216
rect 264756 224204 264762 224256
rect 223482 221416 223488 221468
rect 223540 221456 223546 221468
rect 246298 221456 246304 221468
rect 223540 221428 246304 221456
rect 223540 221416 223546 221428
rect 246298 221416 246304 221428
rect 246356 221416 246362 221468
rect 249702 220056 249708 220108
rect 249760 220096 249766 220108
rect 347038 220096 347044 220108
rect 249760 220068 347044 220096
rect 249760 220056 249766 220068
rect 347038 220056 347044 220068
rect 347096 220056 347102 220108
rect 215202 218016 215208 218068
rect 215260 218056 215266 218068
rect 580166 218056 580172 218068
rect 215260 218028 580172 218056
rect 215260 218016 215266 218028
rect 580166 218016 580172 218028
rect 580224 218016 580230 218068
rect 246942 217268 246948 217320
rect 247000 217308 247006 217320
rect 412634 217308 412640 217320
rect 247000 217280 412640 217308
rect 247000 217268 247006 217280
rect 412634 217268 412640 217280
rect 412692 217268 412698 217320
rect 173158 215908 173164 215960
rect 173216 215948 173222 215960
rect 269022 215948 269028 215960
rect 173216 215920 269028 215948
rect 173216 215908 173222 215920
rect 269022 215908 269028 215920
rect 269080 215908 269086 215960
rect 241422 214548 241428 214600
rect 241480 214588 241486 214600
rect 542354 214588 542360 214600
rect 241480 214560 542360 214588
rect 241480 214548 241486 214560
rect 542354 214548 542360 214560
rect 542412 214548 542418 214600
rect 3142 213936 3148 213988
rect 3200 213976 3206 213988
rect 287054 213976 287060 213988
rect 3200 213948 287060 213976
rect 3200 213936 3206 213948
rect 287054 213936 287060 213948
rect 287112 213936 287118 213988
rect 240778 211828 240784 211880
rect 240836 211868 240842 211880
rect 254302 211868 254308 211880
rect 240836 211840 254308 211868
rect 240836 211828 240842 211840
rect 254302 211828 254308 211840
rect 254360 211828 254366 211880
rect 222102 211760 222108 211812
rect 222160 211800 222166 211812
rect 295978 211800 295984 211812
rect 222160 211772 295984 211800
rect 222160 211760 222166 211772
rect 295978 211760 295984 211772
rect 296036 211760 296042 211812
rect 580902 211080 580908 211132
rect 580960 211120 580966 211132
rect 582374 211120 582380 211132
rect 580960 211092 582380 211120
rect 580960 211080 580966 211092
rect 582374 211080 582380 211092
rect 582432 211080 582438 211132
rect 226242 210808 226248 210860
rect 226300 210848 226306 210860
rect 289078 210848 289084 210860
rect 226300 210820 289084 210848
rect 226300 210808 226306 210820
rect 289078 210808 289084 210820
rect 289136 210808 289142 210860
rect 206278 210740 206284 210792
rect 206336 210780 206342 210792
rect 272518 210780 272524 210792
rect 206336 210752 272524 210780
rect 206336 210740 206342 210752
rect 272518 210740 272524 210752
rect 272576 210740 272582 210792
rect 200758 210672 200764 210724
rect 200816 210712 200822 210724
rect 282914 210712 282920 210724
rect 200816 210684 282920 210712
rect 200816 210672 200822 210684
rect 282914 210672 282920 210684
rect 282972 210672 282978 210724
rect 191098 210604 191104 210656
rect 191156 210644 191162 210656
rect 275094 210644 275100 210656
rect 191156 210616 275100 210644
rect 191156 210604 191162 210616
rect 275094 210604 275100 210616
rect 275152 210604 275158 210656
rect 137278 210536 137284 210588
rect 137336 210576 137342 210588
rect 262122 210576 262128 210588
rect 137336 210548 262128 210576
rect 137336 210536 137342 210548
rect 262122 210536 262128 210548
rect 262180 210536 262186 210588
rect 244182 210468 244188 210520
rect 244240 210508 244246 210520
rect 476758 210508 476764 210520
rect 244240 210480 476764 210508
rect 244240 210468 244246 210480
rect 476758 210468 476764 210480
rect 476816 210468 476822 210520
rect 220630 210400 220636 210452
rect 220688 210440 220694 210452
rect 235258 210440 235264 210452
rect 220688 210412 235264 210440
rect 220688 210400 220694 210412
rect 235258 210400 235264 210412
rect 235316 210400 235322 210452
rect 235902 210400 235908 210452
rect 235960 210440 235966 210452
rect 582558 210440 582564 210452
rect 235960 210412 582564 210440
rect 235960 210400 235966 210412
rect 582558 210400 582564 210412
rect 582616 210400 582622 210452
rect 226978 209448 226984 209500
rect 227036 209488 227042 209500
rect 279510 209488 279516 209500
rect 227036 209460 279516 209488
rect 227036 209448 227042 209460
rect 279510 209448 279516 209460
rect 279568 209448 279574 209500
rect 199378 209380 199384 209432
rect 199436 209420 199442 209432
rect 262950 209420 262956 209432
rect 199436 209392 262956 209420
rect 199436 209380 199442 209392
rect 262950 209380 262956 209392
rect 263008 209380 263014 209432
rect 192478 209312 192484 209364
rect 192536 209352 192542 209364
rect 266446 209352 266452 209364
rect 192536 209324 266452 209352
rect 192536 209312 192542 209324
rect 266446 209312 266452 209324
rect 266504 209312 266510 209364
rect 204898 209244 204904 209296
rect 204956 209284 204962 209296
rect 284662 209284 284668 209296
rect 204956 209256 284668 209284
rect 204956 209244 204962 209256
rect 284662 209244 284668 209256
rect 284720 209244 284726 209296
rect 8202 209176 8208 209228
rect 8260 209216 8266 209228
rect 260742 209216 260748 209228
rect 8260 209188 260748 209216
rect 8260 209176 8266 209188
rect 260742 209176 260748 209188
rect 260800 209176 260806 209228
rect 232958 209108 232964 209160
rect 233016 209148 233022 209160
rect 582834 209148 582840 209160
rect 233016 209120 582840 209148
rect 233016 209108 233022 209120
rect 582834 209108 582840 209120
rect 582892 209108 582898 209160
rect 227622 209040 227628 209092
rect 227680 209080 227686 209092
rect 583294 209080 583300 209092
rect 227680 209052 583300 209080
rect 227680 209040 227686 209052
rect 583294 209040 583300 209052
rect 583352 209040 583358 209092
rect 262858 208836 262864 208888
rect 262916 208876 262922 208888
rect 263870 208876 263876 208888
rect 262916 208848 263876 208876
rect 262916 208836 262922 208848
rect 263870 208836 263876 208848
rect 263928 208836 263934 208888
rect 213178 208020 213184 208072
rect 213236 208060 213242 208072
rect 278590 208060 278596 208072
rect 213236 208032 278596 208060
rect 213236 208020 213242 208032
rect 278590 208020 278596 208032
rect 278648 208020 278654 208072
rect 196618 207952 196624 208004
rect 196676 207992 196682 208004
rect 276014 207992 276020 208004
rect 196676 207964 276020 207992
rect 196676 207952 196682 207964
rect 276014 207952 276020 207964
rect 276072 207952 276078 208004
rect 157978 207884 157984 207936
rect 158036 207924 158042 207936
rect 256878 207924 256884 207936
rect 158036 207896 256884 207924
rect 158036 207884 158042 207896
rect 256878 207884 256884 207896
rect 256936 207884 256942 207936
rect 246022 207816 246028 207868
rect 246080 207856 246086 207868
rect 429194 207856 429200 207868
rect 246080 207828 429200 207856
rect 246080 207816 246086 207828
rect 429194 207816 429200 207828
rect 429252 207816 429258 207868
rect 41322 207748 41328 207800
rect 41380 207788 41386 207800
rect 259178 207788 259184 207800
rect 41380 207760 259184 207788
rect 41380 207748 41386 207760
rect 259178 207748 259184 207760
rect 259236 207748 259242 207800
rect 223850 207680 223856 207732
rect 223908 207720 223914 207732
rect 583386 207720 583392 207732
rect 223908 207692 583392 207720
rect 223908 207680 223914 207692
rect 583386 207680 583392 207692
rect 583444 207680 583450 207732
rect 216398 207612 216404 207664
rect 216456 207652 216462 207664
rect 582926 207652 582932 207664
rect 216456 207624 582932 207652
rect 216456 207612 216462 207624
rect 582926 207612 582932 207624
rect 582984 207612 582990 207664
rect 214282 207000 214288 207052
rect 214340 207040 214346 207052
rect 215938 207040 215944 207052
rect 214340 207012 215944 207040
rect 214340 207000 214346 207012
rect 215938 207000 215944 207012
rect 215996 207000 216002 207052
rect 240318 207000 240324 207052
rect 240376 207040 240382 207052
rect 242158 207040 242164 207052
rect 240376 207012 242164 207040
rect 240376 207000 240382 207012
rect 242158 207000 242164 207012
rect 242216 207000 242222 207052
rect 251174 206592 251180 206644
rect 251232 206632 251238 206644
rect 299474 206632 299480 206644
rect 251232 206604 299480 206632
rect 251232 206592 251238 206604
rect 299474 206592 299480 206604
rect 299532 206592 299538 206644
rect 226426 206524 226432 206576
rect 226484 206564 226490 206576
rect 291838 206564 291844 206576
rect 226484 206536 291844 206564
rect 226484 206524 226490 206536
rect 291838 206524 291844 206536
rect 291896 206524 291902 206576
rect 209038 206456 209044 206508
rect 209096 206496 209102 206508
rect 281258 206496 281264 206508
rect 209096 206468 281264 206496
rect 209096 206456 209102 206468
rect 281258 206456 281264 206468
rect 281316 206456 281322 206508
rect 197998 206388 198004 206440
rect 198056 206428 198062 206440
rect 273346 206428 273352 206440
rect 198056 206400 273352 206428
rect 198056 206388 198062 206400
rect 273346 206388 273352 206400
rect 273404 206388 273410 206440
rect 171042 206320 171048 206372
rect 171100 206360 171106 206372
rect 252646 206360 252652 206372
rect 171100 206332 252652 206360
rect 171100 206320 171106 206332
rect 252646 206320 252652 206332
rect 252704 206320 252710 206372
rect 216858 206252 216864 206304
rect 216916 206292 216922 206304
rect 232498 206292 232504 206304
rect 216916 206264 232504 206292
rect 216916 206252 216922 206264
rect 232498 206252 232504 206264
rect 232556 206252 232562 206304
rect 234430 206252 234436 206304
rect 234488 206292 234494 206304
rect 582742 206292 582748 206304
rect 234488 206264 582748 206292
rect 234488 206252 234494 206264
rect 582742 206252 582748 206264
rect 582800 206252 582806 206304
rect 213822 205640 213828 205692
rect 213880 205680 213886 205692
rect 580166 205680 580172 205692
rect 213880 205652 580172 205680
rect 213880 205640 213886 205652
rect 580166 205640 580172 205652
rect 580224 205640 580230 205692
rect 202782 205164 202788 205216
rect 202840 205204 202846 205216
rect 250622 205204 250628 205216
rect 202840 205176 250628 205204
rect 202840 205164 202846 205176
rect 250622 205164 250628 205176
rect 250680 205164 250686 205216
rect 245562 205096 245568 205148
rect 245620 205136 245626 205148
rect 298738 205136 298744 205148
rect 245620 205108 298744 205136
rect 245620 205096 245626 205108
rect 298738 205096 298744 205108
rect 298796 205096 298802 205148
rect 195238 205028 195244 205080
rect 195296 205068 195302 205080
rect 255498 205068 255504 205080
rect 195296 205040 255504 205068
rect 195296 205028 195302 205040
rect 255498 205028 255504 205040
rect 255556 205028 255562 205080
rect 248506 204960 248512 205012
rect 248564 205000 248570 205012
rect 331214 205000 331220 205012
rect 248564 204972 331220 205000
rect 248564 204960 248570 204972
rect 331214 204960 331220 204972
rect 331272 204960 331278 205012
rect 228910 204892 228916 204944
rect 228968 204932 228974 204944
rect 583202 204932 583208 204944
rect 228968 204904 583208 204932
rect 228968 204892 228974 204904
rect 583202 204892 583208 204904
rect 583260 204892 583266 204944
rect 258718 204824 258724 204876
rect 258776 204864 258782 204876
rect 265526 204864 265532 204876
rect 258776 204836 265532 204864
rect 258776 204824 258782 204836
rect 265526 204824 265532 204836
rect 265584 204824 265590 204876
rect 209038 204348 209044 204400
rect 209096 204388 209102 204400
rect 583386 204388 583392 204400
rect 209096 204360 583392 204388
rect 209096 204348 209102 204360
rect 583386 204348 583392 204360
rect 583444 204348 583450 204400
rect 202046 204280 202052 204332
rect 202104 204320 202110 204332
rect 582466 204320 582472 204332
rect 202104 204292 582472 204320
rect 202104 204280 202110 204292
rect 582466 204280 582472 204292
rect 582524 204280 582530 204332
rect 247310 203600 247316 203652
rect 247368 203640 247374 203652
rect 294598 203640 294604 203652
rect 247368 203612 294604 203640
rect 247368 203600 247374 203612
rect 294598 203600 294604 203612
rect 294656 203600 294662 203652
rect 210418 203532 210424 203584
rect 210476 203572 210482 203584
rect 270770 203572 270776 203584
rect 210476 203544 270776 203572
rect 210476 203532 210482 203544
rect 270770 203532 270776 203544
rect 270828 203532 270834 203584
rect 289078 203232 289084 203244
rect 282886 203204 289084 203232
rect 159358 203124 159364 203176
rect 159416 203164 159422 203176
rect 282886 203164 282914 203204
rect 289078 203192 289084 203204
rect 289136 203192 289142 203244
rect 159416 203136 282914 203164
rect 159416 203124 159422 203136
rect 283834 203124 283840 203176
rect 283892 203164 283898 203176
rect 285674 203164 285680 203176
rect 283892 203136 285680 203164
rect 283892 203124 283898 203136
rect 285674 203124 285680 203136
rect 285732 203124 285738 203176
rect 207290 203056 207296 203108
rect 207348 203096 207354 203108
rect 583018 203096 583024 203108
rect 207348 203068 583024 203096
rect 207348 203056 207354 203068
rect 583018 203056 583024 203068
rect 583076 203056 583082 203108
rect 205542 202988 205548 203040
rect 205600 203028 205606 203040
rect 582650 203028 582656 203040
rect 205600 203000 582656 203028
rect 205600 202988 205606 203000
rect 582650 202988 582656 203000
rect 582708 202988 582714 203040
rect 202966 202920 202972 202972
rect 203024 202960 203030 202972
rect 583570 202960 583576 202972
rect 203024 202932 583576 202960
rect 203024 202920 203030 202932
rect 583570 202920 583576 202932
rect 583628 202920 583634 202972
rect 201218 202852 201224 202904
rect 201276 202892 201282 202904
rect 583846 202892 583852 202904
rect 201276 202864 583852 202892
rect 201276 202852 201282 202864
rect 583846 202852 583852 202864
rect 583904 202852 583910 202904
rect 228174 202784 228180 202836
rect 228232 202824 228238 202836
rect 229002 202824 229008 202836
rect 228232 202796 229008 202824
rect 228232 202784 228238 202796
rect 229002 202784 229008 202796
rect 229060 202784 229066 202836
rect 235166 202444 235172 202496
rect 235224 202484 235230 202496
rect 235902 202484 235908 202496
rect 235224 202456 235908 202484
rect 235224 202444 235230 202456
rect 235902 202444 235908 202456
rect 235960 202444 235966 202496
rect 233418 202308 233424 202360
rect 233476 202348 233482 202360
rect 234522 202348 234528 202360
rect 233476 202320 234528 202348
rect 233476 202308 233482 202320
rect 234522 202308 234528 202320
rect 234580 202308 234586 202360
rect 230750 202240 230756 202292
rect 230808 202280 230814 202292
rect 231762 202280 231768 202292
rect 230808 202252 231768 202280
rect 230808 202240 230814 202252
rect 231762 202240 231768 202252
rect 231820 202240 231826 202292
rect 218606 202104 218612 202156
rect 218664 202144 218670 202156
rect 582374 202144 582380 202156
rect 218664 202116 582380 202144
rect 218664 202104 218670 202116
rect 582374 202104 582380 202116
rect 582432 202104 582438 202156
rect 251634 201968 251640 202020
rect 251692 202008 251698 202020
rect 252462 202008 252468 202020
rect 251692 201980 252468 202008
rect 251692 201968 251698 201980
rect 252462 201968 252468 201980
rect 252520 201968 252526 202020
rect 208210 201900 208216 201952
rect 208268 201940 208274 201952
rect 583202 201940 583208 201952
rect 208268 201912 583208 201940
rect 208268 201900 208274 201912
rect 583202 201900 583208 201912
rect 583260 201900 583266 201952
rect 140038 201832 140044 201884
rect 140096 201872 140102 201884
rect 295978 201872 295984 201884
rect 140096 201844 295984 201872
rect 140096 201832 140102 201844
rect 295978 201832 295984 201844
rect 296036 201832 296042 201884
rect 98638 201764 98644 201816
rect 98696 201804 98702 201816
rect 298646 201804 298652 201816
rect 98696 201776 298652 201804
rect 98696 201764 98702 201776
rect 298646 201764 298652 201776
rect 298704 201764 298710 201816
rect 14458 201696 14464 201748
rect 14516 201736 14522 201748
rect 292482 201736 292488 201748
rect 14516 201708 292488 201736
rect 14516 201696 14522 201708
rect 292482 201696 292488 201708
rect 292540 201696 292546 201748
rect 3234 201628 3240 201680
rect 3292 201668 3298 201680
rect 288158 201668 288164 201680
rect 3292 201640 288164 201668
rect 3292 201628 3298 201640
rect 288158 201628 288164 201640
rect 288216 201628 288222 201680
rect 209866 201560 209872 201612
rect 209924 201600 209930 201612
rect 583294 201600 583300 201612
rect 209924 201572 583300 201600
rect 209924 201560 209930 201572
rect 583294 201560 583300 201572
rect 583352 201560 583358 201612
rect 212534 201492 212540 201544
rect 212592 201532 212598 201544
rect 219342 201532 219348 201544
rect 212592 201504 219348 201532
rect 212592 201492 212598 201504
rect 219342 201492 219348 201504
rect 219400 201492 219406 201544
rect 219434 201492 219440 201544
rect 219492 201532 219498 201544
rect 220630 201532 220636 201544
rect 219492 201504 220636 201532
rect 219492 201492 219498 201504
rect 220630 201492 220636 201504
rect 220688 201492 220694 201544
rect 221182 201424 221188 201476
rect 221240 201464 221246 201476
rect 222102 201464 222108 201476
rect 221240 201436 222108 201464
rect 221240 201424 221246 201436
rect 222102 201424 222108 201436
rect 222160 201424 222166 201476
rect 249886 201356 249892 201408
rect 249944 201396 249950 201408
rect 251174 201396 251180 201408
rect 249944 201368 251180 201396
rect 249944 201356 249950 201368
rect 251174 201356 251180 201368
rect 251232 201356 251238 201408
rect 3418 200812 3424 200864
rect 3476 200852 3482 200864
rect 290826 200852 290832 200864
rect 3476 200824 290832 200852
rect 3476 200812 3482 200824
rect 290826 200812 290832 200824
rect 290884 200812 290890 200864
rect 219342 200744 219348 200796
rect 219400 200784 219406 200796
rect 580258 200784 580264 200796
rect 219400 200756 580264 200784
rect 219400 200744 219406 200756
rect 580258 200744 580264 200756
rect 580316 200744 580322 200796
rect 211614 200404 211620 200456
rect 211672 200444 211678 200456
rect 304258 200444 304264 200456
rect 211672 200416 304264 200444
rect 211672 200404 211678 200416
rect 304258 200404 304264 200416
rect 304316 200404 304322 200456
rect 157242 200336 157248 200388
rect 157300 200376 157306 200388
rect 299474 200376 299480 200388
rect 157300 200348 299480 200376
rect 157300 200336 157306 200348
rect 299474 200336 299480 200348
rect 299532 200336 299538 200388
rect 133138 200268 133144 200320
rect 133196 200308 133202 200320
rect 297726 200308 297732 200320
rect 133196 200280 297732 200308
rect 133196 200268 133202 200280
rect 297726 200268 297732 200280
rect 297784 200268 297790 200320
rect 36538 200200 36544 200252
rect 36596 200240 36602 200252
rect 293402 200240 293408 200252
rect 36596 200212 293408 200240
rect 36596 200200 36602 200212
rect 293402 200200 293408 200212
rect 293460 200200 293466 200252
rect 204714 200132 204720 200184
rect 204772 200172 204778 200184
rect 583662 200172 583668 200184
rect 204772 200144 583668 200172
rect 204772 200132 204778 200144
rect 583662 200132 583668 200144
rect 583720 200132 583726 200184
rect 287606 199860 287612 199912
rect 287664 199900 287670 199912
rect 294782 199900 294788 199912
rect 287664 199872 294788 199900
rect 287664 199860 287670 199872
rect 294782 199860 294788 199872
rect 294840 199860 294846 199912
rect 206738 199792 206744 199844
rect 206796 199832 206802 199844
rect 210418 199832 210424 199844
rect 206796 199804 210424 199832
rect 206796 199792 206802 199804
rect 210418 199792 210424 199804
rect 210476 199792 210482 199844
rect 293144 199804 298094 199832
rect 199930 199724 199936 199776
rect 199988 199764 199994 199776
rect 213178 199764 213184 199776
rect 199988 199736 213184 199764
rect 199988 199724 199994 199736
rect 213178 199724 213184 199736
rect 213236 199724 213242 199776
rect 244182 199724 244188 199776
rect 244240 199764 244246 199776
rect 249242 199764 249248 199776
rect 244240 199736 249248 199764
rect 244240 199724 244246 199736
rect 249242 199724 249248 199736
rect 249300 199724 249306 199776
rect 289630 199764 289636 199776
rect 287164 199736 289636 199764
rect 200022 199656 200028 199708
rect 200080 199696 200086 199708
rect 203518 199696 203524 199708
rect 200080 199668 203524 199696
rect 200080 199656 200086 199668
rect 203518 199656 203524 199668
rect 203576 199656 203582 199708
rect 203702 199656 203708 199708
rect 203760 199696 203766 199708
rect 213270 199696 213276 199708
rect 203760 199668 213276 199696
rect 203760 199656 203766 199668
rect 213270 199656 213276 199668
rect 213328 199656 213334 199708
rect 246298 199696 246304 199708
rect 238726 199668 246304 199696
rect 215018 199628 215024 199640
rect 197326 199600 215024 199628
rect 197326 199288 197354 199600
rect 215018 199588 215024 199600
rect 215076 199588 215082 199640
rect 199378 199520 199384 199572
rect 199436 199560 199442 199572
rect 199436 199532 215294 199560
rect 199436 199520 199442 199532
rect 203702 199492 203708 199504
rect 195946 199260 197354 199288
rect 202846 199464 203708 199492
rect 157978 199044 157984 199096
rect 158036 199084 158042 199096
rect 195946 199084 195974 199260
rect 202846 199084 202874 199464
rect 203702 199452 203708 199464
rect 203760 199452 203766 199504
rect 204070 199452 204076 199504
rect 204128 199492 204134 199504
rect 207658 199492 207664 199504
rect 204128 199464 207664 199492
rect 204128 199452 204134 199464
rect 207658 199452 207664 199464
rect 207716 199452 207722 199504
rect 210326 199452 210332 199504
rect 210384 199452 210390 199504
rect 210418 199452 210424 199504
rect 210476 199452 210482 199504
rect 210510 199452 210516 199504
rect 210568 199492 210574 199504
rect 210568 199464 210648 199492
rect 210568 199452 210574 199464
rect 158036 199056 195974 199084
rect 200408 199056 202874 199084
rect 158036 199044 158042 199056
rect 148318 198976 148324 199028
rect 148376 199016 148382 199028
rect 200408 199016 200436 199056
rect 148376 198988 200436 199016
rect 148376 198976 148382 198988
rect 106918 198908 106924 198960
rect 106976 198948 106982 198960
rect 199930 198948 199936 198960
rect 106976 198920 199936 198948
rect 106976 198908 106982 198920
rect 199930 198908 199936 198920
rect 199988 198908 199994 198960
rect 47578 198772 47584 198824
rect 47636 198812 47642 198824
rect 199838 198812 199844 198824
rect 47636 198784 199844 198812
rect 47636 198772 47642 198784
rect 199838 198772 199844 198784
rect 199896 198772 199902 198824
rect 183002 198704 183008 198756
rect 183060 198744 183066 198756
rect 197998 198744 198004 198756
rect 183060 198716 198004 198744
rect 183060 198704 183066 198716
rect 197998 198704 198004 198716
rect 198056 198704 198062 198756
rect 210344 198268 210372 199452
rect 197326 198240 210372 198268
rect 35158 198092 35164 198144
rect 35216 198132 35222 198144
rect 35216 198104 195974 198132
rect 35216 198092 35222 198104
rect 195946 197996 195974 198104
rect 197326 197996 197354 198240
rect 195946 197968 197354 197996
rect 210436 197860 210464 199452
rect 210620 198404 210648 199464
rect 211154 199452 211160 199504
rect 211212 199452 211218 199504
rect 211246 199452 211252 199504
rect 211304 199452 211310 199504
rect 213178 199452 213184 199504
rect 213236 199452 213242 199504
rect 213270 199452 213276 199504
rect 213328 199452 213334 199504
rect 215018 199452 215024 199504
rect 215076 199492 215082 199504
rect 215076 199464 215156 199492
rect 215076 199452 215082 199464
rect 211172 198540 211200 199452
rect 211264 198880 211292 199452
rect 213196 198948 213224 199452
rect 213288 199016 213316 199452
rect 215128 199152 215156 199464
rect 215266 199220 215294 199532
rect 238018 199452 238024 199504
rect 238076 199452 238082 199504
rect 238036 199288 238064 199452
rect 238726 199288 238754 199668
rect 246298 199656 246304 199668
rect 246356 199656 246362 199708
rect 238036 199260 238754 199288
rect 244016 199600 252554 199628
rect 244016 199220 244044 199600
rect 215266 199192 218054 199220
rect 218026 199152 218054 199192
rect 234586 199192 244044 199220
rect 244108 199532 249380 199560
rect 234586 199152 234614 199192
rect 215128 199124 215340 199152
rect 218026 199124 234614 199152
rect 215312 199084 215340 199124
rect 244108 199084 244136 199532
rect 244182 199452 244188 199504
rect 244240 199452 244246 199504
rect 246206 199452 246212 199504
rect 246264 199452 246270 199504
rect 246298 199452 246304 199504
rect 246356 199452 246362 199504
rect 246482 199452 246488 199504
rect 246540 199452 246546 199504
rect 249242 199452 249248 199504
rect 249300 199452 249306 199504
rect 215312 199056 244136 199084
rect 244200 199016 244228 199452
rect 213288 198988 244228 199016
rect 246224 198948 246252 199452
rect 213196 198920 234614 198948
rect 234586 198880 234614 198920
rect 238128 198920 246252 198948
rect 238128 198880 238156 198920
rect 246316 198880 246344 199452
rect 246500 198948 246528 199452
rect 249260 199288 249288 199452
rect 249168 199260 249288 199288
rect 249168 199016 249196 199260
rect 249352 199084 249380 199532
rect 252526 199492 252554 199600
rect 287054 199560 287060 199572
rect 283116 199532 287060 199560
rect 283116 199492 283144 199532
rect 287054 199520 287060 199532
rect 287112 199520 287118 199572
rect 287164 199492 287192 199736
rect 289630 199724 289636 199736
rect 289688 199724 289694 199776
rect 287698 199656 287704 199708
rect 287756 199696 287762 199708
rect 293144 199696 293172 199804
rect 293218 199724 293224 199776
rect 293276 199764 293282 199776
rect 293276 199736 296760 199764
rect 293276 199724 293282 199736
rect 296622 199696 296628 199708
rect 287756 199668 293172 199696
rect 295306 199668 296628 199696
rect 287756 199656 287762 199668
rect 291286 199628 291292 199640
rect 252526 199464 255314 199492
rect 255286 199152 255314 199464
rect 277366 199464 283144 199492
rect 284266 199464 287192 199492
rect 287256 199600 291292 199628
rect 277366 199152 277394 199464
rect 255286 199124 277394 199152
rect 284266 199084 284294 199464
rect 287256 199424 287284 199600
rect 291286 199588 291292 199600
rect 291344 199588 291350 199640
rect 295306 199560 295334 199668
rect 296622 199656 296628 199668
rect 296680 199656 296686 199708
rect 290476 199532 295334 199560
rect 287606 199452 287612 199504
rect 287664 199452 287670 199504
rect 287698 199452 287704 199504
rect 287756 199452 287762 199504
rect 249352 199056 284294 199084
rect 285968 199396 287284 199424
rect 285968 199016 285996 199396
rect 287624 199016 287652 199452
rect 249168 198988 285996 199016
rect 286336 198988 287652 199016
rect 286336 198948 286364 198988
rect 246500 198920 286364 198948
rect 211264 198852 218054 198880
rect 234586 198852 238156 198880
rect 238864 198852 239076 198880
rect 218026 198812 218054 198852
rect 238864 198812 238892 198852
rect 218026 198784 238892 198812
rect 218026 198716 238984 198744
rect 211172 198512 216536 198540
rect 216508 198404 216536 198512
rect 218026 198472 218054 198716
rect 216646 198444 218054 198472
rect 233206 198580 234614 198608
rect 216646 198404 216674 198444
rect 233206 198404 233234 198580
rect 234586 198540 234614 198580
rect 234586 198512 235994 198540
rect 210620 198376 215294 198404
rect 216508 198376 216674 198404
rect 224926 198376 233234 198404
rect 215266 198268 215294 198376
rect 219406 198308 220814 198336
rect 219406 198268 219434 198308
rect 215266 198240 216674 198268
rect 216646 198064 216674 198240
rect 218026 198240 219434 198268
rect 220786 198268 220814 198308
rect 220786 198240 222194 198268
rect 218026 198064 218054 198240
rect 222166 198132 222194 198240
rect 224926 198132 224954 198376
rect 235966 198200 235994 198512
rect 238956 198404 238984 198716
rect 239048 198676 239076 198852
rect 246224 198852 246344 198880
rect 251146 198852 282408 198880
rect 246224 198744 246252 198852
rect 251146 198744 251174 198852
rect 282380 198812 282408 198852
rect 287716 198812 287744 199452
rect 290476 199220 290504 199532
rect 293218 199452 293224 199504
rect 293276 199452 293282 199504
rect 294138 199452 294144 199504
rect 294196 199452 294202 199504
rect 246224 198716 251174 198744
rect 253906 198784 282224 198812
rect 282380 198784 287744 198812
rect 288406 199192 290504 199220
rect 239048 198648 239444 198676
rect 239416 198540 239444 198648
rect 253906 198540 253934 198784
rect 239416 198512 253934 198540
rect 255286 198716 277394 198744
rect 255286 198404 255314 198716
rect 277366 198540 277394 198716
rect 282196 198676 282224 198784
rect 288406 198676 288434 199192
rect 282196 198648 288434 198676
rect 293236 198608 293264 199452
rect 280126 198580 293264 198608
rect 280126 198540 280154 198580
rect 277366 198512 280154 198540
rect 238956 198376 255314 198404
rect 235966 198172 237374 198200
rect 222166 198104 224954 198132
rect 237346 198132 237374 198172
rect 294156 198132 294184 199452
rect 296732 198948 296760 199736
rect 298066 199016 298094 199804
rect 298066 198988 302234 199016
rect 296732 198920 298094 198948
rect 298066 198608 298094 198920
rect 302206 198880 302234 198988
rect 583754 198880 583760 198892
rect 302206 198852 583760 198880
rect 583754 198840 583760 198852
rect 583812 198840 583818 198892
rect 582374 198744 582380 198756
rect 299446 198716 582380 198744
rect 299446 198608 299474 198716
rect 582374 198704 582380 198716
rect 582432 198704 582438 198756
rect 298066 198580 299474 198608
rect 237346 198104 294184 198132
rect 583110 198064 583116 198076
rect 216646 198036 218054 198064
rect 219406 198036 220814 198064
rect 219406 197996 219434 198036
rect 218026 197968 219434 197996
rect 218026 197928 218054 197968
rect 216646 197900 218054 197928
rect 216646 197860 216674 197900
rect 210436 197832 216674 197860
rect 220786 197860 220814 198036
rect 225984 198036 583116 198064
rect 225984 197928 226012 198036
rect 583110 198024 583116 198036
rect 583168 198024 583174 198076
rect 583754 197996 583760 198008
rect 224926 197900 226012 197928
rect 227686 197968 583760 197996
rect 224926 197860 224954 197900
rect 220786 197832 224954 197860
rect 199930 197752 199936 197804
rect 199988 197792 199994 197804
rect 227686 197792 227714 197968
rect 583754 197956 583760 197968
rect 583812 197956 583818 198008
rect 199988 197764 227714 197792
rect 199988 197752 199994 197764
rect 174538 197344 174544 197396
rect 174596 197384 174602 197396
rect 197998 197384 198004 197396
rect 174596 197356 198004 197384
rect 174596 197344 174602 197356
rect 197998 197344 198004 197356
rect 198056 197344 198062 197396
rect 181530 195984 181536 196036
rect 181588 196024 181594 196036
rect 197998 196024 198004 196036
rect 181588 195996 198004 196024
rect 181588 195984 181594 195996
rect 197998 195984 198004 195996
rect 198056 195984 198062 196036
rect 151722 194556 151728 194608
rect 151780 194596 151786 194608
rect 198090 194596 198096 194608
rect 151780 194568 198096 194596
rect 151780 194556 151786 194568
rect 198090 194556 198096 194568
rect 198148 194556 198154 194608
rect 170490 193196 170496 193248
rect 170548 193236 170554 193248
rect 197722 193236 197728 193248
rect 170548 193208 197728 193236
rect 170548 193196 170554 193208
rect 197722 193196 197728 193208
rect 197780 193196 197786 193248
rect 304258 193128 304264 193180
rect 304316 193168 304322 193180
rect 580166 193168 580172 193180
rect 304316 193140 580172 193168
rect 304316 193128 304322 193140
rect 580166 193128 580172 193140
rect 580224 193128 580230 193180
rect 153102 191836 153108 191888
rect 153160 191876 153166 191888
rect 197630 191876 197636 191888
rect 153160 191848 197636 191876
rect 153160 191836 153166 191848
rect 197630 191836 197636 191848
rect 197688 191836 197694 191888
rect 191190 191020 191196 191072
rect 191248 191060 191254 191072
rect 198090 191060 198096 191072
rect 191248 191032 198096 191060
rect 191248 191020 191254 191032
rect 198090 191020 198096 191032
rect 198148 191020 198154 191072
rect 155862 190476 155868 190528
rect 155920 190516 155926 190528
rect 197354 190516 197360 190528
rect 155920 190488 197360 190516
rect 155920 190476 155926 190488
rect 197354 190476 197360 190488
rect 197412 190476 197418 190528
rect 172422 189116 172428 189168
rect 172480 189156 172486 189168
rect 188430 189156 188436 189168
rect 172480 189128 188436 189156
rect 172480 189116 172486 189128
rect 188430 189116 188436 189128
rect 188488 189116 188494 189168
rect 180150 189048 180156 189100
rect 180208 189088 180214 189100
rect 197906 189088 197912 189100
rect 180208 189060 197912 189088
rect 180208 189048 180214 189060
rect 197906 189048 197912 189060
rect 197964 189048 197970 189100
rect 3510 188980 3516 189032
rect 3568 189020 3574 189032
rect 199378 189020 199384 189032
rect 3568 188992 199384 189020
rect 3568 188980 3574 188992
rect 199378 188980 199384 188992
rect 199436 188980 199442 189032
rect 173158 187688 173164 187740
rect 173216 187728 173222 187740
rect 197354 187728 197360 187740
rect 173216 187700 197360 187728
rect 173216 187688 173222 187700
rect 197354 187688 197360 187700
rect 197412 187688 197418 187740
rect 172422 186396 172428 186448
rect 172480 186436 172486 186448
rect 184382 186436 184388 186448
rect 172480 186408 184388 186436
rect 172480 186396 172486 186408
rect 184382 186396 184388 186408
rect 184440 186396 184446 186448
rect 178770 186328 178776 186380
rect 178828 186368 178834 186380
rect 197538 186368 197544 186380
rect 178828 186340 197544 186368
rect 178828 186328 178834 186340
rect 197538 186328 197544 186340
rect 197596 186328 197602 186380
rect 195330 186192 195336 186244
rect 195388 186232 195394 186244
rect 197630 186232 197636 186244
rect 195388 186204 197636 186232
rect 195388 186192 195394 186204
rect 197630 186192 197636 186204
rect 197688 186192 197694 186244
rect 171778 185580 171784 185632
rect 171836 185620 171842 185632
rect 186958 185620 186964 185632
rect 171836 185592 186964 185620
rect 171836 185580 171842 185592
rect 186958 185580 186964 185592
rect 187016 185580 187022 185632
rect 178862 184152 178868 184204
rect 178920 184192 178926 184204
rect 197354 184192 197360 184204
rect 178920 184164 197360 184192
rect 178920 184152 178926 184164
rect 197354 184152 197360 184164
rect 197412 184152 197418 184204
rect 196710 183744 196716 183796
rect 196768 183784 196774 183796
rect 198366 183784 198372 183796
rect 196768 183756 198372 183784
rect 196768 183744 196774 183756
rect 198366 183744 198372 183756
rect 198424 183744 198430 183796
rect 172422 183608 172428 183660
rect 172480 183648 172486 183660
rect 177298 183648 177304 183660
rect 172480 183620 177304 183648
rect 172480 183608 172486 183620
rect 177298 183608 177304 183620
rect 177356 183608 177362 183660
rect 171686 183540 171692 183592
rect 171744 183580 171750 183592
rect 176010 183580 176016 183592
rect 171744 183552 176016 183580
rect 171744 183540 171750 183552
rect 176010 183540 176016 183552
rect 176068 183540 176074 183592
rect 172422 182248 172428 182300
rect 172480 182288 172486 182300
rect 185578 182288 185584 182300
rect 172480 182260 185584 182288
rect 172480 182248 172486 182260
rect 185578 182248 185584 182260
rect 185636 182248 185642 182300
rect 174630 182180 174636 182232
rect 174688 182220 174694 182232
rect 197722 182220 197728 182232
rect 174688 182192 197728 182220
rect 174688 182180 174694 182192
rect 197722 182180 197728 182192
rect 197780 182180 197786 182232
rect 192478 181432 192484 181484
rect 192536 181472 192542 181484
rect 197354 181472 197360 181484
rect 192536 181444 197360 181472
rect 192536 181432 192542 181444
rect 197354 181432 197360 181444
rect 197412 181432 197418 181484
rect 172422 180820 172428 180872
rect 172480 180860 172486 180872
rect 193858 180860 193864 180872
rect 172480 180832 193864 180860
rect 172480 180820 172486 180832
rect 193858 180820 193864 180832
rect 193916 180820 193922 180872
rect 172054 179460 172060 179512
rect 172112 179500 172118 179512
rect 182910 179500 182916 179512
rect 172112 179472 182916 179500
rect 172112 179460 172118 179472
rect 182910 179460 182916 179472
rect 182968 179460 182974 179512
rect 177390 179392 177396 179444
rect 177448 179432 177454 179444
rect 197354 179432 197360 179444
rect 177448 179404 197360 179432
rect 177448 179392 177454 179404
rect 197354 179392 197360 179404
rect 197412 179392 197418 179444
rect 172146 178100 172152 178152
rect 172204 178140 172210 178152
rect 184290 178140 184296 178152
rect 172204 178112 184296 178140
rect 172204 178100 172210 178112
rect 184290 178100 184296 178112
rect 184348 178100 184354 178152
rect 175918 178032 175924 178084
rect 175976 178072 175982 178084
rect 197906 178072 197912 178084
rect 175976 178044 197912 178072
rect 175976 178032 175982 178044
rect 197906 178032 197912 178044
rect 197964 178032 197970 178084
rect 188522 177352 188528 177404
rect 188580 177392 188586 177404
rect 198090 177392 198096 177404
rect 188580 177364 198096 177392
rect 188580 177352 188586 177364
rect 198090 177352 198096 177364
rect 198148 177352 198154 177404
rect 184382 177284 184388 177336
rect 184440 177324 184446 177336
rect 198182 177324 198188 177336
rect 184440 177296 198188 177324
rect 184440 177284 184446 177296
rect 198182 177284 198188 177296
rect 198240 177284 198246 177336
rect 172422 176740 172428 176792
rect 172480 176780 172486 176792
rect 180058 176780 180064 176792
rect 172480 176752 180064 176780
rect 172480 176740 172486 176752
rect 180058 176740 180064 176752
rect 180116 176740 180122 176792
rect 172238 176672 172244 176724
rect 172296 176712 172302 176724
rect 184198 176712 184204 176724
rect 172296 176684 184204 176712
rect 172296 176672 172302 176684
rect 184198 176672 184204 176684
rect 184256 176672 184262 176724
rect 191282 176332 191288 176384
rect 191340 176372 191346 176384
rect 197814 176372 197820 176384
rect 191340 176344 197820 176372
rect 191340 176332 191346 176344
rect 197814 176332 197820 176344
rect 197872 176332 197878 176384
rect 172422 175244 172428 175296
rect 172480 175284 172486 175296
rect 195422 175284 195428 175296
rect 172480 175256 195428 175284
rect 172480 175244 172486 175256
rect 195422 175244 195428 175256
rect 195480 175244 195486 175296
rect 189718 174496 189724 174548
rect 189776 174536 189782 174548
rect 197354 174536 197360 174548
rect 189776 174508 197360 174536
rect 189776 174496 189782 174508
rect 197354 174496 197360 174508
rect 197412 174496 197418 174548
rect 173434 173884 173440 173936
rect 173492 173924 173498 173936
rect 198550 173924 198556 173936
rect 173492 173896 198556 173924
rect 173492 173884 173498 173896
rect 198550 173884 198556 173896
rect 198608 173884 198614 173936
rect 171778 173204 171784 173256
rect 171836 173244 171842 173256
rect 187050 173244 187056 173256
rect 171836 173216 187056 173244
rect 171836 173204 171842 173216
rect 187050 173204 187056 173216
rect 187108 173204 187114 173256
rect 176010 173136 176016 173188
rect 176068 173176 176074 173188
rect 198090 173176 198096 173188
rect 176068 173148 198096 173176
rect 176068 173136 176074 173148
rect 198090 173136 198096 173148
rect 198148 173136 198154 173188
rect 196802 173000 196808 173052
rect 196860 173040 196866 173052
rect 198458 173040 198464 173052
rect 196860 173012 198464 173040
rect 196860 173000 196866 173012
rect 198458 173000 198464 173012
rect 198516 173000 198522 173052
rect 176010 171776 176016 171828
rect 176068 171816 176074 171828
rect 197354 171816 197360 171828
rect 176068 171788 197360 171816
rect 176068 171776 176074 171788
rect 197354 171776 197360 171788
rect 197412 171776 197418 171828
rect 172238 171096 172244 171148
rect 172296 171136 172302 171148
rect 181438 171136 181444 171148
rect 172296 171108 181444 171136
rect 172296 171096 172302 171108
rect 181438 171096 181444 171108
rect 181496 171096 181502 171148
rect 172238 169736 172244 169788
rect 172296 169776 172302 169788
rect 191098 169776 191104 169788
rect 172296 169748 191104 169776
rect 172296 169736 172302 169748
rect 191098 169736 191104 169748
rect 191156 169736 191162 169788
rect 192570 169736 192576 169788
rect 192628 169776 192634 169788
rect 197722 169776 197728 169788
rect 192628 169748 197728 169776
rect 192628 169736 192634 169748
rect 197722 169736 197728 169748
rect 197780 169736 197786 169788
rect 193950 168512 193956 168564
rect 194008 168552 194014 168564
rect 197722 168552 197728 168564
rect 194008 168524 197728 168552
rect 194008 168512 194014 168524
rect 197722 168512 197728 168524
rect 197780 168512 197786 168564
rect 172422 168376 172428 168428
rect 172480 168416 172486 168428
rect 196618 168416 196624 168428
rect 172480 168388 196624 168416
rect 172480 168376 172486 168388
rect 196618 168376 196624 168388
rect 196676 168376 196682 168428
rect 172422 167084 172428 167136
rect 172480 167124 172486 167136
rect 195238 167124 195244 167136
rect 172480 167096 195244 167124
rect 172480 167084 172486 167096
rect 195238 167084 195244 167096
rect 195296 167084 195302 167136
rect 174722 167016 174728 167068
rect 174780 167056 174786 167068
rect 197906 167056 197912 167068
rect 174780 167028 197912 167056
rect 174780 167016 174786 167028
rect 197906 167016 197912 167028
rect 197964 167016 197970 167068
rect 172054 166268 172060 166320
rect 172112 166308 172118 166320
rect 192478 166308 192484 166320
rect 172112 166280 192484 166308
rect 172112 166268 172118 166280
rect 192478 166268 192484 166280
rect 192536 166268 192542 166320
rect 172422 165656 172428 165708
rect 172480 165696 172486 165708
rect 188338 165696 188344 165708
rect 172480 165668 188344 165696
rect 172480 165656 172486 165668
rect 188338 165656 188344 165668
rect 188396 165656 188402 165708
rect 181622 165588 181628 165640
rect 181680 165628 181686 165640
rect 197354 165628 197360 165640
rect 181680 165600 197360 165628
rect 181680 165588 181686 165600
rect 197354 165588 197360 165600
rect 197412 165588 197418 165640
rect 171134 164296 171140 164348
rect 171192 164336 171198 164348
rect 192478 164336 192484 164348
rect 171192 164308 192484 164336
rect 171192 164296 171198 164308
rect 192478 164296 192484 164308
rect 192536 164296 192542 164348
rect 169202 164228 169208 164280
rect 169260 164268 169266 164280
rect 174538 164268 174544 164280
rect 169260 164240 174544 164268
rect 169260 164228 169266 164240
rect 174538 164228 174544 164240
rect 174596 164228 174602 164280
rect 177482 164228 177488 164280
rect 177540 164268 177546 164280
rect 197630 164268 197636 164280
rect 177540 164240 197636 164268
rect 177540 164228 177546 164240
rect 197630 164228 197636 164240
rect 197688 164228 197694 164280
rect 3234 164160 3240 164212
rect 3292 164200 3298 164212
rect 159358 164200 159364 164212
rect 3292 164172 159364 164200
rect 3292 164160 3298 164172
rect 159358 164160 159364 164172
rect 159416 164160 159422 164212
rect 180242 163480 180248 163532
rect 180300 163520 180306 163532
rect 197354 163520 197360 163532
rect 180300 163492 197360 163520
rect 180300 163480 180306 163492
rect 197354 163480 197360 163492
rect 197412 163480 197418 163532
rect 171870 162936 171876 162988
rect 171928 162976 171934 162988
rect 174538 162976 174544 162988
rect 171928 162948 174544 162976
rect 171928 162936 171934 162948
rect 174538 162936 174544 162948
rect 174596 162936 174602 162988
rect 171686 162868 171692 162920
rect 171744 162908 171750 162920
rect 178678 162908 178684 162920
rect 171744 162880 178684 162908
rect 171744 162868 171750 162880
rect 178678 162868 178684 162880
rect 178736 162868 178742 162920
rect 178954 162188 178960 162240
rect 179012 162228 179018 162240
rect 197630 162228 197636 162240
rect 179012 162200 197636 162228
rect 179012 162188 179018 162200
rect 197630 162188 197636 162200
rect 197688 162188 197694 162240
rect 169386 162120 169392 162172
rect 169444 162160 169450 162172
rect 197446 162160 197452 162172
rect 169444 162132 197452 162160
rect 169444 162120 169450 162132
rect 197446 162120 197452 162132
rect 197504 162120 197510 162172
rect 160002 161440 160008 161492
rect 160060 161480 160066 161492
rect 169294 161480 169300 161492
rect 160060 161452 169300 161480
rect 160060 161440 160066 161452
rect 169294 161440 169300 161452
rect 169352 161440 169358 161492
rect 171686 160828 171692 160880
rect 171744 160868 171750 160880
rect 183002 160868 183008 160880
rect 171744 160840 183008 160868
rect 171744 160828 171750 160840
rect 183002 160828 183008 160840
rect 183060 160828 183066 160880
rect 169294 160760 169300 160812
rect 169352 160800 169358 160812
rect 181530 160800 181536 160812
rect 169352 160772 181536 160800
rect 169352 160760 169358 160772
rect 181530 160760 181536 160772
rect 181588 160760 181594 160812
rect 160830 160692 160836 160744
rect 160888 160732 160894 160744
rect 191190 160732 191196 160744
rect 160888 160704 164234 160732
rect 160888 160692 160894 160704
rect 164206 160664 164234 160704
rect 171888 160704 191196 160732
rect 171888 160664 171916 160704
rect 191190 160692 191196 160704
rect 191248 160692 191254 160744
rect 164206 160636 171916 160664
rect 165154 160488 165160 160540
rect 165212 160528 165218 160540
rect 169294 160528 169300 160540
rect 165212 160500 169300 160528
rect 165212 160488 165218 160500
rect 169294 160488 169300 160500
rect 169352 160488 169358 160540
rect 166810 160420 166816 160472
rect 166868 160460 166874 160472
rect 171686 160460 171692 160472
rect 166868 160432 171692 160460
rect 166868 160420 166874 160432
rect 171686 160420 171692 160432
rect 171744 160420 171750 160472
rect 163130 160352 163136 160404
rect 163188 160392 163194 160404
rect 170490 160392 170496 160404
rect 163188 160364 170496 160392
rect 163188 160352 163194 160364
rect 170490 160352 170496 160364
rect 170548 160352 170554 160404
rect 171870 160080 171876 160132
rect 171928 160120 171934 160132
rect 182818 160120 182824 160132
rect 171928 160092 182824 160120
rect 171928 160080 171934 160092
rect 182818 160080 182824 160092
rect 182876 160080 182882 160132
rect 191374 160080 191380 160132
rect 191432 160120 191438 160132
rect 197354 160120 197360 160132
rect 191432 160092 197360 160120
rect 191432 160080 191438 160092
rect 197354 160080 197360 160092
rect 197412 160080 197418 160132
rect 173342 159332 173348 159384
rect 173400 159372 173406 159384
rect 198458 159372 198464 159384
rect 173400 159344 198464 159372
rect 173400 159332 173406 159344
rect 198458 159332 198464 159344
rect 198516 159332 198522 159384
rect 176102 158720 176108 158772
rect 176160 158760 176166 158772
rect 197538 158760 197544 158772
rect 176160 158732 197544 158760
rect 176160 158720 176166 158732
rect 197538 158720 197544 158732
rect 197596 158720 197602 158772
rect 171962 158652 171968 158704
rect 172020 158692 172026 158704
rect 173250 158692 173256 158704
rect 172020 158664 173256 158692
rect 172020 158652 172026 158664
rect 173250 158652 173256 158664
rect 173308 158652 173314 158704
rect 188430 157972 188436 158024
rect 188488 158012 188494 158024
rect 198458 158012 198464 158024
rect 188488 157984 198464 158012
rect 188488 157972 188494 157984
rect 198458 157972 198464 157984
rect 198516 157972 198522 158024
rect 187142 157360 187148 157412
rect 187200 157400 187206 157412
rect 197354 157400 197360 157412
rect 187200 157372 197360 157400
rect 187200 157360 187206 157372
rect 197354 157360 197360 157372
rect 197412 157360 197418 157412
rect 195422 156884 195428 156936
rect 195480 156924 195486 156936
rect 197998 156924 198004 156936
rect 195480 156896 198004 156924
rect 195480 156884 195486 156896
rect 197998 156884 198004 156896
rect 198056 156884 198062 156936
rect 172238 156000 172244 156052
rect 172296 156040 172302 156052
rect 180150 156040 180156 156052
rect 172296 156012 180156 156040
rect 172296 156000 172302 156012
rect 180150 156000 180156 156012
rect 180208 156000 180214 156052
rect 195514 156000 195520 156052
rect 195572 156040 195578 156052
rect 197906 156040 197912 156052
rect 195572 156012 197912 156040
rect 195572 156000 195578 156012
rect 197906 156000 197912 156012
rect 197964 156000 197970 156052
rect 171962 155320 171968 155372
rect 172020 155360 172026 155372
rect 173434 155360 173440 155372
rect 172020 155332 173440 155360
rect 172020 155320 172026 155332
rect 173434 155320 173440 155332
rect 173492 155320 173498 155372
rect 170490 154572 170496 154624
rect 170548 154612 170554 154624
rect 197722 154612 197728 154624
rect 170548 154584 197728 154612
rect 170548 154572 170554 154584
rect 197722 154572 197728 154584
rect 197780 154572 197786 154624
rect 171686 154504 171692 154556
rect 171744 154544 171750 154556
rect 173158 154544 173164 154556
rect 171744 154516 173164 154544
rect 171744 154504 171750 154516
rect 173158 154504 173164 154516
rect 173216 154504 173222 154556
rect 186958 154504 186964 154556
rect 187016 154544 187022 154556
rect 197354 154544 197360 154556
rect 187016 154516 197360 154544
rect 187016 154504 187022 154516
rect 197354 154504 197360 154516
rect 197412 154504 197418 154556
rect 192662 153212 192668 153264
rect 192720 153252 192726 153264
rect 197354 153252 197360 153264
rect 192720 153224 197360 153252
rect 192720 153212 192726 153224
rect 197354 153212 197360 153224
rect 197412 153212 197418 153264
rect 172330 153144 172336 153196
rect 172388 153184 172394 153196
rect 195330 153184 195336 153196
rect 172388 153156 195336 153184
rect 172388 153144 172394 153156
rect 195330 153144 195336 153156
rect 195388 153144 195394 153196
rect 171502 153076 171508 153128
rect 171560 153116 171566 153128
rect 178770 153116 178776 153128
rect 171560 153088 178776 153116
rect 171560 153076 171566 153088
rect 178770 153076 178776 153088
rect 178828 153076 178834 153128
rect 172330 151648 172336 151700
rect 172388 151688 172394 151700
rect 178862 151688 178868 151700
rect 172388 151660 178868 151688
rect 172388 151648 172394 151660
rect 178862 151648 178868 151660
rect 178920 151648 178926 151700
rect 172422 151580 172428 151632
rect 172480 151620 172486 151632
rect 196710 151620 196716 151632
rect 172480 151592 196716 151620
rect 172480 151580 172486 151592
rect 196710 151580 196716 151592
rect 196768 151580 196774 151632
rect 171318 151172 171324 151224
rect 171376 151212 171382 151224
rect 174630 151212 174636 151224
rect 171376 151184 174636 151212
rect 171376 151172 171382 151184
rect 174630 151172 174636 151184
rect 174688 151172 174694 151224
rect 186958 150424 186964 150476
rect 187016 150464 187022 150476
rect 197446 150464 197452 150476
rect 187016 150436 197452 150464
rect 187016 150424 187022 150436
rect 197446 150424 197452 150436
rect 197504 150424 197510 150476
rect 187050 150356 187056 150408
rect 187108 150396 187114 150408
rect 197354 150396 197360 150408
rect 187108 150368 197360 150396
rect 187108 150356 187114 150368
rect 197354 150356 197360 150368
rect 197412 150356 197418 150408
rect 172238 149676 172244 149728
rect 172296 149716 172302 149728
rect 192570 149716 192576 149728
rect 172296 149688 192576 149716
rect 172296 149676 172302 149688
rect 192570 149676 192576 149688
rect 192628 149676 192634 149728
rect 171502 149608 171508 149660
rect 171560 149648 171566 149660
rect 177390 149648 177396 149660
rect 171560 149620 177396 149648
rect 171560 149608 171566 149620
rect 177390 149608 177396 149620
rect 177448 149608 177454 149660
rect 171686 148996 171692 149048
rect 171744 149036 171750 149048
rect 191282 149036 191288 149048
rect 171744 149008 191288 149036
rect 171744 148996 171750 149008
rect 191282 148996 191288 149008
rect 191340 148996 191346 149048
rect 172422 148928 172428 148980
rect 172480 148968 172486 148980
rect 188522 148968 188528 148980
rect 172480 148940 188528 148968
rect 172480 148928 172486 148940
rect 188522 148928 188528 148940
rect 188580 148928 188586 148980
rect 171318 148316 171324 148368
rect 171376 148356 171382 148368
rect 175918 148356 175924 148368
rect 171376 148328 175924 148356
rect 171376 148316 171382 148328
rect 175918 148316 175924 148328
rect 175976 148316 175982 148368
rect 193858 147704 193864 147756
rect 193916 147744 193922 147756
rect 193916 147716 198136 147744
rect 193916 147704 193922 147716
rect 198108 147688 198136 147716
rect 177390 147636 177396 147688
rect 177448 147676 177454 147688
rect 197538 147676 197544 147688
rect 177448 147648 197544 147676
rect 177448 147636 177454 147648
rect 197538 147636 197544 147648
rect 197596 147636 197602 147688
rect 198090 147636 198096 147688
rect 198148 147636 198154 147688
rect 172422 147568 172428 147620
rect 172480 147608 172486 147620
rect 189718 147608 189724 147620
rect 172480 147580 189724 147608
rect 172480 147568 172486 147580
rect 189718 147568 189724 147580
rect 189776 147568 189782 147620
rect 177298 146888 177304 146940
rect 177356 146928 177362 146940
rect 197354 146928 197360 146940
rect 177356 146900 197360 146928
rect 177356 146888 177362 146900
rect 197354 146888 197360 146900
rect 197412 146888 197418 146940
rect 178770 146276 178776 146328
rect 178828 146316 178834 146328
rect 198182 146316 198188 146328
rect 178828 146288 198188 146316
rect 178828 146276 178834 146288
rect 198182 146276 198188 146288
rect 198240 146276 198246 146328
rect 172330 146208 172336 146260
rect 172388 146248 172394 146260
rect 198734 146248 198740 146260
rect 172388 146220 198740 146248
rect 172388 146208 172394 146220
rect 198734 146208 198740 146220
rect 198792 146208 198798 146260
rect 172422 146140 172428 146192
rect 172480 146180 172486 146192
rect 196802 146180 196808 146192
rect 172480 146152 196808 146180
rect 172480 146140 172486 146152
rect 196802 146140 196808 146152
rect 196860 146140 196866 146192
rect 172146 146072 172152 146124
rect 172204 146112 172210 146124
rect 176010 146112 176016 146124
rect 172204 146084 176016 146112
rect 172204 146072 172210 146084
rect 176010 146072 176016 146084
rect 176068 146072 176074 146124
rect 171318 144848 171324 144900
rect 171376 144888 171382 144900
rect 193950 144888 193956 144900
rect 171376 144860 193956 144888
rect 171376 144848 171382 144860
rect 193950 144848 193956 144860
rect 194008 144848 194014 144900
rect 171962 144168 171968 144220
rect 172020 144208 172026 144220
rect 187142 144208 187148 144220
rect 172020 144180 187148 144208
rect 172020 144168 172026 144180
rect 187142 144168 187148 144180
rect 187200 144168 187206 144220
rect 186314 143556 186320 143608
rect 186372 143596 186378 143608
rect 197446 143596 197452 143608
rect 186372 143568 197452 143596
rect 186372 143556 186378 143568
rect 197446 143556 197452 143568
rect 197504 143556 197510 143608
rect 172422 143488 172428 143540
rect 172480 143528 172486 143540
rect 181622 143528 181628 143540
rect 172480 143500 181628 143528
rect 172480 143488 172486 143500
rect 181622 143488 181628 143500
rect 181680 143488 181686 143540
rect 185578 143488 185584 143540
rect 185636 143528 185642 143540
rect 197354 143528 197360 143540
rect 185636 143500 197360 143528
rect 185636 143488 185642 143500
rect 197354 143488 197360 143500
rect 197412 143488 197418 143540
rect 171686 143352 171692 143404
rect 171744 143392 171750 143404
rect 174722 143392 174728 143404
rect 171744 143364 174728 143392
rect 171744 143352 171750 143364
rect 174722 143352 174728 143364
rect 174780 143352 174786 143404
rect 171870 142808 171876 142860
rect 171928 142848 171934 142860
rect 186314 142848 186320 142860
rect 171928 142820 186320 142848
rect 171928 142808 171934 142820
rect 186314 142808 186320 142820
rect 186372 142808 186378 142860
rect 187050 142128 187056 142180
rect 187108 142168 187114 142180
rect 197354 142168 197360 142180
rect 187108 142140 197360 142168
rect 187108 142128 187114 142140
rect 197354 142128 197360 142140
rect 197412 142128 197418 142180
rect 171502 142060 171508 142112
rect 171560 142100 171566 142112
rect 177482 142100 177488 142112
rect 171560 142072 177488 142100
rect 171560 142060 171566 142072
rect 177482 142060 177488 142072
rect 177540 142060 177546 142112
rect 172422 141516 172428 141568
rect 172480 141556 172486 141568
rect 180242 141556 180248 141568
rect 172480 141528 180248 141556
rect 172480 141516 172486 141528
rect 180242 141516 180248 141528
rect 180300 141516 180306 141568
rect 184290 141380 184296 141432
rect 184348 141420 184354 141432
rect 198458 141420 198464 141432
rect 184348 141392 198464 141420
rect 184348 141380 184354 141392
rect 198458 141380 198464 141392
rect 198516 141380 198522 141432
rect 171502 140972 171508 141024
rect 171560 141012 171566 141024
rect 178954 141012 178960 141024
rect 171560 140984 178960 141012
rect 171560 140972 171566 140984
rect 178954 140972 178960 140984
rect 179012 140972 179018 141024
rect 172422 140700 172428 140752
rect 172480 140740 172486 140752
rect 191374 140740 191380 140752
rect 172480 140712 191380 140740
rect 172480 140700 172486 140712
rect 191374 140700 191380 140712
rect 191432 140700 191438 140752
rect 171686 140632 171692 140684
rect 171744 140672 171750 140684
rect 173342 140672 173348 140684
rect 171744 140644 173348 140672
rect 171744 140632 171750 140644
rect 173342 140632 173348 140644
rect 173400 140632 173406 140684
rect 176010 139408 176016 139460
rect 176068 139448 176074 139460
rect 197354 139448 197360 139460
rect 176068 139420 197360 139448
rect 176068 139408 176074 139420
rect 197354 139408 197360 139420
rect 197412 139408 197418 139460
rect 171318 139340 171324 139392
rect 171376 139380 171382 139392
rect 195514 139380 195520 139392
rect 171376 139352 195520 139380
rect 171376 139340 171382 139352
rect 195514 139340 195520 139352
rect 195572 139340 195578 139392
rect 182910 139272 182916 139324
rect 182968 139312 182974 139324
rect 198182 139312 198188 139324
rect 182968 139284 198188 139312
rect 182968 139272 182974 139284
rect 198182 139272 198188 139284
rect 198240 139272 198246 139324
rect 172422 139204 172428 139256
rect 172480 139244 172486 139256
rect 176102 139244 176108 139256
rect 172480 139216 176108 139244
rect 172480 139204 172486 139216
rect 176102 139204 176108 139216
rect 176160 139204 176166 139256
rect 3234 137912 3240 137964
rect 3292 137952 3298 137964
rect 157978 137952 157984 137964
rect 3292 137924 157984 137952
rect 3292 137912 3298 137924
rect 157978 137912 157984 137924
rect 158036 137912 158042 137964
rect 171502 137912 171508 137964
rect 171560 137952 171566 137964
rect 192662 137952 192668 137964
rect 171560 137924 192668 137952
rect 171560 137912 171566 137924
rect 192662 137912 192668 137924
rect 192720 137912 192726 137964
rect 176654 136620 176660 136672
rect 176712 136660 176718 136672
rect 197538 136660 197544 136672
rect 176712 136632 197544 136660
rect 176712 136620 176718 136632
rect 197538 136620 197544 136632
rect 197596 136620 197602 136672
rect 172422 136552 172428 136604
rect 172480 136592 172486 136604
rect 186958 136592 186964 136604
rect 172480 136564 186964 136592
rect 172480 136552 172486 136564
rect 186958 136552 186964 136564
rect 187016 136552 187022 136604
rect 171686 136484 171692 136536
rect 171744 136524 171750 136536
rect 177390 136524 177396 136536
rect 171744 136496 177396 136524
rect 171744 136484 171750 136496
rect 177390 136484 177396 136496
rect 177448 136484 177454 136536
rect 171502 135600 171508 135652
rect 171560 135640 171566 135652
rect 178770 135640 178776 135652
rect 171560 135612 178776 135640
rect 171560 135600 171566 135612
rect 178770 135600 178776 135612
rect 178828 135600 178834 135652
rect 175274 135260 175280 135312
rect 175332 135300 175338 135312
rect 198182 135300 198188 135312
rect 175332 135272 198188 135300
rect 175332 135260 175338 135272
rect 198182 135260 198188 135272
rect 198240 135260 198246 135312
rect 171502 135192 171508 135244
rect 171560 135232 171566 135244
rect 187050 135232 187056 135244
rect 171560 135204 187056 135232
rect 171560 135192 171566 135204
rect 187050 135192 187056 135204
rect 187108 135192 187114 135244
rect 184198 135124 184204 135176
rect 184256 135164 184262 135176
rect 197354 135164 197360 135176
rect 184256 135136 197360 135164
rect 184256 135124 184262 135136
rect 197354 135124 197360 135136
rect 197412 135124 197418 135176
rect 171870 134716 171876 134768
rect 171928 134756 171934 134768
rect 176010 134756 176016 134768
rect 171928 134728 176016 134756
rect 171928 134716 171934 134728
rect 176010 134716 176016 134728
rect 176068 134716 176074 134768
rect 171686 133832 171692 133884
rect 171744 133872 171750 133884
rect 175274 133872 175280 133884
rect 171744 133844 175280 133872
rect 171744 133832 171750 133844
rect 175274 133832 175280 133844
rect 175332 133832 175338 133884
rect 172422 133356 172428 133408
rect 172480 133396 172486 133408
rect 176654 133396 176660 133408
rect 172480 133368 176660 133396
rect 172480 133356 172486 133368
rect 176654 133356 176660 133368
rect 176712 133356 176718 133408
rect 197446 132512 197452 132524
rect 176304 132484 197452 132512
rect 171686 132404 171692 132456
rect 171744 132444 171750 132456
rect 176304 132444 176332 132484
rect 197446 132472 197452 132484
rect 197504 132472 197510 132524
rect 171744 132416 176332 132444
rect 171744 132404 171750 132416
rect 180058 132404 180064 132456
rect 180116 132444 180122 132456
rect 197354 132444 197360 132456
rect 180116 132416 197360 132444
rect 180116 132404 180122 132416
rect 197354 132404 197360 132416
rect 197412 132404 197418 132456
rect 172422 131724 172428 131776
rect 172480 131764 172486 131776
rect 197906 131764 197912 131776
rect 172480 131736 197912 131764
rect 172480 131724 172486 131736
rect 197906 131724 197912 131736
rect 197964 131724 197970 131776
rect 172422 131112 172428 131164
rect 172480 131152 172486 131164
rect 176654 131152 176660 131164
rect 172480 131124 176660 131152
rect 172480 131112 172486 131124
rect 176654 131112 176660 131124
rect 176712 131112 176718 131164
rect 170398 130364 170404 130416
rect 170456 130404 170462 130416
rect 197446 130404 197452 130416
rect 170456 130376 197452 130404
rect 170456 130364 170462 130376
rect 197446 130364 197452 130376
rect 197504 130364 197510 130416
rect 171686 129820 171692 129872
rect 171744 129860 171750 129872
rect 175918 129860 175924 129872
rect 171744 129832 175924 129860
rect 171744 129820 171750 129832
rect 175918 129820 175924 129832
rect 175976 129820 175982 129872
rect 172054 129752 172060 129804
rect 172112 129792 172118 129804
rect 186314 129792 186320 129804
rect 172112 129764 186320 129792
rect 172112 129752 172118 129764
rect 186314 129752 186320 129764
rect 186372 129752 186378 129804
rect 176654 129684 176660 129736
rect 176712 129724 176718 129736
rect 197354 129724 197360 129736
rect 176712 129696 197360 129724
rect 176712 129684 176718 129696
rect 197354 129684 197360 129696
rect 197412 129684 197418 129736
rect 172422 128392 172428 128444
rect 172480 128432 172486 128444
rect 177298 128432 177304 128444
rect 172480 128404 177304 128432
rect 172480 128392 172486 128404
rect 177298 128392 177304 128404
rect 177356 128392 177362 128444
rect 171594 128324 171600 128376
rect 171652 128364 171658 128376
rect 180150 128364 180156 128376
rect 171652 128336 180156 128364
rect 171652 128324 171658 128336
rect 180150 128324 180156 128336
rect 180208 128324 180214 128376
rect 173250 128256 173256 128308
rect 173308 128296 173314 128308
rect 198090 128296 198096 128308
rect 173308 128268 198096 128296
rect 173308 128256 173314 128268
rect 198090 128256 198096 128268
rect 198148 128256 198154 128308
rect 178678 127576 178684 127628
rect 178736 127616 178742 127628
rect 197998 127616 198004 127628
rect 178736 127588 198004 127616
rect 178736 127576 178742 127588
rect 197998 127576 198004 127588
rect 198056 127576 198062 127628
rect 172054 127032 172060 127084
rect 172112 127072 172118 127084
rect 173158 127072 173164 127084
rect 172112 127044 173164 127072
rect 172112 127032 172118 127044
rect 173158 127032 173164 127044
rect 173216 127032 173222 127084
rect 171686 126964 171692 127016
rect 171744 127004 171750 127016
rect 178034 127004 178040 127016
rect 171744 126976 178040 127004
rect 171744 126964 171750 126976
rect 178034 126964 178040 126976
rect 178092 126964 178098 127016
rect 175918 126896 175924 126948
rect 175976 126936 175982 126948
rect 197354 126936 197360 126948
rect 175976 126908 197360 126936
rect 175976 126896 175982 126908
rect 197354 126896 197360 126908
rect 197412 126896 197418 126948
rect 181438 126216 181444 126268
rect 181496 126256 181502 126268
rect 197906 126256 197912 126268
rect 181496 126228 197912 126256
rect 181496 126216 181502 126228
rect 197906 126216 197912 126228
rect 197964 126216 197970 126268
rect 172422 125672 172428 125724
rect 172480 125712 172486 125724
rect 181530 125712 181536 125724
rect 172480 125684 181536 125712
rect 172480 125672 172486 125684
rect 181530 125672 181536 125684
rect 181588 125672 181594 125724
rect 172146 125604 172152 125656
rect 172204 125644 172210 125656
rect 184198 125644 184204 125656
rect 172204 125616 184204 125644
rect 172204 125604 172210 125616
rect 184198 125604 184204 125616
rect 184256 125604 184262 125656
rect 186314 125536 186320 125588
rect 186372 125576 186378 125588
rect 197630 125576 197636 125588
rect 186372 125548 197636 125576
rect 186372 125536 186378 125548
rect 197630 125536 197636 125548
rect 197688 125536 197694 125588
rect 172330 124856 172336 124908
rect 172388 124896 172394 124908
rect 186958 124896 186964 124908
rect 172388 124868 186964 124896
rect 172388 124856 172394 124868
rect 186958 124856 186964 124868
rect 187016 124856 187022 124908
rect 171870 124312 171876 124364
rect 171928 124352 171934 124364
rect 180058 124352 180064 124364
rect 171928 124324 180064 124352
rect 171928 124312 171934 124324
rect 180058 124312 180064 124324
rect 180116 124312 180122 124364
rect 171686 124244 171692 124296
rect 171744 124284 171750 124296
rect 178678 124284 178684 124296
rect 171744 124256 178684 124284
rect 171744 124244 171750 124256
rect 178678 124244 178684 124256
rect 178736 124244 178742 124296
rect 172422 124176 172428 124228
rect 172480 124216 172486 124228
rect 175918 124216 175924 124228
rect 172480 124188 175924 124216
rect 172480 124176 172486 124188
rect 175918 124176 175924 124188
rect 175976 124176 175982 124228
rect 155862 124108 155868 124160
rect 155920 124148 155926 124160
rect 160646 124148 160652 124160
rect 155920 124120 160652 124148
rect 155920 124108 155926 124120
rect 160646 124108 160652 124120
rect 160704 124108 160710 124160
rect 178034 123428 178040 123480
rect 178092 123468 178098 123480
rect 197630 123468 197636 123480
rect 178092 123440 197636 123468
rect 178092 123428 178098 123440
rect 197630 123428 197636 123440
rect 197688 123428 197694 123480
rect 153102 122816 153108 122868
rect 153160 122856 153166 122868
rect 162854 122856 162860 122868
rect 153160 122828 162860 122856
rect 153160 122816 153166 122828
rect 162854 122816 162860 122828
rect 162912 122816 162918 122868
rect 151722 122748 151728 122800
rect 151780 122788 151786 122800
rect 164878 122788 164884 122800
rect 151780 122760 164884 122788
rect 151780 122748 151786 122760
rect 164878 122748 164884 122760
rect 164936 122748 164942 122800
rect 168926 122748 168932 122800
rect 168984 122788 168990 122800
rect 198826 122788 198832 122800
rect 168984 122760 198832 122788
rect 168984 122748 168990 122760
rect 198826 122748 198832 122760
rect 198884 122748 198890 122800
rect 157242 122680 157248 122732
rect 157300 122720 157306 122732
rect 166902 122720 166908 122732
rect 157300 122692 166908 122720
rect 157300 122680 157306 122692
rect 166902 122680 166908 122692
rect 166960 122680 166966 122732
rect 170398 122680 170404 122732
rect 170456 122720 170462 122732
rect 197354 122720 197360 122732
rect 170456 122692 197360 122720
rect 170456 122680 170462 122692
rect 197354 122680 197360 122692
rect 197412 122680 197418 122732
rect 180150 121388 180156 121440
rect 180208 121428 180214 121440
rect 197538 121428 197544 121440
rect 180208 121400 197544 121428
rect 180208 121388 180214 121400
rect 197538 121388 197544 121400
rect 197596 121388 197602 121440
rect 191098 121320 191104 121372
rect 191156 121360 191162 121372
rect 197354 121360 197360 121372
rect 191156 121332 197360 121360
rect 191156 121320 191162 121332
rect 197354 121320 197360 121332
rect 197412 121320 197418 121372
rect 171778 120708 171784 120760
rect 171836 120748 171842 120760
rect 191742 120748 191748 120760
rect 171836 120720 191748 120748
rect 171836 120708 171842 120720
rect 191742 120708 191748 120720
rect 191800 120708 191806 120760
rect 191742 119960 191748 120012
rect 191800 120000 191806 120012
rect 198274 120000 198280 120012
rect 191800 119972 198280 120000
rect 191800 119960 191806 119972
rect 198274 119960 198280 119972
rect 198332 119960 198338 120012
rect 177298 118600 177304 118652
rect 177356 118640 177362 118652
rect 197354 118640 197360 118652
rect 177356 118612 197360 118640
rect 177356 118600 177362 118612
rect 197354 118600 197360 118612
rect 197412 118600 197418 118652
rect 196618 117172 196624 117224
rect 196676 117212 196682 117224
rect 198458 117212 198464 117224
rect 196676 117184 198464 117212
rect 196676 117172 196682 117184
rect 198458 117172 198464 117184
rect 198516 117172 198522 117224
rect 195238 114860 195244 114912
rect 195296 114900 195302 114912
rect 197906 114900 197912 114912
rect 195296 114872 197912 114900
rect 195296 114860 195302 114872
rect 197906 114860 197912 114872
rect 197964 114860 197970 114912
rect 173158 114452 173164 114504
rect 173216 114492 173222 114504
rect 197354 114492 197360 114504
rect 173216 114464 197360 114492
rect 173216 114452 173222 114464
rect 197354 114452 197360 114464
rect 197412 114452 197418 114504
rect 188338 113092 188344 113144
rect 188396 113132 188402 113144
rect 197354 113132 197360 113144
rect 188396 113104 197360 113132
rect 188396 113092 188402 113104
rect 197354 113092 197360 113104
rect 197412 113092 197418 113144
rect 3418 111732 3424 111784
rect 3476 111772 3482 111784
rect 148318 111772 148324 111784
rect 3476 111744 148324 111772
rect 3476 111732 3482 111744
rect 148318 111732 148324 111744
rect 148376 111732 148382 111784
rect 186958 111732 186964 111784
rect 187016 111772 187022 111784
rect 197354 111772 197360 111784
rect 187016 111744 197360 111772
rect 187016 111732 187022 111744
rect 197354 111732 197360 111744
rect 197412 111732 197418 111784
rect 184198 110372 184204 110424
rect 184256 110412 184262 110424
rect 197538 110412 197544 110424
rect 184256 110384 197544 110412
rect 184256 110372 184262 110384
rect 197538 110372 197544 110384
rect 197596 110372 197602 110424
rect 192478 110304 192484 110356
rect 192536 110344 192542 110356
rect 197354 110344 197360 110356
rect 192536 110316 197360 110344
rect 192536 110304 192542 110316
rect 197354 110304 197360 110316
rect 197412 110304 197418 110356
rect 181530 108264 181536 108316
rect 181588 108304 181594 108316
rect 197538 108304 197544 108316
rect 181588 108276 197544 108304
rect 181588 108264 181594 108276
rect 197538 108264 197544 108276
rect 197596 108264 197602 108316
rect 180058 106904 180064 106956
rect 180116 106944 180122 106956
rect 198090 106944 198096 106956
rect 180116 106916 198096 106944
rect 180116 106904 180122 106916
rect 198090 106904 198096 106916
rect 198148 106904 198154 106956
rect 174538 106224 174544 106276
rect 174596 106264 174602 106276
rect 198550 106264 198556 106276
rect 174596 106236 198556 106264
rect 174596 106224 174602 106236
rect 198550 106224 198556 106236
rect 198608 106224 198614 106276
rect 178678 105544 178684 105596
rect 178736 105584 178742 105596
rect 197446 105584 197452 105596
rect 178736 105556 197452 105584
rect 178736 105544 178742 105556
rect 197446 105544 197452 105556
rect 197504 105544 197510 105596
rect 160002 104796 160008 104848
rect 160060 104836 160066 104848
rect 197538 104836 197544 104848
rect 160060 104808 197544 104836
rect 160060 104796 160066 104808
rect 197538 104796 197544 104808
rect 197596 104796 197602 104848
rect 175918 102756 175924 102808
rect 175976 102796 175982 102808
rect 198090 102796 198096 102808
rect 175976 102768 198096 102796
rect 175976 102756 175982 102768
rect 198090 102756 198096 102768
rect 198148 102756 198154 102808
rect 182818 102076 182824 102128
rect 182876 102116 182882 102128
rect 197906 102116 197912 102128
rect 182876 102088 197912 102116
rect 182876 102076 182882 102088
rect 197906 102076 197912 102088
rect 197964 102076 197970 102128
rect 39298 100716 39304 100768
rect 39356 100756 39362 100768
rect 568574 100756 568580 100768
rect 39356 100728 202276 100756
rect 39356 100716 39362 100728
rect 202248 100700 202276 100728
rect 295536 100728 568580 100756
rect 295536 100700 295564 100728
rect 568574 100716 568580 100728
rect 568632 100716 568638 100768
rect 199930 100648 199936 100700
rect 199988 100688 199994 100700
rect 200574 100688 200580 100700
rect 199988 100660 200580 100688
rect 199988 100648 199994 100660
rect 200574 100648 200580 100660
rect 200632 100648 200638 100700
rect 202230 100648 202236 100700
rect 202288 100648 202294 100700
rect 295518 100648 295524 100700
rect 295576 100648 295582 100700
rect 211522 100104 211528 100156
rect 211580 100144 211586 100156
rect 211706 100144 211712 100156
rect 211580 100116 211712 100144
rect 211580 100104 211586 100116
rect 211706 100104 211712 100116
rect 211764 100104 211770 100156
rect 147582 99764 147588 99816
rect 147640 99804 147646 99816
rect 225138 99804 225144 99816
rect 147640 99776 225144 99804
rect 147640 99764 147646 99776
rect 225138 99764 225144 99776
rect 225196 99764 225202 99816
rect 253198 99764 253204 99816
rect 253256 99804 253262 99816
rect 320174 99804 320180 99816
rect 253256 99776 320180 99804
rect 253256 99764 253262 99776
rect 320174 99764 320180 99776
rect 320232 99764 320238 99816
rect 135162 99696 135168 99748
rect 135220 99736 135226 99748
rect 222838 99736 222844 99748
rect 135220 99708 222844 99736
rect 135220 99696 135226 99708
rect 222838 99696 222844 99708
rect 222896 99696 222902 99748
rect 255682 99696 255688 99748
rect 255740 99736 255746 99748
rect 323578 99736 323584 99748
rect 255740 99708 323584 99736
rect 255740 99696 255746 99708
rect 323578 99696 323584 99708
rect 323636 99696 323642 99748
rect 156598 99628 156604 99680
rect 156656 99668 156662 99680
rect 226058 99668 226064 99680
rect 156656 99640 226064 99668
rect 156656 99628 156662 99640
rect 226058 99628 226064 99640
rect 226116 99628 226122 99680
rect 259914 99628 259920 99680
rect 259972 99668 259978 99680
rect 331858 99668 331864 99680
rect 259972 99640 331864 99668
rect 259972 99628 259978 99640
rect 331858 99628 331864 99640
rect 331916 99628 331922 99680
rect 155862 99560 155868 99612
rect 155920 99600 155926 99612
rect 226610 99600 226616 99612
rect 155920 99572 226616 99600
rect 155920 99560 155926 99572
rect 226610 99560 226616 99572
rect 226668 99560 226674 99612
rect 259270 99560 259276 99612
rect 259328 99600 259334 99612
rect 345014 99600 345020 99612
rect 259328 99572 345020 99600
rect 259328 99560 259334 99572
rect 345014 99560 345020 99572
rect 345072 99560 345078 99612
rect 105538 99492 105544 99544
rect 105596 99532 105602 99544
rect 217962 99532 217968 99544
rect 105596 99504 217968 99532
rect 105596 99492 105602 99504
rect 217962 99492 217968 99504
rect 218020 99492 218026 99544
rect 286686 99492 286692 99544
rect 286744 99532 286750 99544
rect 504358 99532 504364 99544
rect 286744 99504 504364 99532
rect 286744 99492 286750 99504
rect 504358 99492 504364 99504
rect 504416 99492 504422 99544
rect 77202 99424 77208 99476
rect 77260 99464 77266 99476
rect 213086 99464 213092 99476
rect 77260 99436 213092 99464
rect 77260 99424 77266 99436
rect 213086 99424 213092 99436
rect 213144 99424 213150 99476
rect 234982 99424 234988 99476
rect 235040 99424 235046 99476
rect 239214 99424 239220 99476
rect 239272 99424 239278 99476
rect 287882 99424 287888 99476
rect 287940 99464 287946 99476
rect 511994 99464 512000 99476
rect 287940 99436 512000 99464
rect 287940 99424 287946 99436
rect 511994 99424 512000 99436
rect 512052 99424 512058 99476
rect 66162 99356 66168 99408
rect 66220 99396 66226 99408
rect 211246 99396 211252 99408
rect 66220 99368 211252 99396
rect 66220 99356 66226 99368
rect 211246 99356 211252 99368
rect 211304 99356 211310 99408
rect 235000 99272 235028 99424
rect 239232 99272 239260 99424
rect 289078 99356 289084 99408
rect 289136 99396 289142 99408
rect 520366 99396 520372 99408
rect 289136 99368 520372 99396
rect 289136 99356 289142 99368
rect 520366 99356 520372 99368
rect 520424 99356 520430 99408
rect 234982 99220 234988 99272
rect 235040 99220 235046 99272
rect 239214 99220 239220 99272
rect 239272 99220 239278 99272
rect 248322 98948 248328 99000
rect 248380 98988 248386 99000
rect 283374 98988 283380 99000
rect 248380 98960 283380 98988
rect 248380 98948 248386 98960
rect 283374 98948 283380 98960
rect 283432 98948 283438 99000
rect 197262 98880 197268 98932
rect 197320 98920 197326 98932
rect 235534 98920 235540 98932
rect 197320 98892 235540 98920
rect 197320 98880 197326 98892
rect 235534 98880 235540 98892
rect 235592 98880 235598 98932
rect 180058 98812 180064 98864
rect 180116 98852 180122 98864
rect 230658 98852 230664 98864
rect 180116 98824 230664 98852
rect 180116 98812 180122 98824
rect 230658 98812 230664 98824
rect 230716 98812 230722 98864
rect 255038 98812 255044 98864
rect 255096 98852 255102 98864
rect 324406 98852 324412 98864
rect 255096 98824 324412 98852
rect 255096 98812 255102 98824
rect 324406 98812 324412 98824
rect 324464 98812 324470 98864
rect 173158 98744 173164 98796
rect 173216 98784 173222 98796
rect 228910 98784 228916 98796
rect 173216 98756 228916 98784
rect 173216 98744 173222 98756
rect 228910 98744 228916 98756
rect 228968 98744 228974 98796
rect 267826 98744 267832 98796
rect 267884 98784 267890 98796
rect 394694 98784 394700 98796
rect 267884 98756 394700 98784
rect 267884 98744 267890 98756
rect 394694 98744 394700 98756
rect 394752 98744 394758 98796
rect 162118 98676 162124 98728
rect 162176 98716 162182 98728
rect 227622 98716 227628 98728
rect 162176 98688 227628 98716
rect 162176 98676 162182 98688
rect 227622 98676 227628 98688
rect 227680 98676 227686 98728
rect 283650 98676 283656 98728
rect 283708 98716 283714 98728
rect 475378 98716 475384 98728
rect 283708 98688 475384 98716
rect 283708 98676 283714 98688
rect 475378 98676 475384 98688
rect 475436 98676 475442 98728
rect 4798 98608 4804 98660
rect 4856 98648 4862 98660
rect 200298 98648 200304 98660
rect 4856 98620 200304 98648
rect 4856 98608 4862 98620
rect 200298 98608 200304 98620
rect 200356 98608 200362 98660
rect 201402 98608 201408 98660
rect 201460 98648 201466 98660
rect 234338 98648 234344 98660
rect 201460 98620 234344 98648
rect 201460 98608 201466 98620
rect 234338 98608 234344 98620
rect 234396 98608 234402 98660
rect 282454 98608 282460 98660
rect 282512 98648 282518 98660
rect 479518 98648 479524 98660
rect 282512 98620 479524 98648
rect 282512 98608 282518 98620
rect 479518 98608 479524 98620
rect 479576 98608 479582 98660
rect 238938 98268 238944 98320
rect 238996 98308 239002 98320
rect 239398 98308 239404 98320
rect 238996 98280 239404 98308
rect 238996 98268 239002 98280
rect 239398 98268 239404 98280
rect 239456 98268 239462 98320
rect 262858 98132 262864 98184
rect 262916 98172 262922 98184
rect 306374 98172 306380 98184
rect 262916 98144 306380 98172
rect 262916 98132 262922 98144
rect 306374 98132 306380 98144
rect 306432 98132 306438 98184
rect 165522 98064 165528 98116
rect 165580 98104 165586 98116
rect 215294 98104 215300 98116
rect 165580 98076 215300 98104
rect 165580 98064 165586 98076
rect 215294 98064 215300 98076
rect 215352 98064 215358 98116
rect 328454 98104 328460 98116
rect 267706 98076 328460 98104
rect 144822 97996 144828 98048
rect 144880 98036 144886 98048
rect 267706 98036 267734 98076
rect 328454 98064 328460 98076
rect 328512 98064 328518 98116
rect 144880 98008 215294 98036
rect 144880 97996 144886 98008
rect 3418 97928 3424 97980
rect 3476 97968 3482 97980
rect 36538 97968 36544 97980
rect 3476 97940 36544 97968
rect 3476 97928 3482 97940
rect 36538 97928 36544 97940
rect 36596 97928 36602 97980
rect 215266 97968 215294 98008
rect 263612 98008 267734 98036
rect 224586 97968 224592 97980
rect 215266 97940 224592 97968
rect 224586 97928 224592 97940
rect 224644 97928 224650 97980
rect 231210 97928 231216 97980
rect 231268 97968 231274 97980
rect 237374 97968 237380 97980
rect 231268 97940 237380 97968
rect 231268 97928 231274 97940
rect 237374 97928 237380 97940
rect 237432 97928 237438 97980
rect 238662 97928 238668 97980
rect 238720 97968 238726 97980
rect 241422 97968 241428 97980
rect 238720 97940 241428 97968
rect 238720 97928 238726 97940
rect 241422 97928 241428 97940
rect 241480 97928 241486 97980
rect 195330 97860 195336 97912
rect 195388 97900 195394 97912
rect 202138 97900 202144 97912
rect 195388 97872 202144 97900
rect 195388 97860 195394 97872
rect 202138 97860 202144 97872
rect 202196 97860 202202 97912
rect 215294 97792 215300 97844
rect 215352 97832 215358 97844
rect 228266 97832 228272 97844
rect 215352 97804 228272 97832
rect 215352 97792 215358 97804
rect 228266 97792 228272 97804
rect 228324 97792 228330 97844
rect 237374 97792 237380 97844
rect 237432 97832 237438 97844
rect 239030 97832 239036 97844
rect 237432 97804 239036 97832
rect 237432 97792 237438 97804
rect 239030 97792 239036 97804
rect 239088 97792 239094 97844
rect 256418 97792 256424 97844
rect 256476 97832 256482 97844
rect 263612 97832 263640 98008
rect 278774 97996 278780 98048
rect 278832 98036 278838 98048
rect 283558 98036 283564 98048
rect 278832 98008 283564 98036
rect 278832 97996 278838 98008
rect 283558 97996 283564 98008
rect 283616 97996 283622 98048
rect 285766 97996 285772 98048
rect 285824 98036 285830 98048
rect 483014 98036 483020 98048
rect 285824 98008 483020 98036
rect 285824 97996 285830 98008
rect 483014 97996 483020 98008
rect 483072 97996 483078 98048
rect 275738 97860 275744 97912
rect 275796 97900 275802 97912
rect 280706 97900 280712 97912
rect 275796 97872 280712 97900
rect 275796 97860 275802 97872
rect 280706 97860 280712 97872
rect 280764 97860 280770 97912
rect 256476 97804 263640 97832
rect 256476 97792 256482 97804
rect 280982 97792 280988 97844
rect 281040 97832 281046 97844
rect 291654 97832 291660 97844
rect 281040 97804 291660 97832
rect 281040 97792 281046 97804
rect 291654 97792 291660 97804
rect 291712 97792 291718 97844
rect 217318 97724 217324 97776
rect 217376 97764 217382 97776
rect 219710 97764 219716 97776
rect 217376 97736 219716 97764
rect 217376 97724 217382 97736
rect 219710 97724 219716 97736
rect 219768 97724 219774 97776
rect 256878 97724 256884 97776
rect 256936 97764 256942 97776
rect 260190 97764 260196 97776
rect 256936 97736 260196 97764
rect 256936 97724 256942 97736
rect 260190 97724 260196 97736
rect 260248 97724 260254 97776
rect 264974 97724 264980 97776
rect 265032 97764 265038 97776
rect 300578 97764 300584 97776
rect 265032 97736 300584 97764
rect 265032 97724 265038 97736
rect 300578 97724 300584 97736
rect 300636 97724 300642 97776
rect 234522 97656 234528 97708
rect 234580 97696 234586 97708
rect 240226 97696 240232 97708
rect 234580 97668 240232 97696
rect 234580 97656 234586 97668
rect 240226 97656 240232 97668
rect 240284 97656 240290 97708
rect 252646 97656 252652 97708
rect 252704 97696 252710 97708
rect 262858 97696 262864 97708
rect 252704 97668 262864 97696
rect 252704 97656 252710 97668
rect 262858 97656 262864 97668
rect 262916 97656 262922 97708
rect 309870 97696 309876 97708
rect 277366 97668 309876 97696
rect 202138 97588 202144 97640
rect 202196 97628 202202 97640
rect 224034 97628 224040 97640
rect 202196 97600 224040 97628
rect 202196 97588 202202 97600
rect 224034 97588 224040 97600
rect 224092 97588 224098 97640
rect 247310 97588 247316 97640
rect 247368 97628 247374 97640
rect 253198 97628 253204 97640
rect 247368 97600 253204 97628
rect 247368 97588 247374 97600
rect 253198 97588 253204 97600
rect 253256 97588 253262 97640
rect 273070 97588 273076 97640
rect 273128 97628 273134 97640
rect 277366 97628 277394 97668
rect 309870 97656 309876 97668
rect 309928 97656 309934 97708
rect 279326 97628 279332 97640
rect 273128 97600 277394 97628
rect 278424 97600 279332 97628
rect 273128 97588 273134 97600
rect 101398 97520 101404 97572
rect 101456 97560 101462 97572
rect 206186 97560 206192 97572
rect 101456 97532 206192 97560
rect 101456 97520 101462 97532
rect 206186 97520 206192 97532
rect 206244 97520 206250 97572
rect 206462 97520 206468 97572
rect 206520 97560 206526 97572
rect 215478 97560 215484 97572
rect 206520 97532 215484 97560
rect 206520 97520 206526 97532
rect 215478 97520 215484 97532
rect 215536 97520 215542 97572
rect 242710 97520 242716 97572
rect 242768 97560 242774 97572
rect 247678 97560 247684 97572
rect 242768 97532 247684 97560
rect 242768 97520 242774 97532
rect 247678 97520 247684 97532
rect 247736 97520 247742 97572
rect 265342 97520 265348 97572
rect 265400 97560 265406 97572
rect 269758 97560 269764 97572
rect 265400 97532 269764 97560
rect 265400 97520 265406 97532
rect 269758 97520 269764 97532
rect 269816 97520 269822 97572
rect 277118 97520 277124 97572
rect 277176 97560 277182 97572
rect 278424 97560 278452 97600
rect 279326 97588 279332 97600
rect 279384 97588 279390 97640
rect 279418 97588 279424 97640
rect 279476 97628 279482 97640
rect 353938 97628 353944 97640
rect 279476 97600 353944 97628
rect 279476 97588 279482 97600
rect 353938 97588 353944 97600
rect 353996 97588 354002 97640
rect 443638 97560 443644 97572
rect 277176 97532 278452 97560
rect 278792 97532 443644 97560
rect 277176 97520 277182 97532
rect 93118 97452 93124 97504
rect 93176 97492 93182 97504
rect 210234 97492 210240 97504
rect 93176 97464 210240 97492
rect 93176 97452 93182 97464
rect 210234 97452 210240 97464
rect 210292 97452 210298 97504
rect 225874 97492 225880 97504
rect 219406 97464 225880 97492
rect 86310 97384 86316 97436
rect 86368 97424 86374 97436
rect 207934 97424 207940 97436
rect 86368 97396 207940 97424
rect 86368 97384 86374 97396
rect 207934 97384 207940 97396
rect 207992 97384 207998 97436
rect 40678 97316 40684 97368
rect 40736 97356 40742 97368
rect 206646 97356 206652 97368
rect 40736 97328 206652 97356
rect 40736 97316 40742 97328
rect 206646 97316 206652 97328
rect 206704 97316 206710 97368
rect 207658 97316 207664 97368
rect 207716 97356 207722 97368
rect 219406 97356 219434 97464
rect 225874 97452 225880 97464
rect 225932 97452 225938 97504
rect 228450 97452 228456 97504
rect 228508 97492 228514 97504
rect 238202 97492 238208 97504
rect 228508 97464 238208 97492
rect 228508 97452 228514 97464
rect 238202 97452 238208 97464
rect 238260 97452 238266 97504
rect 245746 97452 245752 97504
rect 245804 97492 245810 97504
rect 257338 97492 257344 97504
rect 245804 97464 257344 97492
rect 245804 97452 245810 97464
rect 257338 97452 257344 97464
rect 257396 97452 257402 97504
rect 260282 97452 260288 97504
rect 260340 97492 260346 97504
rect 262858 97492 262864 97504
rect 260340 97464 262864 97492
rect 260340 97452 260346 97464
rect 262858 97452 262864 97464
rect 262916 97452 262922 97504
rect 263778 97452 263784 97504
rect 263836 97492 263842 97504
rect 268378 97492 268384 97504
rect 263836 97464 268384 97492
rect 263836 97452 263842 97464
rect 268378 97452 268384 97464
rect 268436 97452 268442 97504
rect 276750 97452 276756 97504
rect 276808 97492 276814 97504
rect 278792 97492 278820 97532
rect 443638 97520 443644 97532
rect 443696 97520 443702 97572
rect 276808 97464 278820 97492
rect 276808 97452 276814 97464
rect 279786 97452 279792 97504
rect 279844 97492 279850 97504
rect 454678 97492 454684 97504
rect 279844 97464 454684 97492
rect 279844 97452 279850 97464
rect 454678 97452 454684 97464
rect 454736 97452 454742 97504
rect 223482 97384 223488 97436
rect 223540 97424 223546 97436
rect 237006 97424 237012 97436
rect 223540 97396 237012 97424
rect 223540 97384 223546 97396
rect 237006 97384 237012 97396
rect 237064 97384 237070 97436
rect 244458 97384 244464 97436
rect 244516 97424 244522 97436
rect 255958 97424 255964 97436
rect 244516 97396 255964 97424
rect 244516 97384 244522 97396
rect 255958 97384 255964 97396
rect 256016 97384 256022 97436
rect 291654 97384 291660 97436
rect 291712 97424 291718 97436
rect 461578 97424 461584 97436
rect 291712 97396 461584 97424
rect 291712 97384 291718 97396
rect 461578 97384 461584 97396
rect 461636 97384 461642 97436
rect 207716 97328 219434 97356
rect 207716 97316 207722 97328
rect 226058 97316 226064 97368
rect 226116 97356 226122 97368
rect 236178 97356 236184 97368
rect 226116 97328 236184 97356
rect 226116 97316 226122 97328
rect 236178 97316 236184 97328
rect 236236 97316 236242 97368
rect 246298 97316 246304 97368
rect 246356 97356 246362 97368
rect 246356 97328 253244 97356
rect 246356 97316 246362 97328
rect 32398 97248 32404 97300
rect 32456 97288 32462 97300
rect 204898 97288 204904 97300
rect 32456 97260 204904 97288
rect 32456 97248 32462 97260
rect 204898 97248 204904 97260
rect 204956 97248 204962 97300
rect 207474 97248 207480 97300
rect 207532 97288 207538 97300
rect 207750 97288 207756 97300
rect 207532 97260 207756 97288
rect 207532 97248 207538 97260
rect 207750 97248 207756 97260
rect 207808 97248 207814 97300
rect 213730 97248 213736 97300
rect 213788 97288 213794 97300
rect 236822 97288 236828 97300
rect 213788 97260 236828 97288
rect 213788 97248 213794 97260
rect 236822 97248 236828 97260
rect 236880 97248 236886 97300
rect 245102 97248 245108 97300
rect 245160 97288 245166 97300
rect 251818 97288 251824 97300
rect 245160 97260 251824 97288
rect 245160 97248 245166 97260
rect 251818 97248 251824 97260
rect 251876 97248 251882 97300
rect 246114 97180 246120 97232
rect 246172 97220 246178 97232
rect 250438 97220 250444 97232
rect 246172 97192 250444 97220
rect 246172 97180 246178 97192
rect 250438 97180 250444 97192
rect 250496 97180 250502 97232
rect 253216 97220 253244 97328
rect 257890 97316 257896 97368
rect 257948 97356 257954 97368
rect 260282 97356 260288 97368
rect 257948 97328 260288 97356
rect 257948 97316 257954 97328
rect 260282 97316 260288 97328
rect 260340 97316 260346 97368
rect 261110 97316 261116 97368
rect 261168 97356 261174 97368
rect 275278 97356 275284 97368
rect 261168 97328 275284 97356
rect 261168 97316 261174 97328
rect 275278 97316 275284 97328
rect 275336 97316 275342 97368
rect 282362 97316 282368 97368
rect 282420 97356 282426 97368
rect 468478 97356 468484 97368
rect 282420 97328 468484 97356
rect 282420 97316 282426 97328
rect 468478 97316 468484 97328
rect 468536 97316 468542 97368
rect 253842 97248 253848 97300
rect 253900 97288 253906 97300
rect 282178 97288 282184 97300
rect 253900 97260 282184 97288
rect 253900 97248 253906 97260
rect 282178 97248 282184 97260
rect 282236 97248 282242 97300
rect 299658 97248 299664 97300
rect 299716 97288 299722 97300
rect 582926 97288 582932 97300
rect 299716 97260 582932 97288
rect 299716 97248 299722 97260
rect 582926 97248 582932 97260
rect 582984 97248 582990 97300
rect 260006 97220 260012 97232
rect 253216 97192 260012 97220
rect 260006 97180 260012 97192
rect 260064 97180 260070 97232
rect 274726 97180 274732 97232
rect 274784 97220 274790 97232
rect 279418 97220 279424 97232
rect 274784 97192 279424 97220
rect 274784 97180 274790 97192
rect 279418 97180 279424 97192
rect 279476 97180 279482 97232
rect 234890 97112 234896 97164
rect 234948 97152 234954 97164
rect 235166 97152 235172 97164
rect 234948 97124 235172 97152
rect 234948 97112 234954 97124
rect 235166 97112 235172 97124
rect 235224 97112 235230 97164
rect 236638 97112 236644 97164
rect 236696 97152 236702 97164
rect 239582 97152 239588 97164
rect 236696 97124 239588 97152
rect 236696 97112 236702 97124
rect 239582 97112 239588 97124
rect 239640 97112 239646 97164
rect 243262 97112 243268 97164
rect 243320 97152 243326 97164
rect 246298 97152 246304 97164
rect 243320 97124 246304 97152
rect 243320 97112 243326 97124
rect 246298 97112 246304 97124
rect 246356 97112 246362 97164
rect 268010 97112 268016 97164
rect 268068 97152 268074 97164
rect 276750 97152 276756 97164
rect 268068 97124 276756 97152
rect 268068 97112 268074 97124
rect 276750 97112 276756 97124
rect 276808 97112 276814 97164
rect 293402 97112 293408 97164
rect 293460 97152 293466 97164
rect 293862 97152 293868 97164
rect 293460 97124 293868 97152
rect 293460 97112 293466 97124
rect 293862 97112 293868 97124
rect 293920 97112 293926 97164
rect 296070 97112 296076 97164
rect 296128 97152 296134 97164
rect 296438 97152 296444 97164
rect 296128 97124 296444 97152
rect 296128 97112 296134 97124
rect 296438 97112 296444 97124
rect 296496 97112 296502 97164
rect 243446 97044 243452 97096
rect 243504 97084 243510 97096
rect 246390 97084 246396 97096
rect 243504 97056 246396 97084
rect 243504 97044 243510 97056
rect 246390 97044 246396 97056
rect 246448 97044 246454 97096
rect 248966 97044 248972 97096
rect 249024 97084 249030 97096
rect 255774 97084 255780 97096
rect 249024 97056 255780 97084
rect 249024 97044 249030 97056
rect 255774 97044 255780 97056
rect 255832 97044 255838 97096
rect 259546 97044 259552 97096
rect 259604 97084 259610 97096
rect 264238 97084 264244 97096
rect 259604 97056 264244 97084
rect 259604 97044 259610 97056
rect 264238 97044 264244 97056
rect 264296 97044 264302 97096
rect 264606 97044 264612 97096
rect 264664 97084 264670 97096
rect 265894 97084 265900 97096
rect 264664 97056 265900 97084
rect 264664 97044 264670 97056
rect 265894 97044 265900 97056
rect 265952 97044 265958 97096
rect 275370 97044 275376 97096
rect 275428 97084 275434 97096
rect 276658 97084 276664 97096
rect 275428 97056 276664 97084
rect 275428 97044 275434 97056
rect 276658 97044 276664 97056
rect 276716 97044 276722 97096
rect 296254 97044 296260 97096
rect 296312 97084 296318 97096
rect 296622 97084 296628 97096
rect 296312 97056 296628 97084
rect 296312 97044 296318 97056
rect 296622 97044 296628 97056
rect 296680 97044 296686 97096
rect 214558 96976 214564 97028
rect 214616 97016 214622 97028
rect 218146 97016 218152 97028
rect 214616 96988 218152 97016
rect 214616 96976 214622 96988
rect 218146 96976 218152 96988
rect 218204 96976 218210 97028
rect 219802 96976 219808 97028
rect 219860 97016 219866 97028
rect 220630 97016 220636 97028
rect 219860 96988 220636 97016
rect 219860 96976 219866 96988
rect 220630 96976 220636 96988
rect 220688 96976 220694 97028
rect 222286 96976 222292 97028
rect 222344 97016 222350 97028
rect 223114 97016 223120 97028
rect 222344 96988 223120 97016
rect 222344 96976 222350 96988
rect 223114 96976 223120 96988
rect 223172 96976 223178 97028
rect 243906 96976 243912 97028
rect 243964 97016 243970 97028
rect 244182 97016 244188 97028
rect 243964 96988 244188 97016
rect 243964 96976 243970 96988
rect 244182 96976 244188 96988
rect 244240 96976 244246 97028
rect 246758 96976 246764 97028
rect 246816 96976 246822 97028
rect 247126 96976 247132 97028
rect 247184 97016 247190 97028
rect 247184 96988 248414 97016
rect 247184 96976 247190 96988
rect 201954 96908 201960 96960
rect 202012 96948 202018 96960
rect 202598 96948 202604 96960
rect 202012 96920 202604 96948
rect 202012 96908 202018 96920
rect 202598 96908 202604 96920
rect 202656 96908 202662 96960
rect 207750 96908 207756 96960
rect 207808 96948 207814 96960
rect 213638 96948 213644 96960
rect 207808 96920 213644 96948
rect 207808 96908 207814 96920
rect 213638 96908 213644 96920
rect 213696 96908 213702 96960
rect 215386 96908 215392 96960
rect 215444 96948 215450 96960
rect 215938 96948 215944 96960
rect 215444 96920 215944 96948
rect 215444 96908 215450 96920
rect 215938 96908 215944 96920
rect 215996 96908 216002 96960
rect 216858 96908 216864 96960
rect 216916 96948 216922 96960
rect 217502 96948 217508 96960
rect 216916 96920 217508 96948
rect 216916 96908 216922 96920
rect 217502 96908 217508 96920
rect 217560 96908 217566 96960
rect 218238 96908 218244 96960
rect 218296 96948 218302 96960
rect 218606 96948 218612 96960
rect 218296 96920 218612 96948
rect 218296 96908 218302 96920
rect 218606 96908 218612 96920
rect 218664 96908 218670 96960
rect 219894 96908 219900 96960
rect 219952 96948 219958 96960
rect 220262 96948 220268 96960
rect 219952 96920 220268 96948
rect 219952 96908 219958 96920
rect 220262 96908 220268 96920
rect 220320 96908 220326 96960
rect 222654 96908 222660 96960
rect 222712 96948 222718 96960
rect 223298 96948 223304 96960
rect 222712 96920 223304 96948
rect 222712 96908 222718 96920
rect 223298 96908 223304 96920
rect 223356 96908 223362 96960
rect 223666 96908 223672 96960
rect 223724 96948 223730 96960
rect 224678 96948 224684 96960
rect 223724 96920 224684 96948
rect 223724 96908 223730 96920
rect 224678 96908 224684 96920
rect 224736 96908 224742 96960
rect 234706 96908 234712 96960
rect 234764 96948 234770 96960
rect 235626 96948 235632 96960
rect 234764 96920 235632 96948
rect 234764 96908 234770 96920
rect 235626 96908 235632 96920
rect 235684 96908 235690 96960
rect 236270 96908 236276 96960
rect 236328 96948 236334 96960
rect 237098 96948 237104 96960
rect 236328 96920 237104 96948
rect 236328 96908 236334 96920
rect 237098 96908 237104 96920
rect 237156 96908 237162 96960
rect 240502 96908 240508 96960
rect 240560 96948 240566 96960
rect 240962 96948 240968 96960
rect 240560 96920 240968 96948
rect 240560 96908 240566 96920
rect 240962 96908 240968 96920
rect 241020 96908 241026 96960
rect 242066 96908 242072 96960
rect 242124 96948 242130 96960
rect 242526 96948 242532 96960
rect 242124 96920 242532 96948
rect 242124 96908 242130 96920
rect 242526 96908 242532 96920
rect 242584 96908 242590 96960
rect 244918 96908 244924 96960
rect 244976 96948 244982 96960
rect 245470 96948 245476 96960
rect 244976 96920 245476 96948
rect 244976 96908 244982 96920
rect 245470 96908 245476 96920
rect 245528 96908 245534 96960
rect 204254 96840 204260 96892
rect 204312 96880 204318 96892
rect 209406 96880 209412 96892
rect 204312 96852 209412 96880
rect 204312 96840 204318 96852
rect 209406 96840 209412 96852
rect 209464 96840 209470 96892
rect 216766 96840 216772 96892
rect 216824 96880 216830 96892
rect 217594 96880 217600 96892
rect 216824 96852 217600 96880
rect 216824 96840 216830 96852
rect 217594 96840 217600 96852
rect 217652 96840 217658 96892
rect 218422 96840 218428 96892
rect 218480 96880 218486 96892
rect 219250 96880 219256 96892
rect 218480 96852 219256 96880
rect 218480 96840 218486 96852
rect 219250 96840 219256 96852
rect 219308 96840 219314 96892
rect 219618 96840 219624 96892
rect 219676 96880 219682 96892
rect 220078 96880 220084 96892
rect 219676 96852 220084 96880
rect 219676 96840 219682 96852
rect 220078 96840 220084 96852
rect 220136 96840 220142 96892
rect 224218 96840 224224 96892
rect 224276 96880 224282 96892
rect 228634 96880 228640 96892
rect 224276 96852 228640 96880
rect 224276 96840 224282 96852
rect 228634 96840 228640 96852
rect 228692 96840 228698 96892
rect 244274 96840 244280 96892
rect 244332 96880 244338 96892
rect 245378 96880 245384 96892
rect 244332 96852 245384 96880
rect 244332 96840 244338 96852
rect 245378 96840 245384 96852
rect 245436 96840 245442 96892
rect 202598 96772 202604 96824
rect 202656 96812 202662 96824
rect 208210 96812 208216 96824
rect 202656 96784 208216 96812
rect 202656 96772 202662 96784
rect 208210 96772 208216 96784
rect 208268 96772 208274 96824
rect 209222 96772 209228 96824
rect 209280 96812 209286 96824
rect 213822 96812 213828 96824
rect 209280 96784 213828 96812
rect 209280 96772 209286 96784
rect 213822 96772 213828 96784
rect 213880 96772 213886 96824
rect 215294 96812 215300 96824
rect 215266 96772 215300 96812
rect 215352 96772 215358 96824
rect 215938 96772 215944 96824
rect 215996 96812 216002 96824
rect 216950 96812 216956 96824
rect 215996 96784 216956 96812
rect 215996 96772 216002 96784
rect 216950 96772 216956 96784
rect 217008 96772 217014 96824
rect 239122 96772 239128 96824
rect 239180 96812 239186 96824
rect 239950 96812 239956 96824
rect 239180 96784 239956 96812
rect 239180 96772 239186 96784
rect 239950 96772 239956 96784
rect 240008 96772 240014 96824
rect 241882 96772 241888 96824
rect 241940 96812 241946 96824
rect 242618 96812 242624 96824
rect 241940 96784 242624 96812
rect 241940 96772 241946 96784
rect 242618 96772 242624 96784
rect 242676 96772 242682 96824
rect 242894 96772 242900 96824
rect 242952 96812 242958 96824
rect 243814 96812 243820 96824
rect 242952 96784 243820 96812
rect 242952 96772 242958 96784
rect 243814 96772 243820 96784
rect 243872 96772 243878 96824
rect 246776 96812 246804 96976
rect 247770 96908 247776 96960
rect 247828 96948 247834 96960
rect 248138 96948 248144 96960
rect 247828 96920 248144 96948
rect 247828 96908 247834 96920
rect 248138 96908 248144 96920
rect 248196 96908 248202 96960
rect 248386 96948 248414 96988
rect 250806 96976 250812 97028
rect 250864 97016 250870 97028
rect 251082 97016 251088 97028
rect 250864 96988 251088 97016
rect 250864 96976 250870 96988
rect 251082 96976 251088 96988
rect 251140 96976 251146 97028
rect 252186 96976 252192 97028
rect 252244 97016 252250 97028
rect 253290 97016 253296 97028
rect 252244 96988 253296 97016
rect 252244 96976 252250 96988
rect 253290 96976 253296 96988
rect 253348 96976 253354 97028
rect 258258 96976 258264 97028
rect 258316 97016 258322 97028
rect 259270 97016 259276 97028
rect 258316 96988 259276 97016
rect 258316 96976 258322 96988
rect 259270 96976 259276 96988
rect 259328 96976 259334 97028
rect 261294 96976 261300 97028
rect 261352 97016 261358 97028
rect 262950 97016 262956 97028
rect 261352 96988 262956 97016
rect 261352 96976 261358 96988
rect 262950 96976 262956 96988
rect 263008 96976 263014 97028
rect 270862 96976 270868 97028
rect 270920 97016 270926 97028
rect 271506 97016 271512 97028
rect 270920 96988 271512 97016
rect 270920 96976 270926 96988
rect 271506 96976 271512 96988
rect 271564 96976 271570 97028
rect 276106 96976 276112 97028
rect 276164 97016 276170 97028
rect 277302 97016 277308 97028
rect 276164 96988 277308 97016
rect 276164 96976 276170 96988
rect 277302 96976 277308 96988
rect 277360 96976 277366 97028
rect 290734 96976 290740 97028
rect 290792 97016 290798 97028
rect 291102 97016 291108 97028
rect 290792 96988 291108 97016
rect 290792 96976 290798 96988
rect 291102 96976 291108 96988
rect 291160 96976 291166 97028
rect 249058 96948 249064 96960
rect 248386 96920 249064 96948
rect 249058 96908 249064 96920
rect 249116 96908 249122 96960
rect 249150 96908 249156 96960
rect 249208 96948 249214 96960
rect 249702 96948 249708 96960
rect 249208 96920 249708 96948
rect 249208 96908 249214 96920
rect 249702 96908 249708 96920
rect 249760 96908 249766 96960
rect 249978 96908 249984 96960
rect 250036 96948 250042 96960
rect 254578 96948 254584 96960
rect 250036 96920 254584 96948
rect 250036 96908 250042 96920
rect 254578 96908 254584 96920
rect 254636 96908 254642 96960
rect 254670 96908 254676 96960
rect 254728 96948 254734 96960
rect 255038 96948 255044 96960
rect 254728 96920 255044 96948
rect 254728 96908 254734 96920
rect 255038 96908 255044 96920
rect 255096 96908 255102 96960
rect 255866 96908 255872 96960
rect 255924 96948 255930 96960
rect 256510 96948 256516 96960
rect 255924 96920 256516 96948
rect 255924 96908 255930 96920
rect 256510 96908 256516 96920
rect 256568 96908 256574 96960
rect 258534 96908 258540 96960
rect 258592 96948 258598 96960
rect 259086 96948 259092 96960
rect 258592 96920 259092 96948
rect 258592 96908 258598 96920
rect 259086 96908 259092 96920
rect 259144 96908 259150 96960
rect 259730 96908 259736 96960
rect 259788 96948 259794 96960
rect 260742 96948 260748 96960
rect 259788 96920 260748 96948
rect 259788 96908 259794 96920
rect 260742 96908 260748 96920
rect 260800 96908 260806 96960
rect 261662 96908 261668 96960
rect 261720 96948 261726 96960
rect 262122 96948 262128 96960
rect 261720 96920 262128 96948
rect 261720 96908 261726 96920
rect 262122 96908 262128 96920
rect 262180 96908 262186 96960
rect 262582 96908 262588 96960
rect 262640 96948 262646 96960
rect 263502 96948 263508 96960
rect 262640 96920 263508 96948
rect 262640 96908 262646 96920
rect 263502 96908 263508 96920
rect 263560 96908 263566 96960
rect 264146 96908 264152 96960
rect 264204 96948 264210 96960
rect 264698 96948 264704 96960
rect 264204 96920 264704 96948
rect 264204 96908 264210 96920
rect 264698 96908 264704 96920
rect 264756 96908 264762 96960
rect 265618 96908 265624 96960
rect 265676 96948 265682 96960
rect 266078 96948 266084 96960
rect 265676 96920 266084 96948
rect 265676 96908 265682 96920
rect 266078 96908 266084 96920
rect 266136 96908 266142 96960
rect 266630 96908 266636 96960
rect 266688 96948 266694 96960
rect 267366 96948 267372 96960
rect 266688 96920 267372 96948
rect 266688 96908 266694 96920
rect 267366 96908 267372 96920
rect 267424 96908 267430 96960
rect 269482 96908 269488 96960
rect 269540 96948 269546 96960
rect 270402 96948 270408 96960
rect 269540 96920 270408 96948
rect 269540 96908 269546 96920
rect 270402 96908 270408 96920
rect 270460 96908 270466 96960
rect 270678 96908 270684 96960
rect 270736 96948 270742 96960
rect 271414 96948 271420 96960
rect 270736 96920 271420 96948
rect 270736 96908 270742 96920
rect 271414 96908 271420 96920
rect 271472 96908 271478 96960
rect 272242 96908 272248 96960
rect 272300 96948 272306 96960
rect 273070 96948 273076 96960
rect 272300 96920 273076 96948
rect 272300 96908 272306 96920
rect 273070 96908 273076 96920
rect 273128 96908 273134 96960
rect 273898 96908 273904 96960
rect 273956 96948 273962 96960
rect 274542 96948 274548 96960
rect 273956 96920 274548 96948
rect 273956 96908 273962 96920
rect 274542 96908 274548 96920
rect 274600 96908 274606 96960
rect 276566 96908 276572 96960
rect 276624 96948 276630 96960
rect 277118 96948 277124 96960
rect 276624 96920 277124 96948
rect 276624 96908 276630 96920
rect 277118 96908 277124 96920
rect 277176 96908 277182 96960
rect 277762 96908 277768 96960
rect 277820 96948 277826 96960
rect 278406 96948 278412 96960
rect 277820 96920 278412 96948
rect 277820 96908 277826 96920
rect 278406 96908 278412 96920
rect 278464 96908 278470 96960
rect 280154 96908 280160 96960
rect 280212 96948 280218 96960
rect 281350 96948 281356 96960
rect 280212 96920 281356 96948
rect 280212 96908 280218 96920
rect 281350 96908 281356 96920
rect 281408 96908 281414 96960
rect 281810 96908 281816 96960
rect 281868 96948 281874 96960
rect 282454 96948 282460 96960
rect 281868 96920 282460 96948
rect 281868 96908 281874 96920
rect 282454 96908 282460 96920
rect 282512 96908 282518 96960
rect 283190 96908 283196 96960
rect 283248 96948 283254 96960
rect 283834 96948 283840 96960
rect 283248 96920 283840 96948
rect 283248 96908 283254 96920
rect 283834 96908 283840 96920
rect 283892 96908 283898 96960
rect 286318 96908 286324 96960
rect 286376 96948 286382 96960
rect 286686 96948 286692 96960
rect 286376 96920 286692 96948
rect 286376 96908 286382 96920
rect 286686 96908 286692 96920
rect 286744 96908 286750 96960
rect 287514 96908 287520 96960
rect 287572 96948 287578 96960
rect 288066 96948 288072 96960
rect 287572 96920 288072 96948
rect 287572 96908 287578 96920
rect 288066 96908 288072 96920
rect 288124 96908 288130 96960
rect 288710 96908 288716 96960
rect 288768 96948 288774 96960
rect 289446 96948 289452 96960
rect 288768 96920 289452 96948
rect 288768 96908 288774 96920
rect 289446 96908 289452 96920
rect 289504 96908 289510 96960
rect 290090 96908 290096 96960
rect 290148 96948 290154 96960
rect 290826 96948 290832 96960
rect 290148 96920 290832 96948
rect 290148 96908 290154 96920
rect 290826 96908 290832 96920
rect 290884 96908 290890 96960
rect 291746 96908 291752 96960
rect 291804 96948 291810 96960
rect 292482 96948 292488 96960
rect 291804 96920 292488 96948
rect 291804 96908 291810 96920
rect 292482 96908 292488 96920
rect 292540 96908 292546 96960
rect 292758 96908 292764 96960
rect 292816 96948 292822 96960
rect 293494 96948 293500 96960
rect 292816 96920 293500 96948
rect 292816 96908 292822 96920
rect 293494 96908 293500 96920
rect 293552 96908 293558 96960
rect 294598 96908 294604 96960
rect 294656 96948 294662 96960
rect 295058 96948 295064 96960
rect 294656 96920 295064 96948
rect 294656 96908 294662 96920
rect 295058 96908 295064 96920
rect 295116 96908 295122 96960
rect 298830 96908 298836 96960
rect 298888 96948 298894 96960
rect 299382 96948 299388 96960
rect 298888 96920 299388 96948
rect 298888 96908 298894 96920
rect 299382 96908 299388 96920
rect 299440 96908 299446 96960
rect 299842 96908 299848 96960
rect 299900 96948 299906 96960
rect 300762 96948 300768 96960
rect 299900 96920 300768 96948
rect 299900 96908 299906 96920
rect 300762 96908 300768 96920
rect 300820 96908 300826 96960
rect 248782 96840 248788 96892
rect 248840 96880 248846 96892
rect 249610 96880 249616 96892
rect 248840 96852 249616 96880
rect 248840 96840 248846 96852
rect 249610 96840 249616 96852
rect 249668 96840 249674 96892
rect 254026 96840 254032 96892
rect 254084 96880 254090 96892
rect 255130 96880 255136 96892
rect 254084 96852 255136 96880
rect 254084 96840 254090 96852
rect 255130 96840 255136 96852
rect 255188 96840 255194 96892
rect 255406 96840 255412 96892
rect 255464 96880 255470 96892
rect 256602 96880 256608 96892
rect 255464 96852 256608 96880
rect 255464 96840 255470 96852
rect 256602 96840 256608 96852
rect 256660 96840 256666 96892
rect 258718 96840 258724 96892
rect 258776 96880 258782 96892
rect 259178 96880 259184 96892
rect 258776 96852 259184 96880
rect 258776 96840 258782 96852
rect 259178 96840 259184 96852
rect 259236 96840 259242 96892
rect 260098 96840 260104 96892
rect 260156 96880 260162 96892
rect 260650 96880 260656 96892
rect 260156 96852 260656 96880
rect 260156 96840 260162 96852
rect 260650 96840 260656 96852
rect 260708 96840 260714 96892
rect 260926 96840 260932 96892
rect 260984 96880 260990 96892
rect 262030 96880 262036 96892
rect 260984 96852 262036 96880
rect 260984 96840 260990 96852
rect 262030 96840 262036 96852
rect 262088 96840 262094 96892
rect 263134 96840 263140 96892
rect 263192 96840 263198 96892
rect 263962 96840 263968 96892
rect 264020 96880 264026 96892
rect 264790 96880 264796 96892
rect 264020 96852 264796 96880
rect 264020 96840 264026 96852
rect 264790 96840 264796 96852
rect 264848 96840 264854 96892
rect 265802 96840 265808 96892
rect 265860 96880 265866 96892
rect 266262 96880 266268 96892
rect 265860 96852 266268 96880
rect 265860 96840 265866 96852
rect 266262 96840 266268 96852
rect 266320 96840 266326 96892
rect 266814 96840 266820 96892
rect 266872 96880 266878 96892
rect 267550 96880 267556 96892
rect 266872 96852 267556 96880
rect 266872 96840 266878 96852
rect 267550 96840 267556 96852
rect 267608 96840 267614 96892
rect 269666 96840 269672 96892
rect 269724 96880 269730 96892
rect 270310 96880 270316 96892
rect 269724 96852 270316 96880
rect 269724 96840 269730 96852
rect 270310 96840 270316 96852
rect 270368 96840 270374 96892
rect 271046 96840 271052 96892
rect 271104 96880 271110 96892
rect 271598 96880 271604 96892
rect 271104 96852 271604 96880
rect 271104 96840 271110 96852
rect 271598 96840 271604 96852
rect 271656 96840 271662 96892
rect 271874 96840 271880 96892
rect 271932 96880 271938 96892
rect 272978 96880 272984 96892
rect 271932 96852 272984 96880
rect 271932 96840 271938 96852
rect 272978 96840 272984 96852
rect 273036 96840 273042 96892
rect 273254 96840 273260 96892
rect 273312 96880 273318 96892
rect 274082 96880 274088 96892
rect 273312 96852 274088 96880
rect 273312 96840 273318 96852
rect 274082 96840 274088 96852
rect 274140 96840 274146 96892
rect 276382 96840 276388 96892
rect 276440 96880 276446 96892
rect 277210 96880 277216 96892
rect 276440 96852 277216 96880
rect 276440 96840 276446 96852
rect 277210 96840 277216 96852
rect 277268 96840 277274 96892
rect 277946 96840 277952 96892
rect 278004 96880 278010 96892
rect 278682 96880 278688 96892
rect 278004 96852 278688 96880
rect 278004 96840 278010 96852
rect 278682 96840 278688 96852
rect 278740 96840 278746 96892
rect 278958 96840 278964 96892
rect 279016 96880 279022 96892
rect 280062 96880 280068 96892
rect 279016 96852 280068 96880
rect 279016 96840 279022 96852
rect 280062 96840 280068 96852
rect 280120 96840 280126 96892
rect 280798 96840 280804 96892
rect 280856 96880 280862 96892
rect 281258 96880 281264 96892
rect 280856 96852 281264 96880
rect 280856 96840 280862 96852
rect 281258 96840 281264 96852
rect 281316 96840 281322 96892
rect 281994 96840 282000 96892
rect 282052 96880 282058 96892
rect 282638 96880 282644 96892
rect 282052 96852 282644 96880
rect 282052 96840 282058 96852
rect 282638 96840 282644 96852
rect 282696 96840 282702 96892
rect 285674 96840 285680 96892
rect 285732 96880 285738 96892
rect 286778 96880 286784 96892
rect 285732 96852 286784 96880
rect 285732 96840 285738 96852
rect 286778 96840 286784 96852
rect 286836 96840 286842 96892
rect 287054 96840 287060 96892
rect 287112 96880 287118 96892
rect 288158 96880 288164 96892
rect 287112 96852 288164 96880
rect 287112 96840 287118 96852
rect 288158 96840 288164 96852
rect 288216 96840 288222 96892
rect 289906 96840 289912 96892
rect 289964 96880 289970 96892
rect 290734 96880 290740 96892
rect 289964 96852 290740 96880
rect 289964 96840 289970 96852
rect 290734 96840 290740 96852
rect 290792 96840 290798 96892
rect 291930 96840 291936 96892
rect 291988 96880 291994 96892
rect 292298 96880 292304 96892
rect 291988 96852 292304 96880
rect 291988 96840 291994 96852
rect 292298 96840 292304 96852
rect 292356 96840 292362 96892
rect 292942 96840 292948 96892
rect 293000 96880 293006 96892
rect 293586 96880 293592 96892
rect 293000 96852 293592 96880
rect 293000 96840 293006 96852
rect 293586 96840 293592 96852
rect 293644 96840 293650 96892
rect 294230 96840 294236 96892
rect 294288 96880 294294 96892
rect 295150 96880 295156 96892
rect 294288 96852 295156 96880
rect 294288 96840 294294 96852
rect 295150 96840 295156 96852
rect 295208 96840 295214 96892
rect 299474 96840 299480 96892
rect 299532 96880 299538 96892
rect 300670 96880 300676 96892
rect 299532 96852 300676 96880
rect 299532 96840 299538 96852
rect 300670 96840 300676 96852
rect 300728 96840 300734 96892
rect 246942 96812 246948 96824
rect 246776 96784 246948 96812
rect 246942 96772 246948 96784
rect 247000 96772 247006 96824
rect 247494 96772 247500 96824
rect 247552 96812 247558 96824
rect 248230 96812 248236 96824
rect 247552 96784 248236 96812
rect 247552 96772 247558 96784
rect 248230 96772 248236 96784
rect 248288 96772 248294 96824
rect 250162 96772 250168 96824
rect 250220 96812 250226 96824
rect 250806 96812 250812 96824
rect 250220 96784 250812 96812
rect 250220 96772 250226 96784
rect 250806 96772 250812 96784
rect 250864 96772 250870 96824
rect 251174 96772 251180 96824
rect 251232 96812 251238 96824
rect 252186 96812 252192 96824
rect 251232 96784 252192 96812
rect 251232 96772 251238 96784
rect 252186 96772 252192 96784
rect 252244 96772 252250 96824
rect 261570 96772 261576 96824
rect 261628 96812 261634 96824
rect 261938 96812 261944 96824
rect 261628 96784 261944 96812
rect 261628 96772 261634 96784
rect 261938 96772 261944 96784
rect 261996 96772 262002 96824
rect 263152 96812 263180 96840
rect 264330 96812 264336 96824
rect 263152 96784 264336 96812
rect 264330 96772 264336 96784
rect 264388 96772 264394 96824
rect 265158 96772 265164 96824
rect 265216 96812 265222 96824
rect 266170 96812 266176 96824
rect 265216 96784 266176 96812
rect 265216 96772 265222 96784
rect 266170 96772 266176 96784
rect 266228 96772 266234 96824
rect 267182 96772 267188 96824
rect 267240 96812 267246 96824
rect 267642 96812 267648 96824
rect 267240 96784 267648 96812
rect 267240 96772 267246 96784
rect 267642 96772 267648 96784
rect 267700 96772 267706 96824
rect 268194 96772 268200 96824
rect 268252 96812 268258 96824
rect 269022 96812 269028 96824
rect 268252 96784 269028 96812
rect 268252 96772 268258 96784
rect 269022 96772 269028 96784
rect 269080 96772 269086 96824
rect 269206 96772 269212 96824
rect 269264 96812 269270 96824
rect 270218 96812 270224 96824
rect 269264 96784 270224 96812
rect 269264 96772 269270 96784
rect 270218 96772 270224 96784
rect 270276 96772 270282 96824
rect 270494 96772 270500 96824
rect 270552 96812 270558 96824
rect 271690 96812 271696 96824
rect 270552 96784 271696 96812
rect 270552 96772 270558 96784
rect 271690 96772 271696 96784
rect 271748 96772 271754 96824
rect 275094 96772 275100 96824
rect 275152 96812 275158 96824
rect 275738 96812 275744 96824
rect 275152 96784 275744 96812
rect 275152 96772 275158 96784
rect 275738 96772 275744 96784
rect 275796 96772 275802 96824
rect 280614 96772 280620 96824
rect 280672 96812 280678 96824
rect 281166 96812 281172 96824
rect 280672 96784 281172 96812
rect 280672 96772 280678 96784
rect 281166 96772 281172 96784
rect 281224 96772 281230 96824
rect 281626 96772 281632 96824
rect 281684 96812 281690 96824
rect 282822 96812 282828 96824
rect 281684 96784 282828 96812
rect 281684 96772 281690 96784
rect 282822 96772 282828 96784
rect 282880 96772 282886 96824
rect 284478 96772 284484 96824
rect 284536 96812 284542 96824
rect 285214 96812 285220 96824
rect 284536 96784 285220 96812
rect 284536 96772 284542 96784
rect 285214 96772 285220 96784
rect 285272 96772 285278 96824
rect 285858 96772 285864 96824
rect 285916 96812 285922 96824
rect 286870 96812 286876 96824
rect 285916 96784 286876 96812
rect 285916 96772 285922 96784
rect 286870 96772 286876 96784
rect 286928 96772 286934 96824
rect 288894 96772 288900 96824
rect 288952 96812 288958 96824
rect 289630 96812 289636 96824
rect 288952 96784 289636 96812
rect 288952 96772 288958 96784
rect 289630 96772 289636 96784
rect 289688 96772 289694 96824
rect 290550 96772 290556 96824
rect 290608 96812 290614 96824
rect 291010 96812 291016 96824
rect 290608 96784 291016 96812
rect 290608 96772 290614 96784
rect 291010 96772 291016 96784
rect 291068 96772 291074 96824
rect 294414 96772 294420 96824
rect 294472 96812 294478 96824
rect 294966 96812 294972 96824
rect 294472 96784 294972 96812
rect 294472 96772 294478 96784
rect 294966 96772 294972 96784
rect 295024 96772 295030 96824
rect 295610 96772 295616 96824
rect 295668 96812 295674 96824
rect 296254 96812 296260 96824
rect 295668 96784 296260 96812
rect 295668 96772 295674 96784
rect 296254 96772 296260 96784
rect 296312 96772 296318 96824
rect 297266 96772 297272 96824
rect 297324 96812 297330 96824
rect 297818 96812 297824 96824
rect 297324 96784 297824 96812
rect 297324 96772 297330 96784
rect 297818 96772 297824 96784
rect 297876 96772 297882 96824
rect 211798 96704 211804 96756
rect 211856 96744 211862 96756
rect 215110 96744 215116 96756
rect 211856 96716 215116 96744
rect 211856 96704 211862 96716
rect 215110 96704 215116 96716
rect 215168 96704 215174 96756
rect 199378 96636 199384 96688
rect 199436 96676 199442 96688
rect 201862 96676 201868 96688
rect 199436 96648 201868 96676
rect 199436 96636 199442 96648
rect 201862 96636 201868 96648
rect 201920 96636 201926 96688
rect 206922 96636 206928 96688
rect 206980 96676 206986 96688
rect 210602 96676 210608 96688
rect 206980 96648 210608 96676
rect 206980 96636 206986 96648
rect 210602 96636 210608 96648
rect 210660 96636 210666 96688
rect 210786 96636 210792 96688
rect 210844 96676 210850 96688
rect 212074 96676 212080 96688
rect 210844 96648 212080 96676
rect 210844 96636 210850 96648
rect 212074 96636 212080 96648
rect 212132 96636 212138 96688
rect 213362 96636 213368 96688
rect 213420 96676 213426 96688
rect 215266 96676 215294 96772
rect 226978 96704 226984 96756
rect 227036 96744 227042 96756
rect 229278 96744 229284 96756
rect 227036 96716 229284 96744
rect 227036 96704 227042 96716
rect 229278 96704 229284 96716
rect 229336 96704 229342 96756
rect 241606 96704 241612 96756
rect 241664 96744 241670 96756
rect 242710 96744 242716 96756
rect 241664 96716 242716 96744
rect 241664 96704 241670 96716
rect 242710 96704 242716 96716
rect 242768 96704 242774 96756
rect 243078 96704 243084 96756
rect 243136 96744 243142 96756
rect 243906 96744 243912 96756
rect 243136 96716 243912 96744
rect 243136 96704 243142 96716
rect 243906 96704 243912 96716
rect 243964 96704 243970 96756
rect 245930 96704 245936 96756
rect 245988 96744 245994 96756
rect 246758 96744 246764 96756
rect 245988 96716 246764 96744
rect 245988 96704 245994 96716
rect 246758 96704 246764 96716
rect 246816 96704 246822 96756
rect 249794 96704 249800 96756
rect 249852 96744 249858 96756
rect 250990 96744 250996 96756
rect 249852 96716 250996 96744
rect 249852 96704 249858 96716
rect 250990 96704 250996 96716
rect 251048 96704 251054 96756
rect 251634 96704 251640 96756
rect 251692 96744 251698 96756
rect 252370 96744 252376 96756
rect 251692 96716 252376 96744
rect 251692 96704 251698 96716
rect 252370 96704 252376 96716
rect 252428 96704 252434 96756
rect 253014 96704 253020 96756
rect 253072 96744 253078 96756
rect 253842 96744 253848 96756
rect 253072 96716 253848 96744
rect 253072 96704 253078 96716
rect 253842 96704 253848 96716
rect 253900 96704 253906 96756
rect 254394 96704 254400 96756
rect 254452 96744 254458 96756
rect 258718 96744 258724 96756
rect 254452 96716 258724 96744
rect 254452 96704 254458 96716
rect 258718 96704 258724 96716
rect 258776 96704 258782 96756
rect 266354 96704 266360 96756
rect 266412 96744 266418 96756
rect 267458 96744 267464 96756
rect 266412 96716 267464 96744
rect 266412 96704 266418 96716
rect 267458 96704 267464 96716
rect 267516 96704 267522 96756
rect 270034 96704 270040 96756
rect 270092 96744 270098 96756
rect 270092 96716 274864 96744
rect 270092 96704 270098 96716
rect 213420 96648 215294 96676
rect 213420 96636 213426 96648
rect 222838 96636 222844 96688
rect 222896 96676 222902 96688
rect 223482 96676 223488 96688
rect 222896 96648 223488 96676
rect 222896 96636 222902 96648
rect 223482 96636 223488 96648
rect 223540 96636 223546 96688
rect 228542 96636 228548 96688
rect 228600 96676 228606 96688
rect 233786 96676 233792 96688
rect 228600 96648 233792 96676
rect 228600 96636 228606 96648
rect 233786 96636 233792 96648
rect 233844 96636 233850 96688
rect 234798 96636 234804 96688
rect 234856 96676 234862 96688
rect 235258 96676 235264 96688
rect 234856 96648 235264 96676
rect 234856 96636 234862 96648
rect 235258 96636 235264 96648
rect 235316 96636 235322 96688
rect 236086 96636 236092 96688
rect 236144 96676 236150 96688
rect 236730 96676 236736 96688
rect 236144 96648 236736 96676
rect 236144 96636 236150 96648
rect 236730 96636 236736 96648
rect 236788 96636 236794 96688
rect 237650 96636 237656 96688
rect 237708 96676 237714 96688
rect 238478 96676 238484 96688
rect 237708 96648 238484 96676
rect 237708 96636 237714 96648
rect 238478 96636 238484 96648
rect 238536 96636 238542 96688
rect 240134 96636 240140 96688
rect 240192 96676 240198 96688
rect 241238 96676 241244 96688
rect 240192 96648 241244 96676
rect 240192 96636 240198 96648
rect 241238 96636 241244 96648
rect 241296 96636 241302 96688
rect 248506 96636 248512 96688
rect 248564 96676 248570 96688
rect 249426 96676 249432 96688
rect 248564 96648 249432 96676
rect 248564 96636 248570 96648
rect 249426 96636 249432 96648
rect 249484 96636 249490 96688
rect 252830 96636 252836 96688
rect 252888 96676 252894 96688
rect 253658 96676 253664 96688
rect 252888 96648 253664 96676
rect 252888 96636 252894 96648
rect 253658 96636 253664 96648
rect 253716 96636 253722 96688
rect 257246 96636 257252 96688
rect 257304 96676 257310 96688
rect 257798 96676 257804 96688
rect 257304 96648 257804 96676
rect 257304 96636 257310 96648
rect 257798 96636 257804 96648
rect 257856 96636 257862 96688
rect 261754 96636 261760 96688
rect 261812 96676 261818 96688
rect 262122 96676 262128 96688
rect 261812 96648 262128 96676
rect 261812 96636 261818 96648
rect 262122 96636 262128 96648
rect 262180 96636 262186 96688
rect 262306 96636 262312 96688
rect 262364 96676 262370 96688
rect 263318 96676 263324 96688
rect 262364 96648 263324 96676
rect 262364 96636 262370 96648
rect 263318 96636 263324 96648
rect 263376 96636 263382 96688
rect 273530 96636 273536 96688
rect 273588 96676 273594 96688
rect 274358 96676 274364 96688
rect 273588 96648 274364 96676
rect 273588 96636 273594 96648
rect 274358 96636 274364 96648
rect 274416 96636 274422 96688
rect 274836 96676 274864 96716
rect 274910 96704 274916 96756
rect 274968 96744 274974 96756
rect 275830 96744 275836 96756
rect 274968 96716 275836 96744
rect 274968 96704 274974 96716
rect 275830 96704 275836 96716
rect 275888 96704 275894 96756
rect 280430 96704 280436 96756
rect 280488 96744 280494 96756
rect 281442 96744 281448 96756
rect 280488 96716 281448 96744
rect 280488 96704 280494 96716
rect 281442 96704 281448 96716
rect 281500 96704 281506 96756
rect 284662 96704 284668 96756
rect 284720 96744 284726 96756
rect 285398 96744 285404 96756
rect 284720 96716 285404 96744
rect 284720 96704 284726 96716
rect 285398 96704 285404 96716
rect 285456 96704 285462 96756
rect 294782 96704 294788 96756
rect 294840 96744 294846 96756
rect 295242 96744 295248 96756
rect 294840 96716 295248 96744
rect 294840 96704 294846 96716
rect 295242 96704 295248 96716
rect 295300 96704 295306 96756
rect 296806 96704 296812 96756
rect 296864 96744 296870 96756
rect 297726 96744 297732 96756
rect 296864 96716 297732 96744
rect 296864 96704 296870 96716
rect 297726 96704 297732 96716
rect 297784 96704 297790 96756
rect 275278 96676 275284 96688
rect 274836 96648 275284 96676
rect 275278 96636 275284 96648
rect 275336 96636 275342 96688
rect 277578 96636 277584 96688
rect 277636 96676 277642 96688
rect 278498 96676 278504 96688
rect 277636 96648 278504 96676
rect 277636 96636 277642 96648
rect 278498 96636 278504 96648
rect 278556 96636 278562 96688
rect 283466 96636 283472 96688
rect 283524 96676 283530 96688
rect 284110 96676 284116 96688
rect 283524 96648 284116 96676
rect 283524 96636 283530 96648
rect 284110 96636 284116 96648
rect 284168 96636 284174 96688
rect 290366 96636 290372 96688
rect 290424 96676 290430 96688
rect 291194 96676 291200 96688
rect 290424 96648 291200 96676
rect 290424 96636 290430 96648
rect 291194 96636 291200 96648
rect 291252 96636 291258 96688
rect 291378 96636 291384 96688
rect 291436 96676 291442 96688
rect 292390 96676 292396 96688
rect 291436 96648 292396 96676
rect 291436 96636 291442 96648
rect 292390 96636 292396 96648
rect 292448 96636 292454 96688
rect 298646 96636 298652 96688
rect 298704 96676 298710 96688
rect 299198 96676 299204 96688
rect 298704 96648 299204 96676
rect 298704 96636 298710 96648
rect 299198 96636 299204 96648
rect 299256 96636 299262 96688
rect 298002 96568 298008 96620
rect 298060 96608 298066 96620
rect 298738 96608 298744 96620
rect 298060 96580 298744 96608
rect 298060 96568 298066 96580
rect 298738 96568 298744 96580
rect 298796 96568 298802 96620
rect 251358 96296 251364 96348
rect 251416 96336 251422 96348
rect 302326 96336 302332 96348
rect 251416 96308 302332 96336
rect 251416 96296 251422 96308
rect 302326 96296 302332 96308
rect 302384 96296 302390 96348
rect 200022 96228 200028 96280
rect 200080 96268 200086 96280
rect 234982 96268 234988 96280
rect 200080 96240 234988 96268
rect 200080 96228 200086 96240
rect 234982 96228 234988 96240
rect 235040 96228 235046 96280
rect 256694 96228 256700 96280
rect 256752 96268 256758 96280
rect 329834 96268 329840 96280
rect 256752 96240 329840 96268
rect 256752 96228 256758 96240
rect 329834 96228 329840 96240
rect 329892 96228 329898 96280
rect 192478 96160 192484 96212
rect 192536 96200 192542 96212
rect 232498 96200 232504 96212
rect 192536 96172 232504 96200
rect 192536 96160 192542 96172
rect 232498 96160 232504 96172
rect 232556 96160 232562 96212
rect 240318 96160 240324 96212
rect 240376 96200 240382 96212
rect 240686 96200 240692 96212
rect 240376 96172 240692 96200
rect 240376 96160 240382 96172
rect 240686 96160 240692 96172
rect 240744 96160 240750 96212
rect 300578 96160 300584 96212
rect 300636 96200 300642 96212
rect 378134 96200 378140 96212
rect 300636 96172 378140 96200
rect 300636 96160 300642 96172
rect 378134 96160 378140 96172
rect 378192 96160 378198 96212
rect 178678 96092 178684 96144
rect 178736 96132 178742 96144
rect 222010 96132 222016 96144
rect 178736 96104 222016 96132
rect 178736 96092 178742 96104
rect 222010 96092 222016 96104
rect 222068 96092 222074 96144
rect 258074 96092 258080 96144
rect 258132 96132 258138 96144
rect 338114 96132 338120 96144
rect 258132 96104 338120 96132
rect 258132 96092 258138 96104
rect 338114 96092 338120 96104
rect 338172 96092 338178 96144
rect 183462 96024 183468 96076
rect 183520 96064 183526 96076
rect 231302 96064 231308 96076
rect 183520 96036 231308 96064
rect 183520 96024 183526 96036
rect 231302 96024 231308 96036
rect 231360 96024 231366 96076
rect 286042 96024 286048 96076
rect 286100 96064 286106 96076
rect 500954 96064 500960 96076
rect 286100 96036 500960 96064
rect 286100 96024 286106 96036
rect 500954 96024 500960 96036
rect 501012 96024 501018 96076
rect 159358 95956 159364 96008
rect 159416 95996 159422 96008
rect 222746 95996 222752 96008
rect 159416 95968 222752 95996
rect 159416 95956 159422 95968
rect 222746 95956 222752 95968
rect 222804 95956 222810 96008
rect 287330 95956 287336 96008
rect 287388 95996 287394 96008
rect 507854 95996 507860 96008
rect 287388 95968 507860 95996
rect 287388 95956 287394 95968
rect 507854 95956 507860 95968
rect 507912 95956 507918 96008
rect 4062 95888 4068 95940
rect 4120 95928 4126 95940
rect 200482 95928 200488 95940
rect 4120 95900 200488 95928
rect 4120 95888 4126 95900
rect 200482 95888 200488 95900
rect 200540 95888 200546 95940
rect 288526 95888 288532 95940
rect 288584 95928 288590 95940
rect 518894 95928 518900 95940
rect 288584 95900 518900 95928
rect 288584 95888 288590 95900
rect 518894 95888 518900 95900
rect 518952 95888 518958 95940
rect 215570 95412 215576 95464
rect 215628 95452 215634 95464
rect 216214 95452 216220 95464
rect 215628 95424 216220 95452
rect 215628 95412 215634 95424
rect 216214 95412 216220 95424
rect 216272 95412 216278 95464
rect 222930 95208 222936 95260
rect 222988 95248 222994 95260
rect 229370 95248 229376 95260
rect 222988 95220 229376 95248
rect 222988 95208 222994 95220
rect 229370 95208 229376 95220
rect 229428 95208 229434 95260
rect 287974 95072 287980 95124
rect 288032 95112 288038 95124
rect 295978 95112 295984 95124
rect 288032 95084 295984 95112
rect 288032 95072 288038 95084
rect 295978 95072 295984 95084
rect 296036 95072 296042 95124
rect 201586 94868 201592 94920
rect 201644 94908 201650 94920
rect 202414 94908 202420 94920
rect 201644 94880 202420 94908
rect 201644 94868 201650 94880
rect 202414 94868 202420 94880
rect 202472 94868 202478 94920
rect 203334 94868 203340 94920
rect 203392 94908 203398 94920
rect 203518 94908 203524 94920
rect 203392 94880 203524 94908
rect 203392 94868 203398 94880
rect 203518 94868 203524 94880
rect 203576 94868 203582 94920
rect 212718 94868 212724 94920
rect 212776 94908 212782 94920
rect 213178 94908 213184 94920
rect 212776 94880 213184 94908
rect 212776 94868 212782 94880
rect 213178 94868 213184 94880
rect 213236 94868 213242 94920
rect 257062 94868 257068 94920
rect 257120 94908 257126 94920
rect 318058 94908 318064 94920
rect 257120 94880 318064 94908
rect 257120 94868 257126 94880
rect 318058 94868 318064 94880
rect 318116 94868 318122 94920
rect 181438 94800 181444 94852
rect 181496 94840 181502 94852
rect 227898 94840 227904 94852
rect 181496 94812 227904 94840
rect 181496 94800 181502 94812
rect 227898 94800 227904 94812
rect 227956 94800 227962 94852
rect 228358 94800 228364 94852
rect 228416 94800 228422 94852
rect 254210 94800 254216 94852
rect 254268 94840 254274 94852
rect 316034 94840 316040 94852
rect 254268 94812 316040 94840
rect 254268 94800 254274 94812
rect 316034 94800 316040 94812
rect 316092 94800 316098 94852
rect 166902 94732 166908 94784
rect 166960 94772 166966 94784
rect 228376 94772 228404 94800
rect 166960 94744 228404 94772
rect 166960 94732 166966 94744
rect 265894 94732 265900 94784
rect 265952 94772 265958 94784
rect 375374 94772 375380 94784
rect 265952 94744 375380 94772
rect 265952 94732 265958 94744
rect 375374 94732 375380 94744
rect 375432 94732 375438 94784
rect 158622 94664 158628 94716
rect 158680 94704 158686 94716
rect 227070 94704 227076 94716
rect 158680 94676 227076 94704
rect 158680 94664 158686 94676
rect 227070 94664 227076 94676
rect 227128 94664 227134 94716
rect 228358 94664 228364 94716
rect 228416 94704 228422 94716
rect 228416 94676 234568 94704
rect 228416 94664 228422 94676
rect 143442 94596 143448 94648
rect 143500 94636 143506 94648
rect 224402 94636 224408 94648
rect 143500 94608 224408 94636
rect 143500 94596 143506 94608
rect 224402 94596 224408 94608
rect 224460 94596 224466 94648
rect 234540 94636 234568 94676
rect 272058 94664 272064 94716
rect 272116 94704 272122 94716
rect 421006 94704 421012 94716
rect 272116 94676 421012 94704
rect 272116 94664 272122 94676
rect 421006 94664 421012 94676
rect 421064 94664 421070 94716
rect 236362 94636 236368 94648
rect 234540 94608 236368 94636
rect 236362 94596 236368 94608
rect 236420 94596 236426 94648
rect 304994 94596 305000 94648
rect 305052 94636 305058 94648
rect 557534 94636 557540 94648
rect 305052 94608 557540 94636
rect 305052 94596 305058 94608
rect 557534 94596 557540 94608
rect 557592 94596 557598 94648
rect 126882 94528 126888 94580
rect 126940 94568 126946 94580
rect 221734 94568 221740 94580
rect 126940 94540 221740 94568
rect 126940 94528 126946 94540
rect 221734 94528 221740 94540
rect 221792 94528 221798 94580
rect 226702 94528 226708 94580
rect 226760 94568 226766 94580
rect 227346 94568 227352 94580
rect 226760 94540 227352 94568
rect 226760 94528 226766 94540
rect 227346 94528 227352 94540
rect 227404 94528 227410 94580
rect 229002 94528 229008 94580
rect 229060 94568 229066 94580
rect 239214 94568 239220 94580
rect 229060 94540 230428 94568
rect 229060 94528 229066 94540
rect 43438 94460 43444 94512
rect 43496 94500 43502 94512
rect 43496 94472 195974 94500
rect 43496 94460 43502 94472
rect 195946 94432 195974 94472
rect 200390 94460 200396 94512
rect 200448 94500 200454 94512
rect 201218 94500 201224 94512
rect 200448 94472 201224 94500
rect 200448 94460 200454 94472
rect 201218 94460 201224 94472
rect 201276 94460 201282 94512
rect 204438 94460 204444 94512
rect 204496 94500 204502 94512
rect 204622 94500 204628 94512
rect 204496 94472 204628 94500
rect 204496 94460 204502 94472
rect 204622 94460 204628 94472
rect 204680 94460 204686 94512
rect 208486 94460 208492 94512
rect 208544 94500 208550 94512
rect 209498 94500 209504 94512
rect 208544 94472 209504 94500
rect 208544 94460 208550 94472
rect 209498 94460 209504 94472
rect 209556 94460 209562 94512
rect 209866 94460 209872 94512
rect 209924 94500 209930 94512
rect 210878 94500 210884 94512
rect 209924 94472 210884 94500
rect 209924 94460 209930 94472
rect 210878 94460 210884 94472
rect 210936 94460 210942 94512
rect 211522 94460 211528 94512
rect 211580 94500 211586 94512
rect 212166 94500 212172 94512
rect 211580 94472 212172 94500
rect 211580 94460 211586 94472
rect 212166 94460 212172 94472
rect 212224 94460 212230 94512
rect 214006 94460 214012 94512
rect 214064 94500 214070 94512
rect 214374 94500 214380 94512
rect 214064 94472 214380 94500
rect 214064 94460 214070 94472
rect 214374 94460 214380 94472
rect 214432 94460 214438 94512
rect 229370 94460 229376 94512
rect 229428 94500 229434 94512
rect 230198 94500 230204 94512
rect 229428 94472 230204 94500
rect 229428 94460 229434 94472
rect 230198 94460 230204 94472
rect 230256 94460 230262 94512
rect 230400 94500 230428 94540
rect 234448 94540 239220 94568
rect 234448 94500 234476 94540
rect 239214 94528 239220 94540
rect 239272 94528 239278 94580
rect 263594 94528 263600 94580
rect 263652 94568 263658 94580
rect 294598 94568 294604 94580
rect 263652 94540 294604 94568
rect 263652 94528 263658 94540
rect 294598 94528 294604 94540
rect 294656 94528 294662 94580
rect 296070 94528 296076 94580
rect 296128 94568 296134 94580
rect 561674 94568 561680 94580
rect 296128 94540 561680 94568
rect 296128 94528 296134 94540
rect 561674 94528 561680 94540
rect 561732 94528 561738 94580
rect 237374 94500 237380 94512
rect 230400 94472 234476 94500
rect 234586 94472 237380 94500
rect 204162 94432 204168 94444
rect 195946 94404 204168 94432
rect 204162 94392 204168 94404
rect 204220 94392 204226 94444
rect 214190 94392 214196 94444
rect 214248 94432 214254 94444
rect 214834 94432 214840 94444
rect 214248 94404 214840 94432
rect 214248 94392 214254 94404
rect 214834 94392 214840 94404
rect 214892 94392 214898 94444
rect 227622 94392 227628 94444
rect 227680 94432 227686 94444
rect 234586 94432 234614 94472
rect 237374 94460 237380 94472
rect 237432 94460 237438 94512
rect 250346 94460 250352 94512
rect 250404 94500 250410 94512
rect 289078 94500 289084 94512
rect 250404 94472 289084 94500
rect 250404 94460 250410 94472
rect 289078 94460 289084 94472
rect 289136 94460 289142 94512
rect 296990 94460 296996 94512
rect 297048 94500 297054 94512
rect 565814 94500 565820 94512
rect 297048 94472 565820 94500
rect 297048 94460 297054 94472
rect 565814 94460 565820 94472
rect 565872 94460 565878 94512
rect 227680 94404 234614 94432
rect 227680 94392 227686 94404
rect 204622 94324 204628 94376
rect 204680 94364 204686 94376
rect 205450 94364 205456 94376
rect 204680 94336 205456 94364
rect 204680 94324 204686 94336
rect 205450 94324 205456 94336
rect 205508 94324 205514 94376
rect 293862 93848 293868 93900
rect 293920 93888 293926 93900
rect 297358 93888 297364 93900
rect 293920 93860 297364 93888
rect 293920 93848 293926 93860
rect 297358 93848 297364 93860
rect 297416 93848 297422 93900
rect 198642 93508 198648 93560
rect 198700 93548 198706 93560
rect 233878 93548 233884 93560
rect 198700 93520 233884 93548
rect 198700 93508 198706 93520
rect 233878 93508 233884 93520
rect 233936 93508 233942 93560
rect 191742 93440 191748 93492
rect 191800 93480 191806 93492
rect 232590 93480 232596 93492
rect 191800 93452 232596 93480
rect 191800 93440 191806 93452
rect 232590 93440 232596 93452
rect 232648 93440 232654 93492
rect 256326 93440 256332 93492
rect 256384 93480 256390 93492
rect 327074 93480 327080 93492
rect 256384 93452 327080 93480
rect 256384 93440 256390 93452
rect 327074 93440 327080 93452
rect 327132 93440 327138 93492
rect 184842 93372 184848 93424
rect 184900 93412 184906 93424
rect 231394 93412 231400 93424
rect 184900 93384 231400 93412
rect 184900 93372 184906 93384
rect 231394 93372 231400 93384
rect 231452 93372 231458 93424
rect 257890 93372 257896 93424
rect 257948 93412 257954 93424
rect 333974 93412 333980 93424
rect 257948 93384 333980 93412
rect 257948 93372 257954 93384
rect 333974 93372 333980 93384
rect 334032 93372 334038 93424
rect 148962 93304 148968 93356
rect 149020 93344 149026 93356
rect 225230 93344 225236 93356
rect 149020 93316 225236 93344
rect 149020 93304 149026 93316
rect 225230 93304 225236 93316
rect 225288 93304 225294 93356
rect 259178 93304 259184 93356
rect 259236 93344 259242 93356
rect 335998 93344 336004 93356
rect 259236 93316 336004 93344
rect 259236 93304 259242 93316
rect 335998 93304 336004 93316
rect 336056 93304 336062 93356
rect 142062 93236 142068 93288
rect 142120 93276 142126 93288
rect 224126 93276 224132 93288
rect 142120 93248 224132 93276
rect 142120 93236 142126 93248
rect 224126 93236 224132 93248
rect 224184 93236 224190 93288
rect 263318 93236 263324 93288
rect 263376 93276 263382 93288
rect 311158 93276 311164 93288
rect 263376 93248 311164 93276
rect 263376 93236 263382 93248
rect 311158 93236 311164 93248
rect 311216 93236 311222 93288
rect 312538 93236 312544 93288
rect 312596 93276 312602 93288
rect 539594 93276 539600 93288
rect 312596 93248 539600 93276
rect 312596 93236 312602 93248
rect 539594 93236 539600 93248
rect 539652 93236 539658 93288
rect 37182 93168 37188 93220
rect 37240 93208 37246 93220
rect 205910 93208 205916 93220
rect 37240 93180 205916 93208
rect 37240 93168 37246 93180
rect 205910 93168 205916 93180
rect 205968 93168 205974 93220
rect 292482 93168 292488 93220
rect 292540 93208 292546 93220
rect 546586 93208 546592 93220
rect 292540 93180 546592 93208
rect 292540 93168 292546 93180
rect 546586 93168 546592 93180
rect 546644 93168 546650 93220
rect 22002 93100 22008 93152
rect 22060 93140 22066 93152
rect 203610 93140 203616 93152
rect 22060 93112 203616 93140
rect 22060 93100 22066 93112
rect 203610 93100 203616 93112
rect 203668 93100 203674 93152
rect 224862 93100 224868 93152
rect 224920 93140 224926 93152
rect 238294 93140 238300 93152
rect 224920 93112 238300 93140
rect 224920 93100 224926 93112
rect 238294 93100 238300 93112
rect 238352 93100 238358 93152
rect 244182 93100 244188 93152
rect 244240 93140 244246 93152
rect 255314 93140 255320 93152
rect 244240 93112 255320 93140
rect 244240 93100 244246 93112
rect 255314 93100 255320 93112
rect 255372 93100 255378 93152
rect 283558 93100 283564 93152
rect 283616 93140 283622 93152
rect 294690 93140 294696 93152
rect 283616 93112 294696 93140
rect 283616 93100 283622 93112
rect 294690 93100 294696 93112
rect 294748 93100 294754 93152
rect 295242 93100 295248 93152
rect 295300 93140 295306 93152
rect 564434 93140 564440 93152
rect 295300 93112 564440 93140
rect 295300 93100 295306 93112
rect 564434 93100 564440 93112
rect 564492 93100 564498 93152
rect 186222 92148 186228 92200
rect 186280 92188 186286 92200
rect 231578 92188 231584 92200
rect 186280 92160 231584 92188
rect 186280 92148 186286 92160
rect 231578 92148 231584 92160
rect 231636 92148 231642 92200
rect 282178 92148 282184 92200
rect 282236 92188 282242 92200
rect 313274 92188 313280 92200
rect 282236 92160 313280 92188
rect 282236 92148 282242 92160
rect 313274 92148 313280 92160
rect 313332 92148 313338 92200
rect 171042 92080 171048 92132
rect 171100 92120 171106 92132
rect 226978 92120 226984 92132
rect 171100 92092 226984 92120
rect 171100 92080 171106 92092
rect 226978 92080 226984 92092
rect 227036 92080 227042 92132
rect 275370 92080 275376 92132
rect 275428 92120 275434 92132
rect 356054 92120 356060 92132
rect 275428 92092 356060 92120
rect 275428 92080 275434 92092
rect 356054 92080 356060 92092
rect 356112 92080 356118 92132
rect 137278 92012 137284 92064
rect 137336 92052 137342 92064
rect 222562 92052 222568 92064
rect 137336 92024 222568 92052
rect 137336 92012 137342 92024
rect 222562 92012 222568 92024
rect 222620 92012 222626 92064
rect 262122 92012 262128 92064
rect 262180 92052 262186 92064
rect 358814 92052 358820 92064
rect 262180 92024 358820 92052
rect 262180 92012 262186 92024
rect 358814 92012 358820 92024
rect 358872 92012 358878 92064
rect 71038 91944 71044 91996
rect 71096 91984 71102 91996
rect 211430 91984 211436 91996
rect 71096 91956 211436 91984
rect 71096 91944 71102 91956
rect 211430 91944 211436 91956
rect 211488 91944 211494 91996
rect 263410 91944 263416 91996
rect 263468 91984 263474 91996
rect 364978 91984 364984 91996
rect 263468 91956 364984 91984
rect 263468 91944 263474 91956
rect 364978 91944 364984 91956
rect 365036 91944 365042 91996
rect 23382 91876 23388 91928
rect 23440 91916 23446 91928
rect 203794 91916 203800 91928
rect 23440 91888 203800 91916
rect 23440 91876 23446 91888
rect 203794 91876 203800 91888
rect 203852 91876 203858 91928
rect 265986 91876 265992 91928
rect 266044 91916 266050 91928
rect 374638 91916 374644 91928
rect 266044 91888 374644 91916
rect 266044 91876 266050 91888
rect 374638 91876 374644 91888
rect 374696 91876 374702 91928
rect 12342 91808 12348 91860
rect 12400 91848 12406 91860
rect 195330 91848 195336 91860
rect 12400 91820 195336 91848
rect 12400 91808 12406 91820
rect 195330 91808 195336 91820
rect 195388 91808 195394 91860
rect 195882 91808 195888 91860
rect 195940 91848 195946 91860
rect 233418 91848 233424 91860
rect 195940 91820 233424 91848
rect 195940 91808 195946 91820
rect 233418 91808 233424 91820
rect 233476 91808 233482 91860
rect 269758 91808 269764 91860
rect 269816 91848 269822 91860
rect 380894 91848 380900 91860
rect 269816 91820 380900 91848
rect 269816 91808 269822 91820
rect 380894 91808 380900 91820
rect 380952 91808 380958 91860
rect 1302 91740 1308 91792
rect 1360 91780 1366 91792
rect 188338 91780 188344 91792
rect 1360 91752 188344 91780
rect 1360 91740 1366 91752
rect 188338 91740 188344 91752
rect 188396 91740 188402 91792
rect 188982 91740 188988 91792
rect 189040 91780 189046 91792
rect 232222 91780 232228 91792
rect 189040 91752 232228 91780
rect 189040 91740 189046 91752
rect 232222 91740 232228 91752
rect 232280 91740 232286 91792
rect 242802 91740 242808 91792
rect 242860 91780 242866 91792
rect 258074 91780 258080 91792
rect 242860 91752 258080 91780
rect 242860 91740 242866 91752
rect 258074 91740 258080 91752
rect 258132 91740 258138 91792
rect 267642 91740 267648 91792
rect 267700 91780 267706 91792
rect 389818 91780 389824 91792
rect 267700 91752 389824 91780
rect 267700 91740 267706 91752
rect 389818 91740 389824 91752
rect 389876 91740 389882 91792
rect 233142 91332 233148 91384
rect 233200 91372 233206 91384
rect 239674 91372 239680 91384
rect 233200 91344 239680 91372
rect 233200 91332 233206 91344
rect 239674 91332 239680 91344
rect 239732 91332 239738 91384
rect 231762 91060 231768 91112
rect 231820 91100 231826 91112
rect 236638 91100 236644 91112
rect 231820 91072 236644 91100
rect 231820 91060 231826 91072
rect 236638 91060 236644 91072
rect 236696 91060 236702 91112
rect 181530 90720 181536 90772
rect 181588 90760 181594 90772
rect 225506 90760 225512 90772
rect 181588 90732 225512 90760
rect 181588 90720 181594 90732
rect 225506 90720 225512 90732
rect 225564 90720 225570 90772
rect 253658 90720 253664 90772
rect 253716 90760 253722 90772
rect 307018 90760 307024 90772
rect 253716 90732 307024 90760
rect 253716 90720 253722 90732
rect 307018 90720 307024 90732
rect 307076 90720 307082 90772
rect 162210 90652 162216 90704
rect 162268 90692 162274 90704
rect 226610 90692 226616 90704
rect 162268 90664 226616 90692
rect 162268 90652 162274 90664
rect 226610 90652 226616 90664
rect 226668 90652 226674 90704
rect 260650 90652 260656 90704
rect 260708 90692 260714 90704
rect 347038 90692 347044 90704
rect 260708 90664 347044 90692
rect 260708 90652 260714 90664
rect 347038 90652 347044 90664
rect 347096 90652 347102 90704
rect 104158 90584 104164 90636
rect 104216 90624 104222 90636
rect 217410 90624 217416 90636
rect 104216 90596 217416 90624
rect 104216 90584 104222 90596
rect 217410 90584 217416 90596
rect 217468 90584 217474 90636
rect 271506 90584 271512 90636
rect 271564 90624 271570 90636
rect 412634 90624 412640 90636
rect 271564 90596 412640 90624
rect 271564 90584 271570 90596
rect 412634 90584 412640 90596
rect 412692 90584 412698 90636
rect 73062 90516 73068 90568
rect 73120 90556 73126 90568
rect 212350 90556 212356 90568
rect 73120 90528 212356 90556
rect 73120 90516 73126 90528
rect 212350 90516 212356 90528
rect 212408 90516 212414 90568
rect 271782 90516 271788 90568
rect 271840 90556 271846 90568
rect 416866 90556 416872 90568
rect 271840 90528 416872 90556
rect 271840 90516 271846 90528
rect 416866 90516 416872 90528
rect 416924 90516 416930 90568
rect 62022 90448 62028 90500
rect 62080 90488 62086 90500
rect 206922 90488 206928 90500
rect 62080 90460 206928 90488
rect 62080 90448 62086 90460
rect 206922 90448 206928 90460
rect 206980 90448 206986 90500
rect 274266 90448 274272 90500
rect 274324 90488 274330 90500
rect 427906 90488 427912 90500
rect 274324 90460 427912 90488
rect 274324 90448 274330 90460
rect 427906 90448 427912 90460
rect 427964 90448 427970 90500
rect 55122 90380 55128 90432
rect 55180 90420 55186 90432
rect 204254 90420 204260 90432
rect 55180 90392 204260 90420
rect 55180 90380 55186 90392
rect 204254 90380 204260 90392
rect 204312 90380 204318 90432
rect 274542 90380 274548 90432
rect 274600 90420 274606 90432
rect 430574 90420 430580 90432
rect 274600 90392 430580 90420
rect 274600 90380 274606 90392
rect 430574 90380 430580 90392
rect 430632 90380 430638 90432
rect 59262 90312 59268 90364
rect 59320 90352 59326 90364
rect 209774 90352 209780 90364
rect 59320 90324 209780 90352
rect 59320 90312 59326 90324
rect 209774 90312 209780 90324
rect 209832 90312 209838 90364
rect 275738 90312 275744 90364
rect 275796 90352 275802 90364
rect 438946 90352 438952 90364
rect 275796 90324 438952 90352
rect 275796 90312 275802 90324
rect 438946 90312 438952 90324
rect 439004 90312 439010 90364
rect 233602 89904 233608 89956
rect 233660 89944 233666 89956
rect 234430 89944 234436 89956
rect 233660 89916 234436 89944
rect 233660 89904 233666 89916
rect 234430 89904 234436 89916
rect 234488 89904 234494 89956
rect 178770 89360 178776 89412
rect 178828 89400 178834 89412
rect 229370 89400 229376 89412
rect 178828 89372 229376 89400
rect 178828 89360 178834 89372
rect 229370 89360 229376 89372
rect 229428 89360 229434 89412
rect 252278 89360 252284 89412
rect 252336 89400 252342 89412
rect 300854 89400 300860 89412
rect 252336 89372 300860 89400
rect 252336 89360 252342 89372
rect 300854 89360 300860 89372
rect 300912 89360 300918 89412
rect 177298 89292 177304 89344
rect 177356 89332 177362 89344
rect 230014 89332 230020 89344
rect 177356 89304 230020 89332
rect 177356 89292 177362 89304
rect 230014 89292 230020 89304
rect 230072 89292 230078 89344
rect 253290 89292 253296 89344
rect 253348 89332 253354 89344
rect 303614 89332 303620 89344
rect 253348 89304 303620 89332
rect 253348 89292 253354 89304
rect 303614 89292 303620 89304
rect 303672 89292 303678 89344
rect 122098 89224 122104 89276
rect 122156 89264 122162 89276
rect 214282 89264 214288 89276
rect 122156 89236 214288 89264
rect 122156 89224 122162 89236
rect 214282 89224 214288 89236
rect 214340 89224 214346 89276
rect 281166 89224 281172 89276
rect 281224 89264 281230 89276
rect 341518 89264 341524 89276
rect 281224 89236 341524 89264
rect 281224 89224 281230 89236
rect 341518 89224 341524 89236
rect 341576 89224 341582 89276
rect 115198 89156 115204 89208
rect 115256 89196 115262 89208
rect 214190 89196 214196 89208
rect 115256 89168 214196 89196
rect 115256 89156 115262 89168
rect 214190 89156 214196 89168
rect 214248 89156 214254 89208
rect 278314 89156 278320 89208
rect 278372 89196 278378 89208
rect 385678 89196 385684 89208
rect 278372 89168 385684 89196
rect 278372 89156 278378 89168
rect 385678 89156 385684 89168
rect 385736 89156 385742 89208
rect 112438 89088 112444 89140
rect 112496 89128 112502 89140
rect 219066 89128 219072 89140
rect 112496 89100 219072 89128
rect 112496 89088 112502 89100
rect 219066 89088 219072 89100
rect 219124 89088 219130 89140
rect 279878 89088 279884 89140
rect 279936 89128 279942 89140
rect 457438 89128 457444 89140
rect 279936 89100 457444 89128
rect 279936 89088 279942 89100
rect 457438 89088 457444 89100
rect 457496 89088 457502 89140
rect 108942 89020 108948 89072
rect 109000 89060 109006 89072
rect 218514 89060 218520 89072
rect 109000 89032 218520 89060
rect 109000 89020 109006 89032
rect 218514 89020 218520 89032
rect 218572 89020 218578 89072
rect 282454 89020 282460 89072
rect 282512 89060 282518 89072
rect 476114 89060 476120 89072
rect 282512 89032 476120 89060
rect 282512 89020 282518 89032
rect 476114 89020 476120 89032
rect 476172 89020 476178 89072
rect 91002 88952 91008 89004
rect 91060 88992 91066 89004
rect 206278 88992 206284 89004
rect 91060 88964 206284 88992
rect 91060 88952 91066 88964
rect 206278 88952 206284 88964
rect 206336 88952 206342 89004
rect 248046 88952 248052 89004
rect 248104 88992 248110 89004
rect 281534 88992 281540 89004
rect 248104 88964 281540 88992
rect 248104 88952 248110 88964
rect 281534 88952 281540 88964
rect 281592 88952 281598 89004
rect 283834 88952 283840 89004
rect 283892 88992 283898 89004
rect 484394 88992 484400 89004
rect 283892 88964 484400 88992
rect 283892 88952 283898 88964
rect 484394 88952 484400 88964
rect 484452 88952 484458 89004
rect 197170 88000 197176 88052
rect 197228 88040 197234 88052
rect 228542 88040 228548 88052
rect 197228 88012 228548 88040
rect 197228 88000 197234 88012
rect 228542 88000 228548 88012
rect 228600 88000 228606 88052
rect 252370 88000 252376 88052
rect 252428 88040 252434 88052
rect 309134 88040 309140 88052
rect 252428 88012 309140 88040
rect 252428 88000 252434 88012
rect 309134 88000 309140 88012
rect 309192 88000 309198 88052
rect 193122 87932 193128 87984
rect 193180 87972 193186 87984
rect 234890 87972 234896 87984
rect 193180 87944 234896 87972
rect 193180 87932 193186 87944
rect 234890 87932 234896 87944
rect 234948 87932 234954 87984
rect 255038 87932 255044 87984
rect 255096 87972 255102 87984
rect 317414 87972 317420 87984
rect 255096 87944 317420 87972
rect 255096 87932 255102 87944
rect 317414 87932 317420 87944
rect 317472 87932 317478 87984
rect 95142 87864 95148 87916
rect 95200 87904 95206 87916
rect 215570 87904 215576 87916
rect 95200 87876 215576 87904
rect 95200 87864 95206 87876
rect 215570 87864 215576 87876
rect 215628 87864 215634 87916
rect 259270 87864 259276 87916
rect 259328 87904 259334 87916
rect 339494 87904 339500 87916
rect 259328 87876 339500 87904
rect 259328 87864 259334 87876
rect 339494 87864 339500 87876
rect 339552 87864 339558 87916
rect 88978 87796 88984 87848
rect 89036 87836 89042 87848
rect 212718 87836 212724 87848
rect 89036 87808 212724 87836
rect 89036 87796 89042 87808
rect 212718 87796 212724 87808
rect 212776 87796 212782 87848
rect 268562 87796 268568 87848
rect 268620 87836 268626 87848
rect 396718 87836 396724 87848
rect 268620 87808 396724 87836
rect 268620 87796 268626 87808
rect 396718 87796 396724 87808
rect 396776 87796 396782 87848
rect 70302 87728 70308 87780
rect 70360 87768 70366 87780
rect 210418 87768 210424 87780
rect 70360 87740 210424 87768
rect 70360 87728 70366 87740
rect 210418 87728 210424 87740
rect 210476 87728 210482 87780
rect 288066 87728 288072 87780
rect 288124 87768 288130 87780
rect 489178 87768 489184 87780
rect 288124 87740 489184 87768
rect 288124 87728 288130 87740
rect 489178 87728 489184 87740
rect 489236 87728 489242 87780
rect 53742 87660 53748 87712
rect 53800 87700 53806 87712
rect 208670 87700 208676 87712
rect 53800 87672 208676 87700
rect 53800 87660 53806 87672
rect 208670 87660 208676 87672
rect 208728 87660 208734 87712
rect 249426 87660 249432 87712
rect 249484 87700 249490 87712
rect 285674 87700 285680 87712
rect 249484 87672 285680 87700
rect 249484 87660 249490 87672
rect 285674 87660 285680 87672
rect 285732 87660 285738 87712
rect 286686 87660 286692 87712
rect 286744 87700 286750 87712
rect 502334 87700 502340 87712
rect 286744 87672 502340 87700
rect 286744 87660 286750 87672
rect 502334 87660 502340 87672
rect 502392 87660 502398 87712
rect 45462 87592 45468 87644
rect 45520 87632 45526 87644
rect 207566 87632 207572 87644
rect 45520 87604 207572 87632
rect 45520 87592 45526 87604
rect 207566 87592 207572 87604
rect 207624 87592 207630 87644
rect 230382 87592 230388 87644
rect 230440 87632 230446 87644
rect 240410 87632 240416 87644
rect 230440 87604 240416 87632
rect 230440 87592 230446 87604
rect 240410 87592 240416 87604
rect 240468 87592 240474 87644
rect 249518 87592 249524 87644
rect 249576 87632 249582 87644
rect 287054 87632 287060 87644
rect 249576 87604 287060 87632
rect 249576 87592 249582 87604
rect 287054 87592 287060 87604
rect 287112 87592 287118 87644
rect 289446 87592 289452 87644
rect 289504 87632 289510 87644
rect 528646 87632 528652 87644
rect 289504 87604 528652 87632
rect 289504 87592 289510 87604
rect 528646 87592 528652 87604
rect 528704 87592 528710 87644
rect 124122 86640 124128 86692
rect 124180 86680 124186 86692
rect 221182 86680 221188 86692
rect 124180 86652 221188 86680
rect 124180 86640 124186 86652
rect 221182 86640 221188 86652
rect 221240 86640 221246 86692
rect 255130 86640 255136 86692
rect 255188 86680 255194 86692
rect 311250 86680 311256 86692
rect 255188 86652 311256 86680
rect 255188 86640 255194 86652
rect 311250 86640 311256 86652
rect 311308 86640 311314 86692
rect 119982 86572 119988 86624
rect 120040 86612 120046 86624
rect 220446 86612 220452 86624
rect 120040 86584 220452 86612
rect 120040 86572 120046 86584
rect 220446 86572 220452 86584
rect 220504 86572 220510 86624
rect 256510 86572 256516 86624
rect 256568 86612 256574 86624
rect 324498 86612 324504 86624
rect 256568 86584 324504 86612
rect 256568 86572 256574 86584
rect 324498 86572 324504 86584
rect 324556 86572 324562 86624
rect 117222 86504 117228 86556
rect 117280 86544 117286 86556
rect 219986 86544 219992 86556
rect 117280 86516 219992 86544
rect 117280 86504 117286 86516
rect 219986 86504 219992 86516
rect 220044 86504 220050 86556
rect 253750 86504 253756 86556
rect 253808 86544 253814 86556
rect 309778 86544 309784 86556
rect 253808 86516 309784 86544
rect 253808 86504 253814 86516
rect 309778 86504 309784 86516
rect 309836 86504 309842 86556
rect 309870 86504 309876 86556
rect 309928 86544 309934 86556
rect 425054 86544 425060 86556
rect 309928 86516 425060 86544
rect 309928 86504 309934 86516
rect 425054 86504 425060 86516
rect 425112 86504 425118 86556
rect 111058 86436 111064 86488
rect 111116 86476 111122 86488
rect 218238 86476 218244 86488
rect 111116 86448 218244 86476
rect 111116 86436 111122 86448
rect 218238 86436 218244 86448
rect 218296 86436 218302 86488
rect 267366 86436 267372 86488
rect 267424 86476 267430 86488
rect 387794 86476 387800 86488
rect 267424 86448 387800 86476
rect 267424 86436 267430 86448
rect 387794 86436 387800 86448
rect 387852 86436 387858 86488
rect 107010 86368 107016 86420
rect 107068 86408 107074 86420
rect 216858 86408 216864 86420
rect 107068 86380 216864 86408
rect 107068 86368 107074 86380
rect 216858 86368 216864 86380
rect 216916 86368 216922 86420
rect 290826 86368 290832 86420
rect 290884 86408 290890 86420
rect 515398 86408 515404 86420
rect 290884 86380 515404 86408
rect 290884 86368 290890 86380
rect 515398 86368 515404 86380
rect 515456 86368 515462 86420
rect 88242 86300 88248 86352
rect 88300 86340 88306 86352
rect 211798 86340 211804 86352
rect 88300 86312 211804 86340
rect 88300 86300 88306 86312
rect 211798 86300 211804 86312
rect 211856 86300 211862 86352
rect 295150 86300 295156 86352
rect 295208 86340 295214 86352
rect 547874 86340 547880 86352
rect 295208 86312 547880 86340
rect 295208 86300 295214 86312
rect 547874 86300 547880 86312
rect 547932 86300 547938 86352
rect 10962 86232 10968 86284
rect 11020 86272 11026 86284
rect 201678 86272 201684 86284
rect 11020 86244 201684 86272
rect 11020 86232 11026 86244
rect 201678 86232 201684 86244
rect 201736 86232 201742 86284
rect 246390 86232 246396 86284
rect 246448 86272 246454 86284
rect 252554 86272 252560 86284
rect 246448 86244 252560 86272
rect 246448 86232 246454 86244
rect 252554 86232 252560 86244
rect 252612 86232 252618 86284
rect 296346 86232 296352 86284
rect 296404 86272 296410 86284
rect 572714 86272 572720 86284
rect 296404 86244 572720 86272
rect 296404 86232 296410 86244
rect 572714 86232 572720 86244
rect 572772 86232 572778 86284
rect 232498 85552 232504 85604
rect 232556 85592 232562 85604
rect 238846 85592 238852 85604
rect 232556 85564 238852 85592
rect 232556 85552 232562 85564
rect 238846 85552 238852 85564
rect 238904 85552 238910 85604
rect 3142 85484 3148 85536
rect 3200 85524 3206 85536
rect 14458 85524 14464 85536
rect 3200 85496 14464 85524
rect 3200 85484 3206 85496
rect 14458 85484 14464 85496
rect 14516 85484 14522 85536
rect 262950 85212 262956 85264
rect 263008 85252 263014 85264
rect 357434 85252 357440 85264
rect 263008 85224 357440 85252
rect 263008 85212 263014 85224
rect 357434 85212 357440 85224
rect 357492 85212 357498 85264
rect 187050 85144 187056 85196
rect 187108 85184 187114 85196
rect 229186 85184 229192 85196
rect 187108 85156 229192 85184
rect 187108 85144 187114 85156
rect 229186 85144 229192 85156
rect 229244 85144 229250 85196
rect 261846 85144 261852 85196
rect 261904 85184 261910 85196
rect 360194 85184 360200 85196
rect 261904 85156 360200 85184
rect 261904 85144 261910 85156
rect 360194 85144 360200 85156
rect 360252 85144 360258 85196
rect 184198 85076 184204 85128
rect 184256 85116 184262 85128
rect 231026 85116 231032 85128
rect 184256 85088 231032 85116
rect 184256 85076 184262 85088
rect 231026 85076 231032 85088
rect 231084 85076 231090 85128
rect 264330 85076 264336 85128
rect 264388 85116 264394 85128
rect 367094 85116 367100 85128
rect 264388 85088 367100 85116
rect 264388 85076 264394 85088
rect 367094 85076 367100 85088
rect 367152 85076 367158 85128
rect 119338 85008 119344 85060
rect 119396 85048 119402 85060
rect 219618 85048 219624 85060
rect 119396 85020 219624 85048
rect 119396 85008 119402 85020
rect 219618 85008 219624 85020
rect 219676 85008 219682 85060
rect 266078 85008 266084 85060
rect 266136 85048 266142 85060
rect 382274 85048 382280 85060
rect 266136 85020 382280 85048
rect 266136 85008 266142 85020
rect 382274 85008 382280 85020
rect 382332 85008 382338 85060
rect 68922 84940 68928 84992
rect 68980 84980 68986 84992
rect 211890 84980 211896 84992
rect 68980 84952 211896 84980
rect 68980 84940 68986 84952
rect 211890 84940 211896 84952
rect 211948 84940 211954 84992
rect 278406 84940 278412 84992
rect 278464 84980 278470 84992
rect 449158 84980 449164 84992
rect 278464 84952 449164 84980
rect 278464 84940 278470 84952
rect 449158 84940 449164 84952
rect 449216 84940 449222 84992
rect 50982 84872 50988 84924
rect 51040 84912 51046 84924
rect 208578 84912 208584 84924
rect 51040 84884 208584 84912
rect 51040 84872 51046 84884
rect 208578 84872 208584 84884
rect 208636 84872 208642 84924
rect 288158 84872 288164 84924
rect 288216 84912 288222 84924
rect 506474 84912 506480 84924
rect 288216 84884 506480 84912
rect 288216 84872 288222 84884
rect 506474 84872 506480 84884
rect 506532 84872 506538 84924
rect 15102 84804 15108 84856
rect 15160 84844 15166 84856
rect 201586 84844 201592 84856
rect 15160 84816 201592 84844
rect 15160 84804 15166 84816
rect 201586 84804 201592 84816
rect 201644 84804 201650 84856
rect 202230 84804 202236 84856
rect 202288 84844 202294 84856
rect 233050 84844 233056 84856
rect 202288 84816 233056 84844
rect 202288 84804 202294 84816
rect 233050 84804 233056 84816
rect 233108 84804 233114 84856
rect 243906 84804 243912 84856
rect 243964 84844 243970 84856
rect 258166 84844 258172 84856
rect 243964 84816 258172 84844
rect 243964 84804 243970 84816
rect 258166 84804 258172 84816
rect 258224 84804 258230 84856
rect 286778 84804 286784 84856
rect 286836 84844 286842 84856
rect 510706 84844 510712 84856
rect 286836 84816 510712 84844
rect 286836 84804 286842 84816
rect 510706 84804 510712 84816
rect 510764 84804 510770 84856
rect 191650 83784 191656 83836
rect 191708 83824 191714 83836
rect 232222 83824 232228 83836
rect 191708 83796 232228 83824
rect 191708 83784 191714 83796
rect 232222 83784 232228 83796
rect 232280 83784 232286 83836
rect 268838 83784 268844 83836
rect 268896 83824 268902 83836
rect 398926 83824 398932 83836
rect 268896 83796 398932 83824
rect 268896 83784 268902 83796
rect 398926 83784 398932 83796
rect 398984 83784 398990 83836
rect 182818 83716 182824 83768
rect 182876 83756 182882 83768
rect 225046 83756 225052 83768
rect 182876 83728 225052 83756
rect 182876 83716 182882 83728
rect 225046 83716 225052 83728
rect 225104 83716 225110 83768
rect 270126 83716 270132 83768
rect 270184 83756 270190 83768
rect 406378 83756 406384 83768
rect 270184 83728 406384 83756
rect 270184 83716 270190 83728
rect 406378 83716 406384 83728
rect 406436 83716 406442 83768
rect 111702 83648 111708 83700
rect 111760 83688 111766 83700
rect 218790 83688 218796 83700
rect 111760 83660 218796 83688
rect 111760 83648 111766 83660
rect 218790 83648 218796 83660
rect 218848 83648 218854 83700
rect 271598 83648 271604 83700
rect 271656 83688 271662 83700
rect 414014 83688 414020 83700
rect 271656 83660 414020 83688
rect 271656 83648 271662 83660
rect 414014 83648 414020 83660
rect 414072 83648 414078 83700
rect 103422 83580 103428 83632
rect 103480 83620 103486 83632
rect 216766 83620 216772 83632
rect 103480 83592 216772 83620
rect 103480 83580 103486 83592
rect 216766 83580 216772 83592
rect 216824 83580 216830 83632
rect 279510 83580 279516 83632
rect 279568 83620 279574 83632
rect 434714 83620 434720 83632
rect 279568 83592 434720 83620
rect 279568 83580 279574 83592
rect 434714 83580 434720 83592
rect 434772 83580 434778 83632
rect 96522 83512 96528 83564
rect 96580 83552 96586 83564
rect 216398 83552 216404 83564
rect 96580 83524 216404 83552
rect 96580 83512 96586 83524
rect 216398 83512 216404 83524
rect 216456 83512 216462 83564
rect 277118 83512 277124 83564
rect 277176 83552 277182 83564
rect 445754 83552 445760 83564
rect 277176 83524 445760 83552
rect 277176 83512 277182 83524
rect 445754 83512 445760 83524
rect 445812 83512 445818 83564
rect 89622 83444 89628 83496
rect 89680 83484 89686 83496
rect 213178 83484 213184 83496
rect 89680 83456 213184 83484
rect 89680 83444 89686 83456
rect 213178 83444 213184 83456
rect 213236 83444 213242 83496
rect 226978 83444 226984 83496
rect 227036 83484 227042 83496
rect 236546 83484 236552 83496
rect 227036 83456 236552 83484
rect 227036 83444 227042 83456
rect 236546 83444 236552 83456
rect 236604 83444 236610 83496
rect 297818 83444 297824 83496
rect 297876 83484 297882 83496
rect 571334 83484 571340 83496
rect 297876 83456 571340 83484
rect 297876 83444 297882 83456
rect 571334 83444 571340 83456
rect 571392 83444 571398 83496
rect 190362 82492 190368 82544
rect 190420 82532 190426 82544
rect 233878 82532 233884 82544
rect 190420 82504 233884 82532
rect 190420 82492 190426 82504
rect 233878 82492 233884 82504
rect 233936 82492 233942 82544
rect 175182 82424 175188 82476
rect 175240 82464 175246 82476
rect 229554 82464 229560 82476
rect 175240 82436 229560 82464
rect 175240 82424 175246 82436
rect 229554 82424 229560 82436
rect 229612 82424 229618 82476
rect 282638 82424 282644 82476
rect 282696 82464 282702 82476
rect 453298 82464 453304 82476
rect 282696 82436 453304 82464
rect 282696 82424 282702 82436
rect 453298 82424 453304 82436
rect 453356 82424 453362 82476
rect 168282 82356 168288 82408
rect 168340 82396 168346 82408
rect 224218 82396 224224 82408
rect 168340 82368 224224 82396
rect 168340 82356 168346 82368
rect 224218 82356 224224 82368
rect 224276 82356 224282 82408
rect 279970 82356 279976 82408
rect 280028 82396 280034 82408
rect 463694 82396 463700 82408
rect 280028 82368 463700 82396
rect 280028 82356 280034 82368
rect 463694 82356 463700 82368
rect 463752 82356 463758 82408
rect 170398 82288 170404 82340
rect 170456 82328 170462 82340
rect 226794 82328 226800 82340
rect 170456 82300 226800 82328
rect 170456 82288 170462 82300
rect 226794 82288 226800 82300
rect 226852 82288 226858 82340
rect 281258 82288 281264 82340
rect 281316 82328 281322 82340
rect 470594 82328 470600 82340
rect 281316 82300 470600 82328
rect 281316 82288 281322 82300
rect 470594 82288 470600 82300
rect 470652 82288 470658 82340
rect 136542 82220 136548 82272
rect 136600 82260 136606 82272
rect 222286 82260 222292 82272
rect 136600 82232 222292 82260
rect 136600 82220 136606 82232
rect 222286 82220 222292 82232
rect 222344 82220 222350 82272
rect 284110 82220 284116 82272
rect 284168 82260 284174 82272
rect 485774 82260 485780 82272
rect 284168 82232 485780 82260
rect 284168 82220 284174 82232
rect 485774 82220 485780 82232
rect 485832 82220 485838 82272
rect 106182 82152 106188 82204
rect 106240 82192 106246 82204
rect 214558 82192 214564 82204
rect 106240 82164 214564 82192
rect 106240 82152 106246 82164
rect 214558 82152 214564 82164
rect 214616 82152 214622 82204
rect 286870 82152 286876 82204
rect 286928 82192 286934 82204
rect 499574 82192 499580 82204
rect 286928 82164 499580 82192
rect 286928 82152 286934 82164
rect 499574 82152 499580 82164
rect 499632 82152 499638 82204
rect 47670 82084 47676 82136
rect 47728 82124 47734 82136
rect 206646 82124 206652 82136
rect 47728 82096 206652 82124
rect 47728 82084 47734 82096
rect 206646 82084 206652 82096
rect 206704 82084 206710 82136
rect 248138 82084 248144 82136
rect 248196 82124 248202 82136
rect 278774 82124 278780 82136
rect 248196 82096 278780 82124
rect 248196 82084 248202 82096
rect 278774 82084 278780 82096
rect 278832 82084 278838 82136
rect 290918 82084 290924 82136
rect 290976 82124 290982 82136
rect 525058 82124 525064 82136
rect 290976 82096 525064 82124
rect 290976 82084 290982 82096
rect 525058 82084 525064 82096
rect 525116 82084 525122 82136
rect 223482 81404 223488 81456
rect 223540 81444 223546 81456
rect 228450 81444 228456 81456
rect 223540 81416 228456 81444
rect 223540 81404 223546 81416
rect 228450 81404 228456 81416
rect 228508 81404 228514 81456
rect 253842 81064 253848 81116
rect 253900 81104 253906 81116
rect 307846 81104 307852 81116
rect 253900 81076 307852 81104
rect 253900 81064 253906 81076
rect 307846 81064 307852 81076
rect 307904 81064 307910 81116
rect 256602 80996 256608 81048
rect 256660 81036 256666 81048
rect 322934 81036 322940 81048
rect 256660 81008 322940 81036
rect 256660 80996 256666 81008
rect 322934 80996 322940 81008
rect 322992 80996 322998 81048
rect 272886 80928 272892 80980
rect 272944 80968 272950 80980
rect 411898 80968 411904 80980
rect 272944 80940 411904 80968
rect 272944 80928 272950 80940
rect 411898 80928 411904 80940
rect 411956 80928 411962 80980
rect 164142 80860 164148 80912
rect 164200 80900 164206 80912
rect 227990 80900 227996 80912
rect 164200 80872 227996 80900
rect 164200 80860 164206 80872
rect 227990 80860 227996 80872
rect 228048 80860 228054 80912
rect 292298 80860 292304 80912
rect 292356 80900 292362 80912
rect 535454 80900 535460 80912
rect 292356 80872 535460 80900
rect 292356 80860 292362 80872
rect 535454 80860 535460 80872
rect 535512 80860 535518 80912
rect 161382 80792 161388 80844
rect 161440 80832 161446 80844
rect 226702 80832 226708 80844
rect 161440 80804 226708 80832
rect 161440 80792 161446 80804
rect 226702 80792 226708 80804
rect 226760 80792 226766 80844
rect 240502 80792 240508 80844
rect 240560 80832 240566 80844
rect 252646 80832 252652 80844
rect 240560 80804 252652 80832
rect 240560 80792 240566 80804
rect 252646 80792 252652 80804
rect 252704 80792 252710 80844
rect 254578 80792 254584 80844
rect 254636 80832 254642 80844
rect 291194 80832 291200 80844
rect 254636 80804 291200 80832
rect 254636 80792 254642 80804
rect 291194 80792 291200 80804
rect 291252 80792 291258 80844
rect 293678 80792 293684 80844
rect 293736 80832 293742 80844
rect 542354 80832 542360 80844
rect 293736 80804 542360 80832
rect 293736 80792 293742 80804
rect 542354 80792 542360 80804
rect 542412 80792 542418 80844
rect 115842 80724 115848 80776
rect 115900 80764 115906 80776
rect 217318 80764 217324 80776
rect 115900 80736 217324 80764
rect 115900 80724 115906 80736
rect 217318 80724 217324 80736
rect 217376 80724 217382 80776
rect 250898 80724 250904 80776
rect 250956 80764 250962 80776
rect 295334 80764 295340 80776
rect 250956 80736 295340 80764
rect 250956 80724 250962 80736
rect 295334 80724 295340 80736
rect 295392 80724 295398 80776
rect 296530 80724 296536 80776
rect 296588 80764 296594 80776
rect 560294 80764 560300 80776
rect 296588 80736 560300 80764
rect 296588 80724 296594 80736
rect 560294 80724 560300 80736
rect 560352 80724 560358 80776
rect 98730 80656 98736 80708
rect 98788 80696 98794 80708
rect 215386 80696 215392 80708
rect 98788 80668 215392 80696
rect 98788 80656 98794 80668
rect 215386 80656 215392 80668
rect 215444 80656 215450 80708
rect 252186 80656 252192 80708
rect 252244 80696 252250 80708
rect 297450 80696 297456 80708
rect 252244 80668 297456 80696
rect 252244 80656 252250 80668
rect 297450 80656 297456 80668
rect 297508 80656 297514 80708
rect 297726 80656 297732 80708
rect 297784 80696 297790 80708
rect 578234 80696 578240 80708
rect 297784 80668 578240 80696
rect 297784 80656 297790 80668
rect 578234 80656 578240 80668
rect 578292 80656 578298 80708
rect 262858 79568 262864 79620
rect 262916 79608 262922 79620
rect 350534 79608 350540 79620
rect 262916 79580 350540 79608
rect 262916 79568 262922 79580
rect 350534 79568 350540 79580
rect 350592 79568 350598 79620
rect 119890 79500 119896 79552
rect 119948 79540 119954 79552
rect 219894 79540 219900 79552
rect 119948 79512 219900 79540
rect 119948 79500 119954 79512
rect 219894 79500 219900 79512
rect 219952 79500 219958 79552
rect 262030 79500 262036 79552
rect 262088 79540 262094 79552
rect 354674 79540 354680 79552
rect 262088 79512 354680 79540
rect 262088 79500 262094 79512
rect 354674 79500 354680 79512
rect 354732 79500 354738 79552
rect 113082 79432 113088 79484
rect 113140 79472 113146 79484
rect 218422 79472 218428 79484
rect 113140 79444 218428 79472
rect 113140 79432 113146 79444
rect 218422 79432 218428 79444
rect 218480 79432 218486 79484
rect 261938 79432 261944 79484
rect 261996 79472 262002 79484
rect 357526 79472 357532 79484
rect 261996 79444 357532 79472
rect 261996 79432 262002 79444
rect 357526 79432 357532 79444
rect 357584 79432 357590 79484
rect 86218 79364 86224 79416
rect 86276 79404 86282 79416
rect 208486 79404 208492 79416
rect 86276 79376 208492 79404
rect 86276 79364 86282 79376
rect 208486 79364 208492 79376
rect 208544 79364 208550 79416
rect 282546 79364 282552 79416
rect 282604 79404 282610 79416
rect 481634 79404 481640 79416
rect 282604 79376 481640 79404
rect 282604 79364 282610 79376
rect 481634 79364 481640 79376
rect 481692 79364 481698 79416
rect 75822 79296 75828 79348
rect 75880 79336 75886 79348
rect 212810 79336 212816 79348
rect 75880 79308 212816 79336
rect 75880 79296 75886 79308
rect 212810 79296 212816 79308
rect 212868 79296 212874 79348
rect 245194 79296 245200 79348
rect 245252 79336 245258 79348
rect 260834 79336 260840 79348
rect 245252 79308 260840 79336
rect 245252 79296 245258 79308
rect 260834 79296 260840 79308
rect 260892 79296 260898 79348
rect 299198 79296 299204 79348
rect 299256 79336 299262 79348
rect 582834 79336 582840 79348
rect 299256 79308 582840 79336
rect 299256 79296 299262 79308
rect 582834 79296 582840 79308
rect 582892 79296 582898 79348
rect 267458 78140 267464 78192
rect 267516 78180 267522 78192
rect 386414 78180 386420 78192
rect 267516 78152 386420 78180
rect 267516 78140 267522 78152
rect 386414 78140 386420 78152
rect 386472 78140 386478 78192
rect 257338 78072 257344 78124
rect 257396 78112 257402 78124
rect 266354 78112 266360 78124
rect 257396 78084 266360 78112
rect 257396 78072 257402 78084
rect 266354 78072 266360 78084
rect 266412 78072 266418 78124
rect 268930 78072 268936 78124
rect 268988 78112 268994 78124
rect 400214 78112 400220 78124
rect 268988 78084 400220 78112
rect 268988 78072 268994 78084
rect 400214 78072 400220 78084
rect 400272 78072 400278 78124
rect 251818 78004 251824 78056
rect 251876 78044 251882 78056
rect 262214 78044 262220 78056
rect 251876 78016 262220 78044
rect 251876 78004 251882 78016
rect 262214 78004 262220 78016
rect 262272 78004 262278 78056
rect 275278 78004 275284 78056
rect 275336 78044 275342 78056
rect 407206 78044 407212 78056
rect 275336 78016 407212 78044
rect 275336 78004 275342 78016
rect 407206 78004 407212 78016
rect 407264 78004 407270 78056
rect 42702 77936 42708 77988
rect 42760 77976 42766 77988
rect 207106 77976 207112 77988
rect 42760 77948 207112 77976
rect 42760 77936 42766 77948
rect 207106 77936 207112 77948
rect 207164 77936 207170 77988
rect 220722 77936 220728 77988
rect 220780 77976 220786 77988
rect 237466 77976 237472 77988
rect 220780 77948 237472 77976
rect 220780 77936 220786 77948
rect 237466 77936 237472 77948
rect 237524 77936 237530 77988
rect 243998 77936 244004 77988
rect 244056 77976 244062 77988
rect 267826 77976 267832 77988
rect 244056 77948 267832 77976
rect 244056 77936 244062 77948
rect 267826 77936 267832 77948
rect 267884 77936 267890 77988
rect 272978 77936 272984 77988
rect 273036 77976 273042 77988
rect 418154 77976 418160 77988
rect 273036 77948 418160 77976
rect 273036 77936 273042 77948
rect 418154 77936 418160 77948
rect 418212 77936 418218 77988
rect 172422 76916 172428 76968
rect 172480 76956 172486 76968
rect 222930 76956 222936 76968
rect 172480 76928 222936 76956
rect 172480 76916 172486 76928
rect 222930 76916 222936 76928
rect 222988 76916 222994 76968
rect 153010 76848 153016 76900
rect 153068 76888 153074 76900
rect 225322 76888 225328 76900
rect 153068 76860 225328 76888
rect 153068 76848 153074 76860
rect 225322 76848 225328 76860
rect 225380 76848 225386 76900
rect 144730 76780 144736 76832
rect 144788 76820 144794 76832
rect 223666 76820 223672 76832
rect 144788 76792 223672 76820
rect 144788 76780 144794 76792
rect 223666 76780 223672 76792
rect 223724 76780 223730 76832
rect 139302 76712 139308 76764
rect 139360 76752 139366 76764
rect 223850 76752 223856 76764
rect 139360 76724 223856 76752
rect 139360 76712 139366 76724
rect 223850 76712 223856 76724
rect 223908 76712 223914 76764
rect 278498 76712 278504 76764
rect 278556 76752 278562 76764
rect 432598 76752 432604 76764
rect 278556 76724 432604 76752
rect 278556 76712 278562 76724
rect 432598 76712 432604 76724
rect 432656 76712 432662 76764
rect 136450 76644 136456 76696
rect 136508 76684 136514 76696
rect 222654 76684 222660 76696
rect 136508 76656 222660 76684
rect 136508 76644 136514 76656
rect 222654 76644 222660 76656
rect 222712 76644 222718 76696
rect 277210 76644 277216 76696
rect 277268 76684 277274 76696
rect 436738 76684 436744 76696
rect 277268 76656 436744 76684
rect 277268 76644 277274 76656
rect 436738 76644 436744 76656
rect 436796 76644 436802 76696
rect 126790 76576 126796 76628
rect 126848 76616 126854 76628
rect 221458 76616 221464 76628
rect 126848 76588 221464 76616
rect 126848 76576 126854 76588
rect 221458 76576 221464 76588
rect 221516 76576 221522 76628
rect 246298 76576 246304 76628
rect 246356 76616 246362 76628
rect 251174 76616 251180 76628
rect 246356 76588 251180 76616
rect 246356 76576 246362 76588
rect 251174 76576 251180 76588
rect 251232 76576 251238 76628
rect 279418 76576 279424 76628
rect 279476 76616 279482 76628
rect 448606 76616 448612 76628
rect 279476 76588 448612 76616
rect 279476 76576 279482 76588
rect 448606 76576 448612 76588
rect 448664 76576 448670 76628
rect 17862 76508 17868 76560
rect 17920 76548 17926 76560
rect 200942 76548 200948 76560
rect 17920 76520 200948 76548
rect 17920 76508 17926 76520
rect 200942 76508 200948 76520
rect 201000 76508 201006 76560
rect 245286 76508 245292 76560
rect 245344 76548 245350 76560
rect 263594 76548 263600 76560
rect 245344 76520 263600 76548
rect 245344 76508 245350 76520
rect 263594 76508 263600 76520
rect 263652 76508 263658 76560
rect 296254 76508 296260 76560
rect 296312 76548 296318 76560
rect 569954 76548 569960 76560
rect 296312 76520 569960 76548
rect 296312 76508 296318 76520
rect 569954 76508 569960 76520
rect 570012 76508 570018 76560
rect 242526 75828 242532 75880
rect 242584 75868 242590 75880
rect 244274 75868 244280 75880
rect 242584 75840 244280 75868
rect 242584 75828 242590 75840
rect 244274 75828 244280 75840
rect 244332 75828 244338 75880
rect 260282 75420 260288 75472
rect 260340 75460 260346 75472
rect 336734 75460 336740 75472
rect 260340 75432 336740 75460
rect 260340 75420 260346 75432
rect 336734 75420 336740 75432
rect 336792 75420 336798 75472
rect 264238 75352 264244 75404
rect 264296 75392 264302 75404
rect 346394 75392 346400 75404
rect 264296 75364 346400 75392
rect 264296 75352 264302 75364
rect 346394 75352 346400 75364
rect 346452 75352 346458 75404
rect 282730 75284 282736 75336
rect 282788 75324 282794 75336
rect 481726 75324 481732 75336
rect 282788 75296 481732 75324
rect 282788 75284 282794 75296
rect 481726 75284 481732 75296
rect 481784 75284 481790 75336
rect 284202 75216 284208 75268
rect 284260 75256 284266 75268
rect 488534 75256 488540 75268
rect 284260 75228 488540 75256
rect 284260 75216 284266 75228
rect 488534 75216 488540 75228
rect 488592 75216 488598 75268
rect 245378 75148 245384 75200
rect 245436 75188 245442 75200
rect 269206 75188 269212 75200
rect 245436 75160 269212 75188
rect 245436 75148 245442 75160
rect 269206 75148 269212 75160
rect 269264 75148 269270 75200
rect 285214 75148 285220 75200
rect 285272 75188 285278 75200
rect 491294 75188 491300 75200
rect 285272 75160 491300 75188
rect 285272 75148 285278 75160
rect 491294 75148 491300 75160
rect 491352 75148 491358 75200
rect 273070 74128 273076 74180
rect 273128 74168 273134 74180
rect 420914 74168 420920 74180
rect 273128 74140 420920 74168
rect 273128 74128 273134 74140
rect 420914 74128 420920 74140
rect 420972 74128 420978 74180
rect 285306 74060 285312 74112
rect 285364 74100 285370 74112
rect 495434 74100 495440 74112
rect 285364 74072 495440 74100
rect 285364 74060 285370 74072
rect 495434 74060 495440 74072
rect 495492 74060 495498 74112
rect 99282 73992 99288 74044
rect 99340 74032 99346 74044
rect 215938 74032 215944 74044
rect 99340 74004 215944 74032
rect 99340 73992 99346 74004
rect 215938 73992 215944 74004
rect 215996 73992 216002 74044
rect 288250 73992 288256 74044
rect 288308 74032 288314 74044
rect 513374 74032 513380 74044
rect 288308 74004 513380 74032
rect 288308 73992 288314 74004
rect 513374 73992 513380 74004
rect 513432 73992 513438 74044
rect 85482 73924 85488 73976
rect 85540 73964 85546 73976
rect 214006 73964 214012 73976
rect 85540 73936 214012 73964
rect 85540 73924 85546 73936
rect 214006 73924 214012 73936
rect 214064 73924 214070 73976
rect 289538 73924 289544 73976
rect 289596 73964 289602 73976
rect 521654 73964 521660 73976
rect 289596 73936 521660 73964
rect 289596 73924 289602 73936
rect 521654 73924 521660 73936
rect 521712 73924 521718 73976
rect 48222 73856 48228 73908
rect 48280 73896 48286 73908
rect 202322 73896 202328 73908
rect 48280 73868 202328 73896
rect 48280 73856 48286 73868
rect 202322 73856 202328 73868
rect 202380 73856 202386 73908
rect 291010 73856 291016 73908
rect 291068 73896 291074 73908
rect 527174 73896 527180 73908
rect 291068 73868 527180 73896
rect 291068 73856 291074 73868
rect 527174 73856 527180 73868
rect 527232 73856 527238 73908
rect 31662 73788 31668 73840
rect 31720 73828 31726 73840
rect 205082 73828 205088 73840
rect 31720 73800 205088 73828
rect 31720 73788 31726 73800
rect 205082 73788 205088 73800
rect 205140 73788 205146 73840
rect 250990 73788 250996 73840
rect 251048 73828 251054 73840
rect 298094 73828 298100 73840
rect 251048 73800 298100 73828
rect 251048 73788 251054 73800
rect 298094 73788 298100 73800
rect 298152 73788 298158 73840
rect 299290 73788 299296 73840
rect 299348 73828 299354 73840
rect 582742 73828 582748 73840
rect 299348 73800 582748 73828
rect 299348 73788 299354 73800
rect 582742 73788 582748 73800
rect 582800 73788 582806 73840
rect 261754 72700 261760 72752
rect 261812 72740 261818 72752
rect 336090 72740 336096 72752
rect 261812 72712 336096 72740
rect 261812 72700 261818 72712
rect 336090 72700 336096 72712
rect 336148 72700 336154 72752
rect 263502 72632 263508 72684
rect 263560 72672 263566 72684
rect 364334 72672 364340 72684
rect 263560 72644 364340 72672
rect 263560 72632 263566 72644
rect 364334 72632 364340 72644
rect 364392 72632 364398 72684
rect 256050 72564 256056 72616
rect 256108 72604 256114 72616
rect 259454 72604 259460 72616
rect 256108 72576 259460 72604
rect 256108 72564 256114 72576
rect 259454 72564 259460 72576
rect 259512 72564 259518 72616
rect 276750 72564 276756 72616
rect 276808 72604 276814 72616
rect 396074 72604 396080 72616
rect 276808 72576 396080 72604
rect 276808 72564 276814 72576
rect 396074 72564 396080 72576
rect 396132 72564 396138 72616
rect 403618 72564 403624 72616
rect 403676 72604 403682 72616
rect 449894 72604 449900 72616
rect 403676 72576 449900 72604
rect 403676 72564 403682 72576
rect 449894 72564 449900 72576
rect 449952 72564 449958 72616
rect 274358 72496 274364 72548
rect 274416 72536 274422 72548
rect 427814 72536 427820 72548
rect 274416 72508 427820 72536
rect 274416 72496 274422 72508
rect 427814 72496 427820 72508
rect 427872 72496 427878 72548
rect 292390 72428 292396 72480
rect 292448 72468 292454 72480
rect 531406 72468 531412 72480
rect 292448 72440 531412 72468
rect 292448 72428 292454 72440
rect 531406 72428 531412 72440
rect 531464 72428 531470 72480
rect 3418 71680 3424 71732
rect 3476 71720 3482 71732
rect 35158 71720 35164 71732
rect 3476 71692 35164 71720
rect 3476 71680 3482 71692
rect 35158 71680 35164 71692
rect 35216 71680 35222 71732
rect 121362 71340 121368 71392
rect 121420 71380 121426 71392
rect 219802 71380 219808 71392
rect 121420 71352 219808 71380
rect 121420 71340 121426 71352
rect 219802 71340 219808 71352
rect 219860 71340 219866 71392
rect 64782 71272 64788 71324
rect 64840 71312 64846 71324
rect 209866 71312 209872 71324
rect 64840 71284 209872 71312
rect 64840 71272 64846 71284
rect 209866 71272 209872 71284
rect 209924 71272 209930 71324
rect 61930 71204 61936 71256
rect 61988 71244 61994 71256
rect 209958 71244 209964 71256
rect 61988 71216 209964 71244
rect 61988 71204 61994 71216
rect 209958 71204 209964 71216
rect 210016 71204 210022 71256
rect 267550 71204 267556 71256
rect 267608 71244 267614 71256
rect 389174 71244 389180 71256
rect 267608 71216 389180 71244
rect 267608 71204 267614 71216
rect 389174 71204 389180 71216
rect 389232 71204 389238 71256
rect 53650 71136 53656 71188
rect 53708 71176 53714 71188
rect 208854 71176 208860 71188
rect 53708 71148 208860 71176
rect 53708 71136 53714 71148
rect 208854 71136 208860 71148
rect 208912 71136 208918 71188
rect 270218 71136 270224 71188
rect 270276 71176 270282 71188
rect 402974 71176 402980 71188
rect 270276 71148 402980 71176
rect 270276 71136 270282 71148
rect 402974 71136 402980 71148
rect 403032 71136 403038 71188
rect 45370 71068 45376 71120
rect 45428 71108 45434 71120
rect 207290 71108 207296 71120
rect 45428 71080 207296 71108
rect 45428 71068 45434 71080
rect 207290 71068 207296 71080
rect 207348 71068 207354 71120
rect 271690 71068 271696 71120
rect 271748 71108 271754 71120
rect 409874 71108 409880 71120
rect 271748 71080 409880 71108
rect 271748 71068 271754 71080
rect 409874 71068 409880 71080
rect 409932 71068 409938 71120
rect 38562 71000 38568 71052
rect 38620 71040 38626 71052
rect 206002 71040 206008 71052
rect 38620 71012 206008 71040
rect 38620 71000 38626 71012
rect 206002 71000 206008 71012
rect 206060 71000 206066 71052
rect 248230 71000 248236 71052
rect 248288 71040 248294 71052
rect 266998 71040 267004 71052
rect 248288 71012 267004 71040
rect 248288 71000 248294 71012
rect 266998 71000 267004 71012
rect 267056 71000 267062 71052
rect 281350 71000 281356 71052
rect 281408 71040 281414 71052
rect 466454 71040 466460 71052
rect 281408 71012 466460 71040
rect 281408 71000 281414 71012
rect 466454 71000 466460 71012
rect 466512 71000 466518 71052
rect 259086 69980 259092 70032
rect 259144 70020 259150 70032
rect 340966 70020 340972 70032
rect 259144 69992 340972 70020
rect 259144 69980 259150 69992
rect 340966 69980 340972 69992
rect 341024 69980 341030 70032
rect 266170 69912 266176 69964
rect 266228 69952 266234 69964
rect 378778 69952 378784 69964
rect 266228 69924 378784 69952
rect 266228 69912 266234 69924
rect 378778 69912 378784 69924
rect 378836 69912 378842 69964
rect 274450 69844 274456 69896
rect 274508 69884 274514 69896
rect 431218 69884 431224 69896
rect 274508 69856 431224 69884
rect 274508 69844 274514 69856
rect 431218 69844 431224 69856
rect 431276 69844 431282 69896
rect 276658 69776 276664 69828
rect 276716 69816 276722 69828
rect 438854 69816 438860 69828
rect 276716 69788 438860 69816
rect 276716 69776 276722 69788
rect 438854 69776 438860 69788
rect 438912 69776 438918 69828
rect 278590 69708 278596 69760
rect 278648 69748 278654 69760
rect 456886 69748 456892 69760
rect 278648 69720 456892 69748
rect 278648 69708 278654 69720
rect 456886 69708 456892 69720
rect 456944 69708 456950 69760
rect 253198 69640 253204 69692
rect 253256 69680 253262 69692
rect 276106 69680 276112 69692
rect 253256 69652 276112 69680
rect 253256 69640 253262 69652
rect 276106 69640 276112 69652
rect 276164 69640 276170 69692
rect 280062 69640 280068 69692
rect 280120 69680 280126 69692
rect 459554 69680 459560 69692
rect 280120 69652 459560 69680
rect 280120 69640 280126 69652
rect 459554 69640 459560 69652
rect 459612 69640 459618 69692
rect 125410 68416 125416 68468
rect 125468 68456 125474 68468
rect 221274 68456 221280 68468
rect 125468 68428 221280 68456
rect 125468 68416 125474 68428
rect 221274 68416 221280 68428
rect 221332 68416 221338 68468
rect 20622 68348 20628 68400
rect 20680 68388 20686 68400
rect 203334 68388 203340 68400
rect 20680 68360 203340 68388
rect 20680 68348 20686 68360
rect 203334 68348 203340 68360
rect 203392 68348 203398 68400
rect 267274 68348 267280 68400
rect 267332 68388 267338 68400
rect 390646 68388 390652 68400
rect 267332 68360 390652 68388
rect 267332 68348 267338 68360
rect 390646 68348 390652 68360
rect 390704 68348 390710 68400
rect 6822 68280 6828 68332
rect 6880 68320 6886 68332
rect 201034 68320 201040 68332
rect 6880 68292 201040 68320
rect 6880 68280 6886 68292
rect 201034 68280 201040 68292
rect 201092 68280 201098 68332
rect 240318 68280 240324 68332
rect 240376 68320 240382 68332
rect 249886 68320 249892 68332
rect 240376 68292 249892 68320
rect 240376 68280 240382 68292
rect 249886 68280 249892 68292
rect 249944 68280 249950 68332
rect 275830 68280 275836 68332
rect 275888 68320 275894 68332
rect 436094 68320 436100 68332
rect 275888 68292 436100 68320
rect 275888 68280 275894 68292
rect 436094 68280 436100 68292
rect 436152 68280 436158 68332
rect 272794 66852 272800 66904
rect 272852 66892 272858 66904
rect 422294 66892 422300 66904
rect 272852 66864 422300 66892
rect 272852 66852 272858 66864
rect 422294 66852 422300 66864
rect 422352 66852 422358 66904
rect 285398 65492 285404 65544
rect 285456 65532 285462 65544
rect 492674 65532 492680 65544
rect 285456 65504 492680 65532
rect 285456 65492 285462 65504
rect 492674 65492 492680 65504
rect 492732 65492 492738 65544
rect 300670 64132 300676 64184
rect 300728 64172 300734 64184
rect 582650 64172 582656 64184
rect 300728 64144 582656 64172
rect 300728 64132 300734 64144
rect 582650 64132 582656 64144
rect 582708 64132 582714 64184
rect 275922 62772 275928 62824
rect 275980 62812 275986 62824
rect 440326 62812 440332 62824
rect 275980 62784 440332 62812
rect 275980 62772 275986 62784
rect 440326 62772 440332 62784
rect 440384 62772 440390 62824
rect 3050 59304 3056 59356
rect 3108 59344 3114 59356
rect 140038 59344 140044 59356
rect 3108 59316 140044 59344
rect 3108 59304 3114 59316
rect 140038 59304 140044 59316
rect 140096 59304 140102 59356
rect 274174 53048 274180 53100
rect 274232 53088 274238 53100
rect 429194 53088 429200 53100
rect 274232 53060 429200 53088
rect 274232 53048 274238 53060
rect 429194 53048 429200 53060
rect 429252 53048 429258 53100
rect 44082 51688 44088 51740
rect 44140 51728 44146 51740
rect 200758 51728 200764 51740
rect 44140 51700 200764 51728
rect 44140 51688 44146 51700
rect 200758 51688 200764 51700
rect 200816 51688 200822 51740
rect 246758 51688 246764 51740
rect 246816 51728 246822 51740
rect 273254 51728 273260 51740
rect 246816 51700 273260 51728
rect 246816 51688 246822 51700
rect 273254 51688 273260 51700
rect 273312 51688 273318 51740
rect 281442 51688 281448 51740
rect 281500 51728 281506 51740
rect 467834 51728 467840 51740
rect 281500 51700 467840 51728
rect 281500 51688 281506 51700
rect 467834 51688 467840 51700
rect 467892 51688 467898 51740
rect 71682 47540 71688 47592
rect 71740 47580 71746 47592
rect 211522 47580 211528 47592
rect 71740 47552 211528 47580
rect 71740 47540 71746 47552
rect 211522 47540 211528 47552
rect 211580 47540 211586 47592
rect 244090 47540 244096 47592
rect 244148 47580 244154 47592
rect 256694 47580 256700 47592
rect 244148 47552 256700 47580
rect 244148 47540 244154 47552
rect 256694 47540 256700 47552
rect 256752 47540 256758 47592
rect 257798 47540 257804 47592
rect 257856 47580 257862 47592
rect 332686 47580 332692 47592
rect 257856 47552 332692 47580
rect 257856 47540 257862 47552
rect 332686 47540 332692 47552
rect 332744 47540 332750 47592
rect 249610 46180 249616 46232
rect 249668 46220 249674 46232
rect 285766 46220 285772 46232
rect 249668 46192 285772 46220
rect 249668 46180 249674 46192
rect 285766 46180 285772 46192
rect 285824 46180 285830 46232
rect 286594 46180 286600 46232
rect 286652 46220 286658 46232
rect 503714 46220 503720 46232
rect 286652 46192 503720 46220
rect 286652 46180 286658 46192
rect 503714 46180 503720 46192
rect 503772 46180 503778 46232
rect 247678 45772 247684 45824
rect 247736 45812 247742 45824
rect 248414 45812 248420 45824
rect 247736 45784 248420 45812
rect 247736 45772 247742 45784
rect 248414 45772 248420 45784
rect 248472 45772 248478 45824
rect 3418 45500 3424 45552
rect 3476 45540 3482 45552
rect 106918 45540 106924 45552
rect 3476 45512 106924 45540
rect 3476 45500 3482 45512
rect 106918 45500 106924 45512
rect 106976 45500 106982 45552
rect 78582 43392 78588 43444
rect 78640 43432 78646 43444
rect 212902 43432 212908 43444
rect 78640 43404 212908 43432
rect 78640 43392 78646 43404
rect 212902 43392 212908 43404
rect 212960 43392 212966 43444
rect 213178 43392 213184 43444
rect 213236 43432 213242 43444
rect 236730 43432 236736 43444
rect 213236 43404 236736 43432
rect 213236 43392 213242 43404
rect 236730 43392 236736 43404
rect 236788 43392 236794 43444
rect 243814 42712 243820 42764
rect 243872 42752 243878 42764
rect 249794 42752 249800 42764
rect 243872 42724 249800 42752
rect 243872 42712 243878 42724
rect 249794 42712 249800 42724
rect 249852 42712 249858 42764
rect 219342 42032 219348 42084
rect 219400 42072 219406 42084
rect 231210 42072 231216 42084
rect 219400 42044 231216 42072
rect 219400 42032 219406 42044
rect 231210 42032 231216 42044
rect 231268 42032 231274 42084
rect 250438 42032 250444 42084
rect 250496 42072 250502 42084
rect 267734 42072 267740 42084
rect 250496 42044 267740 42072
rect 250496 42032 250502 42044
rect 267734 42032 267740 42044
rect 267792 42032 267798 42084
rect 269022 42032 269028 42084
rect 269080 42072 269086 42084
rect 397454 42072 397460 42084
rect 269080 42044 397460 42072
rect 269080 42032 269086 42044
rect 397454 42032 397460 42044
rect 397512 42032 397518 42084
rect 242618 41420 242624 41472
rect 242676 41460 242682 41472
rect 242894 41460 242900 41472
rect 242676 41432 242900 41460
rect 242676 41420 242682 41432
rect 242894 41420 242900 41432
rect 242952 41420 242958 41472
rect 292206 39312 292212 39364
rect 292264 39352 292270 39364
rect 300118 39352 300124 39364
rect 292264 39324 300124 39352
rect 292264 39312 292270 39324
rect 300118 39312 300124 39324
rect 300176 39312 300182 39364
rect 211798 35164 211804 35216
rect 211856 35204 211862 35216
rect 234706 35204 234712 35216
rect 211856 35176 234712 35204
rect 211856 35164 211862 35176
rect 234706 35164 234712 35176
rect 234764 35164 234770 35216
rect 300762 35164 300768 35216
rect 300820 35204 300826 35216
rect 582558 35204 582564 35216
rect 300820 35176 582564 35204
rect 300820 35164 300826 35176
rect 582558 35164 582564 35176
rect 582616 35164 582622 35216
rect 2866 33056 2872 33108
rect 2924 33096 2930 33108
rect 47578 33096 47584 33108
rect 2924 33068 47584 33096
rect 2924 33056 2930 33068
rect 47578 33056 47584 33068
rect 47636 33056 47642 33108
rect 242710 28908 242716 28960
rect 242768 28948 242774 28960
rect 245654 28948 245660 28960
rect 242768 28920 245660 28948
rect 242768 28908 242774 28920
rect 245654 28908 245660 28920
rect 245712 28908 245718 28960
rect 246850 28228 246856 28280
rect 246908 28268 246914 28280
rect 262858 28268 262864 28280
rect 246908 28240 262864 28268
rect 246908 28228 246914 28240
rect 262858 28228 262864 28240
rect 262916 28228 262922 28280
rect 46842 25508 46848 25560
rect 46900 25548 46906 25560
rect 86310 25548 86316 25560
rect 46900 25520 86316 25548
rect 46900 25508 46906 25520
rect 86310 25508 86316 25520
rect 86368 25508 86374 25560
rect 12250 24080 12256 24132
rect 12308 24120 12314 24132
rect 199378 24120 199384 24132
rect 12308 24092 199384 24120
rect 12308 24080 12314 24092
rect 199378 24080 199384 24092
rect 199436 24080 199442 24132
rect 291102 24080 291108 24132
rect 291160 24120 291166 24132
rect 528554 24120 528560 24132
rect 291160 24092 528560 24120
rect 291160 24080 291166 24092
rect 528554 24080 528560 24092
rect 528612 24080 528618 24132
rect 238938 23536 238944 23588
rect 238996 23576 239002 23588
rect 240226 23576 240232 23588
rect 238996 23548 240232 23576
rect 238996 23536 239002 23548
rect 240226 23536 240232 23548
rect 240284 23536 240290 23588
rect 238662 22720 238668 22772
rect 238720 22760 238726 22772
rect 241514 22760 241520 22772
rect 238720 22732 241520 22760
rect 238720 22720 238726 22732
rect 241514 22720 241520 22732
rect 241572 22720 241578 22772
rect 353938 22720 353944 22772
rect 353996 22760 354002 22772
rect 460934 22760 460940 22772
rect 353996 22732 460940 22760
rect 353996 22720 354002 22732
rect 460934 22720 460940 22732
rect 460992 22720 460998 22772
rect 238018 22040 238024 22092
rect 238076 22080 238082 22092
rect 240594 22080 240600 22092
rect 238076 22052 240600 22080
rect 238076 22040 238082 22052
rect 240594 22040 240600 22052
rect 240652 22040 240658 22092
rect 282822 21360 282828 21412
rect 282880 21400 282886 21412
rect 474734 21400 474740 21412
rect 282880 21372 474740 21400
rect 282880 21360 282886 21372
rect 474734 21360 474740 21372
rect 474792 21360 474798 21412
rect 3418 20612 3424 20664
rect 3476 20652 3482 20664
rect 98638 20652 98644 20664
rect 3476 20624 98644 20652
rect 3476 20612 3482 20624
rect 98638 20612 98644 20624
rect 98696 20612 98702 20664
rect 278682 19932 278688 19984
rect 278740 19972 278746 19984
rect 454034 19972 454040 19984
rect 278740 19944 454040 19972
rect 278740 19932 278746 19944
rect 454034 19932 454040 19944
rect 454092 19932 454098 19984
rect 33042 18572 33048 18624
rect 33100 18612 33106 18624
rect 204622 18612 204628 18624
rect 33100 18584 204628 18612
rect 33100 18572 33106 18584
rect 204622 18572 204628 18584
rect 204680 18572 204686 18624
rect 100662 17212 100668 17264
rect 100720 17252 100726 17264
rect 217042 17252 217048 17264
rect 100720 17224 217048 17252
rect 100720 17212 100726 17224
rect 217042 17212 217048 17224
rect 217100 17212 217106 17264
rect 277302 17212 277308 17264
rect 277360 17252 277366 17264
rect 442994 17252 443000 17264
rect 277360 17224 443000 17252
rect 277360 17212 277366 17224
rect 442994 17212 443000 17224
rect 443052 17212 443058 17264
rect 86862 15852 86868 15904
rect 86920 15892 86926 15904
rect 214742 15892 214748 15904
rect 86920 15864 214748 15892
rect 86920 15852 86926 15864
rect 214742 15852 214748 15864
rect 214800 15852 214806 15904
rect 293770 15852 293776 15904
rect 293828 15892 293834 15904
rect 546494 15892 546500 15904
rect 293828 15864 546500 15892
rect 293828 15852 293834 15864
rect 546494 15852 546500 15864
rect 546552 15852 546558 15904
rect 266262 14492 266268 14544
rect 266320 14532 266326 14544
rect 383562 14532 383568 14544
rect 266320 14504 383568 14532
rect 266320 14492 266326 14504
rect 383562 14492 383568 14504
rect 383620 14492 383626 14544
rect 289630 14424 289636 14476
rect 289688 14464 289694 14476
rect 517514 14464 517520 14476
rect 289688 14436 517520 14464
rect 289688 14424 289694 14436
rect 517514 14424 517520 14436
rect 517572 14424 517578 14476
rect 94498 13064 94504 13116
rect 94556 13104 94562 13116
rect 215754 13104 215760 13116
rect 94556 13076 215760 13104
rect 94556 13064 94562 13076
rect 215754 13064 215760 13076
rect 215812 13064 215818 13116
rect 217962 13064 217968 13116
rect 218020 13104 218026 13116
rect 236270 13104 236276 13116
rect 218020 13076 236276 13104
rect 218020 13064 218026 13076
rect 236270 13064 236276 13076
rect 236328 13064 236334 13116
rect 285490 13064 285496 13116
rect 285548 13104 285554 13116
rect 497090 13104 497096 13116
rect 285548 13076 497096 13104
rect 285548 13064 285554 13076
rect 497090 13064 497096 13076
rect 497148 13064 497154 13116
rect 260742 11840 260748 11892
rect 260800 11880 260806 11892
rect 348050 11880 348056 11892
rect 260800 11852 348056 11880
rect 260800 11840 260806 11852
rect 348050 11840 348056 11852
rect 348108 11840 348114 11892
rect 264790 11772 264796 11824
rect 264848 11812 264854 11824
rect 372890 11812 372896 11824
rect 264848 11784 372896 11812
rect 264848 11772 264854 11784
rect 372890 11772 372896 11784
rect 372948 11772 372954 11824
rect 398926 11772 398932 11824
rect 398984 11812 398990 11824
rect 400122 11812 400128 11824
rect 398984 11784 400128 11812
rect 398984 11772 398990 11784
rect 400122 11772 400128 11784
rect 400180 11772 400186 11824
rect 407206 11772 407212 11824
rect 407264 11812 407270 11824
rect 408402 11812 408408 11824
rect 407264 11784 408408 11812
rect 407264 11772 407270 11784
rect 408402 11772 408408 11784
rect 408460 11772 408466 11824
rect 37090 11704 37096 11756
rect 37148 11744 37154 11756
rect 101398 11744 101404 11756
rect 37148 11716 101404 11744
rect 37148 11704 37154 11716
rect 101398 11704 101404 11716
rect 101456 11704 101462 11756
rect 242894 11704 242900 11756
rect 242952 11744 242958 11756
rect 244090 11744 244096 11756
rect 242952 11716 244096 11744
rect 242952 11704 242958 11716
rect 244090 11704 244096 11716
rect 244148 11704 244154 11756
rect 251174 11704 251180 11756
rect 251232 11744 251238 11756
rect 252370 11744 252376 11756
rect 251232 11716 252376 11744
rect 251232 11704 251238 11716
rect 252370 11704 252376 11716
rect 252428 11704 252434 11756
rect 295978 11704 295984 11756
rect 296036 11744 296042 11756
rect 416774 11744 416780 11756
rect 296036 11716 416780 11744
rect 296036 11704 296042 11716
rect 416774 11704 416780 11716
rect 416832 11704 416838 11756
rect 423766 11704 423772 11756
rect 423824 11744 423830 11756
rect 424962 11744 424968 11756
rect 423824 11716 424968 11744
rect 423824 11704 423830 11716
rect 424962 11704 424968 11716
rect 425020 11704 425026 11756
rect 307846 11636 307852 11688
rect 307904 11676 307910 11688
rect 309042 11676 309048 11688
rect 307904 11648 309048 11676
rect 307904 11636 307910 11648
rect 309042 11636 309048 11648
rect 309100 11636 309106 11688
rect 332686 11636 332692 11688
rect 332744 11676 332750 11688
rect 333882 11676 333888 11688
rect 332744 11648 333888 11676
rect 332744 11636 332750 11648
rect 333882 11636 333888 11648
rect 333940 11636 333946 11688
rect 357526 11636 357532 11688
rect 357584 11676 357590 11688
rect 358722 11676 358728 11688
rect 357584 11648 358728 11676
rect 357584 11636 357590 11648
rect 358722 11636 358728 11648
rect 358780 11636 358786 11688
rect 216582 10276 216588 10328
rect 216640 10316 216646 10328
rect 222838 10316 222844 10328
rect 216640 10288 222844 10316
rect 216640 10276 216646 10288
rect 222838 10276 222844 10288
rect 222896 10276 222902 10328
rect 271414 10276 271420 10328
rect 271472 10316 271478 10328
rect 411806 10316 411812 10328
rect 271472 10288 411812 10316
rect 271472 10276 271478 10288
rect 411806 10276 411812 10288
rect 411864 10276 411870 10328
rect 461578 10276 461584 10328
rect 461636 10316 461642 10328
rect 472250 10316 472256 10328
rect 461636 10288 472256 10316
rect 461636 10276 461642 10288
rect 472250 10276 472256 10288
rect 472308 10276 472314 10328
rect 254854 9324 254860 9376
rect 254912 9364 254918 9376
rect 319714 9364 319720 9376
rect 254912 9336 319720 9364
rect 254912 9324 254918 9336
rect 319714 9324 319720 9336
rect 319772 9324 319778 9376
rect 264698 9256 264704 9308
rect 264756 9296 264762 9308
rect 374086 9296 374092 9308
rect 264756 9268 374092 9296
rect 264756 9256 264762 9268
rect 374086 9256 374092 9268
rect 374144 9256 374150 9308
rect 270310 9188 270316 9240
rect 270368 9228 270374 9240
rect 406010 9228 406016 9240
rect 270368 9200 406016 9228
rect 270368 9188 270374 9200
rect 406010 9188 406016 9200
rect 406068 9188 406074 9240
rect 294690 9120 294696 9172
rect 294748 9160 294754 9172
rect 459186 9160 459192 9172
rect 294748 9132 459192 9160
rect 294748 9120 294754 9132
rect 459186 9120 459192 9132
rect 459244 9120 459250 9172
rect 287974 9052 287980 9104
rect 288032 9092 288038 9104
rect 511258 9092 511264 9104
rect 288032 9064 511264 9092
rect 288032 9052 288038 9064
rect 511258 9052 511264 9064
rect 511316 9052 511322 9104
rect 289354 8984 289360 9036
rect 289412 9024 289418 9036
rect 520734 9024 520740 9036
rect 289412 8996 520740 9024
rect 289412 8984 289418 8996
rect 520734 8984 520740 8996
rect 520792 8984 520798 9036
rect 210970 8916 210976 8968
rect 211028 8956 211034 8968
rect 225598 8956 225604 8968
rect 211028 8928 225604 8956
rect 211028 8916 211034 8928
rect 225598 8916 225604 8928
rect 225656 8916 225662 8968
rect 299382 8916 299388 8968
rect 299440 8956 299446 8968
rect 576302 8956 576308 8968
rect 299440 8928 576308 8956
rect 299440 8916 299446 8928
rect 576302 8916 576308 8928
rect 576360 8916 576366 8968
rect 250806 7692 250812 7744
rect 250864 7732 250870 7744
rect 292574 7732 292580 7744
rect 250864 7704 292580 7732
rect 250864 7692 250870 7704
rect 292574 7692 292580 7704
rect 292632 7692 292638 7744
rect 260190 7624 260196 7676
rect 260248 7664 260254 7676
rect 331582 7664 331588 7676
rect 260248 7636 331588 7664
rect 260248 7624 260254 7636
rect 331582 7624 331588 7636
rect 331640 7624 331646 7676
rect 5258 7556 5264 7608
rect 5316 7596 5322 7608
rect 46198 7596 46204 7608
rect 5316 7568 46204 7596
rect 5316 7556 5322 7568
rect 46198 7556 46204 7568
rect 46256 7556 46262 7608
rect 260098 7556 260104 7608
rect 260156 7596 260162 7608
rect 270034 7596 270040 7608
rect 260156 7568 270040 7596
rect 260156 7556 260162 7568
rect 270034 7556 270040 7568
rect 270092 7556 270098 7608
rect 270402 7556 270408 7608
rect 270460 7596 270466 7608
rect 404814 7596 404820 7608
rect 270460 7568 404820 7596
rect 270460 7556 270466 7568
rect 404814 7556 404820 7568
rect 404872 7556 404878 7608
rect 454678 7556 454684 7608
rect 454736 7596 454742 7608
rect 465166 7596 465172 7608
rect 454736 7568 465172 7596
rect 454736 7556 454742 7568
rect 465166 7556 465172 7568
rect 465224 7556 465230 7608
rect 468478 7556 468484 7608
rect 468536 7596 468542 7608
rect 479334 7596 479340 7608
rect 468536 7568 479340 7596
rect 468536 7556 468542 7568
rect 479334 7556 479340 7568
rect 479392 7556 479398 7608
rect 3418 6808 3424 6860
rect 3476 6848 3482 6860
rect 133138 6848 133144 6860
rect 3476 6820 133144 6848
rect 3476 6808 3482 6820
rect 133138 6808 133144 6820
rect 133196 6808 133202 6860
rect 258718 6468 258724 6520
rect 258776 6508 258782 6520
rect 317322 6508 317328 6520
rect 258776 6480 317328 6508
rect 258776 6468 258782 6480
rect 317322 6468 317328 6480
rect 317380 6468 317386 6520
rect 294598 6400 294604 6452
rect 294656 6440 294662 6452
rect 370590 6440 370596 6452
rect 294656 6412 370596 6440
rect 294656 6400 294662 6412
rect 370590 6400 370596 6412
rect 370648 6400 370654 6452
rect 285582 6332 285588 6384
rect 285640 6372 285646 6384
rect 498194 6372 498200 6384
rect 285640 6344 498200 6372
rect 285640 6332 285646 6344
rect 498194 6332 498200 6344
rect 498252 6332 498258 6384
rect 245470 6264 245476 6316
rect 245528 6304 245534 6316
rect 259822 6304 259828 6316
rect 245528 6276 259828 6304
rect 245528 6264 245534 6276
rect 259822 6264 259828 6276
rect 259880 6264 259886 6316
rect 293494 6264 293500 6316
rect 293552 6304 293558 6316
rect 540790 6304 540796 6316
rect 293552 6276 540796 6304
rect 293552 6264 293558 6276
rect 540790 6264 540796 6276
rect 540848 6264 540854 6316
rect 248322 6196 248328 6248
rect 248380 6236 248386 6248
rect 280706 6236 280712 6248
rect 248380 6208 280712 6236
rect 248380 6196 248386 6208
rect 280706 6196 280712 6208
rect 280764 6196 280770 6248
rect 297358 6196 297364 6248
rect 297416 6236 297422 6248
rect 544378 6236 544384 6248
rect 297416 6208 544384 6236
rect 297416 6196 297422 6208
rect 544378 6196 544384 6208
rect 544436 6196 544442 6248
rect 249702 6128 249708 6180
rect 249760 6168 249766 6180
rect 286594 6168 286600 6180
rect 249760 6140 286600 6168
rect 249760 6128 249766 6140
rect 286594 6128 286600 6140
rect 286652 6128 286658 6180
rect 298738 6128 298744 6180
rect 298796 6168 298802 6180
rect 569126 6168 569132 6180
rect 298796 6140 569132 6168
rect 298796 6128 298802 6140
rect 569126 6128 569132 6140
rect 569184 6128 569190 6180
rect 281902 5516 281908 5568
rect 281960 5556 281966 5568
rect 283466 5556 283472 5568
rect 281960 5528 283472 5556
rect 281960 5516 281966 5528
rect 283466 5516 283472 5528
rect 283524 5516 283530 5568
rect 443638 5516 443644 5568
rect 443696 5556 443702 5568
rect 447410 5556 447416 5568
rect 443696 5528 447416 5556
rect 443696 5516 443702 5528
rect 447410 5516 447416 5528
rect 447468 5516 447474 5568
rect 59630 4836 59636 4888
rect 59688 4876 59694 4888
rect 93118 4876 93124 4888
rect 59688 4848 93124 4876
rect 59688 4836 59694 4848
rect 93118 4836 93124 4848
rect 93176 4836 93182 4888
rect 80882 4768 80888 4820
rect 80940 4808 80946 4820
rect 209038 4808 209044 4820
rect 80940 4780 209044 4808
rect 80940 4768 80946 4780
rect 209038 4768 209044 4780
rect 209096 4768 209102 4820
rect 233418 4428 233424 4480
rect 233476 4468 233482 4480
rect 239122 4468 239128 4480
rect 233476 4440 239128 4468
rect 233476 4428 233482 4440
rect 239122 4428 239128 4440
rect 239180 4428 239186 4480
rect 28902 4156 28908 4208
rect 28960 4196 28966 4208
rect 32398 4196 32404 4208
rect 28960 4168 32404 4196
rect 28960 4156 28966 4168
rect 32398 4156 32404 4168
rect 32456 4156 32462 4208
rect 242434 4156 242440 4208
rect 242492 4196 242498 4208
rect 246390 4196 246396 4208
rect 242492 4168 246396 4196
rect 242492 4156 242498 4168
rect 246390 4156 246396 4168
rect 246448 4156 246454 4208
rect 130562 4088 130568 4140
rect 130620 4128 130626 4140
rect 133230 4128 133236 4140
rect 130620 4100 133236 4128
rect 130620 4088 130626 4100
rect 133230 4088 133236 4100
rect 133288 4088 133294 4140
rect 161290 4088 161296 4140
rect 161348 4128 161354 4140
rect 162118 4128 162124 4140
rect 161348 4100 162124 4128
rect 161348 4088 161354 4100
rect 162118 4088 162124 4100
rect 162176 4088 162182 4140
rect 168374 4088 168380 4140
rect 168432 4128 168438 4140
rect 173158 4128 173164 4140
rect 168432 4100 173164 4128
rect 168432 4088 168438 4100
rect 173158 4088 173164 4100
rect 173216 4088 173222 4140
rect 290182 4088 290188 4140
rect 290240 4128 290246 4140
rect 298094 4128 298100 4140
rect 290240 4100 298100 4128
rect 290240 4088 290246 4100
rect 298094 4088 298100 4100
rect 298152 4088 298158 4140
rect 323578 4088 323584 4140
rect 323636 4128 323642 4140
rect 324406 4128 324412 4140
rect 323636 4100 324412 4128
rect 323636 4088 323642 4100
rect 324406 4088 324412 4100
rect 324464 4088 324470 4140
rect 402514 4088 402520 4140
rect 402572 4128 402578 4140
rect 403066 4128 403072 4140
rect 402572 4100 403072 4128
rect 402572 4088 402578 4100
rect 403066 4088 403072 4100
rect 403124 4088 403130 4140
rect 431218 4088 431224 4140
rect 431276 4128 431282 4140
rect 432046 4128 432052 4140
rect 431276 4100 432052 4128
rect 431276 4088 431282 4100
rect 432046 4088 432052 4100
rect 432104 4088 432110 4140
rect 363598 4020 363604 4072
rect 363656 4060 363662 4072
rect 365806 4060 365812 4072
rect 363656 4032 365812 4060
rect 363656 4020 363662 4032
rect 365806 4020 365812 4032
rect 365864 4020 365870 4072
rect 40770 3952 40776 4004
rect 40828 3992 40834 4004
rect 47670 3992 47676 4004
rect 40828 3964 47676 3992
rect 40828 3952 40834 3964
rect 47670 3952 47676 3964
rect 47728 3952 47734 4004
rect 101030 3952 101036 4004
rect 101088 3992 101094 4004
rect 104158 3992 104164 4004
rect 101088 3964 104164 3992
rect 101088 3952 101094 3964
rect 104158 3952 104164 3964
rect 104216 3952 104222 4004
rect 171778 3952 171784 4004
rect 171836 3992 171842 4004
rect 181530 3992 181536 4004
rect 171836 3964 181536 3992
rect 171836 3952 171842 3964
rect 181530 3952 181536 3964
rect 181588 3952 181594 4004
rect 193214 3952 193220 4004
rect 193272 3992 193278 4004
rect 202230 3992 202236 4004
rect 193272 3964 202236 3992
rect 193272 3952 193278 3964
rect 202230 3952 202236 3964
rect 202288 3952 202294 4004
rect 208578 3952 208584 4004
rect 208636 3992 208642 4004
rect 211798 3992 211804 4004
rect 208636 3964 211804 3992
rect 208636 3952 208642 3964
rect 211798 3952 211804 3964
rect 211856 3952 211862 4004
rect 171870 3884 171876 3936
rect 171928 3924 171934 3936
rect 182818 3924 182824 3936
rect 171928 3896 182824 3924
rect 171928 3884 171934 3896
rect 182818 3884 182824 3896
rect 182876 3884 182882 3936
rect 225138 3884 225144 3936
rect 225196 3924 225202 3936
rect 237650 3924 237656 3936
rect 225196 3896 237656 3924
rect 225196 3884 225202 3896
rect 237650 3884 237656 3896
rect 237708 3884 237714 3936
rect 320174 3924 320180 3936
rect 311866 3896 320180 3924
rect 131758 3816 131764 3868
rect 131816 3856 131822 3868
rect 137278 3856 137284 3868
rect 131816 3828 137284 3856
rect 131816 3816 131822 3828
rect 137278 3816 137284 3828
rect 137336 3816 137342 3868
rect 189718 3816 189724 3868
rect 189776 3856 189782 3868
rect 192478 3856 192484 3868
rect 189776 3828 192484 3856
rect 189776 3816 189782 3828
rect 192478 3816 192484 3828
rect 192536 3816 192542 3868
rect 226334 3816 226340 3868
rect 226392 3856 226398 3868
rect 232498 3856 232504 3868
rect 226392 3828 232504 3856
rect 226392 3816 226398 3828
rect 232498 3816 232504 3828
rect 232556 3816 232562 3868
rect 247586 3816 247592 3868
rect 247644 3856 247650 3868
rect 258074 3856 258080 3868
rect 247644 3828 258080 3856
rect 247644 3816 247650 3828
rect 258074 3816 258080 3828
rect 258132 3816 258138 3868
rect 64846 3760 74534 3788
rect 8754 3680 8760 3732
rect 8812 3720 8818 3732
rect 18598 3720 18604 3732
rect 8812 3692 18604 3720
rect 8812 3680 8818 3692
rect 18598 3680 18604 3692
rect 18656 3680 18662 3732
rect 35894 3680 35900 3732
rect 35952 3720 35958 3732
rect 39298 3720 39304 3732
rect 35952 3692 39304 3720
rect 35952 3680 35958 3692
rect 39298 3680 39304 3692
rect 39356 3680 39362 3732
rect 18230 3612 18236 3664
rect 18288 3652 18294 3664
rect 28258 3652 28264 3664
rect 18288 3624 28264 3652
rect 18288 3612 18294 3624
rect 28258 3612 28264 3624
rect 28316 3612 28322 3664
rect 43438 3652 43444 3664
rect 35866 3624 43444 3652
rect 1670 3544 1676 3596
rect 1728 3584 1734 3596
rect 4798 3584 4804 3596
rect 1728 3556 4804 3584
rect 1728 3544 1734 3556
rect 4798 3544 4804 3556
rect 4856 3544 4862 3596
rect 24210 3544 24216 3596
rect 24268 3584 24274 3596
rect 35866 3584 35894 3624
rect 43438 3612 43444 3624
rect 43496 3612 43502 3664
rect 56042 3612 56048 3664
rect 56100 3652 56106 3664
rect 64846 3652 64874 3760
rect 66714 3680 66720 3732
rect 66772 3720 66778 3732
rect 66772 3692 73292 3720
rect 66772 3680 66778 3692
rect 56100 3624 64874 3652
rect 56100 3612 56106 3624
rect 24268 3556 35894 3584
rect 24268 3544 24274 3556
rect 44266 3544 44272 3596
rect 44324 3584 44330 3596
rect 45370 3584 45376 3596
rect 44324 3556 45376 3584
rect 44324 3544 44330 3556
rect 45370 3544 45376 3556
rect 45428 3544 45434 3596
rect 52546 3544 52552 3596
rect 52604 3584 52610 3596
rect 53650 3584 53656 3596
rect 52604 3556 53656 3584
rect 52604 3544 52610 3556
rect 53650 3544 53656 3556
rect 53708 3544 53714 3596
rect 57238 3544 57244 3596
rect 57296 3584 57302 3596
rect 57882 3584 57888 3596
rect 57296 3556 57888 3584
rect 57296 3544 57302 3556
rect 57882 3544 57888 3556
rect 57940 3544 57946 3596
rect 58434 3544 58440 3596
rect 58492 3584 58498 3596
rect 59262 3584 59268 3596
rect 58492 3556 59268 3584
rect 58492 3544 58498 3556
rect 59262 3544 59268 3556
rect 59320 3544 59326 3596
rect 60826 3544 60832 3596
rect 60884 3584 60890 3596
rect 61930 3584 61936 3596
rect 60884 3556 61936 3584
rect 60884 3544 60890 3556
rect 61930 3544 61936 3556
rect 61988 3544 61994 3596
rect 65518 3544 65524 3596
rect 65576 3584 65582 3596
rect 66162 3584 66168 3596
rect 65576 3556 66168 3584
rect 65576 3544 65582 3556
rect 66162 3544 66168 3556
rect 66220 3544 66226 3596
rect 67910 3544 67916 3596
rect 67968 3584 67974 3596
rect 68922 3584 68928 3596
rect 67968 3556 68928 3584
rect 67968 3544 67974 3556
rect 68922 3544 68928 3556
rect 68980 3544 68986 3596
rect 72602 3544 72608 3596
rect 72660 3584 72666 3596
rect 73062 3584 73068 3596
rect 72660 3556 73068 3584
rect 72660 3544 72666 3556
rect 73062 3544 73068 3556
rect 73120 3544 73126 3596
rect 73264 3584 73292 3692
rect 74506 3652 74534 3760
rect 77386 3748 77392 3800
rect 77444 3788 77450 3800
rect 88978 3788 88984 3800
rect 77444 3760 88984 3788
rect 77444 3748 77450 3760
rect 88978 3748 88984 3760
rect 89036 3748 89042 3800
rect 103514 3748 103520 3800
rect 103572 3788 103578 3800
rect 107010 3788 107016 3800
rect 103572 3760 107016 3788
rect 103572 3748 103578 3760
rect 107010 3748 107016 3760
rect 107068 3748 107074 3800
rect 132954 3748 132960 3800
rect 133012 3788 133018 3800
rect 133012 3760 142154 3788
rect 133012 3748 133018 3760
rect 74902 3680 74908 3732
rect 74960 3720 74966 3732
rect 80698 3720 80704 3732
rect 74960 3692 80704 3720
rect 74960 3680 74966 3692
rect 80698 3680 80704 3692
rect 80756 3680 80762 3732
rect 86218 3720 86224 3732
rect 84166 3692 86224 3720
rect 84166 3652 84194 3692
rect 86218 3680 86224 3692
rect 86276 3680 86282 3732
rect 86770 3680 86776 3732
rect 86828 3720 86834 3732
rect 115106 3720 115112 3732
rect 86828 3692 115112 3720
rect 86828 3680 86834 3692
rect 115106 3680 115112 3692
rect 115164 3680 115170 3732
rect 137646 3720 137652 3732
rect 133984 3692 137652 3720
rect 101490 3652 101496 3664
rect 74506 3624 84194 3652
rect 84396 3624 101496 3652
rect 84396 3584 84424 3624
rect 101490 3612 101496 3624
rect 101548 3612 101554 3664
rect 122098 3652 122104 3664
rect 103716 3624 122104 3652
rect 73264 3556 84424 3584
rect 84470 3544 84476 3596
rect 84528 3584 84534 3596
rect 85482 3584 85488 3596
rect 84528 3556 85488 3584
rect 84528 3544 84534 3556
rect 85482 3544 85488 3556
rect 85540 3544 85546 3596
rect 89162 3544 89168 3596
rect 89220 3584 89226 3596
rect 89622 3584 89628 3596
rect 89220 3556 89628 3584
rect 89220 3544 89226 3556
rect 89622 3544 89628 3556
rect 89680 3544 89686 3596
rect 90358 3544 90364 3596
rect 90416 3584 90422 3596
rect 91002 3584 91008 3596
rect 90416 3556 91008 3584
rect 90416 3544 90422 3556
rect 91002 3544 91008 3556
rect 91060 3544 91066 3596
rect 91554 3544 91560 3596
rect 91612 3584 91618 3596
rect 92382 3584 92388 3596
rect 91612 3556 92388 3584
rect 91612 3544 91618 3556
rect 92382 3544 92388 3556
rect 92440 3544 92446 3596
rect 97442 3544 97448 3596
rect 97500 3584 97506 3596
rect 97902 3584 97908 3596
rect 97500 3556 97908 3584
rect 97500 3544 97506 3556
rect 97902 3544 97908 3556
rect 97960 3544 97966 3596
rect 98638 3544 98644 3596
rect 98696 3584 98702 3596
rect 99282 3584 99288 3596
rect 98696 3556 99288 3584
rect 98696 3544 98702 3556
rect 99282 3544 99288 3556
rect 99340 3544 99346 3596
rect 99834 3544 99840 3596
rect 99892 3584 99898 3596
rect 100662 3584 100668 3596
rect 99892 3556 100668 3584
rect 99892 3544 99898 3556
rect 100662 3544 100668 3556
rect 100720 3544 100726 3596
rect 102226 3544 102232 3596
rect 102284 3584 102290 3596
rect 103514 3584 103520 3596
rect 102284 3556 103520 3584
rect 102284 3544 102290 3556
rect 103514 3544 103520 3556
rect 103572 3544 103578 3596
rect 566 3476 572 3528
rect 624 3516 630 3528
rect 1302 3516 1308 3528
rect 624 3488 1308 3516
rect 624 3476 630 3488
rect 1302 3476 1308 3488
rect 1360 3476 1366 3528
rect 2866 3476 2872 3528
rect 2924 3516 2930 3528
rect 3970 3516 3976 3528
rect 2924 3488 3976 3516
rect 2924 3476 2930 3488
rect 3970 3476 3976 3488
rect 4028 3476 4034 3528
rect 9950 3476 9956 3528
rect 10008 3516 10014 3528
rect 10962 3516 10968 3528
rect 10008 3488 10968 3516
rect 10008 3476 10014 3488
rect 10962 3476 10968 3488
rect 11020 3476 11026 3528
rect 11146 3476 11152 3528
rect 11204 3516 11210 3528
rect 12250 3516 12256 3528
rect 11204 3488 12256 3516
rect 11204 3476 11210 3488
rect 12250 3476 12256 3488
rect 12308 3476 12314 3528
rect 13538 3476 13544 3528
rect 13596 3516 13602 3528
rect 35894 3516 35900 3528
rect 13596 3488 35900 3516
rect 13596 3476 13602 3488
rect 35894 3476 35900 3488
rect 35952 3476 35958 3528
rect 35986 3476 35992 3528
rect 36044 3516 36050 3528
rect 37090 3516 37096 3528
rect 36044 3488 37096 3516
rect 36044 3476 36050 3488
rect 37090 3476 37096 3488
rect 37148 3476 37154 3528
rect 41874 3476 41880 3528
rect 41932 3516 41938 3528
rect 42702 3516 42708 3528
rect 41932 3488 42708 3516
rect 41932 3476 41938 3488
rect 42702 3476 42708 3488
rect 42760 3476 42766 3528
rect 43070 3476 43076 3528
rect 43128 3516 43134 3528
rect 44082 3516 44088 3528
rect 43128 3488 44088 3516
rect 43128 3476 43134 3488
rect 44082 3476 44088 3488
rect 44140 3476 44146 3528
rect 48958 3476 48964 3528
rect 49016 3516 49022 3528
rect 49602 3516 49608 3528
rect 49016 3488 49608 3516
rect 49016 3476 49022 3488
rect 49602 3476 49608 3488
rect 49660 3476 49666 3528
rect 50154 3476 50160 3528
rect 50212 3516 50218 3528
rect 50982 3516 50988 3528
rect 50212 3488 50988 3516
rect 50212 3476 50218 3488
rect 50982 3476 50988 3488
rect 51040 3476 51046 3528
rect 51350 3476 51356 3528
rect 51408 3516 51414 3528
rect 74902 3516 74908 3528
rect 51408 3488 74908 3516
rect 51408 3476 51414 3488
rect 74902 3476 74908 3488
rect 74960 3476 74966 3528
rect 74994 3476 75000 3528
rect 75052 3516 75058 3528
rect 75822 3516 75828 3528
rect 75052 3488 75828 3516
rect 75052 3476 75058 3488
rect 75822 3476 75828 3488
rect 75880 3476 75886 3528
rect 76190 3476 76196 3528
rect 76248 3516 76254 3528
rect 77202 3516 77208 3528
rect 76248 3488 77208 3516
rect 76248 3476 76254 3488
rect 77202 3476 77208 3488
rect 77260 3476 77266 3528
rect 83274 3476 83280 3528
rect 83332 3516 83338 3528
rect 103716 3516 103744 3624
rect 122098 3612 122104 3624
rect 122156 3612 122162 3664
rect 125502 3612 125508 3664
rect 125560 3652 125566 3664
rect 125560 3624 132494 3652
rect 125560 3612 125566 3624
rect 110506 3544 110512 3596
rect 110564 3584 110570 3596
rect 111702 3584 111708 3596
rect 110564 3556 111708 3584
rect 110564 3544 110570 3556
rect 111702 3544 111708 3556
rect 111760 3544 111766 3596
rect 117590 3544 117596 3596
rect 117648 3584 117654 3596
rect 119338 3584 119344 3596
rect 117648 3556 119344 3584
rect 117648 3544 117654 3556
rect 119338 3544 119344 3556
rect 119396 3544 119402 3596
rect 128170 3544 128176 3596
rect 128228 3584 128234 3596
rect 132466 3584 132494 3624
rect 133984 3584 134012 3692
rect 137646 3680 137652 3692
rect 137704 3680 137710 3732
rect 142126 3720 142154 3760
rect 158898 3748 158904 3800
rect 158956 3788 158962 3800
rect 170398 3788 170404 3800
rect 158956 3760 170404 3788
rect 158956 3748 158962 3760
rect 170398 3748 170404 3760
rect 170456 3748 170462 3800
rect 171106 3760 172008 3788
rect 159358 3720 159364 3732
rect 142126 3692 159364 3720
rect 159358 3680 159364 3692
rect 159416 3680 159422 3732
rect 162486 3680 162492 3732
rect 162544 3720 162550 3732
rect 171106 3720 171134 3760
rect 162544 3692 171134 3720
rect 171980 3720 172008 3760
rect 173158 3748 173164 3800
rect 173216 3788 173222 3800
rect 187050 3788 187056 3800
rect 173216 3760 187056 3788
rect 173216 3748 173222 3760
rect 187050 3748 187056 3760
rect 187108 3748 187114 3800
rect 190362 3748 190368 3800
rect 190420 3788 190426 3800
rect 199102 3788 199108 3800
rect 190420 3760 199108 3788
rect 190420 3748 190426 3760
rect 199102 3748 199108 3760
rect 199160 3748 199166 3800
rect 200022 3748 200028 3800
rect 200080 3788 200086 3800
rect 203886 3788 203892 3800
rect 200080 3760 203892 3788
rect 200080 3748 200086 3760
rect 203886 3748 203892 3760
rect 203944 3748 203950 3800
rect 220446 3748 220452 3800
rect 220504 3788 220510 3800
rect 231118 3788 231124 3800
rect 220504 3760 231124 3788
rect 220504 3748 220510 3760
rect 231118 3748 231124 3760
rect 231176 3748 231182 3800
rect 262858 3748 262864 3800
rect 262916 3788 262922 3800
rect 271230 3788 271236 3800
rect 262916 3760 271236 3788
rect 262916 3748 262922 3760
rect 271230 3748 271236 3760
rect 271288 3748 271294 3800
rect 181438 3720 181444 3732
rect 171980 3692 181444 3720
rect 162544 3680 162550 3692
rect 181438 3680 181444 3692
rect 181496 3680 181502 3732
rect 218054 3680 218060 3732
rect 218112 3720 218118 3732
rect 219342 3720 219348 3732
rect 218112 3692 219348 3720
rect 218112 3680 218118 3692
rect 219342 3680 219348 3692
rect 219400 3680 219406 3732
rect 238110 3680 238116 3732
rect 238168 3720 238174 3732
rect 249886 3720 249892 3732
rect 238168 3692 249892 3720
rect 238168 3680 238174 3692
rect 249886 3680 249892 3692
rect 249944 3680 249950 3732
rect 258258 3680 258264 3732
rect 258316 3720 258322 3732
rect 269206 3720 269212 3732
rect 258316 3692 269212 3720
rect 258316 3680 258322 3692
rect 269206 3680 269212 3692
rect 269264 3680 269270 3732
rect 310238 3680 310244 3732
rect 310296 3720 310302 3732
rect 311866 3720 311894 3896
rect 320174 3884 320180 3896
rect 320232 3884 320238 3936
rect 326430 3884 326436 3936
rect 326488 3924 326494 3936
rect 326488 3896 326752 3924
rect 326488 3884 326494 3896
rect 310296 3692 311894 3720
rect 316696 3828 326660 3856
rect 310296 3680 310302 3692
rect 145926 3612 145932 3664
rect 145984 3652 145990 3664
rect 145984 3624 149100 3652
rect 145984 3612 145990 3624
rect 128228 3556 130516 3584
rect 132466 3556 134012 3584
rect 128228 3544 128234 3556
rect 83332 3488 103744 3516
rect 83332 3476 83338 3488
rect 104526 3476 104532 3528
rect 104584 3516 104590 3528
rect 105538 3516 105544 3528
rect 104584 3488 105544 3516
rect 104584 3476 104590 3488
rect 105538 3476 105544 3488
rect 105596 3476 105602 3528
rect 105722 3476 105728 3528
rect 105780 3516 105786 3528
rect 106182 3516 106188 3528
rect 105780 3488 106188 3516
rect 105780 3476 105786 3488
rect 106182 3476 106188 3488
rect 106240 3476 106246 3528
rect 108114 3476 108120 3528
rect 108172 3516 108178 3528
rect 108942 3516 108948 3528
rect 108172 3488 108948 3516
rect 108172 3476 108178 3488
rect 108942 3476 108948 3488
rect 109000 3476 109006 3528
rect 109310 3476 109316 3528
rect 109368 3516 109374 3528
rect 111058 3516 111064 3528
rect 109368 3488 111064 3516
rect 109368 3476 109374 3488
rect 111058 3476 111064 3488
rect 111116 3476 111122 3528
rect 111610 3476 111616 3528
rect 111668 3516 111674 3528
rect 112438 3516 112444 3528
rect 111668 3488 112444 3516
rect 111668 3476 111674 3488
rect 112438 3476 112444 3488
rect 112496 3476 112502 3528
rect 114002 3476 114008 3528
rect 114060 3516 114066 3528
rect 114462 3516 114468 3528
rect 114060 3488 114468 3516
rect 114060 3476 114066 3488
rect 114462 3476 114468 3488
rect 114520 3476 114526 3528
rect 115198 3476 115204 3528
rect 115256 3516 115262 3528
rect 115842 3516 115848 3528
rect 115256 3488 115848 3516
rect 115256 3476 115262 3488
rect 115842 3476 115848 3488
rect 115900 3476 115906 3528
rect 116394 3476 116400 3528
rect 116452 3516 116458 3528
rect 117222 3516 117228 3528
rect 116452 3488 117228 3516
rect 116452 3476 116458 3488
rect 117222 3476 117228 3488
rect 117280 3476 117286 3528
rect 118786 3476 118792 3528
rect 118844 3516 118850 3528
rect 119798 3516 119804 3528
rect 118844 3488 119804 3516
rect 118844 3476 118850 3488
rect 119798 3476 119804 3488
rect 119856 3476 119862 3528
rect 122282 3476 122288 3528
rect 122340 3516 122346 3528
rect 122742 3516 122748 3528
rect 122340 3488 122748 3516
rect 122340 3476 122346 3488
rect 122742 3476 122748 3488
rect 122800 3476 122806 3528
rect 123478 3476 123484 3528
rect 123536 3516 123542 3528
rect 124122 3516 124128 3528
rect 123536 3488 124128 3516
rect 123536 3476 123542 3488
rect 124122 3476 124128 3488
rect 124180 3476 124186 3528
rect 124674 3476 124680 3528
rect 124732 3516 124738 3528
rect 125410 3516 125416 3528
rect 124732 3488 125416 3516
rect 124732 3476 124738 3488
rect 125410 3476 125416 3488
rect 125468 3476 125474 3528
rect 125870 3476 125876 3528
rect 125928 3516 125934 3528
rect 126790 3516 126796 3528
rect 125928 3488 126796 3516
rect 125928 3476 125934 3488
rect 126790 3476 126796 3488
rect 126848 3476 126854 3528
rect 129366 3476 129372 3528
rect 129424 3516 129430 3528
rect 130378 3516 130384 3528
rect 129424 3488 130384 3516
rect 129424 3476 129430 3488
rect 130378 3476 130384 3488
rect 130436 3476 130442 3528
rect 130488 3516 130516 3556
rect 134150 3544 134156 3596
rect 134208 3584 134214 3596
rect 135162 3584 135168 3596
rect 134208 3556 135168 3584
rect 134208 3544 134214 3556
rect 135162 3544 135168 3556
rect 135220 3544 135226 3596
rect 138842 3544 138848 3596
rect 138900 3584 138906 3596
rect 139302 3584 139308 3596
rect 138900 3556 139308 3584
rect 138900 3544 138906 3556
rect 139302 3544 139308 3556
rect 139360 3544 139366 3596
rect 141234 3544 141240 3596
rect 141292 3584 141298 3596
rect 142062 3584 142068 3596
rect 141292 3556 142068 3584
rect 141292 3544 141298 3556
rect 142062 3544 142068 3556
rect 142120 3544 142126 3596
rect 143534 3544 143540 3596
rect 143592 3584 143598 3596
rect 144822 3584 144828 3596
rect 143592 3556 144828 3584
rect 143592 3544 143598 3556
rect 144822 3544 144828 3556
rect 144880 3544 144886 3596
rect 148318 3544 148324 3596
rect 148376 3584 148382 3596
rect 148962 3584 148968 3596
rect 148376 3556 148968 3584
rect 148376 3544 148382 3556
rect 148962 3544 148968 3556
rect 149020 3544 149026 3596
rect 149072 3584 149100 3624
rect 149514 3612 149520 3664
rect 149572 3652 149578 3664
rect 171778 3652 171784 3664
rect 149572 3624 171784 3652
rect 149572 3612 149578 3624
rect 171778 3612 171784 3624
rect 171836 3612 171842 3664
rect 193122 3612 193128 3664
rect 193180 3652 193186 3664
rect 193180 3624 195376 3652
rect 193180 3612 193186 3624
rect 171870 3584 171876 3596
rect 149072 3556 171876 3584
rect 171870 3544 171876 3556
rect 171928 3544 171934 3596
rect 171962 3544 171968 3596
rect 172020 3584 172026 3596
rect 172422 3584 172428 3596
rect 172020 3556 172428 3584
rect 172020 3544 172026 3556
rect 172422 3544 172428 3556
rect 172480 3544 172486 3596
rect 178678 3584 178684 3596
rect 174188 3556 178684 3584
rect 174188 3516 174216 3556
rect 178678 3544 178684 3556
rect 178736 3544 178742 3596
rect 195238 3584 195244 3596
rect 180766 3556 195244 3584
rect 130488 3488 174216 3516
rect 174262 3476 174268 3528
rect 174320 3516 174326 3528
rect 175182 3516 175188 3528
rect 174320 3488 175188 3516
rect 174320 3476 174326 3488
rect 175182 3476 175188 3488
rect 175240 3476 175246 3528
rect 179046 3476 179052 3528
rect 179104 3516 179110 3528
rect 180058 3516 180064 3528
rect 179104 3488 180064 3516
rect 179104 3476 179110 3488
rect 180058 3476 180064 3488
rect 180116 3476 180122 3528
rect 180242 3476 180248 3528
rect 180300 3516 180306 3528
rect 180766 3516 180794 3556
rect 195238 3544 195244 3556
rect 195296 3544 195302 3596
rect 195348 3584 195376 3624
rect 197262 3612 197268 3664
rect 197320 3652 197326 3664
rect 207382 3652 207388 3664
rect 197320 3624 207388 3652
rect 197320 3612 197326 3624
rect 207382 3612 207388 3624
rect 207440 3612 207446 3664
rect 213362 3612 213368 3664
rect 213420 3652 213426 3664
rect 226978 3652 226984 3664
rect 213420 3624 226984 3652
rect 213420 3612 213426 3624
rect 226978 3612 226984 3624
rect 227036 3612 227042 3664
rect 233878 3652 233884 3664
rect 229066 3624 233884 3652
rect 205082 3584 205088 3596
rect 195348 3556 205088 3584
rect 205082 3544 205088 3556
rect 205140 3544 205146 3596
rect 219250 3544 219256 3596
rect 219308 3584 219314 3596
rect 229066 3584 229094 3624
rect 233878 3612 233884 3624
rect 233936 3612 233942 3664
rect 239306 3612 239312 3664
rect 239364 3652 239370 3664
rect 252646 3652 252652 3664
rect 239364 3624 252652 3652
rect 239364 3612 239370 3624
rect 252646 3612 252652 3624
rect 252704 3612 252710 3664
rect 254670 3612 254676 3664
rect 254728 3652 254734 3664
rect 267826 3652 267832 3664
rect 254728 3624 267832 3652
rect 254728 3612 254734 3624
rect 267826 3612 267832 3624
rect 267884 3612 267890 3664
rect 268470 3612 268476 3664
rect 268528 3652 268534 3664
rect 316696 3652 316724 3828
rect 318150 3748 318156 3800
rect 318208 3788 318214 3800
rect 318208 3760 321692 3788
rect 318208 3748 318214 3760
rect 268528 3624 316724 3652
rect 268528 3612 268534 3624
rect 233602 3584 233608 3596
rect 219308 3556 229094 3584
rect 230768 3556 233608 3584
rect 219308 3544 219314 3556
rect 180300 3488 180794 3516
rect 180300 3476 180306 3488
rect 182542 3476 182548 3528
rect 182600 3516 182606 3528
rect 183462 3516 183468 3528
rect 182600 3488 183468 3516
rect 182600 3476 182606 3488
rect 183462 3476 183468 3488
rect 183520 3476 183526 3528
rect 183738 3476 183744 3528
rect 183796 3516 183802 3528
rect 184842 3516 184848 3528
rect 183796 3488 184848 3516
rect 183796 3476 183802 3488
rect 184842 3476 184848 3488
rect 184900 3476 184906 3528
rect 184934 3476 184940 3528
rect 184992 3516 184998 3528
rect 186222 3516 186228 3528
rect 184992 3488 186228 3516
rect 184992 3476 184998 3488
rect 186222 3476 186228 3488
rect 186280 3476 186286 3528
rect 187326 3476 187332 3528
rect 187384 3516 187390 3528
rect 188338 3516 188344 3528
rect 187384 3488 188344 3516
rect 187384 3476 187390 3488
rect 188338 3476 188344 3488
rect 188396 3476 188402 3528
rect 188522 3476 188528 3528
rect 188580 3516 188586 3528
rect 188982 3516 188988 3528
rect 188580 3488 188988 3516
rect 188580 3476 188586 3488
rect 188982 3476 188988 3488
rect 189040 3476 189046 3528
rect 190822 3476 190828 3528
rect 190880 3516 190886 3528
rect 191650 3516 191656 3528
rect 190880 3488 191656 3516
rect 190880 3476 190886 3488
rect 191650 3476 191656 3488
rect 191708 3476 191714 3528
rect 197906 3476 197912 3528
rect 197964 3516 197970 3528
rect 198642 3516 198648 3528
rect 197964 3488 198648 3516
rect 197964 3476 197970 3488
rect 198642 3476 198648 3488
rect 198700 3476 198706 3528
rect 200298 3476 200304 3528
rect 200356 3516 200362 3528
rect 201402 3516 201408 3528
rect 200356 3488 201408 3516
rect 200356 3476 200362 3488
rect 201402 3476 201408 3488
rect 201460 3476 201466 3528
rect 201494 3476 201500 3528
rect 201552 3516 201558 3528
rect 230768 3516 230796 3556
rect 233602 3544 233608 3556
rect 233660 3544 233666 3596
rect 245562 3544 245568 3596
rect 245620 3584 245626 3596
rect 265342 3584 265348 3596
rect 245620 3556 265348 3584
rect 245620 3544 245626 3556
rect 265342 3544 265348 3556
rect 265400 3544 265406 3596
rect 266998 3544 267004 3596
rect 267056 3584 267062 3596
rect 277118 3584 277124 3596
rect 267056 3556 277124 3584
rect 267056 3544 267062 3556
rect 277118 3544 277124 3556
rect 277176 3544 277182 3596
rect 296070 3544 296076 3596
rect 296128 3584 296134 3596
rect 303706 3584 303712 3596
rect 296128 3556 303712 3584
rect 296128 3544 296134 3556
rect 303706 3544 303712 3556
rect 303764 3544 303770 3596
rect 311158 3544 311164 3596
rect 311216 3584 311222 3596
rect 321664 3584 321692 3760
rect 326632 3652 326660 3828
rect 326724 3720 326752 3896
rect 331858 3884 331864 3936
rect 331916 3924 331922 3936
rect 517606 3924 517612 3936
rect 331916 3896 345014 3924
rect 331916 3884 331922 3896
rect 327718 3816 327724 3868
rect 327776 3856 327782 3868
rect 344554 3856 344560 3868
rect 327776 3828 344560 3856
rect 327776 3816 327782 3828
rect 344554 3816 344560 3828
rect 344612 3816 344618 3868
rect 336090 3748 336096 3800
rect 336148 3788 336154 3800
rect 344986 3788 345014 3896
rect 509206 3896 517612 3924
rect 449158 3816 449164 3868
rect 449216 3856 449222 3868
rect 453298 3856 453304 3868
rect 449216 3828 453304 3856
rect 449216 3816 449222 3828
rect 453298 3816 453304 3828
rect 453356 3816 453362 3868
rect 349246 3788 349252 3800
rect 336148 3760 336412 3788
rect 344986 3760 349252 3788
rect 336148 3748 336154 3760
rect 336274 3720 336280 3732
rect 326724 3692 336280 3720
rect 336274 3680 336280 3692
rect 336332 3680 336338 3732
rect 336384 3720 336412 3760
rect 349246 3748 349252 3760
rect 349304 3748 349310 3800
rect 416774 3748 416780 3800
rect 416832 3788 416838 3800
rect 417878 3788 417884 3800
rect 416832 3760 417884 3788
rect 416832 3748 416838 3760
rect 417878 3748 417884 3760
rect 417936 3748 417942 3800
rect 436738 3748 436744 3800
rect 436796 3788 436802 3800
rect 445018 3788 445024 3800
rect 436796 3760 445024 3788
rect 436796 3748 436802 3760
rect 445018 3748 445024 3760
rect 445076 3748 445082 3800
rect 450630 3748 450636 3800
rect 450688 3788 450694 3800
rect 458082 3788 458088 3800
rect 450688 3760 458088 3788
rect 450688 3748 450694 3760
rect 458082 3748 458088 3760
rect 458140 3748 458146 3800
rect 506474 3748 506480 3800
rect 506532 3788 506538 3800
rect 509206 3788 509234 3896
rect 517606 3884 517612 3896
rect 517664 3884 517670 3936
rect 575106 3884 575112 3936
rect 575164 3924 575170 3936
rect 582834 3924 582840 3936
rect 575164 3896 582840 3924
rect 575164 3884 575170 3896
rect 582834 3884 582840 3896
rect 582892 3884 582898 3936
rect 515398 3816 515404 3868
rect 515456 3856 515462 3868
rect 525426 3856 525432 3868
rect 515456 3828 525432 3856
rect 515456 3816 515462 3828
rect 525426 3816 525432 3828
rect 525484 3816 525490 3868
rect 566826 3816 566832 3868
rect 566884 3856 566890 3868
rect 571334 3856 571340 3868
rect 566884 3828 571340 3856
rect 566884 3816 566890 3828
rect 571334 3816 571340 3828
rect 571392 3816 571398 3868
rect 572714 3816 572720 3868
rect 572772 3856 572778 3868
rect 583294 3856 583300 3868
rect 572772 3828 583300 3856
rect 572772 3816 572778 3828
rect 583294 3816 583300 3828
rect 583352 3816 583358 3868
rect 506532 3760 509234 3788
rect 506532 3748 506538 3760
rect 517146 3748 517152 3800
rect 517204 3788 517210 3800
rect 517204 3760 523724 3788
rect 517204 3748 517210 3760
rect 362310 3720 362316 3732
rect 336384 3692 362316 3720
rect 362310 3680 362316 3692
rect 362368 3680 362374 3732
rect 409874 3680 409880 3732
rect 409932 3720 409938 3732
rect 410794 3720 410800 3732
rect 409932 3692 410800 3720
rect 409932 3680 409938 3692
rect 410794 3680 410800 3692
rect 410852 3680 410858 3732
rect 411898 3680 411904 3732
rect 411956 3720 411962 3732
rect 423766 3720 423772 3732
rect 411956 3692 423772 3720
rect 411956 3680 411962 3692
rect 423766 3680 423772 3692
rect 423824 3680 423830 3732
rect 432598 3680 432604 3732
rect 432656 3720 432662 3732
rect 452102 3720 452108 3732
rect 432656 3692 452108 3720
rect 432656 3680 432662 3692
rect 452102 3680 452108 3692
rect 452160 3680 452166 3732
rect 453390 3680 453396 3732
rect 453448 3720 453454 3732
rect 478138 3720 478144 3732
rect 453448 3692 478144 3720
rect 453448 3680 453454 3692
rect 478138 3680 478144 3692
rect 478196 3680 478202 3732
rect 499390 3680 499396 3732
rect 499448 3720 499454 3732
rect 510706 3720 510712 3732
rect 499448 3692 510712 3720
rect 499448 3680 499454 3692
rect 510706 3680 510712 3692
rect 510764 3680 510770 3732
rect 515950 3680 515956 3732
rect 516008 3720 516014 3732
rect 518894 3720 518900 3732
rect 516008 3692 518900 3720
rect 516008 3680 516014 3692
rect 518894 3680 518900 3692
rect 518952 3680 518958 3732
rect 523696 3720 523724 3760
rect 525058 3748 525064 3800
rect 525116 3788 525122 3800
rect 531314 3788 531320 3800
rect 525116 3760 531320 3788
rect 525116 3748 525122 3760
rect 531314 3748 531320 3760
rect 531372 3748 531378 3800
rect 556154 3748 556160 3800
rect 556212 3788 556218 3800
rect 568574 3788 568580 3800
rect 556212 3760 568580 3788
rect 556212 3748 556218 3760
rect 568574 3748 568580 3760
rect 568632 3748 568638 3800
rect 570322 3748 570328 3800
rect 570380 3788 570386 3800
rect 583202 3788 583208 3800
rect 570380 3760 583208 3788
rect 570380 3748 570386 3760
rect 583202 3748 583208 3760
rect 583260 3748 583266 3800
rect 528646 3720 528652 3732
rect 523696 3692 528652 3720
rect 528646 3680 528652 3692
rect 528704 3680 528710 3732
rect 534902 3680 534908 3732
rect 534960 3720 534966 3732
rect 546586 3720 546592 3732
rect 534960 3692 546592 3720
rect 534960 3680 534966 3692
rect 546586 3680 546592 3692
rect 546644 3680 546650 3732
rect 563238 3680 563244 3732
rect 563296 3720 563302 3732
rect 575566 3720 575572 3732
rect 563296 3692 575572 3720
rect 563296 3680 563302 3692
rect 575566 3680 575572 3692
rect 575624 3680 575630 3732
rect 371694 3652 371700 3664
rect 326632 3624 371700 3652
rect 371694 3612 371700 3624
rect 371752 3612 371758 3664
rect 374638 3612 374644 3664
rect 374696 3652 374702 3664
rect 384758 3652 384764 3664
rect 374696 3624 384764 3652
rect 374696 3612 374702 3624
rect 384758 3612 384764 3624
rect 384816 3612 384822 3664
rect 385678 3612 385684 3664
rect 385736 3652 385742 3664
rect 455690 3652 455696 3664
rect 385736 3624 455696 3652
rect 385736 3612 385742 3624
rect 455690 3612 455696 3624
rect 455748 3612 455754 3664
rect 475470 3612 475476 3664
rect 475528 3652 475534 3664
rect 487614 3652 487620 3664
rect 475528 3624 487620 3652
rect 475528 3612 475534 3624
rect 487614 3612 487620 3624
rect 487672 3612 487678 3664
rect 491110 3612 491116 3664
rect 491168 3652 491174 3664
rect 494054 3652 494060 3664
rect 491168 3624 494060 3652
rect 491168 3612 491174 3624
rect 494054 3612 494060 3624
rect 494112 3612 494118 3664
rect 497458 3612 497464 3664
rect 497516 3652 497522 3664
rect 523034 3652 523040 3664
rect 497516 3624 523040 3652
rect 497516 3612 497522 3624
rect 523034 3612 523040 3624
rect 523092 3612 523098 3664
rect 524230 3612 524236 3664
rect 524288 3652 524294 3664
rect 536834 3652 536840 3664
rect 524288 3624 536840 3652
rect 524288 3612 524294 3624
rect 536834 3612 536840 3624
rect 536892 3612 536898 3664
rect 541986 3612 541992 3664
rect 542044 3652 542050 3664
rect 554774 3652 554780 3664
rect 542044 3624 554780 3652
rect 542044 3612 542050 3624
rect 554774 3612 554780 3624
rect 554832 3612 554838 3664
rect 557350 3612 557356 3664
rect 557408 3652 557414 3664
rect 569954 3652 569960 3664
rect 557408 3624 569960 3652
rect 557408 3612 557414 3624
rect 569954 3612 569960 3624
rect 570012 3612 570018 3664
rect 571518 3612 571524 3664
rect 571576 3652 571582 3664
rect 583478 3652 583484 3664
rect 571576 3624 583484 3652
rect 571576 3612 571582 3624
rect 583478 3612 583484 3624
rect 583536 3612 583542 3664
rect 332686 3584 332692 3596
rect 311216 3556 311894 3584
rect 321664 3556 332692 3584
rect 311216 3544 311222 3556
rect 201552 3488 230796 3516
rect 201552 3476 201558 3488
rect 231026 3476 231032 3528
rect 231084 3516 231090 3528
rect 231762 3516 231768 3528
rect 231084 3488 231768 3516
rect 231084 3476 231090 3488
rect 231762 3476 231768 3488
rect 231820 3476 231826 3528
rect 232222 3476 232228 3528
rect 232280 3516 232286 3528
rect 233142 3516 233148 3528
rect 232280 3488 233148 3516
rect 232280 3476 232286 3488
rect 233142 3476 233148 3488
rect 233200 3476 233206 3528
rect 237006 3476 237012 3528
rect 237064 3516 237070 3528
rect 238018 3516 238024 3528
rect 237064 3488 238024 3516
rect 237064 3476 237070 3488
rect 238018 3476 238024 3488
rect 238076 3476 238082 3528
rect 246942 3476 246948 3528
rect 247000 3516 247006 3528
rect 272426 3516 272432 3528
rect 247000 3488 272432 3516
rect 247000 3476 247006 3488
rect 272426 3476 272432 3488
rect 272484 3476 272490 3528
rect 278314 3476 278320 3528
rect 278372 3516 278378 3528
rect 278774 3516 278780 3528
rect 278372 3488 278780 3516
rect 278372 3476 278378 3488
rect 278774 3476 278780 3488
rect 278832 3476 278838 3528
rect 279510 3476 279516 3528
rect 279568 3516 279574 3528
rect 281534 3516 281540 3528
rect 279568 3488 281540 3516
rect 279568 3476 279574 3488
rect 281534 3476 281540 3488
rect 281592 3476 281598 3528
rect 284294 3476 284300 3528
rect 284352 3516 284358 3528
rect 285766 3516 285772 3528
rect 284352 3488 285772 3516
rect 284352 3476 284358 3488
rect 285766 3476 285772 3488
rect 285824 3476 285830 3528
rect 294874 3476 294880 3528
rect 294932 3516 294938 3528
rect 295334 3516 295340 3528
rect 294932 3488 295340 3516
rect 294932 3476 294938 3488
rect 295334 3476 295340 3488
rect 295392 3476 295398 3528
rect 297450 3476 297456 3528
rect 297508 3516 297514 3528
rect 298462 3516 298468 3528
rect 297508 3488 298468 3516
rect 297508 3476 297514 3488
rect 298462 3476 298468 3488
rect 298520 3476 298526 3528
rect 300762 3476 300768 3528
rect 300820 3516 300826 3528
rect 309134 3516 309140 3528
rect 300820 3488 309140 3516
rect 300820 3476 300826 3488
rect 309134 3476 309140 3488
rect 309192 3476 309198 3528
rect 309778 3476 309784 3528
rect 309836 3516 309842 3528
rect 311434 3516 311440 3528
rect 309836 3488 311440 3516
rect 309836 3476 309842 3488
rect 311434 3476 311440 3488
rect 311492 3476 311498 3528
rect 311866 3516 311894 3556
rect 332686 3544 332692 3556
rect 332744 3544 332750 3596
rect 341518 3544 341524 3596
rect 341576 3584 341582 3596
rect 469858 3584 469864 3596
rect 341576 3556 469864 3584
rect 341576 3544 341582 3556
rect 469858 3544 469864 3556
rect 469916 3544 469922 3596
rect 472618 3544 472624 3596
rect 472676 3584 472682 3596
rect 473446 3584 473452 3596
rect 472676 3556 473452 3584
rect 472676 3544 472682 3556
rect 473446 3544 473452 3556
rect 473504 3544 473510 3596
rect 481634 3544 481640 3596
rect 481692 3584 481698 3596
rect 482830 3584 482836 3596
rect 481692 3556 482836 3584
rect 481692 3544 481698 3556
rect 482830 3544 482836 3556
rect 482888 3544 482894 3596
rect 489178 3544 489184 3596
rect 489236 3584 489242 3596
rect 510062 3584 510068 3596
rect 489236 3556 510068 3584
rect 489236 3544 489242 3556
rect 510062 3544 510068 3556
rect 510120 3544 510126 3596
rect 519538 3544 519544 3596
rect 519596 3584 519602 3596
rect 520366 3584 520372 3596
rect 519596 3556 520372 3584
rect 519596 3544 519602 3556
rect 520366 3544 520372 3556
rect 520424 3544 520430 3596
rect 522298 3544 522304 3596
rect 522356 3584 522362 3596
rect 550266 3584 550272 3596
rect 522356 3556 550272 3584
rect 522356 3544 522362 3556
rect 550266 3544 550272 3556
rect 550324 3544 550330 3596
rect 552658 3544 552664 3596
rect 552716 3584 552722 3596
rect 564342 3584 564348 3596
rect 552716 3556 564348 3584
rect 552716 3544 552722 3556
rect 564342 3544 564348 3556
rect 564400 3544 564406 3596
rect 564434 3544 564440 3596
rect 564492 3584 564498 3596
rect 578234 3584 578240 3596
rect 564492 3556 578240 3584
rect 564492 3544 564498 3556
rect 578234 3544 578240 3556
rect 578292 3544 578298 3596
rect 363506 3516 363512 3528
rect 311866 3488 363512 3516
rect 363506 3476 363512 3488
rect 363564 3476 363570 3528
rect 364978 3476 364984 3528
rect 365036 3516 365042 3528
rect 367002 3516 367008 3528
rect 365036 3488 367008 3516
rect 365036 3476 365042 3488
rect 367002 3476 367008 3488
rect 367060 3476 367066 3528
rect 370498 3476 370504 3528
rect 370556 3516 370562 3528
rect 551462 3516 551468 3528
rect 370556 3488 551468 3516
rect 370556 3476 370562 3488
rect 551462 3476 551468 3488
rect 551520 3476 551526 3528
rect 559742 3476 559748 3528
rect 559800 3516 559806 3528
rect 572806 3516 572812 3528
rect 559800 3488 572812 3516
rect 559800 3476 559806 3488
rect 572806 3476 572812 3488
rect 572864 3476 572870 3528
rect 574094 3516 574100 3528
rect 572916 3488 574100 3516
rect 4062 3408 4068 3460
rect 4120 3448 4126 3460
rect 15838 3448 15844 3460
rect 4120 3420 15844 3448
rect 4120 3408 4126 3420
rect 15838 3408 15844 3420
rect 15896 3408 15902 3460
rect 17034 3408 17040 3460
rect 17092 3448 17098 3460
rect 17862 3448 17868 3460
rect 17092 3420 17868 3448
rect 17092 3408 17098 3420
rect 17862 3408 17868 3420
rect 17920 3408 17926 3460
rect 19426 3408 19432 3460
rect 19484 3448 19490 3460
rect 20622 3448 20628 3460
rect 19484 3420 20628 3448
rect 19484 3408 19490 3420
rect 20622 3408 20628 3420
rect 20680 3408 20686 3460
rect 25314 3408 25320 3460
rect 25372 3448 25378 3460
rect 26142 3448 26148 3460
rect 25372 3420 26148 3448
rect 25372 3408 25378 3420
rect 26142 3408 26148 3420
rect 26200 3408 26206 3460
rect 26510 3408 26516 3460
rect 26568 3448 26574 3460
rect 27522 3448 27528 3460
rect 26568 3420 27528 3448
rect 26568 3408 26574 3420
rect 27522 3408 27528 3420
rect 27580 3408 27586 3460
rect 32398 3408 32404 3460
rect 32456 3448 32462 3460
rect 33042 3448 33048 3460
rect 32456 3420 33048 3448
rect 32456 3408 32462 3420
rect 33042 3408 33048 3420
rect 33100 3408 33106 3460
rect 33594 3408 33600 3460
rect 33652 3448 33658 3460
rect 34422 3448 34428 3460
rect 33652 3420 34428 3448
rect 33652 3408 33658 3420
rect 34422 3408 34428 3420
rect 34480 3408 34486 3460
rect 203242 3448 203248 3460
rect 35866 3420 203248 3448
rect 35866 3380 35894 3420
rect 203242 3408 203248 3420
rect 203300 3408 203306 3460
rect 213914 3408 213920 3460
rect 213972 3448 213978 3460
rect 214466 3448 214472 3460
rect 213972 3420 214472 3448
rect 213972 3408 213978 3420
rect 214466 3408 214472 3420
rect 214524 3408 214530 3460
rect 216858 3408 216864 3460
rect 216916 3448 216922 3460
rect 217962 3448 217968 3460
rect 216916 3420 217968 3448
rect 216916 3408 216922 3420
rect 217962 3408 217968 3420
rect 218020 3408 218026 3460
rect 218072 3420 219434 3448
rect 20640 3352 35894 3380
rect 20640 3324 20668 3352
rect 92750 3340 92756 3392
rect 92808 3380 92814 3392
rect 94498 3380 94504 3392
rect 92808 3352 94504 3380
rect 92808 3340 92814 3352
rect 94498 3340 94504 3352
rect 94556 3340 94562 3392
rect 153102 3340 153108 3392
rect 153160 3380 153166 3392
rect 154206 3380 154212 3392
rect 153160 3352 154212 3380
rect 153160 3340 153166 3352
rect 154206 3340 154212 3352
rect 154264 3340 154270 3392
rect 155402 3340 155408 3392
rect 155460 3380 155466 3392
rect 155862 3380 155868 3392
rect 155460 3352 155868 3380
rect 155460 3340 155466 3352
rect 155862 3340 155868 3352
rect 155920 3340 155926 3392
rect 157794 3340 157800 3392
rect 157852 3380 157858 3392
rect 158622 3380 158628 3392
rect 157852 3352 158628 3380
rect 157852 3340 157858 3352
rect 158622 3340 158628 3352
rect 158680 3340 158686 3392
rect 163682 3340 163688 3392
rect 163740 3380 163746 3392
rect 164142 3380 164148 3392
rect 163740 3352 164148 3380
rect 163740 3340 163746 3352
rect 164142 3340 164148 3352
rect 164200 3340 164206 3392
rect 164878 3340 164884 3392
rect 164936 3380 164942 3392
rect 165522 3380 165528 3392
rect 164936 3352 165528 3380
rect 164936 3340 164942 3352
rect 165522 3340 165528 3352
rect 165580 3340 165586 3392
rect 166074 3340 166080 3392
rect 166132 3380 166138 3392
rect 166902 3380 166908 3392
rect 166132 3352 166908 3380
rect 166132 3340 166138 3352
rect 166902 3340 166908 3352
rect 166960 3340 166966 3392
rect 167178 3340 167184 3392
rect 167236 3380 167242 3392
rect 168282 3380 168288 3392
rect 167236 3352 168288 3380
rect 167236 3340 167242 3352
rect 168282 3340 168288 3352
rect 168340 3340 168346 3392
rect 181438 3340 181444 3392
rect 181496 3380 181502 3392
rect 184198 3380 184204 3392
rect 181496 3352 184204 3380
rect 181496 3340 181502 3352
rect 184198 3340 184204 3352
rect 184256 3340 184262 3392
rect 212166 3340 212172 3392
rect 212224 3380 212230 3392
rect 218072 3380 218100 3420
rect 212224 3352 218100 3380
rect 219406 3380 219434 3420
rect 220722 3408 220728 3460
rect 220780 3448 220786 3460
rect 221550 3448 221556 3460
rect 220780 3420 221556 3448
rect 220780 3408 220786 3420
rect 221550 3408 221556 3420
rect 221608 3408 221614 3460
rect 222746 3408 222752 3460
rect 222804 3448 222810 3460
rect 223482 3448 223488 3460
rect 222804 3420 223488 3448
rect 222804 3408 222810 3420
rect 223482 3408 223488 3420
rect 223540 3408 223546 3460
rect 223942 3408 223948 3460
rect 224000 3448 224006 3460
rect 224862 3448 224868 3460
rect 224000 3420 224868 3448
rect 224000 3408 224006 3420
rect 224862 3408 224868 3420
rect 224920 3408 224926 3460
rect 229830 3408 229836 3460
rect 229888 3448 229894 3460
rect 240226 3448 240232 3460
rect 229888 3420 240232 3448
rect 229888 3408 229894 3420
rect 240226 3408 240232 3420
rect 240284 3408 240290 3460
rect 242894 3408 242900 3460
rect 242952 3448 242958 3460
rect 245654 3448 245660 3460
rect 242952 3420 245660 3448
rect 242952 3408 242958 3420
rect 245654 3408 245660 3420
rect 245712 3408 245718 3460
rect 249058 3408 249064 3460
rect 249116 3448 249122 3460
rect 274818 3448 274824 3460
rect 249116 3420 274824 3448
rect 249116 3408 249122 3420
rect 274818 3408 274824 3420
rect 274876 3408 274882 3460
rect 275278 3408 275284 3460
rect 275336 3448 275342 3460
rect 288986 3448 288992 3460
rect 275336 3420 288992 3448
rect 275336 3408 275342 3420
rect 288986 3408 288992 3420
rect 289044 3408 289050 3460
rect 300118 3408 300124 3460
rect 300176 3448 300182 3460
rect 537202 3448 537208 3460
rect 300176 3420 537208 3448
rect 300176 3408 300182 3420
rect 537202 3408 537208 3420
rect 537260 3408 537266 3460
rect 554958 3408 554964 3460
rect 555016 3448 555022 3460
rect 572916 3448 572944 3488
rect 574094 3476 574100 3488
rect 574152 3476 574158 3528
rect 577406 3476 577412 3528
rect 577464 3516 577470 3528
rect 582742 3516 582748 3528
rect 577464 3488 582748 3516
rect 577464 3476 577470 3488
rect 582742 3476 582748 3488
rect 582800 3476 582806 3528
rect 555016 3420 572944 3448
rect 555016 3408 555022 3420
rect 573910 3408 573916 3460
rect 573968 3448 573974 3460
rect 583110 3448 583116 3460
rect 573968 3420 583116 3448
rect 573968 3408 573974 3420
rect 583110 3408 583116 3420
rect 583168 3408 583174 3460
rect 228358 3380 228364 3392
rect 219406 3352 228364 3380
rect 212224 3340 212230 3352
rect 228358 3340 228364 3352
rect 228416 3340 228422 3392
rect 267826 3340 267832 3392
rect 267884 3380 267890 3392
rect 273254 3380 273260 3392
rect 267884 3352 273260 3380
rect 267884 3340 267890 3352
rect 273254 3340 273260 3352
rect 273312 3340 273318 3392
rect 299658 3340 299664 3392
rect 299716 3380 299722 3392
rect 302326 3380 302332 3392
rect 299716 3352 302332 3380
rect 299716 3340 299722 3352
rect 302326 3340 302332 3352
rect 302384 3340 302390 3392
rect 373994 3340 374000 3392
rect 374052 3380 374058 3392
rect 375282 3380 375288 3392
rect 374052 3352 375288 3380
rect 374052 3340 374058 3352
rect 375282 3340 375288 3352
rect 375340 3340 375346 3392
rect 378778 3340 378784 3392
rect 378836 3380 378842 3392
rect 379974 3380 379980 3392
rect 378836 3352 379980 3380
rect 378836 3340 378842 3352
rect 379974 3340 379980 3352
rect 380032 3340 380038 3392
rect 396718 3340 396724 3392
rect 396776 3380 396782 3392
rect 398926 3380 398932 3392
rect 396776 3352 398932 3380
rect 396776 3340 396782 3352
rect 398926 3340 398932 3352
rect 398984 3340 398990 3392
rect 406378 3340 406384 3392
rect 406436 3380 406442 3392
rect 407206 3380 407212 3392
rect 406436 3352 407212 3380
rect 406436 3340 406442 3352
rect 407206 3340 407212 3352
rect 407264 3340 407270 3392
rect 420178 3340 420184 3392
rect 420236 3380 420242 3392
rect 421006 3380 421012 3392
rect 420236 3352 421012 3380
rect 420236 3340 420242 3352
rect 421006 3340 421012 3352
rect 421064 3340 421070 3392
rect 427262 3340 427268 3392
rect 427320 3380 427326 3392
rect 427906 3380 427912 3392
rect 427320 3352 427912 3380
rect 427320 3340 427326 3352
rect 427906 3340 427912 3352
rect 427964 3340 427970 3392
rect 440234 3340 440240 3392
rect 440292 3380 440298 3392
rect 441522 3380 441528 3392
rect 440292 3352 441528 3380
rect 440292 3340 440298 3352
rect 441522 3340 441528 3352
rect 441580 3340 441586 3392
rect 493318 3340 493324 3392
rect 493376 3380 493382 3392
rect 494698 3380 494704 3392
rect 493376 3352 494704 3380
rect 493376 3340 493382 3352
rect 494698 3340 494704 3352
rect 494756 3340 494762 3392
rect 504358 3340 504364 3392
rect 504416 3380 504422 3392
rect 505370 3380 505376 3392
rect 504416 3352 505376 3380
rect 504416 3340 504422 3352
rect 505370 3340 505376 3352
rect 505428 3340 505434 3392
rect 20622 3272 20628 3324
rect 20680 3272 20686 3324
rect 34790 3272 34796 3324
rect 34848 3312 34854 3324
rect 35802 3312 35808 3324
rect 34848 3284 35808 3312
rect 34848 3272 34854 3284
rect 35802 3272 35808 3284
rect 35860 3272 35866 3324
rect 64322 3272 64328 3324
rect 64380 3312 64386 3324
rect 64782 3312 64788 3324
rect 64380 3284 64788 3312
rect 64380 3272 64386 3284
rect 64782 3272 64788 3284
rect 64840 3272 64846 3324
rect 106918 3272 106924 3324
rect 106976 3312 106982 3324
rect 107562 3312 107568 3324
rect 106976 3284 107568 3312
rect 106976 3272 106982 3284
rect 107562 3272 107568 3284
rect 107620 3272 107626 3324
rect 135254 3272 135260 3324
rect 135312 3312 135318 3324
rect 136542 3312 136548 3324
rect 135312 3284 136548 3312
rect 135312 3272 135318 3284
rect 136542 3272 136548 3284
rect 136600 3272 136606 3324
rect 151814 3272 151820 3324
rect 151872 3312 151878 3324
rect 156598 3312 156604 3324
rect 151872 3284 156604 3312
rect 151872 3272 151878 3284
rect 156598 3272 156604 3284
rect 156656 3272 156662 3324
rect 156690 3272 156696 3324
rect 156748 3312 156754 3324
rect 162210 3312 162216 3324
rect 156748 3284 162216 3312
rect 156748 3272 156754 3284
rect 162210 3272 162216 3284
rect 162268 3272 162274 3324
rect 335998 3272 336004 3324
rect 336056 3312 336062 3324
rect 342162 3312 342168 3324
rect 336056 3284 342168 3312
rect 336056 3272 336062 3284
rect 342162 3272 342168 3284
rect 342220 3272 342226 3324
rect 367830 3272 367836 3324
rect 367888 3312 367894 3324
rect 369394 3312 369400 3324
rect 367888 3284 369400 3312
rect 367888 3272 367894 3284
rect 369394 3272 369400 3284
rect 369452 3272 369458 3324
rect 93946 3204 93952 3256
rect 94004 3244 94010 3256
rect 98730 3244 98736 3256
rect 94004 3216 98736 3244
rect 94004 3204 94010 3216
rect 98730 3204 98736 3216
rect 98788 3204 98794 3256
rect 209774 3204 209780 3256
rect 209832 3244 209838 3256
rect 213178 3244 213184 3256
rect 209832 3216 213184 3244
rect 209832 3204 209838 3216
rect 213178 3204 213184 3216
rect 213236 3204 213242 3256
rect 215662 3204 215668 3256
rect 215720 3244 215726 3256
rect 216582 3244 216588 3256
rect 215720 3216 216588 3244
rect 215720 3204 215726 3216
rect 216582 3204 216588 3216
rect 216640 3204 216646 3256
rect 259822 3204 259828 3256
rect 259880 3244 259886 3256
rect 261754 3244 261760 3256
rect 259880 3216 261760 3244
rect 259880 3204 259886 3216
rect 261754 3204 261760 3216
rect 261812 3204 261818 3256
rect 296162 3204 296168 3256
rect 296220 3244 296226 3256
rect 297266 3244 297272 3256
rect 296220 3216 297272 3244
rect 296220 3204 296226 3216
rect 297266 3204 297272 3216
rect 297324 3204 297330 3256
rect 39574 3136 39580 3188
rect 39632 3176 39638 3188
rect 40678 3176 40684 3188
rect 39632 3148 40684 3176
rect 39632 3136 39638 3148
rect 40678 3136 40684 3148
rect 40736 3136 40742 3188
rect 73798 3136 73804 3188
rect 73856 3176 73862 3188
rect 75178 3176 75184 3188
rect 73856 3148 75184 3176
rect 73856 3136 73862 3148
rect 75178 3136 75184 3148
rect 75236 3136 75242 3188
rect 147122 3136 147128 3188
rect 147180 3176 147186 3188
rect 147582 3176 147588 3188
rect 147180 3148 147588 3176
rect 147180 3136 147186 3148
rect 147582 3136 147588 3148
rect 147640 3136 147646 3188
rect 160094 3136 160100 3188
rect 160152 3176 160158 3188
rect 161382 3176 161388 3188
rect 160152 3148 161388 3176
rect 160152 3136 160158 3148
rect 161382 3136 161388 3148
rect 161440 3136 161446 3188
rect 230382 3136 230388 3188
rect 230440 3176 230446 3188
rect 235810 3176 235816 3188
rect 230440 3148 235816 3176
rect 230440 3136 230446 3148
rect 235810 3136 235816 3148
rect 235868 3136 235874 3188
rect 251174 3136 251180 3188
rect 251232 3176 251238 3188
rect 258166 3176 258172 3188
rect 251232 3148 258172 3176
rect 251232 3136 251238 3148
rect 258166 3136 258172 3148
rect 258224 3136 258230 3188
rect 311250 3136 311256 3188
rect 311308 3176 311314 3188
rect 315022 3176 315028 3188
rect 311308 3148 315028 3176
rect 311308 3136 311314 3148
rect 315022 3136 315028 3148
rect 315080 3136 315086 3188
rect 320910 3068 320916 3120
rect 320968 3108 320974 3120
rect 324314 3108 324320 3120
rect 320968 3080 324320 3108
rect 320968 3068 320974 3080
rect 324314 3068 324320 3080
rect 324372 3068 324378 3120
rect 347038 3068 347044 3120
rect 347096 3108 347102 3120
rect 350442 3108 350448 3120
rect 347096 3080 350448 3108
rect 347096 3068 347102 3080
rect 350442 3068 350448 3080
rect 350500 3068 350506 3120
rect 457438 3068 457444 3120
rect 457496 3108 457502 3120
rect 462774 3108 462780 3120
rect 457496 3080 462780 3108
rect 457496 3068 457502 3080
rect 462774 3068 462780 3080
rect 462832 3068 462838 3120
rect 547874 3068 547880 3120
rect 547932 3108 547938 3120
rect 550634 3108 550640 3120
rect 547932 3080 550640 3108
rect 547932 3068 547938 3080
rect 550634 3068 550640 3080
rect 550692 3068 550698 3120
rect 27706 3000 27712 3052
rect 27764 3040 27770 3052
rect 35250 3040 35256 3052
rect 27764 3012 35256 3040
rect 27764 3000 27770 3012
rect 35250 3000 35256 3012
rect 35308 3000 35314 3052
rect 69106 3000 69112 3052
rect 69164 3040 69170 3052
rect 71038 3040 71044 3052
rect 69164 3012 71044 3040
rect 69164 3000 69170 3012
rect 71038 3000 71044 3012
rect 71096 3000 71102 3052
rect 85666 3000 85672 3052
rect 85724 3040 85730 3052
rect 86862 3040 86868 3052
rect 85724 3012 86868 3040
rect 85724 3000 85730 3012
rect 86862 3000 86868 3012
rect 86920 3000 86926 3052
rect 176654 3000 176660 3052
rect 176712 3040 176718 3052
rect 178770 3040 178776 3052
rect 176712 3012 178776 3040
rect 176712 3000 176718 3012
rect 178770 3000 178776 3012
rect 178828 3000 178834 3052
rect 191558 3000 191564 3052
rect 191616 3040 191622 3052
rect 192018 3040 192024 3052
rect 191616 3012 192024 3040
rect 191616 3000 191622 3012
rect 192018 3000 192024 3012
rect 192076 3000 192082 3052
rect 389818 3000 389824 3052
rect 389876 3040 389882 3052
rect 391842 3040 391848 3052
rect 389876 3012 391848 3040
rect 389876 3000 389882 3012
rect 391842 3000 391848 3012
rect 391900 3000 391906 3052
rect 437934 3000 437940 3052
rect 437992 3040 437998 3052
rect 438946 3040 438952 3052
rect 437992 3012 438952 3040
rect 437992 3000 437998 3012
rect 438946 3000 438952 3012
rect 439004 3000 439010 3052
rect 447778 3000 447784 3052
rect 447836 3040 447842 3052
rect 448606 3040 448612 3052
rect 447836 3012 448612 3040
rect 447836 3000 447842 3012
rect 448606 3000 448612 3012
rect 448664 3000 448670 3052
rect 479518 3000 479524 3052
rect 479576 3040 479582 3052
rect 480530 3040 480536 3052
rect 479576 3012 480536 3040
rect 479576 3000 479582 3012
rect 480530 3000 480536 3012
rect 480588 3000 480594 3052
rect 578602 3000 578608 3052
rect 578660 3040 578666 3052
rect 582374 3040 582380 3052
rect 578660 3012 582380 3040
rect 578660 3000 578666 3012
rect 582374 3000 582380 3012
rect 582432 3000 582438 3052
rect 175458 2932 175464 2984
rect 175516 2972 175522 2984
rect 177298 2972 177304 2984
rect 175516 2944 177304 2972
rect 175516 2932 175522 2944
rect 177298 2932 177304 2944
rect 177356 2932 177362 2984
rect 283098 2932 283104 2984
rect 283156 2972 283162 2984
rect 285674 2972 285680 2984
rect 283156 2944 285680 2972
rect 283156 2932 283162 2944
rect 285674 2932 285680 2944
rect 285732 2932 285738 2984
rect 316678 2932 316684 2984
rect 316736 2972 316742 2984
rect 322106 2972 322112 2984
rect 316736 2944 322112 2972
rect 316736 2932 316742 2944
rect 322106 2932 322112 2944
rect 322164 2932 322170 2984
rect 82078 2864 82084 2916
rect 82136 2904 82142 2916
rect 83458 2904 83464 2916
rect 82136 2876 83464 2904
rect 82136 2864 82142 2876
rect 83458 2864 83464 2876
rect 83516 2864 83522 2916
rect 142430 2864 142436 2916
rect 142488 2904 142494 2916
rect 143442 2904 143448 2916
rect 142488 2876 143448 2904
rect 142488 2864 142494 2876
rect 143442 2864 143448 2876
rect 143500 2864 143506 2916
rect 186130 2864 186136 2916
rect 186188 2904 186194 2916
rect 186958 2904 186964 2916
rect 186188 2876 186964 2904
rect 186188 2864 186194 2876
rect 186958 2864 186964 2876
rect 187016 2864 187022 2916
rect 289078 2864 289084 2916
rect 289136 2904 289142 2916
rect 293678 2904 293684 2916
rect 289136 2876 293684 2904
rect 289136 2864 289142 2876
rect 293678 2864 293684 2876
rect 293736 2864 293742 2916
rect 307018 2864 307024 2916
rect 307076 2904 307082 2916
rect 307938 2904 307944 2916
rect 307076 2876 307944 2904
rect 307076 2864 307082 2876
rect 307938 2864 307944 2876
rect 307996 2864 308002 2916
rect 429838 2864 429844 2916
rect 429896 2904 429902 2916
rect 434438 2904 434444 2916
rect 429896 2876 434444 2904
rect 429896 2864 429902 2876
rect 434438 2864 434444 2876
rect 434496 2864 434502 2916
rect 150618 2252 150624 2304
rect 150676 2292 150682 2304
rect 207658 2292 207664 2304
rect 150676 2264 207664 2292
rect 150676 2252 150682 2264
rect 207658 2252 207664 2264
rect 207716 2252 207722 2304
rect 140038 2184 140044 2236
rect 140096 2224 140102 2236
rect 202138 2224 202144 2236
rect 140096 2196 202144 2224
rect 140096 2184 140102 2196
rect 202138 2184 202144 2196
rect 202196 2184 202202 2236
rect 63218 2116 63224 2168
rect 63276 2156 63282 2168
rect 210142 2156 210148 2168
rect 63276 2128 210148 2156
rect 63276 2116 63282 2128
rect 210142 2116 210148 2128
rect 210200 2116 210206 2168
rect 7650 2048 7656 2100
rect 7708 2088 7714 2100
rect 200390 2088 200396 2100
rect 7708 2060 200396 2088
rect 7708 2048 7714 2060
rect 200390 2048 200396 2060
rect 200448 2048 200454 2100
rect 206186 2048 206192 2100
rect 206244 2088 206250 2100
rect 235074 2088 235080 2100
rect 206244 2060 235080 2088
rect 206244 2048 206250 2060
rect 235074 2048 235080 2060
rect 235132 2048 235138 2100
<< via1 >>
rect 331220 702992 331272 703044
rect 332508 702992 332560 703044
rect 294604 700544 294656 700596
rect 364984 700544 365036 700596
rect 298744 700476 298796 700528
rect 397460 700476 397512 700528
rect 40500 700408 40552 700460
rect 41328 700408 41380 700460
rect 305644 700408 305696 700460
rect 494796 700408 494848 700460
rect 137836 700340 137888 700392
rect 195244 700340 195296 700392
rect 244924 700340 244976 700392
rect 462320 700340 462372 700392
rect 24308 700272 24360 700324
rect 137284 700272 137336 700324
rect 218980 700272 219032 700324
rect 240784 700272 240836 700324
rect 242164 700272 242216 700324
rect 527180 700272 527232 700324
rect 559656 700272 559708 700324
rect 582932 700272 582984 700324
rect 154120 699728 154172 699780
rect 157984 699728 158036 699780
rect 105452 699660 105504 699712
rect 106188 699660 106240 699712
rect 170312 699660 170364 699712
rect 171048 699660 171100 699712
rect 235172 699660 235224 699712
rect 235908 699660 235960 699712
rect 282184 699660 282236 699712
rect 283840 699660 283892 699712
rect 347044 699660 347096 699712
rect 348792 699660 348844 699712
rect 476764 699660 476816 699712
rect 478512 699660 478564 699712
rect 266360 697552 266412 697604
rect 267648 697552 267700 697604
rect 3424 683136 3476 683188
rect 199384 683136 199436 683188
rect 3516 670692 3568 670744
rect 260104 670692 260156 670744
rect 3424 656888 3476 656940
rect 262864 656888 262916 656940
rect 251088 649272 251140 649324
rect 266360 649272 266412 649324
rect 3424 632068 3476 632120
rect 258724 632068 258776 632120
rect 3148 618264 3200 618316
rect 231124 618264 231176 618316
rect 235908 606432 235960 606484
rect 252560 606432 252612 606484
rect 3240 605820 3292 605872
rect 192484 605820 192536 605872
rect 3332 579640 3384 579692
rect 255964 579640 256016 579692
rect 3424 565836 3476 565888
rect 39304 565836 39356 565888
rect 3424 553392 3476 553444
rect 173164 553392 173216 553444
rect 3424 527144 3476 527196
rect 210424 527144 210476 527196
rect 3424 514768 3476 514820
rect 206284 514768 206336 514820
rect 3056 474716 3108 474768
rect 198004 474716 198056 474768
rect 3516 462340 3568 462392
rect 191104 462340 191156 462392
rect 238668 458804 238720 458856
rect 583392 458804 583444 458856
rect 291844 456764 291896 456816
rect 580172 456764 580224 456816
rect 3148 448536 3200 448588
rect 166264 448536 166316 448588
rect 224868 430584 224920 430636
rect 580172 430584 580224 430636
rect 3516 422288 3568 422340
rect 196624 422288 196676 422340
rect 289084 418140 289136 418192
rect 580172 418140 580224 418192
rect 2872 409844 2924 409896
rect 249064 409844 249116 409896
rect 234528 403588 234580 403640
rect 583484 403588 583536 403640
rect 3516 397468 3568 397520
rect 177304 397468 177356 397520
rect 3516 371220 3568 371272
rect 213184 371220 213236 371272
rect 246304 364352 246356 364404
rect 580172 364352 580224 364404
rect 3148 357416 3200 357468
rect 280344 357416 280396 357468
rect 231124 355308 231176 355360
rect 267280 355308 267332 355360
rect 231768 353948 231820 354000
rect 583668 353948 583720 354000
rect 295984 351908 296036 351960
rect 579896 351908 579948 351960
rect 3332 345040 3384 345092
rect 226984 345040 227036 345092
rect 39304 344292 39356 344344
rect 269948 344292 270000 344344
rect 580908 343204 580960 343256
rect 583484 343204 583536 343256
rect 235264 324300 235316 324352
rect 580172 324300 580224 324352
rect 3332 318792 3384 318844
rect 209044 318792 209096 318844
rect 249064 318044 249116 318096
rect 277768 318044 277820 318096
rect 220728 311856 220780 311908
rect 580172 311856 580224 311908
rect 3516 304988 3568 305040
rect 200764 304988 200816 305040
rect 229008 300092 229060 300144
rect 583576 300092 583628 300144
rect 252468 294584 252520 294636
rect 282184 294584 282236 294636
rect 3516 292544 3568 292596
rect 282092 292544 282144 292596
rect 177304 286288 177356 286340
rect 276848 286288 276900 286340
rect 232504 271872 232556 271924
rect 580172 271872 580224 271924
rect 3056 266364 3108 266416
rect 285680 266364 285732 266416
rect 217968 258068 218020 258120
rect 580172 258068 580224 258120
rect 3516 253920 3568 253972
rect 285588 253920 285640 253972
rect 240048 246304 240100 246356
rect 582932 246304 582984 246356
rect 3056 240116 3108 240168
rect 204904 240116 204956 240168
rect 215944 231820 215996 231872
rect 580172 231820 580224 231872
rect 166264 228352 166316 228404
rect 274272 228352 274324 228404
rect 3424 226992 3476 227044
rect 271696 226992 271748 227044
rect 89628 224204 89680 224256
rect 259460 224204 259512 224256
rect 260104 224204 260156 224256
rect 264704 224204 264756 224256
rect 223488 221416 223540 221468
rect 246304 221416 246356 221468
rect 249708 220056 249760 220108
rect 347044 220056 347096 220108
rect 215208 218016 215260 218068
rect 580172 218016 580224 218068
rect 246948 217268 247000 217320
rect 412640 217268 412692 217320
rect 173164 215908 173216 215960
rect 269028 215908 269080 215960
rect 241428 214548 241480 214600
rect 542360 214548 542412 214600
rect 3148 213936 3200 213988
rect 287060 213936 287112 213988
rect 240784 211828 240836 211880
rect 254308 211828 254360 211880
rect 222108 211760 222160 211812
rect 295984 211760 296036 211812
rect 580908 211080 580960 211132
rect 582380 211080 582432 211132
rect 226248 210808 226300 210860
rect 289084 210808 289136 210860
rect 206284 210740 206336 210792
rect 272524 210740 272576 210792
rect 200764 210672 200816 210724
rect 282920 210672 282972 210724
rect 191104 210604 191156 210656
rect 275100 210604 275152 210656
rect 137284 210536 137336 210588
rect 262128 210536 262180 210588
rect 244188 210468 244240 210520
rect 476764 210468 476816 210520
rect 220636 210400 220688 210452
rect 235264 210400 235316 210452
rect 235908 210400 235960 210452
rect 582564 210400 582616 210452
rect 226984 209448 227036 209500
rect 279516 209448 279568 209500
rect 199384 209380 199436 209432
rect 262956 209380 263008 209432
rect 192484 209312 192536 209364
rect 266452 209312 266504 209364
rect 204904 209244 204956 209296
rect 284668 209244 284720 209296
rect 8208 209176 8260 209228
rect 260748 209176 260800 209228
rect 232964 209108 233016 209160
rect 582840 209108 582892 209160
rect 227628 209040 227680 209092
rect 583300 209040 583352 209092
rect 262864 208836 262916 208888
rect 263876 208836 263928 208888
rect 213184 208020 213236 208072
rect 278596 208020 278648 208072
rect 196624 207952 196676 208004
rect 276020 207952 276072 208004
rect 157984 207884 158036 207936
rect 256884 207884 256936 207936
rect 246028 207816 246080 207868
rect 429200 207816 429252 207868
rect 41328 207748 41380 207800
rect 259184 207748 259236 207800
rect 223856 207680 223908 207732
rect 583392 207680 583444 207732
rect 216404 207612 216456 207664
rect 582932 207612 582984 207664
rect 214288 207000 214340 207052
rect 215944 207000 215996 207052
rect 240324 207000 240376 207052
rect 242164 207000 242216 207052
rect 251180 206592 251232 206644
rect 299480 206592 299532 206644
rect 226432 206524 226484 206576
rect 291844 206524 291896 206576
rect 209044 206456 209096 206508
rect 281264 206456 281316 206508
rect 198004 206388 198056 206440
rect 273352 206388 273404 206440
rect 171048 206320 171100 206372
rect 252652 206320 252704 206372
rect 216864 206252 216916 206304
rect 232504 206252 232556 206304
rect 234436 206252 234488 206304
rect 582748 206252 582800 206304
rect 213828 205640 213880 205692
rect 580172 205640 580224 205692
rect 202788 205164 202840 205216
rect 250628 205164 250680 205216
rect 245568 205096 245620 205148
rect 298744 205096 298796 205148
rect 195244 205028 195296 205080
rect 255504 205028 255556 205080
rect 248512 204960 248564 205012
rect 331220 204960 331272 205012
rect 228916 204892 228968 204944
rect 583208 204892 583260 204944
rect 258724 204824 258776 204876
rect 265532 204824 265584 204876
rect 209044 204348 209096 204400
rect 583392 204348 583444 204400
rect 202052 204280 202104 204332
rect 582472 204280 582524 204332
rect 247316 203600 247368 203652
rect 294604 203600 294656 203652
rect 210424 203532 210476 203584
rect 270776 203532 270828 203584
rect 159364 203124 159416 203176
rect 289084 203192 289136 203244
rect 283840 203124 283892 203176
rect 285680 203124 285732 203176
rect 207296 203056 207348 203108
rect 583024 203056 583076 203108
rect 205548 202988 205600 203040
rect 582656 202988 582708 203040
rect 202972 202920 203024 202972
rect 583576 202920 583628 202972
rect 201224 202852 201276 202904
rect 583852 202852 583904 202904
rect 228180 202784 228232 202836
rect 229008 202784 229060 202836
rect 235172 202444 235224 202496
rect 235908 202444 235960 202496
rect 233424 202308 233476 202360
rect 234528 202308 234580 202360
rect 230756 202240 230808 202292
rect 231768 202240 231820 202292
rect 218612 202104 218664 202156
rect 582380 202104 582432 202156
rect 251640 201968 251692 202020
rect 252468 201968 252520 202020
rect 208216 201900 208268 201952
rect 583208 201900 583260 201952
rect 140044 201832 140096 201884
rect 295984 201832 296036 201884
rect 98644 201764 98696 201816
rect 298652 201764 298704 201816
rect 14464 201696 14516 201748
rect 292488 201696 292540 201748
rect 3240 201628 3292 201680
rect 288164 201628 288216 201680
rect 209872 201560 209924 201612
rect 583300 201560 583352 201612
rect 212540 201492 212592 201544
rect 219348 201492 219400 201544
rect 219440 201492 219492 201544
rect 220636 201492 220688 201544
rect 221188 201424 221240 201476
rect 222108 201424 222160 201476
rect 249892 201356 249944 201408
rect 251180 201356 251232 201408
rect 3424 200812 3476 200864
rect 290832 200812 290884 200864
rect 219348 200744 219400 200796
rect 580264 200744 580316 200796
rect 211620 200404 211672 200456
rect 304264 200404 304316 200456
rect 157248 200336 157300 200388
rect 299480 200336 299532 200388
rect 133144 200268 133196 200320
rect 297732 200268 297784 200320
rect 36544 200200 36596 200252
rect 293408 200200 293460 200252
rect 204720 200132 204772 200184
rect 583668 200132 583720 200184
rect 287612 199860 287664 199912
rect 294788 199860 294840 199912
rect 206744 199792 206796 199844
rect 210424 199792 210476 199844
rect 199936 199724 199988 199776
rect 213184 199724 213236 199776
rect 244188 199724 244240 199776
rect 249248 199724 249300 199776
rect 200028 199656 200080 199708
rect 203524 199656 203576 199708
rect 203708 199656 203760 199708
rect 213276 199656 213328 199708
rect 215024 199588 215076 199640
rect 199384 199520 199436 199572
rect 157984 199044 158036 199096
rect 203708 199452 203760 199504
rect 204076 199452 204128 199504
rect 207664 199452 207716 199504
rect 210332 199452 210384 199504
rect 210424 199452 210476 199504
rect 210516 199452 210568 199504
rect 148324 198976 148376 199028
rect 106924 198908 106976 198960
rect 199936 198908 199988 198960
rect 47584 198772 47636 198824
rect 199844 198772 199896 198824
rect 183008 198704 183060 198756
rect 198004 198704 198056 198756
rect 35164 198092 35216 198144
rect 211160 199452 211212 199504
rect 211252 199452 211304 199504
rect 213184 199452 213236 199504
rect 213276 199452 213328 199504
rect 215024 199452 215076 199504
rect 238024 199452 238076 199504
rect 246304 199656 246356 199708
rect 244188 199452 244240 199504
rect 246212 199452 246264 199504
rect 246304 199452 246356 199504
rect 246488 199452 246540 199504
rect 249248 199452 249300 199504
rect 287060 199520 287112 199572
rect 289636 199724 289688 199776
rect 287704 199656 287756 199708
rect 293224 199724 293276 199776
rect 291292 199588 291344 199640
rect 296628 199656 296680 199708
rect 287612 199452 287664 199504
rect 287704 199452 287756 199504
rect 293224 199452 293276 199504
rect 294144 199452 294196 199504
rect 583760 198840 583812 198892
rect 582380 198704 582432 198756
rect 583116 198024 583168 198076
rect 199936 197752 199988 197804
rect 583760 197956 583812 198008
rect 174544 197344 174596 197396
rect 198004 197344 198056 197396
rect 181536 195984 181588 196036
rect 198004 195984 198056 196036
rect 151728 194556 151780 194608
rect 198096 194556 198148 194608
rect 170496 193196 170548 193248
rect 197728 193196 197780 193248
rect 304264 193128 304316 193180
rect 580172 193128 580224 193180
rect 153108 191836 153160 191888
rect 197636 191836 197688 191888
rect 191196 191020 191248 191072
rect 198096 191020 198148 191072
rect 155868 190476 155920 190528
rect 197360 190476 197412 190528
rect 172428 189116 172480 189168
rect 188436 189116 188488 189168
rect 180156 189048 180208 189100
rect 197912 189048 197964 189100
rect 3516 188980 3568 189032
rect 199384 188980 199436 189032
rect 173164 187688 173216 187740
rect 197360 187688 197412 187740
rect 172428 186396 172480 186448
rect 184388 186396 184440 186448
rect 178776 186328 178828 186380
rect 197544 186328 197596 186380
rect 195336 186192 195388 186244
rect 197636 186192 197688 186244
rect 171784 185580 171836 185632
rect 186964 185580 187016 185632
rect 178868 184152 178920 184204
rect 197360 184152 197412 184204
rect 196716 183744 196768 183796
rect 198372 183744 198424 183796
rect 172428 183608 172480 183660
rect 177304 183608 177356 183660
rect 171692 183540 171744 183592
rect 176016 183540 176068 183592
rect 172428 182248 172480 182300
rect 185584 182248 185636 182300
rect 174636 182180 174688 182232
rect 197728 182180 197780 182232
rect 192484 181432 192536 181484
rect 197360 181432 197412 181484
rect 172428 180820 172480 180872
rect 193864 180820 193916 180872
rect 172060 179460 172112 179512
rect 182916 179460 182968 179512
rect 177396 179392 177448 179444
rect 197360 179392 197412 179444
rect 172152 178100 172204 178152
rect 184296 178100 184348 178152
rect 175924 178032 175976 178084
rect 197912 178032 197964 178084
rect 188528 177352 188580 177404
rect 198096 177352 198148 177404
rect 184388 177284 184440 177336
rect 198188 177284 198240 177336
rect 172428 176740 172480 176792
rect 180064 176740 180116 176792
rect 172244 176672 172296 176724
rect 184204 176672 184256 176724
rect 191288 176332 191340 176384
rect 197820 176332 197872 176384
rect 172428 175244 172480 175296
rect 195428 175244 195480 175296
rect 189724 174496 189776 174548
rect 197360 174496 197412 174548
rect 173440 173884 173492 173936
rect 198556 173884 198608 173936
rect 171784 173204 171836 173256
rect 187056 173204 187108 173256
rect 176016 173136 176068 173188
rect 198096 173136 198148 173188
rect 196808 173000 196860 173052
rect 198464 173000 198516 173052
rect 176016 171776 176068 171828
rect 197360 171776 197412 171828
rect 172244 171096 172296 171148
rect 181444 171096 181496 171148
rect 172244 169736 172296 169788
rect 191104 169736 191156 169788
rect 192576 169736 192628 169788
rect 197728 169736 197780 169788
rect 193956 168512 194008 168564
rect 197728 168512 197780 168564
rect 172428 168376 172480 168428
rect 196624 168376 196676 168428
rect 172428 167084 172480 167136
rect 195244 167084 195296 167136
rect 174728 167016 174780 167068
rect 197912 167016 197964 167068
rect 172060 166268 172112 166320
rect 192484 166268 192536 166320
rect 172428 165656 172480 165708
rect 188344 165656 188396 165708
rect 181628 165588 181680 165640
rect 197360 165588 197412 165640
rect 171140 164296 171192 164348
rect 192484 164296 192536 164348
rect 169208 164228 169260 164280
rect 174544 164228 174596 164280
rect 177488 164228 177540 164280
rect 197636 164228 197688 164280
rect 3240 164160 3292 164212
rect 159364 164160 159416 164212
rect 180248 163480 180300 163532
rect 197360 163480 197412 163532
rect 171876 162936 171928 162988
rect 174544 162936 174596 162988
rect 171692 162868 171744 162920
rect 178684 162868 178736 162920
rect 178960 162188 179012 162240
rect 197636 162188 197688 162240
rect 169392 162120 169444 162172
rect 197452 162120 197504 162172
rect 160008 161440 160060 161492
rect 169300 161440 169352 161492
rect 171692 160828 171744 160880
rect 183008 160828 183060 160880
rect 169300 160760 169352 160812
rect 181536 160760 181588 160812
rect 160836 160692 160888 160744
rect 191196 160692 191248 160744
rect 165160 160488 165212 160540
rect 169300 160488 169352 160540
rect 166816 160420 166868 160472
rect 171692 160420 171744 160472
rect 163136 160352 163188 160404
rect 170496 160352 170548 160404
rect 171876 160080 171928 160132
rect 182824 160080 182876 160132
rect 191380 160080 191432 160132
rect 197360 160080 197412 160132
rect 173348 159332 173400 159384
rect 198464 159332 198516 159384
rect 176108 158720 176160 158772
rect 197544 158720 197596 158772
rect 171968 158652 172020 158704
rect 173256 158652 173308 158704
rect 188436 157972 188488 158024
rect 198464 157972 198516 158024
rect 187148 157360 187200 157412
rect 197360 157360 197412 157412
rect 195428 156884 195480 156936
rect 198004 156884 198056 156936
rect 172244 156000 172296 156052
rect 180156 156000 180208 156052
rect 195520 156000 195572 156052
rect 197912 156000 197964 156052
rect 171968 155320 172020 155372
rect 173440 155320 173492 155372
rect 170496 154572 170548 154624
rect 197728 154572 197780 154624
rect 171692 154504 171744 154556
rect 173164 154504 173216 154556
rect 186964 154504 187016 154556
rect 197360 154504 197412 154556
rect 192668 153212 192720 153264
rect 197360 153212 197412 153264
rect 172336 153144 172388 153196
rect 195336 153144 195388 153196
rect 171508 153076 171560 153128
rect 178776 153076 178828 153128
rect 172336 151648 172388 151700
rect 178868 151648 178920 151700
rect 172428 151580 172480 151632
rect 196716 151580 196768 151632
rect 171324 151172 171376 151224
rect 174636 151172 174688 151224
rect 186964 150424 187016 150476
rect 197452 150424 197504 150476
rect 187056 150356 187108 150408
rect 197360 150356 197412 150408
rect 172244 149676 172296 149728
rect 192576 149676 192628 149728
rect 171508 149608 171560 149660
rect 177396 149608 177448 149660
rect 171692 148996 171744 149048
rect 191288 148996 191340 149048
rect 172428 148928 172480 148980
rect 188528 148928 188580 148980
rect 171324 148316 171376 148368
rect 175924 148316 175976 148368
rect 193864 147704 193916 147756
rect 177396 147636 177448 147688
rect 197544 147636 197596 147688
rect 198096 147636 198148 147688
rect 172428 147568 172480 147620
rect 189724 147568 189776 147620
rect 177304 146888 177356 146940
rect 197360 146888 197412 146940
rect 178776 146276 178828 146328
rect 198188 146276 198240 146328
rect 172336 146208 172388 146260
rect 198740 146208 198792 146260
rect 172428 146140 172480 146192
rect 196808 146140 196860 146192
rect 172152 146072 172204 146124
rect 176016 146072 176068 146124
rect 171324 144848 171376 144900
rect 193956 144848 194008 144900
rect 171968 144168 172020 144220
rect 187148 144168 187200 144220
rect 186320 143556 186372 143608
rect 197452 143556 197504 143608
rect 172428 143488 172480 143540
rect 181628 143488 181680 143540
rect 185584 143488 185636 143540
rect 197360 143488 197412 143540
rect 171692 143352 171744 143404
rect 174728 143352 174780 143404
rect 171876 142808 171928 142860
rect 186320 142808 186372 142860
rect 187056 142128 187108 142180
rect 197360 142128 197412 142180
rect 171508 142060 171560 142112
rect 177488 142060 177540 142112
rect 172428 141516 172480 141568
rect 180248 141516 180300 141568
rect 184296 141380 184348 141432
rect 198464 141380 198516 141432
rect 171508 140972 171560 141024
rect 178960 140972 179012 141024
rect 172428 140700 172480 140752
rect 191380 140700 191432 140752
rect 171692 140632 171744 140684
rect 173348 140632 173400 140684
rect 176016 139408 176068 139460
rect 197360 139408 197412 139460
rect 171324 139340 171376 139392
rect 195520 139340 195572 139392
rect 182916 139272 182968 139324
rect 198188 139272 198240 139324
rect 172428 139204 172480 139256
rect 176108 139204 176160 139256
rect 3240 137912 3292 137964
rect 157984 137912 158036 137964
rect 171508 137912 171560 137964
rect 192668 137912 192720 137964
rect 176660 136620 176712 136672
rect 197544 136620 197596 136672
rect 172428 136552 172480 136604
rect 186964 136552 187016 136604
rect 171692 136484 171744 136536
rect 177396 136484 177448 136536
rect 171508 135600 171560 135652
rect 178776 135600 178828 135652
rect 175280 135260 175332 135312
rect 198188 135260 198240 135312
rect 171508 135192 171560 135244
rect 187056 135192 187108 135244
rect 184204 135124 184256 135176
rect 197360 135124 197412 135176
rect 171876 134716 171928 134768
rect 176016 134716 176068 134768
rect 171692 133832 171744 133884
rect 175280 133832 175332 133884
rect 172428 133356 172480 133408
rect 176660 133356 176712 133408
rect 171692 132404 171744 132456
rect 197452 132472 197504 132524
rect 180064 132404 180116 132456
rect 197360 132404 197412 132456
rect 172428 131724 172480 131776
rect 197912 131724 197964 131776
rect 172428 131112 172480 131164
rect 176660 131112 176712 131164
rect 170404 130364 170456 130416
rect 197452 130364 197504 130416
rect 171692 129820 171744 129872
rect 175924 129820 175976 129872
rect 172060 129752 172112 129804
rect 186320 129752 186372 129804
rect 176660 129684 176712 129736
rect 197360 129684 197412 129736
rect 172428 128392 172480 128444
rect 177304 128392 177356 128444
rect 171600 128324 171652 128376
rect 180156 128324 180208 128376
rect 173256 128256 173308 128308
rect 198096 128256 198148 128308
rect 178684 127576 178736 127628
rect 198004 127576 198056 127628
rect 172060 127032 172112 127084
rect 173164 127032 173216 127084
rect 171692 126964 171744 127016
rect 178040 126964 178092 127016
rect 175924 126896 175976 126948
rect 197360 126896 197412 126948
rect 181444 126216 181496 126268
rect 197912 126216 197964 126268
rect 172428 125672 172480 125724
rect 181536 125672 181588 125724
rect 172152 125604 172204 125656
rect 184204 125604 184256 125656
rect 186320 125536 186372 125588
rect 197636 125536 197688 125588
rect 172336 124856 172388 124908
rect 186964 124856 187016 124908
rect 171876 124312 171928 124364
rect 180064 124312 180116 124364
rect 171692 124244 171744 124296
rect 178684 124244 178736 124296
rect 172428 124176 172480 124228
rect 175924 124176 175976 124228
rect 155868 124108 155920 124160
rect 160652 124108 160704 124160
rect 178040 123428 178092 123480
rect 197636 123428 197688 123480
rect 153108 122816 153160 122868
rect 162860 122816 162912 122868
rect 151728 122748 151780 122800
rect 164884 122748 164936 122800
rect 168932 122748 168984 122800
rect 198832 122748 198884 122800
rect 157248 122680 157300 122732
rect 166908 122680 166960 122732
rect 170404 122680 170456 122732
rect 197360 122680 197412 122732
rect 180156 121388 180208 121440
rect 197544 121388 197596 121440
rect 191104 121320 191156 121372
rect 197360 121320 197412 121372
rect 171784 120708 171836 120760
rect 191748 120708 191800 120760
rect 191748 119960 191800 120012
rect 198280 119960 198332 120012
rect 177304 118600 177356 118652
rect 197360 118600 197412 118652
rect 196624 117172 196676 117224
rect 198464 117172 198516 117224
rect 195244 114860 195296 114912
rect 197912 114860 197964 114912
rect 173164 114452 173216 114504
rect 197360 114452 197412 114504
rect 188344 113092 188396 113144
rect 197360 113092 197412 113144
rect 3424 111732 3476 111784
rect 148324 111732 148376 111784
rect 186964 111732 187016 111784
rect 197360 111732 197412 111784
rect 184204 110372 184256 110424
rect 197544 110372 197596 110424
rect 192484 110304 192536 110356
rect 197360 110304 197412 110356
rect 181536 108264 181588 108316
rect 197544 108264 197596 108316
rect 180064 106904 180116 106956
rect 198096 106904 198148 106956
rect 174544 106224 174596 106276
rect 198556 106224 198608 106276
rect 178684 105544 178736 105596
rect 197452 105544 197504 105596
rect 160008 104796 160060 104848
rect 197544 104796 197596 104848
rect 175924 102756 175976 102808
rect 198096 102756 198148 102808
rect 182824 102076 182876 102128
rect 197912 102076 197964 102128
rect 39304 100716 39356 100768
rect 568580 100716 568632 100768
rect 199936 100648 199988 100700
rect 200580 100648 200632 100700
rect 202236 100648 202288 100700
rect 295524 100648 295576 100700
rect 211528 100104 211580 100156
rect 211712 100104 211764 100156
rect 147588 99764 147640 99816
rect 225144 99764 225196 99816
rect 253204 99764 253256 99816
rect 320180 99764 320232 99816
rect 135168 99696 135220 99748
rect 222844 99696 222896 99748
rect 255688 99696 255740 99748
rect 323584 99696 323636 99748
rect 156604 99628 156656 99680
rect 226064 99628 226116 99680
rect 259920 99628 259972 99680
rect 331864 99628 331916 99680
rect 155868 99560 155920 99612
rect 226616 99560 226668 99612
rect 259276 99560 259328 99612
rect 345020 99560 345072 99612
rect 105544 99492 105596 99544
rect 217968 99492 218020 99544
rect 286692 99492 286744 99544
rect 504364 99492 504416 99544
rect 77208 99424 77260 99476
rect 213092 99424 213144 99476
rect 234988 99424 235040 99476
rect 239220 99424 239272 99476
rect 287888 99424 287940 99476
rect 512000 99424 512052 99476
rect 66168 99356 66220 99408
rect 211252 99356 211304 99408
rect 289084 99356 289136 99408
rect 520372 99356 520424 99408
rect 234988 99220 235040 99272
rect 239220 99220 239272 99272
rect 248328 98948 248380 99000
rect 283380 98948 283432 99000
rect 197268 98880 197320 98932
rect 235540 98880 235592 98932
rect 180064 98812 180116 98864
rect 230664 98812 230716 98864
rect 255044 98812 255096 98864
rect 324412 98812 324464 98864
rect 173164 98744 173216 98796
rect 228916 98744 228968 98796
rect 267832 98744 267884 98796
rect 394700 98744 394752 98796
rect 162124 98676 162176 98728
rect 227628 98676 227680 98728
rect 283656 98676 283708 98728
rect 475384 98676 475436 98728
rect 4804 98608 4856 98660
rect 200304 98608 200356 98660
rect 201408 98608 201460 98660
rect 234344 98608 234396 98660
rect 282460 98608 282512 98660
rect 479524 98608 479576 98660
rect 238944 98268 238996 98320
rect 239404 98268 239456 98320
rect 262864 98132 262916 98184
rect 306380 98132 306432 98184
rect 165528 98064 165580 98116
rect 215300 98064 215352 98116
rect 144828 97996 144880 98048
rect 328460 98064 328512 98116
rect 3424 97928 3476 97980
rect 36544 97928 36596 97980
rect 224592 97928 224644 97980
rect 231216 97928 231268 97980
rect 237380 97928 237432 97980
rect 238668 97928 238720 97980
rect 241428 97928 241480 97980
rect 195336 97860 195388 97912
rect 202144 97860 202196 97912
rect 215300 97792 215352 97844
rect 228272 97792 228324 97844
rect 237380 97792 237432 97844
rect 239036 97792 239088 97844
rect 256424 97792 256476 97844
rect 278780 97996 278832 98048
rect 283564 97996 283616 98048
rect 285772 97996 285824 98048
rect 483020 97996 483072 98048
rect 275744 97860 275796 97912
rect 280712 97860 280764 97912
rect 280988 97792 281040 97844
rect 291660 97792 291712 97844
rect 217324 97724 217376 97776
rect 219716 97724 219768 97776
rect 256884 97724 256936 97776
rect 260196 97724 260248 97776
rect 264980 97724 265032 97776
rect 300584 97724 300636 97776
rect 234528 97656 234580 97708
rect 240232 97656 240284 97708
rect 252652 97656 252704 97708
rect 262864 97656 262916 97708
rect 202144 97588 202196 97640
rect 224040 97588 224092 97640
rect 247316 97588 247368 97640
rect 253204 97588 253256 97640
rect 273076 97588 273128 97640
rect 309876 97656 309928 97708
rect 101404 97520 101456 97572
rect 206192 97520 206244 97572
rect 206468 97520 206520 97572
rect 215484 97520 215536 97572
rect 242716 97520 242768 97572
rect 247684 97520 247736 97572
rect 265348 97520 265400 97572
rect 269764 97520 269816 97572
rect 277124 97520 277176 97572
rect 279332 97588 279384 97640
rect 279424 97588 279476 97640
rect 353944 97588 353996 97640
rect 93124 97452 93176 97504
rect 210240 97452 210292 97504
rect 86316 97384 86368 97436
rect 207940 97384 207992 97436
rect 40684 97316 40736 97368
rect 206652 97316 206704 97368
rect 207664 97316 207716 97368
rect 225880 97452 225932 97504
rect 228456 97452 228508 97504
rect 238208 97452 238260 97504
rect 245752 97452 245804 97504
rect 257344 97452 257396 97504
rect 260288 97452 260340 97504
rect 262864 97452 262916 97504
rect 263784 97452 263836 97504
rect 268384 97452 268436 97504
rect 276756 97452 276808 97504
rect 443644 97520 443696 97572
rect 279792 97452 279844 97504
rect 454684 97452 454736 97504
rect 223488 97384 223540 97436
rect 237012 97384 237064 97436
rect 244464 97384 244516 97436
rect 255964 97384 256016 97436
rect 291660 97384 291712 97436
rect 461584 97384 461636 97436
rect 226064 97316 226116 97368
rect 236184 97316 236236 97368
rect 246304 97316 246356 97368
rect 32404 97248 32456 97300
rect 204904 97248 204956 97300
rect 207480 97248 207532 97300
rect 207756 97248 207808 97300
rect 213736 97248 213788 97300
rect 236828 97248 236880 97300
rect 245108 97248 245160 97300
rect 251824 97248 251876 97300
rect 246120 97180 246172 97232
rect 250444 97180 250496 97232
rect 257896 97316 257948 97368
rect 260288 97316 260340 97368
rect 261116 97316 261168 97368
rect 275284 97316 275336 97368
rect 282368 97316 282420 97368
rect 468484 97316 468536 97368
rect 253848 97248 253900 97300
rect 282184 97248 282236 97300
rect 299664 97248 299716 97300
rect 582932 97248 582984 97300
rect 260012 97180 260064 97232
rect 274732 97180 274784 97232
rect 279424 97180 279476 97232
rect 234896 97112 234948 97164
rect 235172 97112 235224 97164
rect 236644 97112 236696 97164
rect 239588 97112 239640 97164
rect 243268 97112 243320 97164
rect 246304 97112 246356 97164
rect 268016 97112 268068 97164
rect 276756 97112 276808 97164
rect 293408 97112 293460 97164
rect 293868 97112 293920 97164
rect 296076 97112 296128 97164
rect 296444 97112 296496 97164
rect 243452 97044 243504 97096
rect 246396 97044 246448 97096
rect 248972 97044 249024 97096
rect 255780 97044 255832 97096
rect 259552 97044 259604 97096
rect 264244 97044 264296 97096
rect 264612 97044 264664 97096
rect 265900 97044 265952 97096
rect 275376 97044 275428 97096
rect 276664 97044 276716 97096
rect 296260 97044 296312 97096
rect 296628 97044 296680 97096
rect 214564 96976 214616 97028
rect 218152 96976 218204 97028
rect 219808 96976 219860 97028
rect 220636 96976 220688 97028
rect 222292 96976 222344 97028
rect 223120 96976 223172 97028
rect 243912 96976 243964 97028
rect 244188 96976 244240 97028
rect 246764 96976 246816 97028
rect 247132 96976 247184 97028
rect 201960 96908 202012 96960
rect 202604 96908 202656 96960
rect 207756 96908 207808 96960
rect 213644 96908 213696 96960
rect 215392 96908 215444 96960
rect 215944 96908 215996 96960
rect 216864 96908 216916 96960
rect 217508 96908 217560 96960
rect 218244 96908 218296 96960
rect 218612 96908 218664 96960
rect 219900 96908 219952 96960
rect 220268 96908 220320 96960
rect 222660 96908 222712 96960
rect 223304 96908 223356 96960
rect 223672 96908 223724 96960
rect 224684 96908 224736 96960
rect 234712 96908 234764 96960
rect 235632 96908 235684 96960
rect 236276 96908 236328 96960
rect 237104 96908 237156 96960
rect 240508 96908 240560 96960
rect 240968 96908 241020 96960
rect 242072 96908 242124 96960
rect 242532 96908 242584 96960
rect 244924 96908 244976 96960
rect 245476 96908 245528 96960
rect 204260 96840 204312 96892
rect 209412 96840 209464 96892
rect 216772 96840 216824 96892
rect 217600 96840 217652 96892
rect 218428 96840 218480 96892
rect 219256 96840 219308 96892
rect 219624 96840 219676 96892
rect 220084 96840 220136 96892
rect 224224 96840 224276 96892
rect 228640 96840 228692 96892
rect 244280 96840 244332 96892
rect 245384 96840 245436 96892
rect 202604 96772 202656 96824
rect 208216 96772 208268 96824
rect 209228 96772 209280 96824
rect 213828 96772 213880 96824
rect 215300 96772 215352 96824
rect 215944 96772 215996 96824
rect 216956 96772 217008 96824
rect 239128 96772 239180 96824
rect 239956 96772 240008 96824
rect 241888 96772 241940 96824
rect 242624 96772 242676 96824
rect 242900 96772 242952 96824
rect 243820 96772 243872 96824
rect 247776 96908 247828 96960
rect 248144 96908 248196 96960
rect 250812 96976 250864 97028
rect 251088 96976 251140 97028
rect 252192 96976 252244 97028
rect 253296 96976 253348 97028
rect 258264 96976 258316 97028
rect 259276 96976 259328 97028
rect 261300 96976 261352 97028
rect 262956 96976 263008 97028
rect 270868 96976 270920 97028
rect 271512 96976 271564 97028
rect 276112 96976 276164 97028
rect 277308 96976 277360 97028
rect 290740 96976 290792 97028
rect 291108 96976 291160 97028
rect 249064 96908 249116 96960
rect 249156 96908 249208 96960
rect 249708 96908 249760 96960
rect 249984 96908 250036 96960
rect 254584 96908 254636 96960
rect 254676 96908 254728 96960
rect 255044 96908 255096 96960
rect 255872 96908 255924 96960
rect 256516 96908 256568 96960
rect 258540 96908 258592 96960
rect 259092 96908 259144 96960
rect 259736 96908 259788 96960
rect 260748 96908 260800 96960
rect 261668 96908 261720 96960
rect 262128 96908 262180 96960
rect 262588 96908 262640 96960
rect 263508 96908 263560 96960
rect 264152 96908 264204 96960
rect 264704 96908 264756 96960
rect 265624 96908 265676 96960
rect 266084 96908 266136 96960
rect 266636 96908 266688 96960
rect 267372 96908 267424 96960
rect 269488 96908 269540 96960
rect 270408 96908 270460 96960
rect 270684 96908 270736 96960
rect 271420 96908 271472 96960
rect 272248 96908 272300 96960
rect 273076 96908 273128 96960
rect 273904 96908 273956 96960
rect 274548 96908 274600 96960
rect 276572 96908 276624 96960
rect 277124 96908 277176 96960
rect 277768 96908 277820 96960
rect 278412 96908 278464 96960
rect 280160 96908 280212 96960
rect 281356 96908 281408 96960
rect 281816 96908 281868 96960
rect 282460 96908 282512 96960
rect 283196 96908 283248 96960
rect 283840 96908 283892 96960
rect 286324 96908 286376 96960
rect 286692 96908 286744 96960
rect 287520 96908 287572 96960
rect 288072 96908 288124 96960
rect 288716 96908 288768 96960
rect 289452 96908 289504 96960
rect 290096 96908 290148 96960
rect 290832 96908 290884 96960
rect 291752 96908 291804 96960
rect 292488 96908 292540 96960
rect 292764 96908 292816 96960
rect 293500 96908 293552 96960
rect 294604 96908 294656 96960
rect 295064 96908 295116 96960
rect 298836 96908 298888 96960
rect 299388 96908 299440 96960
rect 299848 96908 299900 96960
rect 300768 96908 300820 96960
rect 248788 96840 248840 96892
rect 249616 96840 249668 96892
rect 254032 96840 254084 96892
rect 255136 96840 255188 96892
rect 255412 96840 255464 96892
rect 256608 96840 256660 96892
rect 258724 96840 258776 96892
rect 259184 96840 259236 96892
rect 260104 96840 260156 96892
rect 260656 96840 260708 96892
rect 260932 96840 260984 96892
rect 262036 96840 262088 96892
rect 263140 96840 263192 96892
rect 263968 96840 264020 96892
rect 264796 96840 264848 96892
rect 265808 96840 265860 96892
rect 266268 96840 266320 96892
rect 266820 96840 266872 96892
rect 267556 96840 267608 96892
rect 269672 96840 269724 96892
rect 270316 96840 270368 96892
rect 271052 96840 271104 96892
rect 271604 96840 271656 96892
rect 271880 96840 271932 96892
rect 272984 96840 273036 96892
rect 273260 96840 273312 96892
rect 274088 96840 274140 96892
rect 276388 96840 276440 96892
rect 277216 96840 277268 96892
rect 277952 96840 278004 96892
rect 278688 96840 278740 96892
rect 278964 96840 279016 96892
rect 280068 96840 280120 96892
rect 280804 96840 280856 96892
rect 281264 96840 281316 96892
rect 282000 96840 282052 96892
rect 282644 96840 282696 96892
rect 285680 96840 285732 96892
rect 286784 96840 286836 96892
rect 287060 96840 287112 96892
rect 288164 96840 288216 96892
rect 289912 96840 289964 96892
rect 290740 96840 290792 96892
rect 291936 96840 291988 96892
rect 292304 96840 292356 96892
rect 292948 96840 293000 96892
rect 293592 96840 293644 96892
rect 294236 96840 294288 96892
rect 295156 96840 295208 96892
rect 299480 96840 299532 96892
rect 300676 96840 300728 96892
rect 246948 96772 247000 96824
rect 247500 96772 247552 96824
rect 248236 96772 248288 96824
rect 250168 96772 250220 96824
rect 250812 96772 250864 96824
rect 251180 96772 251232 96824
rect 252192 96772 252244 96824
rect 261576 96772 261628 96824
rect 261944 96772 261996 96824
rect 264336 96772 264388 96824
rect 265164 96772 265216 96824
rect 266176 96772 266228 96824
rect 267188 96772 267240 96824
rect 267648 96772 267700 96824
rect 268200 96772 268252 96824
rect 269028 96772 269080 96824
rect 269212 96772 269264 96824
rect 270224 96772 270276 96824
rect 270500 96772 270552 96824
rect 271696 96772 271748 96824
rect 275100 96772 275152 96824
rect 275744 96772 275796 96824
rect 280620 96772 280672 96824
rect 281172 96772 281224 96824
rect 281632 96772 281684 96824
rect 282828 96772 282880 96824
rect 284484 96772 284536 96824
rect 285220 96772 285272 96824
rect 285864 96772 285916 96824
rect 286876 96772 286928 96824
rect 288900 96772 288952 96824
rect 289636 96772 289688 96824
rect 290556 96772 290608 96824
rect 291016 96772 291068 96824
rect 294420 96772 294472 96824
rect 294972 96772 295024 96824
rect 295616 96772 295668 96824
rect 296260 96772 296312 96824
rect 297272 96772 297324 96824
rect 297824 96772 297876 96824
rect 211804 96704 211856 96756
rect 215116 96704 215168 96756
rect 199384 96636 199436 96688
rect 201868 96636 201920 96688
rect 206928 96636 206980 96688
rect 210608 96636 210660 96688
rect 210792 96636 210844 96688
rect 212080 96636 212132 96688
rect 213368 96636 213420 96688
rect 226984 96704 227036 96756
rect 229284 96704 229336 96756
rect 241612 96704 241664 96756
rect 242716 96704 242768 96756
rect 243084 96704 243136 96756
rect 243912 96704 243964 96756
rect 245936 96704 245988 96756
rect 246764 96704 246816 96756
rect 249800 96704 249852 96756
rect 250996 96704 251048 96756
rect 251640 96704 251692 96756
rect 252376 96704 252428 96756
rect 253020 96704 253072 96756
rect 253848 96704 253900 96756
rect 254400 96704 254452 96756
rect 258724 96704 258776 96756
rect 266360 96704 266412 96756
rect 267464 96704 267516 96756
rect 270040 96704 270092 96756
rect 222844 96636 222896 96688
rect 223488 96636 223540 96688
rect 228548 96636 228600 96688
rect 233792 96636 233844 96688
rect 234804 96636 234856 96688
rect 235264 96636 235316 96688
rect 236092 96636 236144 96688
rect 236736 96636 236788 96688
rect 237656 96636 237708 96688
rect 238484 96636 238536 96688
rect 240140 96636 240192 96688
rect 241244 96636 241296 96688
rect 248512 96636 248564 96688
rect 249432 96636 249484 96688
rect 252836 96636 252888 96688
rect 253664 96636 253716 96688
rect 257252 96636 257304 96688
rect 257804 96636 257856 96688
rect 261760 96636 261812 96688
rect 262128 96636 262180 96688
rect 262312 96636 262364 96688
rect 263324 96636 263376 96688
rect 273536 96636 273588 96688
rect 274364 96636 274416 96688
rect 274916 96704 274968 96756
rect 275836 96704 275888 96756
rect 280436 96704 280488 96756
rect 281448 96704 281500 96756
rect 284668 96704 284720 96756
rect 285404 96704 285456 96756
rect 294788 96704 294840 96756
rect 295248 96704 295300 96756
rect 296812 96704 296864 96756
rect 297732 96704 297784 96756
rect 275284 96636 275336 96688
rect 277584 96636 277636 96688
rect 278504 96636 278556 96688
rect 283472 96636 283524 96688
rect 284116 96636 284168 96688
rect 290372 96636 290424 96688
rect 291200 96636 291252 96688
rect 291384 96636 291436 96688
rect 292396 96636 292448 96688
rect 298652 96636 298704 96688
rect 299204 96636 299256 96688
rect 298008 96568 298060 96620
rect 298744 96568 298796 96620
rect 251364 96296 251416 96348
rect 302332 96296 302384 96348
rect 200028 96228 200080 96280
rect 234988 96228 235040 96280
rect 256700 96228 256752 96280
rect 329840 96228 329892 96280
rect 192484 96160 192536 96212
rect 232504 96160 232556 96212
rect 240324 96160 240376 96212
rect 240692 96160 240744 96212
rect 300584 96160 300636 96212
rect 378140 96160 378192 96212
rect 178684 96092 178736 96144
rect 222016 96092 222068 96144
rect 258080 96092 258132 96144
rect 338120 96092 338172 96144
rect 183468 96024 183520 96076
rect 231308 96024 231360 96076
rect 286048 96024 286100 96076
rect 500960 96024 501012 96076
rect 159364 95956 159416 96008
rect 222752 95956 222804 96008
rect 287336 95956 287388 96008
rect 507860 95956 507912 96008
rect 4068 95888 4120 95940
rect 200488 95888 200540 95940
rect 288532 95888 288584 95940
rect 518900 95888 518952 95940
rect 215576 95412 215628 95464
rect 216220 95412 216272 95464
rect 222936 95208 222988 95260
rect 229376 95208 229428 95260
rect 287980 95072 288032 95124
rect 295984 95072 296036 95124
rect 201592 94868 201644 94920
rect 202420 94868 202472 94920
rect 203340 94868 203392 94920
rect 203524 94868 203576 94920
rect 212724 94868 212776 94920
rect 213184 94868 213236 94920
rect 257068 94868 257120 94920
rect 318064 94868 318116 94920
rect 181444 94800 181496 94852
rect 227904 94800 227956 94852
rect 228364 94800 228416 94852
rect 254216 94800 254268 94852
rect 316040 94800 316092 94852
rect 166908 94732 166960 94784
rect 265900 94732 265952 94784
rect 375380 94732 375432 94784
rect 158628 94664 158680 94716
rect 227076 94664 227128 94716
rect 228364 94664 228416 94716
rect 143448 94596 143500 94648
rect 224408 94596 224460 94648
rect 272064 94664 272116 94716
rect 421012 94664 421064 94716
rect 236368 94596 236420 94648
rect 305000 94596 305052 94648
rect 557540 94596 557592 94648
rect 126888 94528 126940 94580
rect 221740 94528 221792 94580
rect 226708 94528 226760 94580
rect 227352 94528 227404 94580
rect 229008 94528 229060 94580
rect 43444 94460 43496 94512
rect 200396 94460 200448 94512
rect 201224 94460 201276 94512
rect 204444 94460 204496 94512
rect 204628 94460 204680 94512
rect 208492 94460 208544 94512
rect 209504 94460 209556 94512
rect 209872 94460 209924 94512
rect 210884 94460 210936 94512
rect 211528 94460 211580 94512
rect 212172 94460 212224 94512
rect 214012 94460 214064 94512
rect 214380 94460 214432 94512
rect 229376 94460 229428 94512
rect 230204 94460 230256 94512
rect 239220 94528 239272 94580
rect 263600 94528 263652 94580
rect 294604 94528 294656 94580
rect 296076 94528 296128 94580
rect 561680 94528 561732 94580
rect 204168 94392 204220 94444
rect 214196 94392 214248 94444
rect 214840 94392 214892 94444
rect 227628 94392 227680 94444
rect 237380 94460 237432 94512
rect 250352 94460 250404 94512
rect 289084 94460 289136 94512
rect 296996 94460 297048 94512
rect 565820 94460 565872 94512
rect 204628 94324 204680 94376
rect 205456 94324 205508 94376
rect 293868 93848 293920 93900
rect 297364 93848 297416 93900
rect 198648 93508 198700 93560
rect 233884 93508 233936 93560
rect 191748 93440 191800 93492
rect 232596 93440 232648 93492
rect 256332 93440 256384 93492
rect 327080 93440 327132 93492
rect 184848 93372 184900 93424
rect 231400 93372 231452 93424
rect 257896 93372 257948 93424
rect 333980 93372 334032 93424
rect 148968 93304 149020 93356
rect 225236 93304 225288 93356
rect 259184 93304 259236 93356
rect 336004 93304 336056 93356
rect 142068 93236 142120 93288
rect 224132 93236 224184 93288
rect 263324 93236 263376 93288
rect 311164 93236 311216 93288
rect 312544 93236 312596 93288
rect 539600 93236 539652 93288
rect 37188 93168 37240 93220
rect 205916 93168 205968 93220
rect 292488 93168 292540 93220
rect 546592 93168 546644 93220
rect 22008 93100 22060 93152
rect 203616 93100 203668 93152
rect 224868 93100 224920 93152
rect 238300 93100 238352 93152
rect 244188 93100 244240 93152
rect 255320 93100 255372 93152
rect 283564 93100 283616 93152
rect 294696 93100 294748 93152
rect 295248 93100 295300 93152
rect 564440 93100 564492 93152
rect 186228 92148 186280 92200
rect 231584 92148 231636 92200
rect 282184 92148 282236 92200
rect 313280 92148 313332 92200
rect 171048 92080 171100 92132
rect 226984 92080 227036 92132
rect 275376 92080 275428 92132
rect 356060 92080 356112 92132
rect 137284 92012 137336 92064
rect 222568 92012 222620 92064
rect 262128 92012 262180 92064
rect 358820 92012 358872 92064
rect 71044 91944 71096 91996
rect 211436 91944 211488 91996
rect 263416 91944 263468 91996
rect 364984 91944 365036 91996
rect 23388 91876 23440 91928
rect 203800 91876 203852 91928
rect 265992 91876 266044 91928
rect 374644 91876 374696 91928
rect 12348 91808 12400 91860
rect 195336 91808 195388 91860
rect 195888 91808 195940 91860
rect 233424 91808 233476 91860
rect 269764 91808 269816 91860
rect 380900 91808 380952 91860
rect 1308 91740 1360 91792
rect 188344 91740 188396 91792
rect 188988 91740 189040 91792
rect 232228 91740 232280 91792
rect 242808 91740 242860 91792
rect 258080 91740 258132 91792
rect 267648 91740 267700 91792
rect 389824 91740 389876 91792
rect 233148 91332 233200 91384
rect 239680 91332 239732 91384
rect 231768 91060 231820 91112
rect 236644 91060 236696 91112
rect 181536 90720 181588 90772
rect 225512 90720 225564 90772
rect 253664 90720 253716 90772
rect 307024 90720 307076 90772
rect 162216 90652 162268 90704
rect 226616 90652 226668 90704
rect 260656 90652 260708 90704
rect 347044 90652 347096 90704
rect 104164 90584 104216 90636
rect 217416 90584 217468 90636
rect 271512 90584 271564 90636
rect 412640 90584 412692 90636
rect 73068 90516 73120 90568
rect 212356 90516 212408 90568
rect 271788 90516 271840 90568
rect 416872 90516 416924 90568
rect 62028 90448 62080 90500
rect 206928 90448 206980 90500
rect 274272 90448 274324 90500
rect 427912 90448 427964 90500
rect 55128 90380 55180 90432
rect 204260 90380 204312 90432
rect 274548 90380 274600 90432
rect 430580 90380 430632 90432
rect 59268 90312 59320 90364
rect 209780 90312 209832 90364
rect 275744 90312 275796 90364
rect 438952 90312 439004 90364
rect 233608 89904 233660 89956
rect 234436 89904 234488 89956
rect 178776 89360 178828 89412
rect 229376 89360 229428 89412
rect 252284 89360 252336 89412
rect 300860 89360 300912 89412
rect 177304 89292 177356 89344
rect 230020 89292 230072 89344
rect 253296 89292 253348 89344
rect 303620 89292 303672 89344
rect 122104 89224 122156 89276
rect 214288 89224 214340 89276
rect 281172 89224 281224 89276
rect 341524 89224 341576 89276
rect 115204 89156 115256 89208
rect 214196 89156 214248 89208
rect 278320 89156 278372 89208
rect 385684 89156 385736 89208
rect 112444 89088 112496 89140
rect 219072 89088 219124 89140
rect 279884 89088 279936 89140
rect 457444 89088 457496 89140
rect 108948 89020 109000 89072
rect 218520 89020 218572 89072
rect 282460 89020 282512 89072
rect 476120 89020 476172 89072
rect 91008 88952 91060 89004
rect 206284 88952 206336 89004
rect 248052 88952 248104 89004
rect 281540 88952 281592 89004
rect 283840 88952 283892 89004
rect 484400 88952 484452 89004
rect 197176 88000 197228 88052
rect 228548 88000 228600 88052
rect 252376 88000 252428 88052
rect 309140 88000 309192 88052
rect 193128 87932 193180 87984
rect 234896 87932 234948 87984
rect 255044 87932 255096 87984
rect 317420 87932 317472 87984
rect 95148 87864 95200 87916
rect 215576 87864 215628 87916
rect 259276 87864 259328 87916
rect 339500 87864 339552 87916
rect 88984 87796 89036 87848
rect 212724 87796 212776 87848
rect 268568 87796 268620 87848
rect 396724 87796 396776 87848
rect 70308 87728 70360 87780
rect 210424 87728 210476 87780
rect 288072 87728 288124 87780
rect 489184 87728 489236 87780
rect 53748 87660 53800 87712
rect 208676 87660 208728 87712
rect 249432 87660 249484 87712
rect 285680 87660 285732 87712
rect 286692 87660 286744 87712
rect 502340 87660 502392 87712
rect 45468 87592 45520 87644
rect 207572 87592 207624 87644
rect 230388 87592 230440 87644
rect 240416 87592 240468 87644
rect 249524 87592 249576 87644
rect 287060 87592 287112 87644
rect 289452 87592 289504 87644
rect 528652 87592 528704 87644
rect 124128 86640 124180 86692
rect 221188 86640 221240 86692
rect 255136 86640 255188 86692
rect 311256 86640 311308 86692
rect 119988 86572 120040 86624
rect 220452 86572 220504 86624
rect 256516 86572 256568 86624
rect 324504 86572 324556 86624
rect 117228 86504 117280 86556
rect 219992 86504 220044 86556
rect 253756 86504 253808 86556
rect 309784 86504 309836 86556
rect 309876 86504 309928 86556
rect 425060 86504 425112 86556
rect 111064 86436 111116 86488
rect 218244 86436 218296 86488
rect 267372 86436 267424 86488
rect 387800 86436 387852 86488
rect 107016 86368 107068 86420
rect 216864 86368 216916 86420
rect 290832 86368 290884 86420
rect 515404 86368 515456 86420
rect 88248 86300 88300 86352
rect 211804 86300 211856 86352
rect 295156 86300 295208 86352
rect 547880 86300 547932 86352
rect 10968 86232 11020 86284
rect 201684 86232 201736 86284
rect 246396 86232 246448 86284
rect 252560 86232 252612 86284
rect 296352 86232 296404 86284
rect 572720 86232 572772 86284
rect 232504 85552 232556 85604
rect 238852 85552 238904 85604
rect 3148 85484 3200 85536
rect 14464 85484 14516 85536
rect 262956 85212 263008 85264
rect 357440 85212 357492 85264
rect 187056 85144 187108 85196
rect 229192 85144 229244 85196
rect 261852 85144 261904 85196
rect 360200 85144 360252 85196
rect 184204 85076 184256 85128
rect 231032 85076 231084 85128
rect 264336 85076 264388 85128
rect 367100 85076 367152 85128
rect 119344 85008 119396 85060
rect 219624 85008 219676 85060
rect 266084 85008 266136 85060
rect 382280 85008 382332 85060
rect 68928 84940 68980 84992
rect 211896 84940 211948 84992
rect 278412 84940 278464 84992
rect 449164 84940 449216 84992
rect 50988 84872 51040 84924
rect 208584 84872 208636 84924
rect 288164 84872 288216 84924
rect 506480 84872 506532 84924
rect 15108 84804 15160 84856
rect 201592 84804 201644 84856
rect 202236 84804 202288 84856
rect 233056 84804 233108 84856
rect 243912 84804 243964 84856
rect 258172 84804 258224 84856
rect 286784 84804 286836 84856
rect 510712 84804 510764 84856
rect 191656 83784 191708 83836
rect 232228 83784 232280 83836
rect 268844 83784 268896 83836
rect 398932 83784 398984 83836
rect 182824 83716 182876 83768
rect 225052 83716 225104 83768
rect 270132 83716 270184 83768
rect 406384 83716 406436 83768
rect 111708 83648 111760 83700
rect 218796 83648 218848 83700
rect 271604 83648 271656 83700
rect 414020 83648 414072 83700
rect 103428 83580 103480 83632
rect 216772 83580 216824 83632
rect 279516 83580 279568 83632
rect 434720 83580 434772 83632
rect 96528 83512 96580 83564
rect 216404 83512 216456 83564
rect 277124 83512 277176 83564
rect 445760 83512 445812 83564
rect 89628 83444 89680 83496
rect 213184 83444 213236 83496
rect 226984 83444 227036 83496
rect 236552 83444 236604 83496
rect 297824 83444 297876 83496
rect 571340 83444 571392 83496
rect 190368 82492 190420 82544
rect 233884 82492 233936 82544
rect 175188 82424 175240 82476
rect 229560 82424 229612 82476
rect 282644 82424 282696 82476
rect 453304 82424 453356 82476
rect 168288 82356 168340 82408
rect 224224 82356 224276 82408
rect 279976 82356 280028 82408
rect 463700 82356 463752 82408
rect 170404 82288 170456 82340
rect 226800 82288 226852 82340
rect 281264 82288 281316 82340
rect 470600 82288 470652 82340
rect 136548 82220 136600 82272
rect 222292 82220 222344 82272
rect 284116 82220 284168 82272
rect 485780 82220 485832 82272
rect 106188 82152 106240 82204
rect 214564 82152 214616 82204
rect 286876 82152 286928 82204
rect 499580 82152 499632 82204
rect 47676 82084 47728 82136
rect 206652 82084 206704 82136
rect 248144 82084 248196 82136
rect 278780 82084 278832 82136
rect 290924 82084 290976 82136
rect 525064 82084 525116 82136
rect 223488 81404 223540 81456
rect 228456 81404 228508 81456
rect 253848 81064 253900 81116
rect 307852 81064 307904 81116
rect 256608 80996 256660 81048
rect 322940 80996 322992 81048
rect 272892 80928 272944 80980
rect 411904 80928 411956 80980
rect 164148 80860 164200 80912
rect 227996 80860 228048 80912
rect 292304 80860 292356 80912
rect 535460 80860 535512 80912
rect 161388 80792 161440 80844
rect 226708 80792 226760 80844
rect 240508 80792 240560 80844
rect 252652 80792 252704 80844
rect 254584 80792 254636 80844
rect 291200 80792 291252 80844
rect 293684 80792 293736 80844
rect 542360 80792 542412 80844
rect 115848 80724 115900 80776
rect 217324 80724 217376 80776
rect 250904 80724 250956 80776
rect 295340 80724 295392 80776
rect 296536 80724 296588 80776
rect 560300 80724 560352 80776
rect 98736 80656 98788 80708
rect 215392 80656 215444 80708
rect 252192 80656 252244 80708
rect 297456 80656 297508 80708
rect 297732 80656 297784 80708
rect 578240 80656 578292 80708
rect 262864 79568 262916 79620
rect 350540 79568 350592 79620
rect 119896 79500 119948 79552
rect 219900 79500 219952 79552
rect 262036 79500 262088 79552
rect 354680 79500 354732 79552
rect 113088 79432 113140 79484
rect 218428 79432 218480 79484
rect 261944 79432 261996 79484
rect 357532 79432 357584 79484
rect 86224 79364 86276 79416
rect 208492 79364 208544 79416
rect 282552 79364 282604 79416
rect 481640 79364 481692 79416
rect 75828 79296 75880 79348
rect 212816 79296 212868 79348
rect 245200 79296 245252 79348
rect 260840 79296 260892 79348
rect 299204 79296 299256 79348
rect 582840 79296 582892 79348
rect 267464 78140 267516 78192
rect 386420 78140 386472 78192
rect 257344 78072 257396 78124
rect 266360 78072 266412 78124
rect 268936 78072 268988 78124
rect 400220 78072 400272 78124
rect 251824 78004 251876 78056
rect 262220 78004 262272 78056
rect 275284 78004 275336 78056
rect 407212 78004 407264 78056
rect 42708 77936 42760 77988
rect 207112 77936 207164 77988
rect 220728 77936 220780 77988
rect 237472 77936 237524 77988
rect 244004 77936 244056 77988
rect 267832 77936 267884 77988
rect 272984 77936 273036 77988
rect 418160 77936 418212 77988
rect 172428 76916 172480 76968
rect 222936 76916 222988 76968
rect 153016 76848 153068 76900
rect 225328 76848 225380 76900
rect 144736 76780 144788 76832
rect 223672 76780 223724 76832
rect 139308 76712 139360 76764
rect 223856 76712 223908 76764
rect 278504 76712 278556 76764
rect 432604 76712 432656 76764
rect 136456 76644 136508 76696
rect 222660 76644 222712 76696
rect 277216 76644 277268 76696
rect 436744 76644 436796 76696
rect 126796 76576 126848 76628
rect 221464 76576 221516 76628
rect 246304 76576 246356 76628
rect 251180 76576 251232 76628
rect 279424 76576 279476 76628
rect 448612 76576 448664 76628
rect 17868 76508 17920 76560
rect 200948 76508 201000 76560
rect 245292 76508 245344 76560
rect 263600 76508 263652 76560
rect 296260 76508 296312 76560
rect 569960 76508 570012 76560
rect 242532 75828 242584 75880
rect 244280 75828 244332 75880
rect 260288 75420 260340 75472
rect 336740 75420 336792 75472
rect 264244 75352 264296 75404
rect 346400 75352 346452 75404
rect 282736 75284 282788 75336
rect 481732 75284 481784 75336
rect 284208 75216 284260 75268
rect 488540 75216 488592 75268
rect 245384 75148 245436 75200
rect 269212 75148 269264 75200
rect 285220 75148 285272 75200
rect 491300 75148 491352 75200
rect 273076 74128 273128 74180
rect 420920 74128 420972 74180
rect 285312 74060 285364 74112
rect 495440 74060 495492 74112
rect 99288 73992 99340 74044
rect 215944 73992 215996 74044
rect 288256 73992 288308 74044
rect 513380 73992 513432 74044
rect 85488 73924 85540 73976
rect 214012 73924 214064 73976
rect 289544 73924 289596 73976
rect 521660 73924 521712 73976
rect 48228 73856 48280 73908
rect 202328 73856 202380 73908
rect 291016 73856 291068 73908
rect 527180 73856 527232 73908
rect 31668 73788 31720 73840
rect 205088 73788 205140 73840
rect 250996 73788 251048 73840
rect 298100 73788 298152 73840
rect 299296 73788 299348 73840
rect 582748 73788 582800 73840
rect 261760 72700 261812 72752
rect 336096 72700 336148 72752
rect 263508 72632 263560 72684
rect 364340 72632 364392 72684
rect 256056 72564 256108 72616
rect 259460 72564 259512 72616
rect 276756 72564 276808 72616
rect 396080 72564 396132 72616
rect 403624 72564 403676 72616
rect 449900 72564 449952 72616
rect 274364 72496 274416 72548
rect 427820 72496 427872 72548
rect 292396 72428 292448 72480
rect 531412 72428 531464 72480
rect 3424 71680 3476 71732
rect 35164 71680 35216 71732
rect 121368 71340 121420 71392
rect 219808 71340 219860 71392
rect 64788 71272 64840 71324
rect 209872 71272 209924 71324
rect 61936 71204 61988 71256
rect 209964 71204 210016 71256
rect 267556 71204 267608 71256
rect 389180 71204 389232 71256
rect 53656 71136 53708 71188
rect 208860 71136 208912 71188
rect 270224 71136 270276 71188
rect 402980 71136 403032 71188
rect 45376 71068 45428 71120
rect 207296 71068 207348 71120
rect 271696 71068 271748 71120
rect 409880 71068 409932 71120
rect 38568 71000 38620 71052
rect 206008 71000 206060 71052
rect 248236 71000 248288 71052
rect 267004 71000 267056 71052
rect 281356 71000 281408 71052
rect 466460 71000 466512 71052
rect 259092 69980 259144 70032
rect 340972 69980 341024 70032
rect 266176 69912 266228 69964
rect 378784 69912 378836 69964
rect 274456 69844 274508 69896
rect 431224 69844 431276 69896
rect 276664 69776 276716 69828
rect 438860 69776 438912 69828
rect 278596 69708 278648 69760
rect 456892 69708 456944 69760
rect 253204 69640 253256 69692
rect 276112 69640 276164 69692
rect 280068 69640 280120 69692
rect 459560 69640 459612 69692
rect 125416 68416 125468 68468
rect 221280 68416 221332 68468
rect 20628 68348 20680 68400
rect 203340 68348 203392 68400
rect 267280 68348 267332 68400
rect 390652 68348 390704 68400
rect 6828 68280 6880 68332
rect 201040 68280 201092 68332
rect 240324 68280 240376 68332
rect 249892 68280 249944 68332
rect 275836 68280 275888 68332
rect 436100 68280 436152 68332
rect 272800 66852 272852 66904
rect 422300 66852 422352 66904
rect 285404 65492 285456 65544
rect 492680 65492 492732 65544
rect 300676 64132 300728 64184
rect 582656 64132 582708 64184
rect 275928 62772 275980 62824
rect 440332 62772 440384 62824
rect 3056 59304 3108 59356
rect 140044 59304 140096 59356
rect 274180 53048 274232 53100
rect 429200 53048 429252 53100
rect 44088 51688 44140 51740
rect 200764 51688 200816 51740
rect 246764 51688 246816 51740
rect 273260 51688 273312 51740
rect 281448 51688 281500 51740
rect 467840 51688 467892 51740
rect 71688 47540 71740 47592
rect 211528 47540 211580 47592
rect 244096 47540 244148 47592
rect 256700 47540 256752 47592
rect 257804 47540 257856 47592
rect 332692 47540 332744 47592
rect 249616 46180 249668 46232
rect 285772 46180 285824 46232
rect 286600 46180 286652 46232
rect 503720 46180 503772 46232
rect 247684 45772 247736 45824
rect 248420 45772 248472 45824
rect 3424 45500 3476 45552
rect 106924 45500 106976 45552
rect 78588 43392 78640 43444
rect 212908 43392 212960 43444
rect 213184 43392 213236 43444
rect 236736 43392 236788 43444
rect 243820 42712 243872 42764
rect 249800 42712 249852 42764
rect 219348 42032 219400 42084
rect 231216 42032 231268 42084
rect 250444 42032 250496 42084
rect 267740 42032 267792 42084
rect 269028 42032 269080 42084
rect 397460 42032 397512 42084
rect 242624 41420 242676 41472
rect 242900 41420 242952 41472
rect 292212 39312 292264 39364
rect 300124 39312 300176 39364
rect 211804 35164 211856 35216
rect 234712 35164 234764 35216
rect 300768 35164 300820 35216
rect 582564 35164 582616 35216
rect 2872 33056 2924 33108
rect 47584 33056 47636 33108
rect 242716 28908 242768 28960
rect 245660 28908 245712 28960
rect 246856 28228 246908 28280
rect 262864 28228 262916 28280
rect 46848 25508 46900 25560
rect 86316 25508 86368 25560
rect 12256 24080 12308 24132
rect 199384 24080 199436 24132
rect 291108 24080 291160 24132
rect 528560 24080 528612 24132
rect 238944 23536 238996 23588
rect 240232 23536 240284 23588
rect 238668 22720 238720 22772
rect 241520 22720 241572 22772
rect 353944 22720 353996 22772
rect 460940 22720 460992 22772
rect 238024 22040 238076 22092
rect 240600 22040 240652 22092
rect 282828 21360 282880 21412
rect 474740 21360 474792 21412
rect 3424 20612 3476 20664
rect 98644 20612 98696 20664
rect 278688 19932 278740 19984
rect 454040 19932 454092 19984
rect 33048 18572 33100 18624
rect 204628 18572 204680 18624
rect 100668 17212 100720 17264
rect 217048 17212 217100 17264
rect 277308 17212 277360 17264
rect 443000 17212 443052 17264
rect 86868 15852 86920 15904
rect 214748 15852 214800 15904
rect 293776 15852 293828 15904
rect 546500 15852 546552 15904
rect 266268 14492 266320 14544
rect 383568 14492 383620 14544
rect 289636 14424 289688 14476
rect 517520 14424 517572 14476
rect 94504 13064 94556 13116
rect 215760 13064 215812 13116
rect 217968 13064 218020 13116
rect 236276 13064 236328 13116
rect 285496 13064 285548 13116
rect 497096 13064 497148 13116
rect 260748 11840 260800 11892
rect 348056 11840 348108 11892
rect 264796 11772 264848 11824
rect 372896 11772 372948 11824
rect 398932 11772 398984 11824
rect 400128 11772 400180 11824
rect 407212 11772 407264 11824
rect 408408 11772 408460 11824
rect 37096 11704 37148 11756
rect 101404 11704 101456 11756
rect 242900 11704 242952 11756
rect 244096 11704 244148 11756
rect 251180 11704 251232 11756
rect 252376 11704 252428 11756
rect 295984 11704 296036 11756
rect 416780 11704 416832 11756
rect 423772 11704 423824 11756
rect 424968 11704 425020 11756
rect 307852 11636 307904 11688
rect 309048 11636 309100 11688
rect 332692 11636 332744 11688
rect 333888 11636 333940 11688
rect 357532 11636 357584 11688
rect 358728 11636 358780 11688
rect 216588 10276 216640 10328
rect 222844 10276 222896 10328
rect 271420 10276 271472 10328
rect 411812 10276 411864 10328
rect 461584 10276 461636 10328
rect 472256 10276 472308 10328
rect 254860 9324 254912 9376
rect 319720 9324 319772 9376
rect 264704 9256 264756 9308
rect 374092 9256 374144 9308
rect 270316 9188 270368 9240
rect 406016 9188 406068 9240
rect 294696 9120 294748 9172
rect 459192 9120 459244 9172
rect 287980 9052 288032 9104
rect 511264 9052 511316 9104
rect 289360 8984 289412 9036
rect 520740 8984 520792 9036
rect 210976 8916 211028 8968
rect 225604 8916 225656 8968
rect 299388 8916 299440 8968
rect 576308 8916 576360 8968
rect 250812 7692 250864 7744
rect 292580 7692 292632 7744
rect 260196 7624 260248 7676
rect 331588 7624 331640 7676
rect 5264 7556 5316 7608
rect 46204 7556 46256 7608
rect 260104 7556 260156 7608
rect 270040 7556 270092 7608
rect 270408 7556 270460 7608
rect 404820 7556 404872 7608
rect 454684 7556 454736 7608
rect 465172 7556 465224 7608
rect 468484 7556 468536 7608
rect 479340 7556 479392 7608
rect 3424 6808 3476 6860
rect 133144 6808 133196 6860
rect 258724 6468 258776 6520
rect 317328 6468 317380 6520
rect 294604 6400 294656 6452
rect 370596 6400 370648 6452
rect 285588 6332 285640 6384
rect 498200 6332 498252 6384
rect 245476 6264 245528 6316
rect 259828 6264 259880 6316
rect 293500 6264 293552 6316
rect 540796 6264 540848 6316
rect 248328 6196 248380 6248
rect 280712 6196 280764 6248
rect 297364 6196 297416 6248
rect 544384 6196 544436 6248
rect 249708 6128 249760 6180
rect 286600 6128 286652 6180
rect 298744 6128 298796 6180
rect 569132 6128 569184 6180
rect 281908 5516 281960 5568
rect 283472 5516 283524 5568
rect 443644 5516 443696 5568
rect 447416 5516 447468 5568
rect 59636 4836 59688 4888
rect 93124 4836 93176 4888
rect 80888 4768 80940 4820
rect 209044 4768 209096 4820
rect 233424 4428 233476 4480
rect 239128 4428 239180 4480
rect 28908 4156 28960 4208
rect 32404 4156 32456 4208
rect 242440 4156 242492 4208
rect 246396 4156 246448 4208
rect 130568 4088 130620 4140
rect 133236 4088 133288 4140
rect 161296 4088 161348 4140
rect 162124 4088 162176 4140
rect 168380 4088 168432 4140
rect 173164 4088 173216 4140
rect 290188 4088 290240 4140
rect 298100 4088 298152 4140
rect 323584 4088 323636 4140
rect 324412 4088 324464 4140
rect 402520 4088 402572 4140
rect 403072 4088 403124 4140
rect 431224 4088 431276 4140
rect 432052 4088 432104 4140
rect 363604 4020 363656 4072
rect 365812 4020 365864 4072
rect 40776 3952 40828 4004
rect 47676 3952 47728 4004
rect 101036 3952 101088 4004
rect 104164 3952 104216 4004
rect 171784 3952 171836 4004
rect 181536 3952 181588 4004
rect 193220 3952 193272 4004
rect 202236 3952 202288 4004
rect 208584 3952 208636 4004
rect 211804 3952 211856 4004
rect 171876 3884 171928 3936
rect 182824 3884 182876 3936
rect 225144 3884 225196 3936
rect 237656 3884 237708 3936
rect 131764 3816 131816 3868
rect 137284 3816 137336 3868
rect 189724 3816 189776 3868
rect 192484 3816 192536 3868
rect 226340 3816 226392 3868
rect 232504 3816 232556 3868
rect 247592 3816 247644 3868
rect 258080 3816 258132 3868
rect 8760 3680 8812 3732
rect 18604 3680 18656 3732
rect 35900 3680 35952 3732
rect 39304 3680 39356 3732
rect 18236 3612 18288 3664
rect 28264 3612 28316 3664
rect 1676 3544 1728 3596
rect 4804 3544 4856 3596
rect 24216 3544 24268 3596
rect 43444 3612 43496 3664
rect 56048 3612 56100 3664
rect 66720 3680 66772 3732
rect 44272 3544 44324 3596
rect 45376 3544 45428 3596
rect 52552 3544 52604 3596
rect 53656 3544 53708 3596
rect 57244 3544 57296 3596
rect 57888 3544 57940 3596
rect 58440 3544 58492 3596
rect 59268 3544 59320 3596
rect 60832 3544 60884 3596
rect 61936 3544 61988 3596
rect 65524 3544 65576 3596
rect 66168 3544 66220 3596
rect 67916 3544 67968 3596
rect 68928 3544 68980 3596
rect 72608 3544 72660 3596
rect 73068 3544 73120 3596
rect 77392 3748 77444 3800
rect 88984 3748 89036 3800
rect 103520 3748 103572 3800
rect 107016 3748 107068 3800
rect 132960 3748 133012 3800
rect 74908 3680 74960 3732
rect 80704 3680 80756 3732
rect 86224 3680 86276 3732
rect 86776 3680 86828 3732
rect 115112 3680 115164 3732
rect 101496 3612 101548 3664
rect 84476 3544 84528 3596
rect 85488 3544 85540 3596
rect 89168 3544 89220 3596
rect 89628 3544 89680 3596
rect 90364 3544 90416 3596
rect 91008 3544 91060 3596
rect 91560 3544 91612 3596
rect 92388 3544 92440 3596
rect 97448 3544 97500 3596
rect 97908 3544 97960 3596
rect 98644 3544 98696 3596
rect 99288 3544 99340 3596
rect 99840 3544 99892 3596
rect 100668 3544 100720 3596
rect 102232 3544 102284 3596
rect 103520 3544 103572 3596
rect 572 3476 624 3528
rect 1308 3476 1360 3528
rect 2872 3476 2924 3528
rect 3976 3476 4028 3528
rect 9956 3476 10008 3528
rect 10968 3476 11020 3528
rect 11152 3476 11204 3528
rect 12256 3476 12308 3528
rect 13544 3476 13596 3528
rect 35900 3476 35952 3528
rect 35992 3476 36044 3528
rect 37096 3476 37148 3528
rect 41880 3476 41932 3528
rect 42708 3476 42760 3528
rect 43076 3476 43128 3528
rect 44088 3476 44140 3528
rect 48964 3476 49016 3528
rect 49608 3476 49660 3528
rect 50160 3476 50212 3528
rect 50988 3476 51040 3528
rect 51356 3476 51408 3528
rect 74908 3476 74960 3528
rect 75000 3476 75052 3528
rect 75828 3476 75880 3528
rect 76196 3476 76248 3528
rect 77208 3476 77260 3528
rect 83280 3476 83332 3528
rect 122104 3612 122156 3664
rect 125508 3612 125560 3664
rect 110512 3544 110564 3596
rect 111708 3544 111760 3596
rect 117596 3544 117648 3596
rect 119344 3544 119396 3596
rect 128176 3544 128228 3596
rect 137652 3680 137704 3732
rect 158904 3748 158956 3800
rect 170404 3748 170456 3800
rect 159364 3680 159416 3732
rect 162492 3680 162544 3732
rect 173164 3748 173216 3800
rect 187056 3748 187108 3800
rect 190368 3748 190420 3800
rect 199108 3748 199160 3800
rect 200028 3748 200080 3800
rect 203892 3748 203944 3800
rect 220452 3748 220504 3800
rect 231124 3748 231176 3800
rect 262864 3748 262916 3800
rect 271236 3748 271288 3800
rect 181444 3680 181496 3732
rect 218060 3680 218112 3732
rect 219348 3680 219400 3732
rect 238116 3680 238168 3732
rect 249892 3680 249944 3732
rect 258264 3680 258316 3732
rect 269212 3680 269264 3732
rect 310244 3680 310296 3732
rect 320180 3884 320232 3936
rect 326436 3884 326488 3936
rect 145932 3612 145984 3664
rect 104532 3476 104584 3528
rect 105544 3476 105596 3528
rect 105728 3476 105780 3528
rect 106188 3476 106240 3528
rect 108120 3476 108172 3528
rect 108948 3476 109000 3528
rect 109316 3476 109368 3528
rect 111064 3476 111116 3528
rect 111616 3476 111668 3528
rect 112444 3476 112496 3528
rect 114008 3476 114060 3528
rect 114468 3476 114520 3528
rect 115204 3476 115256 3528
rect 115848 3476 115900 3528
rect 116400 3476 116452 3528
rect 117228 3476 117280 3528
rect 118792 3476 118844 3528
rect 119804 3476 119856 3528
rect 122288 3476 122340 3528
rect 122748 3476 122800 3528
rect 123484 3476 123536 3528
rect 124128 3476 124180 3528
rect 124680 3476 124732 3528
rect 125416 3476 125468 3528
rect 125876 3476 125928 3528
rect 126796 3476 126848 3528
rect 129372 3476 129424 3528
rect 130384 3476 130436 3528
rect 134156 3544 134208 3596
rect 135168 3544 135220 3596
rect 138848 3544 138900 3596
rect 139308 3544 139360 3596
rect 141240 3544 141292 3596
rect 142068 3544 142120 3596
rect 143540 3544 143592 3596
rect 144828 3544 144880 3596
rect 148324 3544 148376 3596
rect 148968 3544 149020 3596
rect 149520 3612 149572 3664
rect 171784 3612 171836 3664
rect 193128 3612 193180 3664
rect 171876 3544 171928 3596
rect 171968 3544 172020 3596
rect 172428 3544 172480 3596
rect 178684 3544 178736 3596
rect 174268 3476 174320 3528
rect 175188 3476 175240 3528
rect 179052 3476 179104 3528
rect 180064 3476 180116 3528
rect 180248 3476 180300 3528
rect 195244 3544 195296 3596
rect 197268 3612 197320 3664
rect 207388 3612 207440 3664
rect 213368 3612 213420 3664
rect 226984 3612 227036 3664
rect 205088 3544 205140 3596
rect 219256 3544 219308 3596
rect 233884 3612 233936 3664
rect 239312 3612 239364 3664
rect 252652 3612 252704 3664
rect 254676 3612 254728 3664
rect 267832 3612 267884 3664
rect 268476 3612 268528 3664
rect 318156 3748 318208 3800
rect 182548 3476 182600 3528
rect 183468 3476 183520 3528
rect 183744 3476 183796 3528
rect 184848 3476 184900 3528
rect 184940 3476 184992 3528
rect 186228 3476 186280 3528
rect 187332 3476 187384 3528
rect 188344 3476 188396 3528
rect 188528 3476 188580 3528
rect 188988 3476 189040 3528
rect 190828 3476 190880 3528
rect 191656 3476 191708 3528
rect 197912 3476 197964 3528
rect 198648 3476 198700 3528
rect 200304 3476 200356 3528
rect 201408 3476 201460 3528
rect 201500 3476 201552 3528
rect 233608 3544 233660 3596
rect 245568 3544 245620 3596
rect 265348 3544 265400 3596
rect 267004 3544 267056 3596
rect 277124 3544 277176 3596
rect 296076 3544 296128 3596
rect 303712 3544 303764 3596
rect 311164 3544 311216 3596
rect 331864 3884 331916 3936
rect 327724 3816 327776 3868
rect 344560 3816 344612 3868
rect 336096 3748 336148 3800
rect 449164 3816 449216 3868
rect 453304 3816 453356 3868
rect 336280 3680 336332 3732
rect 349252 3748 349304 3800
rect 416780 3748 416832 3800
rect 417884 3748 417936 3800
rect 436744 3748 436796 3800
rect 445024 3748 445076 3800
rect 450636 3748 450688 3800
rect 458088 3748 458140 3800
rect 506480 3748 506532 3800
rect 517612 3884 517664 3936
rect 575112 3884 575164 3936
rect 582840 3884 582892 3936
rect 515404 3816 515456 3868
rect 525432 3816 525484 3868
rect 566832 3816 566884 3868
rect 571340 3816 571392 3868
rect 572720 3816 572772 3868
rect 583300 3816 583352 3868
rect 517152 3748 517204 3800
rect 362316 3680 362368 3732
rect 409880 3680 409932 3732
rect 410800 3680 410852 3732
rect 411904 3680 411956 3732
rect 423772 3680 423824 3732
rect 432604 3680 432656 3732
rect 452108 3680 452160 3732
rect 453396 3680 453448 3732
rect 478144 3680 478196 3732
rect 499396 3680 499448 3732
rect 510712 3680 510764 3732
rect 515956 3680 516008 3732
rect 518900 3680 518952 3732
rect 525064 3748 525116 3800
rect 531320 3748 531372 3800
rect 556160 3748 556212 3800
rect 568580 3748 568632 3800
rect 570328 3748 570380 3800
rect 583208 3748 583260 3800
rect 528652 3680 528704 3732
rect 534908 3680 534960 3732
rect 546592 3680 546644 3732
rect 563244 3680 563296 3732
rect 575572 3680 575624 3732
rect 371700 3612 371752 3664
rect 374644 3612 374696 3664
rect 384764 3612 384816 3664
rect 385684 3612 385736 3664
rect 455696 3612 455748 3664
rect 475476 3612 475528 3664
rect 487620 3612 487672 3664
rect 491116 3612 491168 3664
rect 494060 3612 494112 3664
rect 497464 3612 497516 3664
rect 523040 3612 523092 3664
rect 524236 3612 524288 3664
rect 536840 3612 536892 3664
rect 541992 3612 542044 3664
rect 554780 3612 554832 3664
rect 557356 3612 557408 3664
rect 569960 3612 570012 3664
rect 571524 3612 571576 3664
rect 583484 3612 583536 3664
rect 231032 3476 231084 3528
rect 231768 3476 231820 3528
rect 232228 3476 232280 3528
rect 233148 3476 233200 3528
rect 237012 3476 237064 3528
rect 238024 3476 238076 3528
rect 246948 3476 247000 3528
rect 272432 3476 272484 3528
rect 278320 3476 278372 3528
rect 278780 3476 278832 3528
rect 279516 3476 279568 3528
rect 281540 3476 281592 3528
rect 284300 3476 284352 3528
rect 285772 3476 285824 3528
rect 294880 3476 294932 3528
rect 295340 3476 295392 3528
rect 297456 3476 297508 3528
rect 298468 3476 298520 3528
rect 300768 3476 300820 3528
rect 309140 3476 309192 3528
rect 309784 3476 309836 3528
rect 311440 3476 311492 3528
rect 332692 3544 332744 3596
rect 341524 3544 341576 3596
rect 469864 3544 469916 3596
rect 472624 3544 472676 3596
rect 473452 3544 473504 3596
rect 481640 3544 481692 3596
rect 482836 3544 482888 3596
rect 489184 3544 489236 3596
rect 510068 3544 510120 3596
rect 519544 3544 519596 3596
rect 520372 3544 520424 3596
rect 522304 3544 522356 3596
rect 550272 3544 550324 3596
rect 552664 3544 552716 3596
rect 564348 3544 564400 3596
rect 564440 3544 564492 3596
rect 578240 3544 578292 3596
rect 363512 3476 363564 3528
rect 364984 3476 365036 3528
rect 367008 3476 367060 3528
rect 370504 3476 370556 3528
rect 551468 3476 551520 3528
rect 559748 3476 559800 3528
rect 572812 3476 572864 3528
rect 4068 3408 4120 3460
rect 15844 3408 15896 3460
rect 17040 3408 17092 3460
rect 17868 3408 17920 3460
rect 19432 3408 19484 3460
rect 20628 3408 20680 3460
rect 25320 3408 25372 3460
rect 26148 3408 26200 3460
rect 26516 3408 26568 3460
rect 27528 3408 27580 3460
rect 32404 3408 32456 3460
rect 33048 3408 33100 3460
rect 33600 3408 33652 3460
rect 34428 3408 34480 3460
rect 203248 3408 203300 3460
rect 213920 3408 213972 3460
rect 214472 3408 214524 3460
rect 216864 3408 216916 3460
rect 217968 3408 218020 3460
rect 92756 3340 92808 3392
rect 94504 3340 94556 3392
rect 153108 3340 153160 3392
rect 154212 3340 154264 3392
rect 155408 3340 155460 3392
rect 155868 3340 155920 3392
rect 157800 3340 157852 3392
rect 158628 3340 158680 3392
rect 163688 3340 163740 3392
rect 164148 3340 164200 3392
rect 164884 3340 164936 3392
rect 165528 3340 165580 3392
rect 166080 3340 166132 3392
rect 166908 3340 166960 3392
rect 167184 3340 167236 3392
rect 168288 3340 168340 3392
rect 181444 3340 181496 3392
rect 184204 3340 184256 3392
rect 212172 3340 212224 3392
rect 220728 3408 220780 3460
rect 221556 3408 221608 3460
rect 222752 3408 222804 3460
rect 223488 3408 223540 3460
rect 223948 3408 224000 3460
rect 224868 3408 224920 3460
rect 229836 3408 229888 3460
rect 240232 3408 240284 3460
rect 242900 3408 242952 3460
rect 245660 3408 245712 3460
rect 249064 3408 249116 3460
rect 274824 3408 274876 3460
rect 275284 3408 275336 3460
rect 288992 3408 289044 3460
rect 300124 3408 300176 3460
rect 537208 3408 537260 3460
rect 554964 3408 555016 3460
rect 574100 3476 574152 3528
rect 577412 3476 577464 3528
rect 582748 3476 582800 3528
rect 573916 3408 573968 3460
rect 583116 3408 583168 3460
rect 228364 3340 228416 3392
rect 267832 3340 267884 3392
rect 273260 3340 273312 3392
rect 299664 3340 299716 3392
rect 302332 3340 302384 3392
rect 374000 3340 374052 3392
rect 375288 3340 375340 3392
rect 378784 3340 378836 3392
rect 379980 3340 380032 3392
rect 396724 3340 396776 3392
rect 398932 3340 398984 3392
rect 406384 3340 406436 3392
rect 407212 3340 407264 3392
rect 420184 3340 420236 3392
rect 421012 3340 421064 3392
rect 427268 3340 427320 3392
rect 427912 3340 427964 3392
rect 440240 3340 440292 3392
rect 441528 3340 441580 3392
rect 493324 3340 493376 3392
rect 494704 3340 494756 3392
rect 504364 3340 504416 3392
rect 505376 3340 505428 3392
rect 20628 3272 20680 3324
rect 34796 3272 34848 3324
rect 35808 3272 35860 3324
rect 64328 3272 64380 3324
rect 64788 3272 64840 3324
rect 106924 3272 106976 3324
rect 107568 3272 107620 3324
rect 135260 3272 135312 3324
rect 136548 3272 136600 3324
rect 151820 3272 151872 3324
rect 156604 3272 156656 3324
rect 156696 3272 156748 3324
rect 162216 3272 162268 3324
rect 336004 3272 336056 3324
rect 342168 3272 342220 3324
rect 367836 3272 367888 3324
rect 369400 3272 369452 3324
rect 93952 3204 94004 3256
rect 98736 3204 98788 3256
rect 209780 3204 209832 3256
rect 213184 3204 213236 3256
rect 215668 3204 215720 3256
rect 216588 3204 216640 3256
rect 259828 3204 259880 3256
rect 261760 3204 261812 3256
rect 296168 3204 296220 3256
rect 297272 3204 297324 3256
rect 39580 3136 39632 3188
rect 40684 3136 40736 3188
rect 73804 3136 73856 3188
rect 75184 3136 75236 3188
rect 147128 3136 147180 3188
rect 147588 3136 147640 3188
rect 160100 3136 160152 3188
rect 161388 3136 161440 3188
rect 230388 3136 230440 3188
rect 235816 3136 235868 3188
rect 251180 3136 251232 3188
rect 258172 3136 258224 3188
rect 311256 3136 311308 3188
rect 315028 3136 315080 3188
rect 320916 3068 320968 3120
rect 324320 3068 324372 3120
rect 347044 3068 347096 3120
rect 350448 3068 350500 3120
rect 457444 3068 457496 3120
rect 462780 3068 462832 3120
rect 547880 3068 547932 3120
rect 550640 3068 550692 3120
rect 27712 3000 27764 3052
rect 35256 3000 35308 3052
rect 69112 3000 69164 3052
rect 71044 3000 71096 3052
rect 85672 3000 85724 3052
rect 86868 3000 86920 3052
rect 176660 3000 176712 3052
rect 178776 3000 178828 3052
rect 191564 3000 191616 3052
rect 192024 3000 192076 3052
rect 389824 3000 389876 3052
rect 391848 3000 391900 3052
rect 437940 3000 437992 3052
rect 438952 3000 439004 3052
rect 447784 3000 447836 3052
rect 448612 3000 448664 3052
rect 479524 3000 479576 3052
rect 480536 3000 480588 3052
rect 578608 3000 578660 3052
rect 582380 3000 582432 3052
rect 175464 2932 175516 2984
rect 177304 2932 177356 2984
rect 283104 2932 283156 2984
rect 285680 2932 285732 2984
rect 316684 2932 316736 2984
rect 322112 2932 322164 2984
rect 82084 2864 82136 2916
rect 83464 2864 83516 2916
rect 142436 2864 142488 2916
rect 143448 2864 143500 2916
rect 186136 2864 186188 2916
rect 186964 2864 187016 2916
rect 289084 2864 289136 2916
rect 293684 2864 293736 2916
rect 307024 2864 307076 2916
rect 307944 2864 307996 2916
rect 429844 2864 429896 2916
rect 434444 2864 434496 2916
rect 150624 2252 150676 2304
rect 207664 2252 207716 2304
rect 140044 2184 140096 2236
rect 202144 2184 202196 2236
rect 63224 2116 63276 2168
rect 210148 2116 210200 2168
rect 7656 2048 7708 2100
rect 200396 2048 200448 2100
rect 206192 2048 206244 2100
rect 235080 2048 235132 2100
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 89364 703582 89668 703610
rect 8128 702434 8156 703520
rect 8128 702406 8248 702434
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 3436 683194 3464 684247
rect 3424 683188 3476 683194
rect 3424 683130 3476 683136
rect 3514 671256 3570 671265
rect 3514 671191 3570 671200
rect 3528 670750 3556 671191
rect 3516 670744 3568 670750
rect 3516 670686 3568 670692
rect 3422 658200 3478 658209
rect 3422 658135 3478 658144
rect 3436 656946 3464 658135
rect 3424 656940 3476 656946
rect 3424 656882 3476 656888
rect 3424 632120 3476 632126
rect 3422 632088 3424 632097
rect 3476 632088 3478 632097
rect 3422 632023 3478 632032
rect 3146 619168 3202 619177
rect 3146 619103 3202 619112
rect 3160 618322 3188 619103
rect 3148 618316 3200 618322
rect 3148 618258 3200 618264
rect 3238 606112 3294 606121
rect 3238 606047 3294 606056
rect 3252 605878 3280 606047
rect 3240 605872 3292 605878
rect 3240 605814 3292 605820
rect 3330 580000 3386 580009
rect 3330 579935 3386 579944
rect 3344 579698 3372 579935
rect 3332 579692 3384 579698
rect 3332 579634 3384 579640
rect 3422 566944 3478 566953
rect 3422 566879 3478 566888
rect 3436 565894 3464 566879
rect 3424 565888 3476 565894
rect 3424 565830 3476 565836
rect 3422 553888 3478 553897
rect 3422 553823 3478 553832
rect 3436 553450 3464 553823
rect 3424 553444 3476 553450
rect 3424 553386 3476 553392
rect 3422 527912 3478 527921
rect 3422 527847 3478 527856
rect 3436 527202 3464 527847
rect 3424 527196 3476 527202
rect 3424 527138 3476 527144
rect 3422 514856 3478 514865
rect 3422 514791 3424 514800
rect 3476 514791 3478 514800
rect 3424 514762 3476 514768
rect 3422 501800 3478 501809
rect 3422 501735 3478 501744
rect 3054 475688 3110 475697
rect 3054 475623 3110 475632
rect 3068 474774 3096 475623
rect 3056 474768 3108 474774
rect 3056 474710 3108 474716
rect 3146 449576 3202 449585
rect 3146 449511 3202 449520
rect 3160 448594 3188 449511
rect 3148 448588 3200 448594
rect 3148 448530 3200 448536
rect 2870 410544 2926 410553
rect 2870 410479 2926 410488
rect 2884 409902 2912 410479
rect 2872 409896 2924 409902
rect 2872 409838 2924 409844
rect 3146 358456 3202 358465
rect 3146 358391 3202 358400
rect 3160 357474 3188 358391
rect 3148 357468 3200 357474
rect 3148 357410 3200 357416
rect 3330 345400 3386 345409
rect 3330 345335 3386 345344
rect 3344 345098 3372 345335
rect 3332 345092 3384 345098
rect 3332 345034 3384 345040
rect 3330 319288 3386 319297
rect 3330 319223 3386 319232
rect 3344 318850 3372 319223
rect 3332 318844 3384 318850
rect 3332 318786 3384 318792
rect 3054 267200 3110 267209
rect 3054 267135 3110 267144
rect 3068 266422 3096 267135
rect 3056 266416 3108 266422
rect 3056 266358 3108 266364
rect 3054 241088 3110 241097
rect 3054 241023 3110 241032
rect 3068 240174 3096 241023
rect 3056 240168 3108 240174
rect 3056 240110 3108 240116
rect 3436 227050 3464 501735
rect 3514 462632 3570 462641
rect 3514 462567 3570 462576
rect 3528 462398 3556 462567
rect 3516 462392 3568 462398
rect 3516 462334 3568 462340
rect 3514 423600 3570 423609
rect 3514 423535 3570 423544
rect 3528 422346 3556 423535
rect 3516 422340 3568 422346
rect 3516 422282 3568 422288
rect 3516 397520 3568 397526
rect 3514 397488 3516 397497
rect 3568 397488 3570 397497
rect 3514 397423 3570 397432
rect 3514 371376 3570 371385
rect 3514 371311 3570 371320
rect 3528 371278 3556 371311
rect 3516 371272 3568 371278
rect 3516 371214 3568 371220
rect 3514 306232 3570 306241
rect 3514 306167 3570 306176
rect 3528 305046 3556 306167
rect 3516 305040 3568 305046
rect 3516 304982 3568 304988
rect 3514 293176 3570 293185
rect 3514 293111 3570 293120
rect 3528 292602 3556 293111
rect 3516 292596 3568 292602
rect 3516 292538 3568 292544
rect 3514 254144 3570 254153
rect 3514 254079 3570 254088
rect 3528 253978 3556 254079
rect 3516 253972 3568 253978
rect 3516 253914 3568 253920
rect 3424 227044 3476 227050
rect 3424 226986 3476 226992
rect 3146 214976 3202 214985
rect 3146 214911 3202 214920
rect 3160 213994 3188 214911
rect 3148 213988 3200 213994
rect 3148 213930 3200 213936
rect 8220 209234 8248 702406
rect 24320 700330 24348 703520
rect 40512 700466 40540 703520
rect 72988 702434 73016 703520
rect 89180 703474 89208 703520
rect 89364 703474 89392 703582
rect 89180 703446 89392 703474
rect 72988 702406 73108 702434
rect 40500 700460 40552 700466
rect 40500 700402 40552 700408
rect 41328 700460 41380 700466
rect 41328 700402 41380 700408
rect 24308 700324 24360 700330
rect 24308 700266 24360 700272
rect 39304 565888 39356 565894
rect 39304 565830 39356 565836
rect 39316 344350 39344 565830
rect 39304 344344 39356 344350
rect 39304 344286 39356 344292
rect 8208 209228 8260 209234
rect 8208 209170 8260 209176
rect 41340 207806 41368 700402
rect 41328 207800 41380 207806
rect 41328 207742 41380 207748
rect 73080 205193 73108 702406
rect 89640 224262 89668 703582
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 299492 703582 299980 703610
rect 105464 699718 105492 703520
rect 137848 700398 137876 703520
rect 137836 700392 137888 700398
rect 137836 700334 137888 700340
rect 137284 700324 137336 700330
rect 137284 700266 137336 700272
rect 105452 699712 105504 699718
rect 105452 699654 105504 699660
rect 106188 699712 106240 699718
rect 106188 699654 106240 699660
rect 89628 224256 89680 224262
rect 89628 224198 89680 224204
rect 73066 205184 73122 205193
rect 73066 205119 73122 205128
rect 106200 203697 106228 699654
rect 137296 210594 137324 700266
rect 154132 699786 154160 703520
rect 154120 699780 154172 699786
rect 154120 699722 154172 699728
rect 157984 699780 158036 699786
rect 157984 699722 158036 699728
rect 137284 210588 137336 210594
rect 137284 210530 137336 210536
rect 157996 207942 158024 699722
rect 170324 699718 170352 703520
rect 195244 700392 195296 700398
rect 195244 700334 195296 700340
rect 170312 699712 170364 699718
rect 170312 699654 170364 699660
rect 171048 699712 171100 699718
rect 171048 699654 171100 699660
rect 166264 448588 166316 448594
rect 166264 448530 166316 448536
rect 166276 228410 166304 448530
rect 166264 228404 166316 228410
rect 166264 228346 166316 228352
rect 157984 207936 158036 207942
rect 157984 207878 158036 207884
rect 171060 206378 171088 699654
rect 192484 605872 192536 605878
rect 192484 605814 192536 605820
rect 173164 553444 173216 553450
rect 173164 553386 173216 553392
rect 173176 215966 173204 553386
rect 191104 462392 191156 462398
rect 191104 462334 191156 462340
rect 177304 397520 177356 397526
rect 177304 397462 177356 397468
rect 177316 286346 177344 397462
rect 177304 286340 177356 286346
rect 177304 286282 177356 286288
rect 173164 215960 173216 215966
rect 173164 215902 173216 215908
rect 191116 210662 191144 462334
rect 191104 210656 191156 210662
rect 191104 210598 191156 210604
rect 192496 209370 192524 605814
rect 192484 209364 192536 209370
rect 192484 209306 192536 209312
rect 171048 206372 171100 206378
rect 171048 206314 171100 206320
rect 195256 205086 195284 700334
rect 199384 683188 199436 683194
rect 199384 683130 199436 683136
rect 198004 474768 198056 474774
rect 198004 474710 198056 474716
rect 196624 422340 196676 422346
rect 196624 422282 196676 422288
rect 196636 208010 196664 422282
rect 196624 208004 196676 208010
rect 196624 207946 196676 207952
rect 198016 206446 198044 474710
rect 199396 209438 199424 683130
rect 200764 305040 200816 305046
rect 200764 304982 200816 304988
rect 200776 210730 200804 304982
rect 200764 210724 200816 210730
rect 200764 210666 200816 210672
rect 199384 209432 199436 209438
rect 199384 209374 199436 209380
rect 198004 206440 198056 206446
rect 198004 206382 198056 206388
rect 202800 205222 202828 703520
rect 218992 700330 219020 703520
rect 218980 700324 219032 700330
rect 218980 700266 219032 700272
rect 235184 699718 235212 703520
rect 244924 700392 244976 700398
rect 244924 700334 244976 700340
rect 240784 700324 240836 700330
rect 240784 700266 240836 700272
rect 242164 700324 242216 700330
rect 242164 700266 242216 700272
rect 235172 699712 235224 699718
rect 235172 699654 235224 699660
rect 235908 699712 235960 699718
rect 235908 699654 235960 699660
rect 231124 618316 231176 618322
rect 231124 618258 231176 618264
rect 210424 527196 210476 527202
rect 210424 527138 210476 527144
rect 206284 514820 206336 514826
rect 206284 514762 206336 514768
rect 204904 240168 204956 240174
rect 204904 240110 204956 240116
rect 204916 209302 204944 240110
rect 206296 210798 206324 514762
rect 209044 318844 209096 318850
rect 209044 318786 209096 318792
rect 206284 210792 206336 210798
rect 206284 210734 206336 210740
rect 204904 209296 204956 209302
rect 204904 209238 204956 209244
rect 209056 206514 209084 318786
rect 209044 206508 209096 206514
rect 209044 206450 209096 206456
rect 202788 205216 202840 205222
rect 202788 205158 202840 205164
rect 195244 205080 195296 205086
rect 195244 205022 195296 205028
rect 209044 204400 209096 204406
rect 209044 204342 209096 204348
rect 202052 204332 202104 204338
rect 202052 204274 202104 204280
rect 106186 203688 106242 203697
rect 106186 203623 106242 203632
rect 159364 203176 159416 203182
rect 159364 203118 159416 203124
rect 3238 201920 3294 201929
rect 3238 201855 3294 201864
rect 140044 201884 140096 201890
rect 3252 201686 3280 201855
rect 140044 201826 140096 201832
rect 98644 201816 98696 201822
rect 98644 201758 98696 201764
rect 14464 201748 14516 201754
rect 14464 201690 14516 201696
rect 3240 201680 3292 201686
rect 3240 201622 3292 201628
rect 3424 200864 3476 200870
rect 3424 200806 3476 200812
rect 3240 164212 3292 164218
rect 3240 164154 3292 164160
rect 3252 162897 3280 164154
rect 3238 162888 3294 162897
rect 3238 162823 3294 162832
rect 3436 149841 3464 200806
rect 3516 189032 3568 189038
rect 3516 188974 3568 188980
rect 3528 188873 3556 188974
rect 3514 188864 3570 188873
rect 3514 188799 3570 188808
rect 3422 149832 3478 149841
rect 3422 149767 3478 149776
rect 3240 137964 3292 137970
rect 3240 137906 3292 137912
rect 3252 136785 3280 137906
rect 3238 136776 3294 136785
rect 3238 136711 3294 136720
rect 3424 111784 3476 111790
rect 3424 111726 3476 111732
rect 3436 110673 3464 111726
rect 3422 110664 3478 110673
rect 3422 110599 3478 110608
rect 4804 98660 4856 98666
rect 4804 98602 4856 98608
rect 3424 97980 3476 97986
rect 3424 97922 3476 97928
rect 3436 97617 3464 97922
rect 3422 97608 3478 97617
rect 3422 97543 3478 97552
rect 4068 95940 4120 95946
rect 4068 95882 4120 95888
rect 1308 91792 1360 91798
rect 1308 91734 1360 91740
rect 1320 3534 1348 91734
rect 3148 85536 3200 85542
rect 3148 85478 3200 85484
rect 3160 84697 3188 85478
rect 3146 84688 3202 84697
rect 3146 84623 3202 84632
rect 3424 71732 3476 71738
rect 3424 71674 3476 71680
rect 3436 71641 3464 71674
rect 3422 71632 3478 71641
rect 3422 71567 3478 71576
rect 3056 59356 3108 59362
rect 3056 59298 3108 59304
rect 3068 58585 3096 59298
rect 3054 58576 3110 58585
rect 3054 58511 3110 58520
rect 3424 45552 3476 45558
rect 3422 45520 3424 45529
rect 3476 45520 3478 45529
rect 3422 45455 3478 45464
rect 2872 33108 2924 33114
rect 2872 33050 2924 33056
rect 2884 32473 2912 33050
rect 2870 32464 2926 32473
rect 2870 32399 2926 32408
rect 3424 20664 3476 20670
rect 3424 20606 3476 20612
rect 3436 19417 3464 20606
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 4080 6914 4108 95882
rect 3988 6886 4108 6914
rect 3424 6860 3476 6866
rect 3424 6802 3476 6808
rect 3436 6497 3464 6802
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 1676 3596 1728 3602
rect 1676 3538 1728 3544
rect 572 3528 624 3534
rect 572 3470 624 3476
rect 1308 3528 1360 3534
rect 1308 3470 1360 3476
rect 584 480 612 3470
rect 1688 480 1716 3538
rect 3988 3534 4016 6886
rect 4816 3602 4844 98602
rect 12348 91860 12400 91866
rect 12348 91802 12400 91808
rect 10968 86284 11020 86290
rect 10968 86226 11020 86232
rect 6828 68332 6880 68338
rect 6828 68274 6880 68280
rect 5264 7608 5316 7614
rect 5264 7550 5316 7556
rect 4804 3596 4856 3602
rect 4804 3538 4856 3544
rect 2872 3528 2924 3534
rect 2872 3470 2924 3476
rect 3976 3528 4028 3534
rect 3976 3470 4028 3476
rect 2884 480 2912 3470
rect 4068 3460 4120 3466
rect 4068 3402 4120 3408
rect 4080 480 4108 3402
rect 5276 480 5304 7550
rect 6840 6914 6868 68274
rect 6472 6886 6868 6914
rect 6472 480 6500 6886
rect 8760 3732 8812 3738
rect 8760 3674 8812 3680
rect 7656 2100 7708 2106
rect 7656 2042 7708 2048
rect 7668 480 7696 2042
rect 8772 480 8800 3674
rect 10980 3534 11008 86226
rect 12256 24132 12308 24138
rect 12256 24074 12308 24080
rect 12268 3534 12296 24074
rect 9956 3528 10008 3534
rect 9956 3470 10008 3476
rect 10968 3528 11020 3534
rect 10968 3470 11020 3476
rect 11152 3528 11204 3534
rect 11152 3470 11204 3476
rect 12256 3528 12308 3534
rect 12256 3470 12308 3476
rect 9968 480 9996 3470
rect 11164 480 11192 3470
rect 12360 480 12388 91802
rect 14476 85542 14504 201690
rect 36544 200252 36596 200258
rect 36544 200194 36596 200200
rect 35164 198144 35216 198150
rect 35164 198086 35216 198092
rect 15842 101008 15898 101017
rect 15842 100943 15898 100952
rect 14464 85536 14516 85542
rect 14464 85478 14516 85484
rect 15108 84856 15160 84862
rect 15108 84798 15160 84804
rect 15120 6914 15148 84798
rect 14752 6886 15148 6914
rect 13544 3528 13596 3534
rect 13544 3470 13596 3476
rect 13556 480 13584 3470
rect 14752 480 14780 6886
rect 15856 3466 15884 100943
rect 30286 98696 30342 98705
rect 30286 98631 30342 98640
rect 18602 95840 18658 95849
rect 18602 95775 18658 95784
rect 17868 76560 17920 76566
rect 17868 76502 17920 76508
rect 15934 3496 15990 3505
rect 15844 3460 15896 3466
rect 17880 3466 17908 76502
rect 18616 3738 18644 95775
rect 22008 93152 22060 93158
rect 22008 93094 22060 93100
rect 26146 93120 26202 93129
rect 20628 68400 20680 68406
rect 20628 68342 20680 68348
rect 18604 3732 18656 3738
rect 18604 3674 18656 3680
rect 18236 3664 18288 3670
rect 18236 3606 18288 3612
rect 15934 3431 15990 3440
rect 17040 3460 17092 3466
rect 15844 3402 15896 3408
rect 15948 480 15976 3431
rect 17040 3402 17092 3408
rect 17868 3460 17920 3466
rect 17868 3402 17920 3408
rect 17052 480 17080 3402
rect 18248 480 18276 3606
rect 20640 3466 20668 68342
rect 22020 6914 22048 93094
rect 26146 93055 26202 93064
rect 23388 91928 23440 91934
rect 23388 91870 23440 91876
rect 23400 6914 23428 91870
rect 21836 6886 22048 6914
rect 23032 6886 23428 6914
rect 19432 3460 19484 3466
rect 19432 3402 19484 3408
rect 20628 3460 20680 3466
rect 20628 3402 20680 3408
rect 19444 480 19472 3402
rect 20628 3324 20680 3330
rect 20628 3266 20680 3272
rect 20640 480 20668 3266
rect 21836 480 21864 6886
rect 23032 480 23060 6886
rect 24216 3596 24268 3602
rect 24216 3538 24268 3544
rect 24228 480 24256 3538
rect 26160 3466 26188 93055
rect 28262 91760 28318 91769
rect 28262 91695 28318 91704
rect 27526 87544 27582 87553
rect 27526 87479 27582 87488
rect 27540 3466 27568 87479
rect 28276 3670 28304 91695
rect 30300 6914 30328 98631
rect 32404 97300 32456 97306
rect 32404 97242 32456 97248
rect 31668 73840 31720 73846
rect 31668 73782 31720 73788
rect 31680 6914 31708 73782
rect 30116 6886 30328 6914
rect 31312 6886 31708 6914
rect 28908 4208 28960 4214
rect 28908 4150 28960 4156
rect 28264 3664 28316 3670
rect 28264 3606 28316 3612
rect 25320 3460 25372 3466
rect 25320 3402 25372 3408
rect 26148 3460 26200 3466
rect 26148 3402 26200 3408
rect 26516 3460 26568 3466
rect 26516 3402 26568 3408
rect 27528 3460 27580 3466
rect 27528 3402 27580 3408
rect 25332 480 25360 3402
rect 26528 480 26556 3402
rect 27712 3052 27764 3058
rect 27712 2994 27764 3000
rect 27724 480 27752 2994
rect 28920 480 28948 4150
rect 30116 480 30144 6886
rect 31312 480 31340 6886
rect 32416 4214 32444 97242
rect 34426 93256 34482 93265
rect 34426 93191 34482 93200
rect 33048 18624 33100 18630
rect 33048 18566 33100 18572
rect 32404 4208 32456 4214
rect 32404 4150 32456 4156
rect 33060 3466 33088 18566
rect 34440 3466 34468 93191
rect 35176 71738 35204 198086
rect 36556 97986 36584 200194
rect 47584 198824 47636 198830
rect 47584 198766 47636 198772
rect 39304 100768 39356 100774
rect 39304 100710 39356 100716
rect 36544 97980 36596 97986
rect 36544 97922 36596 97928
rect 37188 93220 37240 93226
rect 37188 93162 37240 93168
rect 35254 82104 35310 82113
rect 35254 82039 35310 82048
rect 35164 71732 35216 71738
rect 35164 71674 35216 71680
rect 32404 3460 32456 3466
rect 32404 3402 32456 3408
rect 33048 3460 33100 3466
rect 33048 3402 33100 3408
rect 33600 3460 33652 3466
rect 33600 3402 33652 3408
rect 34428 3460 34480 3466
rect 34428 3402 34480 3408
rect 32416 480 32444 3402
rect 33612 480 33640 3402
rect 34796 3324 34848 3330
rect 34796 3266 34848 3272
rect 34808 480 34836 3266
rect 35268 3058 35296 82039
rect 35806 73808 35862 73817
rect 35806 73743 35862 73752
rect 35820 3330 35848 73743
rect 37096 11756 37148 11762
rect 37096 11698 37148 11704
rect 35900 3732 35952 3738
rect 35900 3674 35952 3680
rect 35912 3534 35940 3674
rect 37108 3534 37136 11698
rect 35900 3528 35952 3534
rect 35900 3470 35952 3476
rect 35992 3528 36044 3534
rect 35992 3470 36044 3476
rect 37096 3528 37148 3534
rect 37096 3470 37148 3476
rect 35808 3324 35860 3330
rect 35808 3266 35860 3272
rect 35256 3052 35308 3058
rect 35256 2994 35308 3000
rect 36004 480 36032 3470
rect 37200 480 37228 93162
rect 38568 71052 38620 71058
rect 38568 70994 38620 71000
rect 38580 6914 38608 70994
rect 38396 6886 38608 6914
rect 38396 480 38424 6886
rect 39316 3738 39344 100710
rect 40684 97368 40736 97374
rect 40684 97310 40736 97316
rect 39304 3732 39356 3738
rect 39304 3674 39356 3680
rect 40696 3194 40724 97310
rect 46202 97200 46258 97209
rect 46202 97135 46258 97144
rect 43444 94512 43496 94518
rect 43444 94454 43496 94460
rect 42708 77988 42760 77994
rect 42708 77930 42760 77936
rect 40776 4004 40828 4010
rect 40776 3946 40828 3952
rect 39580 3188 39632 3194
rect 39580 3130 39632 3136
rect 40684 3188 40736 3194
rect 40684 3130 40736 3136
rect 39592 480 39620 3130
rect 40788 1986 40816 3946
rect 42720 3534 42748 77930
rect 43456 3670 43484 94454
rect 45468 87644 45520 87650
rect 45468 87586 45520 87592
rect 45376 71120 45428 71126
rect 45376 71062 45428 71068
rect 44088 51740 44140 51746
rect 44088 51682 44140 51688
rect 43444 3664 43496 3670
rect 43444 3606 43496 3612
rect 44100 3534 44128 51682
rect 45388 16574 45416 71062
rect 45296 16546 45416 16574
rect 44272 3596 44324 3602
rect 44272 3538 44324 3544
rect 41880 3528 41932 3534
rect 41880 3470 41932 3476
rect 42708 3528 42760 3534
rect 42708 3470 42760 3476
rect 43076 3528 43128 3534
rect 43076 3470 43128 3476
rect 44088 3528 44140 3534
rect 44088 3470 44140 3476
rect 40696 1958 40816 1986
rect 40696 480 40724 1958
rect 41892 480 41920 3470
rect 43088 480 43116 3470
rect 44284 480 44312 3538
rect 45296 3482 45324 16546
rect 45480 6914 45508 87586
rect 46216 7614 46244 97135
rect 47596 33114 47624 198766
rect 77208 99476 77260 99482
rect 77208 99418 77260 99424
rect 66168 99408 66220 99414
rect 66168 99350 66220 99356
rect 62028 90500 62080 90506
rect 62028 90442 62080 90448
rect 55128 90432 55180 90438
rect 55128 90374 55180 90380
rect 53748 87712 53800 87718
rect 53748 87654 53800 87660
rect 50988 84924 51040 84930
rect 50988 84866 51040 84872
rect 47676 82136 47728 82142
rect 47676 82078 47728 82084
rect 47584 33108 47636 33114
rect 47584 33050 47636 33056
rect 46848 25560 46900 25566
rect 46848 25502 46900 25508
rect 46204 7608 46256 7614
rect 46204 7550 46256 7556
rect 46860 6914 46888 25502
rect 45388 6886 45508 6914
rect 46676 6886 46888 6914
rect 45388 3602 45416 6886
rect 45376 3596 45428 3602
rect 45376 3538 45428 3544
rect 45296 3454 45508 3482
rect 45480 480 45508 3454
rect 46676 480 46704 6886
rect 47688 4010 47716 82078
rect 49606 80744 49662 80753
rect 49606 80679 49662 80688
rect 48228 73908 48280 73914
rect 48228 73850 48280 73856
rect 48240 6914 48268 73850
rect 47872 6886 48268 6914
rect 47676 4004 47728 4010
rect 47676 3946 47728 3952
rect 47872 480 47900 6886
rect 49620 3534 49648 80679
rect 51000 3534 51028 84866
rect 53656 71188 53708 71194
rect 53656 71130 53708 71136
rect 53668 16574 53696 71130
rect 53576 16546 53696 16574
rect 52552 3596 52604 3602
rect 52552 3538 52604 3544
rect 48964 3528 49016 3534
rect 48964 3470 49016 3476
rect 49608 3528 49660 3534
rect 49608 3470 49660 3476
rect 50160 3528 50212 3534
rect 50160 3470 50212 3476
rect 50988 3528 51040 3534
rect 50988 3470 51040 3476
rect 51356 3528 51408 3534
rect 51356 3470 51408 3476
rect 48976 480 49004 3470
rect 50172 480 50200 3470
rect 51368 480 51396 3470
rect 52564 480 52592 3538
rect 53576 3482 53604 16546
rect 53760 6914 53788 87654
rect 55140 6914 55168 90374
rect 59268 90364 59320 90370
rect 59268 90306 59320 90312
rect 57886 84824 57942 84833
rect 57886 84759 57942 84768
rect 53668 6886 53788 6914
rect 54956 6886 55168 6914
rect 53668 3602 53696 6886
rect 53656 3596 53708 3602
rect 53656 3538 53708 3544
rect 53576 3454 53788 3482
rect 53760 480 53788 3454
rect 54956 480 54984 6886
rect 56048 3664 56100 3670
rect 56048 3606 56100 3612
rect 56060 480 56088 3606
rect 57900 3602 57928 84759
rect 59280 3602 59308 90306
rect 61936 71256 61988 71262
rect 61936 71198 61988 71204
rect 59636 4888 59688 4894
rect 59636 4830 59688 4836
rect 57244 3596 57296 3602
rect 57244 3538 57296 3544
rect 57888 3596 57940 3602
rect 57888 3538 57940 3544
rect 58440 3596 58492 3602
rect 58440 3538 58492 3544
rect 59268 3596 59320 3602
rect 59268 3538 59320 3544
rect 57256 480 57284 3538
rect 58452 480 58480 3538
rect 59648 480 59676 4830
rect 61948 3602 61976 71198
rect 60832 3596 60884 3602
rect 60832 3538 60884 3544
rect 61936 3596 61988 3602
rect 61936 3538 61988 3544
rect 60844 480 60872 3538
rect 62040 480 62068 90442
rect 64788 71324 64840 71330
rect 64788 71266 64840 71272
rect 64800 3330 64828 71266
rect 66180 3602 66208 99350
rect 71044 91996 71096 92002
rect 71044 91938 71096 91944
rect 70308 87780 70360 87786
rect 70308 87722 70360 87728
rect 68928 84992 68980 84998
rect 68928 84934 68980 84940
rect 66720 3732 66772 3738
rect 66720 3674 66772 3680
rect 65524 3596 65576 3602
rect 65524 3538 65576 3544
rect 66168 3596 66220 3602
rect 66168 3538 66220 3544
rect 64328 3324 64380 3330
rect 64328 3266 64380 3272
rect 64788 3324 64840 3330
rect 64788 3266 64840 3272
rect 63224 2168 63276 2174
rect 63224 2110 63276 2116
rect 63236 480 63264 2110
rect 64340 480 64368 3266
rect 65536 480 65564 3538
rect 66732 480 66760 3674
rect 68940 3602 68968 84934
rect 67916 3596 67968 3602
rect 67916 3538 67968 3544
rect 68928 3596 68980 3602
rect 68928 3538 68980 3544
rect 67928 480 67956 3538
rect 69112 3052 69164 3058
rect 69112 2994 69164 3000
rect 69124 480 69152 2994
rect 70320 480 70348 87722
rect 71056 3058 71084 91938
rect 73068 90568 73120 90574
rect 73068 90510 73120 90516
rect 71688 47592 71740 47598
rect 71688 47534 71740 47540
rect 71700 6914 71728 47534
rect 71516 6886 71728 6914
rect 71044 3052 71096 3058
rect 71044 2994 71096 3000
rect 71516 480 71544 6886
rect 73080 3602 73108 90510
rect 75182 87680 75238 87689
rect 75182 87615 75238 87624
rect 74908 3732 74960 3738
rect 74908 3674 74960 3680
rect 72608 3596 72660 3602
rect 72608 3538 72660 3544
rect 73068 3596 73120 3602
rect 73068 3538 73120 3544
rect 72620 480 72648 3538
rect 74920 3534 74948 3674
rect 74908 3528 74960 3534
rect 74908 3470 74960 3476
rect 75000 3528 75052 3534
rect 75000 3470 75052 3476
rect 73804 3188 73856 3194
rect 73804 3130 73856 3136
rect 73816 480 73844 3130
rect 75012 480 75040 3470
rect 75196 3194 75224 87615
rect 75828 79348 75880 79354
rect 75828 79290 75880 79296
rect 75840 3534 75868 79290
rect 77220 3534 77248 99418
rect 80702 98832 80758 98841
rect 80702 98767 80758 98776
rect 79966 89040 80022 89049
rect 79966 88975 80022 88984
rect 78588 43444 78640 43450
rect 78588 43386 78640 43392
rect 77392 3800 77444 3806
rect 77392 3742 77444 3748
rect 75828 3528 75880 3534
rect 75828 3470 75880 3476
rect 76196 3528 76248 3534
rect 76196 3470 76248 3476
rect 77208 3528 77260 3534
rect 77208 3470 77260 3476
rect 75184 3188 75236 3194
rect 75184 3130 75236 3136
rect 76208 480 76236 3470
rect 77404 480 77432 3742
rect 78600 480 78628 43386
rect 79980 6914 80008 88975
rect 79704 6886 80008 6914
rect 79704 480 79732 6886
rect 80716 3738 80744 98767
rect 93124 97504 93176 97510
rect 93124 97446 93176 97452
rect 86316 97436 86368 97442
rect 86316 97378 86368 97384
rect 83462 84960 83518 84969
rect 83462 84895 83518 84904
rect 80888 4820 80940 4826
rect 80888 4762 80940 4768
rect 80704 3732 80756 3738
rect 80704 3674 80756 3680
rect 80900 480 80928 4762
rect 83280 3528 83332 3534
rect 83280 3470 83332 3476
rect 82084 2916 82136 2922
rect 82084 2858 82136 2864
rect 82096 480 82124 2858
rect 83292 480 83320 3470
rect 83476 2922 83504 84895
rect 86224 79416 86276 79422
rect 86224 79358 86276 79364
rect 85488 73976 85540 73982
rect 85488 73918 85540 73924
rect 85500 3602 85528 73918
rect 86236 3738 86264 79358
rect 86328 25566 86356 97378
rect 91008 89004 91060 89010
rect 91008 88946 91060 88952
rect 88984 87848 89036 87854
rect 88984 87790 89036 87796
rect 88248 86352 88300 86358
rect 88248 86294 88300 86300
rect 86316 25560 86368 25566
rect 86316 25502 86368 25508
rect 86868 15904 86920 15910
rect 86868 15846 86920 15852
rect 86224 3732 86276 3738
rect 86224 3674 86276 3680
rect 86776 3732 86828 3738
rect 86776 3674 86828 3680
rect 84476 3596 84528 3602
rect 84476 3538 84528 3544
rect 85488 3596 85540 3602
rect 85488 3538 85540 3544
rect 83464 2916 83516 2922
rect 83464 2858 83516 2864
rect 84488 480 84516 3538
rect 85672 3052 85724 3058
rect 85672 2994 85724 3000
rect 85684 480 85712 2994
rect 86788 1850 86816 3674
rect 86880 3058 86908 15846
rect 88260 6914 88288 86294
rect 87984 6886 88288 6914
rect 86868 3052 86920 3058
rect 86868 2994 86920 3000
rect 86788 1822 86908 1850
rect 86880 480 86908 1822
rect 87984 480 88012 6886
rect 88996 3806 89024 87790
rect 89628 83496 89680 83502
rect 89628 83438 89680 83444
rect 88984 3800 89036 3806
rect 88984 3742 89036 3748
rect 89640 3602 89668 83438
rect 91020 3602 91048 88946
rect 92386 73944 92442 73953
rect 92386 73879 92442 73888
rect 92400 3602 92428 73879
rect 93136 4894 93164 97446
rect 97906 89176 97962 89185
rect 97906 89111 97962 89120
rect 95148 87916 95200 87922
rect 95148 87858 95200 87864
rect 94504 13116 94556 13122
rect 94504 13058 94556 13064
rect 93124 4888 93176 4894
rect 93124 4830 93176 4836
rect 89168 3596 89220 3602
rect 89168 3538 89220 3544
rect 89628 3596 89680 3602
rect 89628 3538 89680 3544
rect 90364 3596 90416 3602
rect 90364 3538 90416 3544
rect 91008 3596 91060 3602
rect 91008 3538 91060 3544
rect 91560 3596 91612 3602
rect 91560 3538 91612 3544
rect 92388 3596 92440 3602
rect 92388 3538 92440 3544
rect 89180 480 89208 3538
rect 90376 480 90404 3538
rect 91572 480 91600 3538
rect 94516 3398 94544 13058
rect 92756 3392 92808 3398
rect 92756 3334 92808 3340
rect 94504 3392 94556 3398
rect 94504 3334 94556 3340
rect 92768 480 92796 3334
rect 93952 3256 94004 3262
rect 93952 3198 94004 3204
rect 93964 480 93992 3198
rect 95160 480 95188 87858
rect 96528 83564 96580 83570
rect 96528 83506 96580 83512
rect 96540 6914 96568 83506
rect 96264 6886 96568 6914
rect 96264 480 96292 6886
rect 97920 3602 97948 89111
rect 98656 20670 98684 201758
rect 133144 200320 133196 200326
rect 133144 200262 133196 200268
rect 106924 198960 106976 198966
rect 106924 198902 106976 198908
rect 105544 99544 105596 99550
rect 105544 99486 105596 99492
rect 101404 97572 101456 97578
rect 101404 97514 101456 97520
rect 98736 80708 98788 80714
rect 98736 80650 98788 80656
rect 98644 20664 98696 20670
rect 98644 20606 98696 20612
rect 97448 3596 97500 3602
rect 97448 3538 97500 3544
rect 97908 3596 97960 3602
rect 97908 3538 97960 3544
rect 98644 3596 98696 3602
rect 98644 3538 98696 3544
rect 97460 480 97488 3538
rect 98656 480 98684 3538
rect 98748 3262 98776 80650
rect 99288 74044 99340 74050
rect 99288 73986 99340 73992
rect 99300 3602 99328 73986
rect 100668 17264 100720 17270
rect 100668 17206 100720 17212
rect 100680 3602 100708 17206
rect 101416 11762 101444 97514
rect 104164 90636 104216 90642
rect 104164 90578 104216 90584
rect 103428 83632 103480 83638
rect 103428 83574 103480 83580
rect 101494 79384 101550 79393
rect 101494 79319 101550 79328
rect 101404 11756 101456 11762
rect 101404 11698 101456 11704
rect 101036 4004 101088 4010
rect 101036 3946 101088 3952
rect 99288 3596 99340 3602
rect 99288 3538 99340 3544
rect 99840 3596 99892 3602
rect 99840 3538 99892 3544
rect 100668 3596 100720 3602
rect 100668 3538 100720 3544
rect 98736 3256 98788 3262
rect 98736 3198 98788 3204
rect 99852 480 99880 3538
rect 101048 480 101076 3946
rect 101508 3670 101536 79319
rect 103440 6914 103468 83574
rect 103348 6886 103468 6914
rect 101496 3664 101548 3670
rect 101496 3606 101548 3612
rect 102232 3596 102284 3602
rect 102232 3538 102284 3544
rect 102244 480 102272 3538
rect 103348 480 103376 6886
rect 104176 4010 104204 90578
rect 104164 4004 104216 4010
rect 104164 3946 104216 3952
rect 103520 3800 103572 3806
rect 103520 3742 103572 3748
rect 103532 3602 103560 3742
rect 103520 3596 103572 3602
rect 103520 3538 103572 3544
rect 105556 3534 105584 99486
rect 106188 82204 106240 82210
rect 106188 82146 106240 82152
rect 106200 3534 106228 82146
rect 106936 45558 106964 198902
rect 130382 95976 130438 95985
rect 130382 95911 130438 95920
rect 126888 94580 126940 94586
rect 126888 94522 126940 94528
rect 125506 93392 125562 93401
rect 125506 93327 125562 93336
rect 122104 89276 122156 89282
rect 122104 89218 122156 89224
rect 115204 89208 115256 89214
rect 115204 89150 115256 89156
rect 112444 89140 112496 89146
rect 112444 89082 112496 89088
rect 108948 89072 109000 89078
rect 108948 89014 109000 89020
rect 107016 86420 107068 86426
rect 107016 86362 107068 86368
rect 106924 45552 106976 45558
rect 106924 45494 106976 45500
rect 107028 3806 107056 86362
rect 107566 44840 107622 44849
rect 107566 44775 107622 44784
rect 107016 3800 107068 3806
rect 107016 3742 107068 3748
rect 104532 3528 104584 3534
rect 104532 3470 104584 3476
rect 105544 3528 105596 3534
rect 105544 3470 105596 3476
rect 105728 3528 105780 3534
rect 105728 3470 105780 3476
rect 106188 3528 106240 3534
rect 106188 3470 106240 3476
rect 104544 480 104572 3470
rect 105740 480 105768 3470
rect 107580 3330 107608 44775
rect 108960 3534 108988 89014
rect 111064 86488 111116 86494
rect 111064 86430 111116 86436
rect 110512 3596 110564 3602
rect 110512 3538 110564 3544
rect 108120 3528 108172 3534
rect 108120 3470 108172 3476
rect 108948 3528 109000 3534
rect 108948 3470 109000 3476
rect 109316 3528 109368 3534
rect 109316 3470 109368 3476
rect 106924 3324 106976 3330
rect 106924 3266 106976 3272
rect 107568 3324 107620 3330
rect 107568 3266 107620 3272
rect 106936 480 106964 3266
rect 108132 480 108160 3470
rect 109328 480 109356 3470
rect 110524 480 110552 3538
rect 111076 3534 111104 86430
rect 111708 83700 111760 83706
rect 111708 83642 111760 83648
rect 111720 3602 111748 83642
rect 111708 3596 111760 3602
rect 111708 3538 111760 3544
rect 112456 3534 112484 89082
rect 113088 79484 113140 79490
rect 113088 79426 113140 79432
rect 113100 6914 113128 79426
rect 114466 77888 114522 77897
rect 114466 77823 114522 77832
rect 112824 6886 113128 6914
rect 111064 3528 111116 3534
rect 111064 3470 111116 3476
rect 111616 3528 111668 3534
rect 111616 3470 111668 3476
rect 112444 3528 112496 3534
rect 112444 3470 112496 3476
rect 111628 480 111656 3470
rect 112824 480 112852 6886
rect 114480 3534 114508 77823
rect 115216 6914 115244 89150
rect 119988 86624 120040 86630
rect 119988 86566 120040 86572
rect 117228 86556 117280 86562
rect 117228 86498 117280 86504
rect 115848 80776 115900 80782
rect 115848 80718 115900 80724
rect 115124 6886 115244 6914
rect 115124 3738 115152 6886
rect 115112 3732 115164 3738
rect 115112 3674 115164 3680
rect 115860 3534 115888 80718
rect 117240 3534 117268 86498
rect 119344 85060 119396 85066
rect 119344 85002 119396 85008
rect 119356 3602 119384 85002
rect 119896 79552 119948 79558
rect 119896 79494 119948 79500
rect 119908 16574 119936 79494
rect 119816 16546 119936 16574
rect 117596 3596 117648 3602
rect 117596 3538 117648 3544
rect 119344 3596 119396 3602
rect 119344 3538 119396 3544
rect 114008 3528 114060 3534
rect 114008 3470 114060 3476
rect 114468 3528 114520 3534
rect 114468 3470 114520 3476
rect 115204 3528 115256 3534
rect 115204 3470 115256 3476
rect 115848 3528 115900 3534
rect 115848 3470 115900 3476
rect 116400 3528 116452 3534
rect 116400 3470 116452 3476
rect 117228 3528 117280 3534
rect 117228 3470 117280 3476
rect 114020 480 114048 3470
rect 115216 480 115244 3470
rect 116412 480 116440 3470
rect 117608 480 117636 3538
rect 119816 3534 119844 16546
rect 120000 6914 120028 86566
rect 121368 71392 121420 71398
rect 121368 71334 121420 71340
rect 121380 6914 121408 71334
rect 119908 6886 120028 6914
rect 121104 6886 121408 6914
rect 118792 3528 118844 3534
rect 118792 3470 118844 3476
rect 119804 3528 119856 3534
rect 119804 3470 119856 3476
rect 118804 480 118832 3470
rect 119908 480 119936 6886
rect 121104 480 121132 6886
rect 122116 3670 122144 89218
rect 124128 86692 124180 86698
rect 124128 86634 124180 86640
rect 122746 79520 122802 79529
rect 122746 79455 122802 79464
rect 122104 3664 122156 3670
rect 122104 3606 122156 3612
rect 122760 3534 122788 79455
rect 124140 3534 124168 86634
rect 125416 68468 125468 68474
rect 125416 68410 125468 68416
rect 125428 3534 125456 68410
rect 125520 3670 125548 93327
rect 126796 76628 126848 76634
rect 126796 76570 126848 76576
rect 125508 3664 125560 3670
rect 125508 3606 125560 3612
rect 126808 3534 126836 76570
rect 122288 3528 122340 3534
rect 122288 3470 122340 3476
rect 122748 3528 122800 3534
rect 122748 3470 122800 3476
rect 123484 3528 123536 3534
rect 123484 3470 123536 3476
rect 124128 3528 124180 3534
rect 124128 3470 124180 3476
rect 124680 3528 124732 3534
rect 124680 3470 124732 3476
rect 125416 3528 125468 3534
rect 125416 3470 125468 3476
rect 125876 3528 125928 3534
rect 125876 3470 125928 3476
rect 126796 3528 126848 3534
rect 126796 3470 126848 3476
rect 126900 3482 126928 94522
rect 128176 3596 128228 3602
rect 128176 3538 128228 3544
rect 122300 480 122328 3470
rect 123496 480 123524 3470
rect 124692 480 124720 3470
rect 125888 480 125916 3470
rect 126900 3454 127020 3482
rect 126992 480 127020 3454
rect 128188 480 128216 3538
rect 130396 3534 130424 95911
rect 133156 6866 133184 200262
rect 135168 99748 135220 99754
rect 135168 99690 135220 99696
rect 133234 83464 133290 83473
rect 133234 83399 133290 83408
rect 133144 6860 133196 6866
rect 133144 6802 133196 6808
rect 133248 4146 133276 83399
rect 130568 4140 130620 4146
rect 130568 4082 130620 4088
rect 133236 4140 133288 4146
rect 133236 4082 133288 4088
rect 129372 3528 129424 3534
rect 129372 3470 129424 3476
rect 130384 3528 130436 3534
rect 130384 3470 130436 3476
rect 129384 480 129412 3470
rect 130580 480 130608 4082
rect 131764 3868 131816 3874
rect 131764 3810 131816 3816
rect 131776 480 131804 3810
rect 132960 3800 133012 3806
rect 132960 3742 133012 3748
rect 132972 480 133000 3742
rect 135180 3602 135208 99690
rect 137284 92064 137336 92070
rect 137284 92006 137336 92012
rect 136548 82272 136600 82278
rect 136548 82214 136600 82220
rect 136456 76696 136508 76702
rect 136456 76638 136508 76644
rect 134156 3596 134208 3602
rect 134156 3538 134208 3544
rect 135168 3596 135220 3602
rect 135168 3538 135220 3544
rect 134168 480 134196 3538
rect 135260 3324 135312 3330
rect 135260 3266 135312 3272
rect 135272 480 135300 3266
rect 136468 480 136496 76638
rect 136560 3330 136588 82214
rect 137296 3874 137324 92006
rect 139308 76764 139360 76770
rect 139308 76706 139360 76712
rect 137284 3868 137336 3874
rect 137284 3810 137336 3816
rect 137652 3732 137704 3738
rect 137652 3674 137704 3680
rect 136548 3324 136600 3330
rect 136548 3266 136600 3272
rect 137664 480 137692 3674
rect 139320 3602 139348 76706
rect 140056 59362 140084 201826
rect 157248 200388 157300 200394
rect 157248 200330 157300 200336
rect 148324 199028 148376 199034
rect 148324 198970 148376 198976
rect 148336 111790 148364 198970
rect 151728 194608 151780 194614
rect 151728 194550 151780 194556
rect 151740 122806 151768 194550
rect 153108 191888 153160 191894
rect 153108 191830 153160 191836
rect 153120 122874 153148 191830
rect 155868 190528 155920 190534
rect 155868 190470 155920 190476
rect 155880 124166 155908 190470
rect 155868 124160 155920 124166
rect 155868 124102 155920 124108
rect 153108 122868 153160 122874
rect 153108 122810 153160 122816
rect 151728 122800 151780 122806
rect 151728 122742 151780 122748
rect 157260 122738 157288 200330
rect 157984 199096 158036 199102
rect 157984 199038 158036 199044
rect 157996 137970 158024 199038
rect 159376 164218 159404 203118
rect 201224 202904 201276 202910
rect 201224 202846 201276 202852
rect 200394 200152 200450 200161
rect 200394 200087 200450 200096
rect 200408 199988 200436 200087
rect 201236 199988 201264 202846
rect 202064 199988 202092 204274
rect 207296 203108 207348 203114
rect 207296 203050 207348 203056
rect 205548 203040 205600 203046
rect 205548 202982 205600 202988
rect 202972 202972 203024 202978
rect 202972 202914 203024 202920
rect 202984 199988 203012 202914
rect 204720 200184 204772 200190
rect 204720 200126 204772 200132
rect 204732 199988 204760 200126
rect 205560 199988 205588 202982
rect 207308 199988 207336 203050
rect 208216 201952 208268 201958
rect 208216 201894 208268 201900
rect 208228 199988 208256 201894
rect 209056 199988 209084 204342
rect 210436 203590 210464 527138
rect 224868 430636 224920 430642
rect 224868 430578 224920 430584
rect 213184 371272 213236 371278
rect 213184 371214 213236 371220
rect 213196 208078 213224 371214
rect 220728 311908 220780 311914
rect 220728 311850 220780 311856
rect 217968 258120 218020 258126
rect 217968 258062 218020 258068
rect 215944 231872 215996 231878
rect 215944 231814 215996 231820
rect 215208 218068 215260 218074
rect 215208 218010 215260 218016
rect 213184 208072 213236 208078
rect 213184 208014 213236 208020
rect 214288 207052 214340 207058
rect 214288 206994 214340 207000
rect 213828 205692 213880 205698
rect 213828 205634 213880 205640
rect 210424 203584 210476 203590
rect 210424 203526 210476 203532
rect 209872 201612 209924 201618
rect 209872 201554 209924 201560
rect 209884 199988 209912 201554
rect 212540 201544 212592 201550
rect 212540 201486 212592 201492
rect 211620 200456 211672 200462
rect 211620 200398 211672 200404
rect 210344 199974 210556 200002
rect 211632 199988 211660 200398
rect 212552 199988 212580 201486
rect 213840 200002 213868 205634
rect 213394 199974 213868 200002
rect 214300 199988 214328 206994
rect 215220 200002 215248 218010
rect 215956 207058 215984 231814
rect 216404 207664 216456 207670
rect 216404 207606 216456 207612
rect 215944 207052 215996 207058
rect 215944 206994 215996 207000
rect 216416 200002 216444 207606
rect 216864 206304 216916 206310
rect 216864 206246 216916 206252
rect 215142 199974 215248 200002
rect 216062 199974 216444 200002
rect 216876 199988 216904 206246
rect 217980 200002 218008 258062
rect 220636 210452 220688 210458
rect 220636 210394 220688 210400
rect 218612 202156 218664 202162
rect 218612 202098 218664 202104
rect 217810 199974 218008 200002
rect 218624 199988 218652 202098
rect 220648 201550 220676 210394
rect 219348 201544 219400 201550
rect 219348 201486 219400 201492
rect 219440 201544 219492 201550
rect 219440 201486 219492 201492
rect 220636 201544 220688 201550
rect 220636 201486 220688 201492
rect 219360 200802 219388 201486
rect 219348 200796 219400 200802
rect 219348 200738 219400 200744
rect 219452 199988 219480 201486
rect 220740 200002 220768 311850
rect 223488 221468 223540 221474
rect 223488 221410 223540 221416
rect 222108 211812 222160 211818
rect 222108 211754 222160 211760
rect 222120 201482 222148 211754
rect 223500 204254 223528 221410
rect 223856 207732 223908 207738
rect 223856 207674 223908 207680
rect 223408 204226 223528 204254
rect 222382 202192 222438 202201
rect 222382 202127 222438 202136
rect 221188 201476 221240 201482
rect 221188 201418 221240 201424
rect 222108 201476 222160 201482
rect 222108 201418 222160 201424
rect 220386 199974 220768 200002
rect 221200 199988 221228 201418
rect 222396 200002 222424 202127
rect 223408 200002 223436 204226
rect 222134 199974 222424 200002
rect 222962 199974 223436 200002
rect 223868 199988 223896 207674
rect 224880 200002 224908 430578
rect 231136 355366 231164 618258
rect 235920 606490 235948 699654
rect 235908 606484 235960 606490
rect 235908 606426 235960 606432
rect 238668 458856 238720 458862
rect 238668 458798 238720 458804
rect 234528 403640 234580 403646
rect 234528 403582 234580 403588
rect 231124 355360 231176 355366
rect 231124 355302 231176 355308
rect 231768 354000 231820 354006
rect 231768 353942 231820 353948
rect 226984 345092 227036 345098
rect 226984 345034 227036 345040
rect 226248 210860 226300 210866
rect 226248 210802 226300 210808
rect 226260 200114 226288 210802
rect 226996 209506 227024 345034
rect 229008 300144 229060 300150
rect 229008 300086 229060 300092
rect 226984 209500 227036 209506
rect 226984 209442 227036 209448
rect 227628 209092 227680 209098
rect 227628 209034 227680 209040
rect 226432 206576 226484 206582
rect 226432 206518 226484 206524
rect 225984 200086 226288 200114
rect 225984 200002 226012 200086
rect 224710 199974 224908 200002
rect 225630 199974 226012 200002
rect 226444 199988 226472 206518
rect 227640 200002 227668 209034
rect 228916 204944 228968 204950
rect 228916 204886 228968 204892
rect 228180 202836 228232 202842
rect 228180 202778 228232 202784
rect 227378 199974 227668 200002
rect 228192 199988 228220 202778
rect 228928 200002 228956 204886
rect 229020 202842 229048 300086
rect 231674 204912 231730 204921
rect 231674 204847 231730 204856
rect 230386 203552 230442 203561
rect 230386 203487 230442 203496
rect 229008 202836 229060 202842
rect 229008 202778 229060 202784
rect 230400 200002 230428 203487
rect 230756 202292 230808 202298
rect 230756 202234 230808 202240
rect 228928 199974 229034 200002
rect 229954 199974 230428 200002
rect 230768 199988 230796 202234
rect 231688 199988 231716 204847
rect 231780 202298 231808 353942
rect 232504 271924 232556 271930
rect 232504 271866 232556 271872
rect 232516 206310 232544 271866
rect 232964 209160 233016 209166
rect 232964 209102 233016 209108
rect 232504 206304 232556 206310
rect 232504 206246 232556 206252
rect 231768 202292 231820 202298
rect 231768 202234 231820 202240
rect 232976 200002 233004 209102
rect 234436 206304 234488 206310
rect 234436 206246 234488 206252
rect 233424 202360 233476 202366
rect 233424 202302 233476 202308
rect 232530 199974 233004 200002
rect 233436 199988 233464 202302
rect 234448 200002 234476 206246
rect 234540 202366 234568 403582
rect 235264 324352 235316 324358
rect 235264 324294 235316 324300
rect 235276 210458 235304 324294
rect 235264 210452 235316 210458
rect 235264 210394 235316 210400
rect 235908 210452 235960 210458
rect 235908 210394 235960 210400
rect 235920 202502 235948 210394
rect 237194 206272 237250 206281
rect 237194 206207 237250 206216
rect 235998 205048 236054 205057
rect 235998 204983 236054 204992
rect 235172 202496 235224 202502
rect 235172 202438 235224 202444
rect 235908 202496 235960 202502
rect 235908 202438 235960 202444
rect 234528 202360 234580 202366
rect 234528 202302 234580 202308
rect 234278 199974 234476 200002
rect 235184 199988 235212 202438
rect 236012 199988 236040 204983
rect 237208 200002 237236 206207
rect 238680 200002 238708 458798
rect 240048 246356 240100 246362
rect 240048 246298 240100 246304
rect 240060 205634 240088 246298
rect 240796 211886 240824 700266
rect 241428 214600 241480 214606
rect 241428 214542 241480 214548
rect 240784 211880 240836 211886
rect 240784 211822 240836 211828
rect 240324 207052 240376 207058
rect 240324 206994 240376 207000
rect 239968 205606 240088 205634
rect 239968 200002 239996 205606
rect 236854 199974 237236 200002
rect 238602 199974 238708 200002
rect 239522 199974 239996 200002
rect 240336 199988 240364 206994
rect 241440 200002 241468 214542
rect 242176 207058 242204 700266
rect 244188 210520 244240 210526
rect 244188 210462 244240 210468
rect 242530 207632 242586 207641
rect 242530 207567 242586 207576
rect 242164 207052 242216 207058
rect 242164 206994 242216 207000
rect 242544 200002 242572 207567
rect 242990 202872 243046 202881
rect 242990 202807 243046 202816
rect 241270 199974 241468 200002
rect 242098 199974 242572 200002
rect 243004 199988 243032 202807
rect 244200 200002 244228 210462
rect 244936 202881 244964 700334
rect 267660 697610 267688 703520
rect 283852 699718 283880 703520
rect 294604 700596 294656 700602
rect 294604 700538 294656 700544
rect 282184 699712 282236 699718
rect 282184 699654 282236 699660
rect 283840 699712 283892 699718
rect 283840 699654 283892 699660
rect 266360 697604 266412 697610
rect 266360 697546 266412 697552
rect 267648 697604 267700 697610
rect 267648 697546 267700 697552
rect 260104 670744 260156 670750
rect 260104 670686 260156 670692
rect 251088 649324 251140 649330
rect 251088 649266 251140 649272
rect 249064 409896 249116 409902
rect 249064 409838 249116 409844
rect 246304 364404 246356 364410
rect 246304 364346 246356 364352
rect 246316 221474 246344 364346
rect 249076 318102 249104 409838
rect 249064 318096 249116 318102
rect 249064 318038 249116 318044
rect 246304 221468 246356 221474
rect 246304 221410 246356 221416
rect 249708 220108 249760 220114
rect 249708 220050 249760 220056
rect 246948 217320 247000 217326
rect 246948 217262 247000 217268
rect 246028 207868 246080 207874
rect 246028 207810 246080 207816
rect 245568 205148 245620 205154
rect 245568 205090 245620 205096
rect 244922 202872 244978 202881
rect 244922 202807 244978 202816
rect 244738 202736 244794 202745
rect 244738 202671 244794 202680
rect 243846 199974 244228 200002
rect 244752 199988 244780 202671
rect 245580 199988 245608 205090
rect 246040 202745 246068 207810
rect 246960 204254 246988 217262
rect 248512 205012 248564 205018
rect 248512 204954 248564 204960
rect 246776 204226 246988 204254
rect 246026 202736 246082 202745
rect 246026 202671 246082 202680
rect 246776 200002 246804 204226
rect 247316 203652 247368 203658
rect 247316 203594 247368 203600
rect 246422 199974 246804 200002
rect 247328 199988 247356 203594
rect 248524 200002 248552 204954
rect 249720 204254 249748 220050
rect 250628 205216 250680 205222
rect 250628 205158 250680 205164
rect 249536 204226 249748 204254
rect 249536 200002 249564 204226
rect 250640 202609 250668 205158
rect 250626 202600 250682 202609
rect 250626 202535 250682 202544
rect 249892 201408 249944 201414
rect 249892 201350 249944 201356
rect 248170 199974 248552 200002
rect 249090 199974 249564 200002
rect 249904 199988 249932 201350
rect 251100 200002 251128 649266
rect 258724 632120 258776 632126
rect 258724 632062 258776 632068
rect 252560 606484 252612 606490
rect 252560 606426 252612 606432
rect 252468 294636 252520 294642
rect 252468 294578 252520 294584
rect 251180 206644 251232 206650
rect 251180 206586 251232 206592
rect 251192 201414 251220 206586
rect 252480 202026 252508 294578
rect 251640 202020 251692 202026
rect 251640 201962 251692 201968
rect 252468 202020 252520 202026
rect 252468 201962 252520 201968
rect 251180 201408 251232 201414
rect 251180 201350 251232 201356
rect 250838 199974 251128 200002
rect 251652 199988 251680 201962
rect 252572 199988 252600 606426
rect 255964 579692 256016 579698
rect 255964 579634 256016 579640
rect 254308 211880 254360 211886
rect 254308 211822 254360 211828
rect 252652 206372 252704 206378
rect 252652 206314 252704 206320
rect 252664 202881 252692 206314
rect 252650 202872 252706 202881
rect 252650 202807 252706 202816
rect 253386 202600 253442 202609
rect 253386 202535 253442 202544
rect 253400 199988 253428 202535
rect 254320 199988 254348 211822
rect 255504 205080 255556 205086
rect 255504 205022 255556 205028
rect 255318 203688 255374 203697
rect 255318 203623 255374 203632
rect 255134 202872 255190 202881
rect 255134 202807 255190 202816
rect 255148 199988 255176 202807
rect 255332 201929 255360 203623
rect 255318 201920 255374 201929
rect 255318 201855 255374 201864
rect 255516 200002 255544 205022
rect 255976 203833 256004 579634
rect 256884 207936 256936 207942
rect 256884 207878 256936 207884
rect 255962 203824 256018 203833
rect 255962 203759 256018 203768
rect 255516 199974 255990 200002
rect 256896 199988 256924 207878
rect 258630 205184 258686 205193
rect 258630 205119 258686 205128
rect 257710 201920 257766 201929
rect 257710 201855 257766 201864
rect 257724 199988 257752 201855
rect 258644 199988 258672 205119
rect 258736 204882 258764 632062
rect 260116 224262 260144 670686
rect 262864 656940 262916 656946
rect 262864 656882 262916 656888
rect 259460 224256 259512 224262
rect 259460 224198 259512 224204
rect 260104 224256 260156 224262
rect 260104 224198 260156 224204
rect 259184 207800 259236 207806
rect 259184 207742 259236 207748
rect 258724 204876 258776 204882
rect 258724 204818 258776 204824
rect 259196 202881 259224 207742
rect 259182 202872 259238 202881
rect 259182 202807 259238 202816
rect 259472 199988 259500 224198
rect 262128 210588 262180 210594
rect 262128 210530 262180 210536
rect 260748 209228 260800 209234
rect 260748 209170 260800 209176
rect 260378 202872 260434 202881
rect 260760 202858 260788 209170
rect 260760 202830 260880 202858
rect 260378 202807 260434 202816
rect 260392 199988 260420 202807
rect 260852 200114 260880 202830
rect 260852 200086 261248 200114
rect 261220 199988 261248 200086
rect 262140 199988 262168 210530
rect 262876 208894 262904 656882
rect 266372 649330 266400 697546
rect 266360 649324 266412 649330
rect 266360 649266 266412 649272
rect 280344 357468 280396 357474
rect 280344 357410 280396 357416
rect 267280 355360 267332 355366
rect 267280 355302 267332 355308
rect 264704 224256 264756 224262
rect 264704 224198 264756 224204
rect 262956 209432 263008 209438
rect 262956 209374 263008 209380
rect 262864 208888 262916 208894
rect 262864 208830 262916 208836
rect 262968 199988 262996 209374
rect 263876 208888 263928 208894
rect 263876 208830 263928 208836
rect 263888 199988 263916 208830
rect 264716 199988 264744 224198
rect 266452 209364 266504 209370
rect 266452 209306 266504 209312
rect 265532 204876 265584 204882
rect 265532 204818 265584 204824
rect 265544 199988 265572 204818
rect 266464 199988 266492 209306
rect 267292 199988 267320 355302
rect 269948 344344 270000 344350
rect 269948 344286 270000 344292
rect 269028 215960 269080 215966
rect 269028 215902 269080 215908
rect 268198 203824 268254 203833
rect 268198 203759 268254 203768
rect 268212 199988 268240 203759
rect 269040 199988 269068 215902
rect 269960 199988 269988 344286
rect 277768 318096 277820 318102
rect 277768 318038 277820 318044
rect 276848 286340 276900 286346
rect 276848 286282 276900 286288
rect 274272 228404 274324 228410
rect 274272 228346 274324 228352
rect 271696 227044 271748 227050
rect 271696 226986 271748 226992
rect 270776 203584 270828 203590
rect 270776 203526 270828 203532
rect 270788 199988 270816 203526
rect 271708 199988 271736 226986
rect 272524 210792 272576 210798
rect 272524 210734 272576 210740
rect 272536 199988 272564 210734
rect 273352 206440 273404 206446
rect 273352 206382 273404 206388
rect 273364 199988 273392 206382
rect 274284 199988 274312 228346
rect 275100 210656 275152 210662
rect 275100 210598 275152 210604
rect 275112 199988 275140 210598
rect 276020 208004 276072 208010
rect 276020 207946 276072 207952
rect 276032 199988 276060 207946
rect 276860 199988 276888 286282
rect 277780 199988 277808 318038
rect 279516 209500 279568 209506
rect 279516 209442 279568 209448
rect 278596 208072 278648 208078
rect 278596 208014 278648 208020
rect 278608 199988 278636 208014
rect 279528 199988 279556 209442
rect 280356 199988 280384 357410
rect 282196 294642 282224 699654
rect 291844 456816 291896 456822
rect 291844 456758 291896 456764
rect 289084 418192 289136 418198
rect 289084 418134 289136 418140
rect 282184 294636 282236 294642
rect 282184 294578 282236 294584
rect 282092 292596 282144 292602
rect 282092 292538 282144 292544
rect 281264 206508 281316 206514
rect 281264 206450 281316 206456
rect 281276 199988 281304 206450
rect 282104 199988 282132 292538
rect 285680 266416 285732 266422
rect 285680 266358 285732 266364
rect 285588 253972 285640 253978
rect 285588 253914 285640 253920
rect 282920 210724 282972 210730
rect 282920 210666 282972 210672
rect 282932 199988 282960 210666
rect 284668 209296 284720 209302
rect 284668 209238 284720 209244
rect 283840 203176 283892 203182
rect 283840 203118 283892 203124
rect 283852 199988 283880 203118
rect 284680 199988 284708 209238
rect 285600 199988 285628 253914
rect 285692 203182 285720 266358
rect 287060 213988 287112 213994
rect 287060 213930 287112 213936
rect 285680 203176 285732 203182
rect 285680 203118 285732 203124
rect 287072 202994 287100 213930
rect 289096 210866 289124 418134
rect 289084 210860 289136 210866
rect 289084 210802 289136 210808
rect 291856 206582 291884 456758
rect 291844 206576 291896 206582
rect 291844 206518 291896 206524
rect 294616 203658 294644 700538
rect 298744 700528 298796 700534
rect 298744 700470 298796 700476
rect 295984 351960 296036 351966
rect 295984 351902 296036 351908
rect 295996 211818 296024 351902
rect 295984 211812 296036 211818
rect 295984 211754 296036 211760
rect 298756 205154 298784 700470
rect 299492 206650 299520 703582
rect 299952 703474 299980 703582
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 412652 703582 413508 703610
rect 300136 703474 300164 703520
rect 299952 703446 300164 703474
rect 332520 703050 332548 703520
rect 331220 703044 331272 703050
rect 331220 702986 331272 702992
rect 332508 703044 332560 703050
rect 332508 702986 332560 702992
rect 305644 700460 305696 700466
rect 305644 700402 305696 700408
rect 305656 207641 305684 700402
rect 305642 207632 305698 207641
rect 305642 207567 305698 207576
rect 299480 206644 299532 206650
rect 299480 206586 299532 206592
rect 298744 205148 298796 205154
rect 298744 205090 298796 205096
rect 331232 205018 331260 702986
rect 348804 699718 348832 703520
rect 364996 700602 365024 703520
rect 364984 700596 365036 700602
rect 364984 700538 365036 700544
rect 397472 700534 397500 703520
rect 397460 700528 397512 700534
rect 397460 700470 397512 700476
rect 347044 699712 347096 699718
rect 347044 699654 347096 699660
rect 348792 699712 348844 699718
rect 348792 699654 348844 699660
rect 347056 220114 347084 699654
rect 347044 220108 347096 220114
rect 347044 220050 347096 220056
rect 412652 217326 412680 703582
rect 413480 703474 413508 703582
rect 413622 703520 413734 704960
rect 429212 703582 429700 703610
rect 413664 703474 413692 703520
rect 413480 703446 413692 703474
rect 412640 217320 412692 217326
rect 412640 217262 412692 217268
rect 429212 207874 429240 703582
rect 429672 703474 429700 703582
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 429856 703474 429884 703520
rect 429672 703446 429884 703474
rect 462332 700398 462360 703520
rect 462320 700392 462372 700398
rect 462320 700334 462372 700340
rect 478524 699718 478552 703520
rect 494808 700466 494836 703520
rect 494796 700460 494848 700466
rect 494796 700402 494848 700408
rect 527192 700330 527220 703520
rect 543476 702434 543504 703520
rect 542372 702406 543504 702434
rect 527180 700324 527232 700330
rect 527180 700266 527232 700272
rect 476764 699712 476816 699718
rect 476764 699654 476816 699660
rect 478512 699712 478564 699718
rect 478512 699654 478564 699660
rect 476776 210526 476804 699654
rect 542372 214606 542400 702406
rect 559668 700330 559696 703520
rect 559656 700324 559708 700330
rect 559656 700266 559708 700272
rect 582932 700324 582984 700330
rect 582932 700266 582984 700272
rect 582470 670712 582526 670721
rect 582470 670647 582526 670656
rect 580170 458144 580226 458153
rect 580170 458079 580226 458088
rect 580184 456822 580212 458079
rect 580172 456816 580224 456822
rect 580172 456758 580224 456764
rect 580170 431624 580226 431633
rect 580170 431559 580226 431568
rect 580184 430642 580212 431559
rect 580172 430636 580224 430642
rect 580172 430578 580224 430584
rect 580170 418296 580226 418305
rect 580170 418231 580226 418240
rect 580184 418198 580212 418231
rect 580172 418192 580224 418198
rect 580172 418134 580224 418140
rect 580906 378448 580962 378457
rect 580906 378383 580962 378392
rect 580170 365120 580226 365129
rect 580170 365055 580226 365064
rect 580184 364410 580212 365055
rect 580172 364404 580224 364410
rect 580172 364346 580224 364352
rect 579896 351960 579948 351966
rect 579894 351928 579896 351937
rect 579948 351928 579950 351937
rect 579894 351863 579950 351872
rect 580920 343262 580948 378383
rect 580908 343256 580960 343262
rect 580908 343198 580960 343204
rect 580170 325272 580226 325281
rect 580170 325207 580226 325216
rect 580184 324358 580212 325207
rect 580172 324352 580224 324358
rect 580172 324294 580224 324300
rect 580170 312080 580226 312089
rect 580170 312015 580226 312024
rect 580184 311914 580212 312015
rect 580172 311908 580224 311914
rect 580172 311850 580224 311856
rect 580906 298752 580962 298761
rect 580906 298687 580962 298696
rect 580170 272232 580226 272241
rect 580170 272167 580226 272176
rect 580184 271930 580212 272167
rect 580172 271924 580224 271930
rect 580172 271866 580224 271872
rect 580170 258904 580226 258913
rect 580170 258839 580226 258848
rect 580184 258126 580212 258839
rect 580172 258120 580224 258126
rect 580172 258062 580224 258068
rect 580170 232384 580226 232393
rect 580170 232319 580226 232328
rect 580184 231878 580212 232319
rect 580172 231872 580224 231878
rect 580172 231814 580224 231820
rect 580170 219056 580226 219065
rect 580170 218991 580226 219000
rect 580184 218074 580212 218991
rect 580172 218068 580224 218074
rect 580172 218010 580224 218016
rect 542360 214600 542412 214606
rect 542360 214542 542412 214548
rect 580920 211138 580948 298687
rect 580908 211132 580960 211138
rect 580908 211074 580960 211080
rect 582380 211132 582432 211138
rect 582380 211074 582432 211080
rect 476764 210520 476816 210526
rect 476764 210462 476816 210468
rect 429200 207868 429252 207874
rect 429200 207810 429252 207816
rect 580170 205728 580226 205737
rect 580170 205663 580172 205672
rect 580224 205663 580226 205672
rect 580172 205634 580224 205640
rect 331220 205012 331272 205018
rect 331220 204954 331272 204960
rect 294604 203652 294656 203658
rect 294604 203594 294656 203600
rect 289084 203244 289136 203250
rect 289084 203186 289136 203192
rect 286888 202966 287100 202994
rect 286888 200002 286916 202966
rect 288164 201680 288216 201686
rect 288164 201622 288216 201628
rect 286442 199974 286916 200002
rect 288176 199988 288204 201622
rect 289096 199988 289124 203186
rect 582392 202162 582420 211074
rect 582484 206281 582512 670647
rect 582562 644056 582618 644065
rect 582562 643991 582618 644000
rect 582576 210458 582604 643991
rect 582654 630864 582710 630873
rect 582654 630799 582710 630808
rect 582564 210452 582616 210458
rect 582564 210394 582616 210400
rect 582470 206272 582526 206281
rect 582470 206207 582526 206216
rect 582668 205057 582696 630799
rect 582746 617536 582802 617545
rect 582746 617471 582802 617480
rect 582760 206310 582788 617471
rect 582838 591016 582894 591025
rect 582838 590951 582894 590960
rect 582852 209166 582880 590951
rect 582944 246362 582972 700266
rect 583758 696960 583814 696969
rect 583758 696895 583814 696904
rect 583390 683904 583446 683913
rect 583390 683839 583446 683848
rect 583022 564360 583078 564369
rect 583022 564295 583078 564304
rect 582932 246356 582984 246362
rect 582932 246298 582984 246304
rect 582930 245576 582986 245585
rect 582930 245511 582986 245520
rect 582840 209160 582892 209166
rect 582840 209102 582892 209108
rect 582944 207670 582972 245511
rect 582932 207664 582984 207670
rect 582932 207606 582984 207612
rect 582748 206304 582800 206310
rect 582748 206246 582800 206252
rect 582654 205048 582710 205057
rect 582654 204983 582710 204992
rect 583036 204921 583064 564295
rect 583114 537840 583170 537849
rect 583114 537775 583170 537784
rect 583022 204912 583078 204921
rect 583022 204847 583078 204856
rect 582472 204332 582524 204338
rect 582472 204274 582524 204280
rect 582380 202156 582432 202162
rect 582380 202098 582432 202104
rect 295984 201884 296036 201890
rect 295984 201826 296036 201832
rect 292488 201748 292540 201754
rect 292488 201690 292540 201696
rect 290832 200864 290884 200870
rect 290832 200806 290884 200812
rect 290844 199988 290872 200806
rect 292500 199988 292528 201690
rect 293408 200252 293460 200258
rect 293408 200194 293460 200200
rect 293420 199988 293448 200194
rect 295996 199988 296024 201826
rect 298652 201816 298704 201822
rect 298652 201758 298704 201764
rect 297732 200320 297784 200326
rect 297732 200262 297784 200268
rect 297744 199988 297772 200262
rect 298664 199988 298692 201758
rect 580264 200796 580316 200802
rect 580264 200738 580316 200744
rect 304264 200456 304316 200462
rect 304264 200398 304316 200404
rect 299480 200388 299532 200394
rect 299480 200330 299532 200336
rect 299492 199988 299520 200330
rect 203536 199838 203826 199866
rect 206494 199850 206784 199866
rect 206494 199844 206796 199850
rect 206494 199838 206744 199844
rect 199936 199776 199988 199782
rect 199936 199718 199988 199724
rect 199842 199608 199898 199617
rect 199384 199572 199436 199578
rect 199842 199543 199898 199552
rect 199384 199514 199436 199520
rect 198002 199336 198058 199345
rect 198002 199271 198058 199280
rect 198016 198762 198044 199271
rect 183008 198756 183060 198762
rect 183008 198698 183060 198704
rect 198004 198756 198056 198762
rect 198004 198698 198056 198704
rect 174544 197396 174596 197402
rect 174544 197338 174596 197344
rect 170496 193248 170548 193254
rect 170496 193190 170548 193196
rect 170402 173292 170458 173301
rect 170402 173227 170458 173236
rect 169208 164280 169260 164286
rect 169208 164222 169260 164228
rect 159364 164212 159416 164218
rect 159364 164154 159416 164160
rect 160008 161492 160060 161498
rect 160008 161434 160060 161440
rect 157984 137964 158036 137970
rect 157984 137906 158036 137912
rect 157248 122732 157300 122738
rect 157248 122674 157300 122680
rect 148324 111784 148376 111790
rect 148324 111726 148376 111732
rect 160020 104854 160048 161434
rect 160836 160744 160888 160750
rect 169220 160698 169248 164222
rect 169392 162172 169444 162178
rect 169392 162114 169444 162120
rect 169298 161528 169354 161537
rect 169298 161463 169300 161472
rect 169352 161463 169354 161472
rect 169300 161434 169352 161440
rect 169300 160812 169352 160818
rect 169300 160754 169352 160760
rect 160888 160692 160954 160698
rect 160836 160686 160954 160692
rect 160848 160670 160954 160686
rect 168958 160670 169248 160698
rect 169312 160546 169340 160754
rect 165160 160540 165212 160546
rect 165160 160482 165212 160488
rect 169300 160540 169352 160546
rect 169300 160482 169352 160488
rect 165172 160426 165200 160482
rect 162886 160410 163176 160426
rect 162886 160404 163188 160410
rect 162886 160398 163136 160404
rect 164910 160398 165200 160426
rect 166816 160472 166868 160478
rect 166868 160420 166934 160426
rect 166816 160414 166934 160420
rect 166828 160398 166934 160414
rect 163136 160346 163188 160352
rect 169404 144265 169432 162114
rect 169390 144256 169446 144265
rect 169390 144191 169446 144200
rect 170416 130422 170444 173227
rect 170508 160410 170536 193190
rect 172426 189272 172482 189281
rect 172426 189207 172482 189216
rect 172440 189174 172468 189207
rect 172428 189168 172480 189174
rect 172428 189110 172480 189116
rect 171782 187776 171838 187785
rect 171782 187711 171838 187720
rect 173164 187740 173216 187746
rect 171796 185638 171824 187711
rect 173164 187682 173216 187688
rect 172426 186824 172482 186833
rect 172426 186759 172482 186768
rect 172440 186454 172468 186759
rect 172428 186448 172480 186454
rect 172428 186390 172480 186396
rect 171784 185632 171836 185638
rect 171784 185574 171836 185580
rect 171782 185464 171838 185473
rect 171782 185399 171838 185408
rect 171690 184240 171746 184249
rect 171690 184175 171746 184184
rect 171704 183598 171732 184175
rect 171692 183592 171744 183598
rect 171692 183534 171744 183540
rect 171796 173262 171824 185399
rect 172426 183696 172482 183705
rect 172426 183631 172428 183640
rect 172480 183631 172482 183640
rect 172428 183602 172480 183608
rect 172426 182472 172482 182481
rect 172426 182407 172482 182416
rect 172440 182306 172468 182407
rect 172428 182300 172480 182306
rect 172428 182242 172480 182248
rect 172426 181112 172482 181121
rect 172426 181047 172482 181056
rect 172440 180878 172468 181047
rect 172428 180872 172480 180878
rect 172428 180814 172480 180820
rect 172058 179888 172114 179897
rect 172058 179823 172114 179832
rect 172072 179518 172100 179823
rect 172060 179512 172112 179518
rect 172060 179454 172112 179460
rect 172150 178664 172206 178673
rect 172150 178599 172206 178608
rect 172164 178158 172192 178599
rect 172152 178152 172204 178158
rect 172152 178094 172204 178100
rect 172242 177304 172298 177313
rect 172242 177239 172298 177248
rect 172256 176730 172284 177239
rect 172428 176792 172480 176798
rect 172426 176760 172428 176769
rect 172480 176760 172482 176769
rect 172244 176724 172296 176730
rect 172426 176695 172482 176704
rect 172244 176666 172296 176672
rect 172426 175400 172482 175409
rect 172426 175335 172482 175344
rect 172440 175302 172468 175335
rect 172428 175296 172480 175302
rect 172428 175238 172480 175244
rect 171966 174176 172022 174185
rect 171966 174111 172022 174120
rect 171784 173256 171836 173262
rect 171784 173198 171836 173204
rect 171782 169824 171838 169833
rect 171782 169759 171838 169768
rect 171138 164792 171194 164801
rect 171138 164727 171194 164736
rect 171152 164354 171180 164727
rect 171140 164348 171192 164354
rect 171140 164290 171192 164296
rect 171690 163432 171746 163441
rect 171690 163367 171746 163376
rect 171704 162926 171732 163367
rect 171692 162920 171744 162926
rect 171692 162862 171744 162868
rect 171692 160880 171744 160886
rect 171692 160822 171744 160828
rect 171704 160478 171732 160822
rect 171692 160472 171744 160478
rect 171692 160414 171744 160420
rect 170496 160404 170548 160410
rect 170496 160346 170548 160352
rect 170496 154624 170548 154630
rect 170496 154566 170548 154572
rect 170508 137601 170536 154566
rect 171692 154556 171744 154562
rect 171692 154498 171744 154504
rect 171704 153241 171732 154498
rect 171690 153232 171746 153241
rect 171690 153167 171746 153176
rect 171508 153128 171560 153134
rect 171508 153070 171560 153076
rect 171520 152697 171548 153070
rect 171506 152688 171562 152697
rect 171506 152623 171562 152632
rect 171324 151224 171376 151230
rect 171324 151166 171376 151172
rect 171336 150521 171364 151166
rect 171322 150512 171378 150521
rect 171322 150447 171378 150456
rect 171508 149660 171560 149666
rect 171508 149602 171560 149608
rect 171520 149433 171548 149602
rect 171506 149424 171562 149433
rect 171506 149359 171562 149368
rect 171692 149048 171744 149054
rect 171692 148990 171744 148996
rect 171324 148368 171376 148374
rect 171322 148336 171324 148345
rect 171376 148336 171378 148345
rect 171322 148271 171378 148280
rect 171704 147801 171732 148990
rect 171690 147792 171746 147801
rect 171690 147727 171746 147736
rect 171324 144900 171376 144906
rect 171324 144842 171376 144848
rect 171336 143585 171364 144842
rect 171322 143576 171378 143585
rect 171322 143511 171378 143520
rect 171692 143404 171744 143410
rect 171692 143346 171744 143352
rect 171704 143041 171732 143346
rect 171690 143032 171746 143041
rect 171690 142967 171746 142976
rect 171508 142112 171560 142118
rect 171508 142054 171560 142060
rect 171520 141953 171548 142054
rect 171506 141944 171562 141953
rect 171506 141879 171562 141888
rect 171508 141024 171560 141030
rect 171508 140966 171560 140972
rect 171520 140865 171548 140966
rect 171506 140856 171562 140865
rect 171506 140791 171562 140800
rect 171692 140684 171744 140690
rect 171692 140626 171744 140632
rect 171704 139777 171732 140626
rect 171690 139768 171746 139777
rect 171690 139703 171746 139712
rect 171324 139392 171376 139398
rect 171324 139334 171376 139340
rect 171336 138689 171364 139334
rect 171322 138680 171378 138689
rect 171322 138615 171378 138624
rect 171508 137964 171560 137970
rect 171508 137906 171560 137912
rect 170494 137592 170550 137601
rect 170494 137527 170550 137536
rect 171520 137057 171548 137906
rect 171506 137048 171562 137057
rect 171506 136983 171562 136992
rect 171692 136536 171744 136542
rect 171692 136478 171744 136484
rect 171704 135969 171732 136478
rect 171690 135960 171746 135969
rect 171690 135895 171746 135904
rect 171508 135652 171560 135658
rect 171508 135594 171560 135600
rect 171520 135425 171548 135594
rect 171506 135416 171562 135425
rect 171506 135351 171562 135360
rect 171508 135244 171560 135250
rect 171508 135186 171560 135192
rect 171520 134337 171548 135186
rect 171506 134328 171562 134337
rect 171506 134263 171562 134272
rect 171692 133884 171744 133890
rect 171692 133826 171744 133832
rect 171704 132841 171732 133826
rect 171690 132832 171746 132841
rect 171690 132767 171746 132776
rect 171692 132456 171744 132462
rect 171692 132398 171744 132404
rect 171704 132297 171732 132398
rect 171690 132288 171746 132297
rect 171690 132223 171746 132232
rect 171690 130656 171746 130665
rect 171690 130591 171746 130600
rect 170404 130416 170456 130422
rect 170404 130358 170456 130364
rect 171704 129878 171732 130591
rect 171692 129872 171744 129878
rect 171692 129814 171744 129820
rect 170402 129568 170458 129577
rect 170402 129503 170458 129512
rect 160652 124160 160704 124166
rect 160704 124108 160954 124114
rect 160652 124102 160954 124108
rect 160664 124086 160954 124102
rect 162872 122874 162900 124100
rect 162860 122868 162912 122874
rect 162860 122810 162912 122816
rect 164896 122806 164924 124100
rect 164884 122800 164936 122806
rect 164884 122742 164936 122748
rect 166920 122738 166948 124100
rect 168944 122806 168972 124100
rect 168932 122800 168984 122806
rect 168932 122742 168984 122748
rect 170416 122738 170444 129503
rect 171598 129024 171654 129033
rect 171598 128959 171654 128968
rect 171612 128382 171640 128959
rect 171600 128376 171652 128382
rect 171600 128318 171652 128324
rect 171690 127936 171746 127945
rect 171690 127871 171746 127880
rect 171704 127022 171732 127871
rect 171692 127016 171744 127022
rect 171692 126958 171744 126964
rect 171690 124672 171746 124681
rect 171690 124607 171746 124616
rect 171704 124302 171732 124607
rect 171692 124296 171744 124302
rect 171692 124238 171744 124244
rect 166908 122732 166960 122738
rect 166908 122674 166960 122680
rect 170404 122732 170456 122738
rect 170404 122674 170456 122680
rect 171796 120766 171824 169759
rect 171874 163024 171930 163033
rect 171874 162959 171876 162968
rect 171928 162959 171930 162968
rect 171876 162930 171928 162936
rect 171874 160440 171930 160449
rect 171874 160375 171930 160384
rect 171888 160138 171916 160375
rect 171876 160132 171928 160138
rect 171876 160074 171928 160080
rect 171980 158710 172008 174111
rect 172242 171728 172298 171737
rect 172242 171663 172298 171672
rect 172256 171154 172284 171663
rect 172244 171148 172296 171154
rect 172244 171090 172296 171096
rect 172242 170368 172298 170377
rect 172242 170303 172298 170312
rect 172256 169794 172284 170303
rect 172244 169788 172296 169794
rect 172244 169730 172296 169736
rect 172426 168600 172482 168609
rect 172426 168535 172482 168544
rect 172440 168434 172468 168535
rect 172428 168428 172480 168434
rect 172428 168370 172480 168376
rect 172426 167376 172482 167385
rect 172426 167311 172482 167320
rect 172440 167142 172468 167311
rect 172428 167136 172480 167142
rect 172428 167078 172480 167084
rect 172060 166320 172112 166326
rect 172060 166262 172112 166268
rect 171968 158704 172020 158710
rect 171968 158646 172020 158652
rect 172072 157334 172100 166262
rect 172426 166016 172482 166025
rect 172426 165951 172482 165960
rect 172440 165714 172468 165951
rect 172428 165708 172480 165714
rect 172428 165650 172480 165656
rect 171888 157306 172100 157334
rect 171888 149977 171916 157306
rect 172244 156052 172296 156058
rect 172244 155994 172296 156000
rect 171968 155372 172020 155378
rect 171968 155314 172020 155320
rect 171874 149968 171930 149977
rect 171874 149903 171930 149912
rect 171980 146713 172008 155314
rect 172256 153785 172284 155994
rect 173176 154562 173204 187682
rect 173440 173936 173492 173942
rect 173440 173878 173492 173884
rect 173348 159384 173400 159390
rect 173348 159326 173400 159332
rect 173256 158704 173308 158710
rect 173256 158646 173308 158652
rect 173164 154556 173216 154562
rect 173164 154498 173216 154504
rect 172242 153776 172298 153785
rect 172242 153711 172298 153720
rect 172336 153196 172388 153202
rect 172336 153138 172388 153144
rect 172348 152153 172376 153138
rect 172334 152144 172390 152153
rect 172334 152079 172390 152088
rect 172336 151700 172388 151706
rect 172336 151642 172388 151648
rect 172348 151609 172376 151642
rect 172428 151632 172480 151638
rect 172334 151600 172390 151609
rect 172428 151574 172480 151580
rect 172334 151535 172390 151544
rect 172440 151065 172468 151574
rect 172426 151056 172482 151065
rect 172426 150991 172482 151000
rect 172244 149728 172296 149734
rect 172244 149670 172296 149676
rect 171966 146704 172022 146713
rect 171966 146639 172022 146648
rect 172150 146160 172206 146169
rect 172150 146095 172152 146104
rect 172204 146095 172206 146104
rect 172152 146066 172204 146072
rect 172256 144537 172284 149670
rect 172428 148980 172480 148986
rect 172428 148922 172480 148928
rect 172440 148889 172468 148922
rect 172426 148880 172482 148889
rect 172426 148815 172482 148824
rect 172428 147620 172480 147626
rect 172428 147562 172480 147568
rect 172440 147257 172468 147562
rect 172426 147248 172482 147257
rect 172426 147183 172482 147192
rect 172336 146260 172388 146266
rect 172336 146202 172388 146208
rect 172348 145081 172376 146202
rect 172428 146192 172480 146198
rect 172428 146134 172480 146140
rect 172440 145625 172468 146134
rect 172426 145616 172482 145625
rect 172426 145551 172482 145560
rect 172334 145072 172390 145081
rect 172334 145007 172390 145016
rect 172242 144528 172298 144537
rect 172242 144463 172298 144472
rect 171968 144220 172020 144226
rect 171968 144162 172020 144168
rect 171876 142860 171928 142866
rect 171876 142802 171928 142808
rect 171888 134881 171916 142802
rect 171980 138145 172008 144162
rect 172428 143540 172480 143546
rect 172428 143482 172480 143488
rect 172440 142497 172468 143482
rect 172426 142488 172482 142497
rect 172426 142423 172482 142432
rect 172428 141568 172480 141574
rect 172428 141510 172480 141516
rect 172440 141409 172468 141510
rect 172426 141400 172482 141409
rect 172426 141335 172482 141344
rect 172428 140752 172480 140758
rect 172428 140694 172480 140700
rect 172440 140321 172468 140694
rect 172426 140312 172482 140321
rect 172426 140247 172482 140256
rect 172428 139256 172480 139262
rect 172426 139224 172428 139233
rect 172480 139224 172482 139233
rect 172426 139159 172482 139168
rect 171966 138136 172022 138145
rect 171966 138071 172022 138080
rect 172428 136604 172480 136610
rect 172428 136546 172480 136552
rect 172440 136513 172468 136546
rect 172426 136504 172482 136513
rect 172426 136439 172482 136448
rect 171874 134872 171930 134881
rect 171874 134807 171930 134816
rect 171876 134768 171928 134774
rect 171876 134710 171928 134716
rect 171888 133929 171916 134710
rect 171874 133920 171930 133929
rect 171874 133855 171930 133864
rect 172428 133408 172480 133414
rect 172426 133376 172428 133385
rect 172480 133376 172482 133385
rect 172426 133311 172482 133320
rect 172428 131776 172480 131782
rect 172426 131744 172428 131753
rect 172480 131744 172482 131753
rect 172426 131679 172482 131688
rect 172426 131200 172482 131209
rect 172426 131135 172428 131144
rect 172480 131135 172482 131144
rect 172428 131106 172480 131112
rect 172058 130112 172114 130121
rect 172058 130047 172114 130056
rect 172072 129810 172100 130047
rect 172060 129804 172112 129810
rect 172060 129746 172112 129752
rect 172426 128480 172482 128489
rect 172426 128415 172428 128424
rect 172480 128415 172482 128424
rect 172428 128386 172480 128392
rect 173268 128314 173296 158646
rect 173360 140690 173388 159326
rect 173452 155378 173480 173878
rect 174556 164286 174584 197338
rect 181536 196036 181588 196042
rect 181536 195978 181588 195984
rect 180156 189100 180208 189106
rect 180156 189042 180208 189048
rect 178776 186380 178828 186386
rect 178776 186322 178828 186328
rect 177304 183660 177356 183666
rect 177304 183602 177356 183608
rect 176016 183592 176068 183598
rect 176016 183534 176068 183540
rect 174636 182232 174688 182238
rect 174636 182174 174688 182180
rect 174544 164280 174596 164286
rect 174544 164222 174596 164228
rect 174544 162988 174596 162994
rect 174544 162930 174596 162936
rect 173440 155372 173492 155378
rect 173440 155314 173492 155320
rect 173348 140684 173400 140690
rect 173348 140626 173400 140632
rect 173256 128308 173308 128314
rect 173256 128250 173308 128256
rect 172058 127392 172114 127401
rect 172058 127327 172114 127336
rect 172072 127090 172100 127327
rect 172060 127084 172112 127090
rect 172060 127026 172112 127032
rect 173164 127084 173216 127090
rect 173164 127026 173216 127032
rect 172334 126848 172390 126857
rect 172334 126783 172390 126792
rect 172150 126304 172206 126313
rect 172150 126239 172206 126248
rect 172164 125662 172192 126239
rect 172152 125656 172204 125662
rect 172152 125598 172204 125604
rect 171874 125216 171930 125225
rect 171874 125151 171930 125160
rect 171888 124370 171916 125151
rect 172348 124914 172376 126783
rect 172426 125760 172482 125769
rect 172426 125695 172428 125704
rect 172480 125695 172482 125704
rect 172428 125666 172480 125672
rect 172336 124908 172388 124914
rect 172336 124850 172388 124856
rect 171876 124364 171928 124370
rect 171876 124306 171928 124312
rect 172426 124264 172482 124273
rect 172426 124199 172428 124208
rect 172480 124199 172482 124208
rect 172428 124170 172480 124176
rect 171784 120760 171836 120766
rect 171784 120702 171836 120708
rect 173176 114510 173204 127026
rect 173164 114504 173216 114510
rect 173164 114446 173216 114452
rect 174556 106282 174584 162930
rect 174648 151230 174676 182174
rect 175924 178084 175976 178090
rect 175924 178026 175976 178032
rect 174728 167068 174780 167074
rect 174728 167010 174780 167016
rect 174636 151224 174688 151230
rect 174636 151166 174688 151172
rect 174740 143410 174768 167010
rect 175936 148374 175964 178026
rect 176028 173194 176056 183534
rect 176016 173188 176068 173194
rect 176016 173130 176068 173136
rect 176016 171828 176068 171834
rect 176016 171770 176068 171776
rect 175924 148368 175976 148374
rect 175924 148310 175976 148316
rect 176028 146130 176056 171770
rect 176108 158772 176160 158778
rect 176108 158714 176160 158720
rect 176016 146124 176068 146130
rect 176016 146066 176068 146072
rect 174728 143404 174780 143410
rect 174728 143346 174780 143352
rect 176016 139460 176068 139466
rect 176016 139402 176068 139408
rect 175280 135312 175332 135318
rect 175280 135254 175332 135260
rect 175292 133890 175320 135254
rect 176028 134774 176056 139402
rect 176120 139262 176148 158714
rect 177316 146946 177344 183602
rect 177396 179444 177448 179450
rect 177396 179386 177448 179392
rect 177408 149666 177436 179386
rect 177488 164280 177540 164286
rect 177488 164222 177540 164228
rect 177396 149660 177448 149666
rect 177396 149602 177448 149608
rect 177396 147688 177448 147694
rect 177396 147630 177448 147636
rect 177304 146940 177356 146946
rect 177304 146882 177356 146888
rect 176108 139256 176160 139262
rect 176108 139198 176160 139204
rect 176660 136672 176712 136678
rect 176660 136614 176712 136620
rect 176016 134768 176068 134774
rect 176016 134710 176068 134716
rect 175280 133884 175332 133890
rect 175280 133826 175332 133832
rect 176672 133414 176700 136614
rect 177408 136542 177436 147630
rect 177500 142118 177528 164222
rect 178684 162920 178736 162926
rect 178684 162862 178736 162868
rect 177488 142112 177540 142118
rect 177488 142054 177540 142060
rect 177396 136536 177448 136542
rect 177396 136478 177448 136484
rect 176660 133408 176712 133414
rect 176660 133350 176712 133356
rect 176660 131164 176712 131170
rect 176660 131106 176712 131112
rect 175924 129872 175976 129878
rect 175924 129814 175976 129820
rect 175936 126954 175964 129814
rect 176672 129742 176700 131106
rect 176660 129736 176712 129742
rect 176660 129678 176712 129684
rect 177304 128444 177356 128450
rect 177304 128386 177356 128392
rect 175924 126948 175976 126954
rect 175924 126890 175976 126896
rect 175924 124228 175976 124234
rect 175924 124170 175976 124176
rect 174544 106276 174596 106282
rect 174544 106218 174596 106224
rect 160008 104848 160060 104854
rect 160008 104790 160060 104796
rect 175936 102814 175964 124170
rect 177316 118658 177344 128386
rect 178696 127634 178724 162862
rect 178788 153134 178816 186322
rect 178868 184204 178920 184210
rect 178868 184146 178920 184152
rect 178776 153128 178828 153134
rect 178776 153070 178828 153076
rect 178880 151706 178908 184146
rect 180064 176792 180116 176798
rect 180064 176734 180116 176740
rect 178960 162240 179012 162246
rect 178960 162182 179012 162188
rect 178868 151700 178920 151706
rect 178868 151642 178920 151648
rect 178776 146328 178828 146334
rect 178776 146270 178828 146276
rect 178788 135658 178816 146270
rect 178972 141030 179000 162182
rect 178960 141024 179012 141030
rect 178960 140966 179012 140972
rect 178776 135652 178828 135658
rect 178776 135594 178828 135600
rect 180076 132462 180104 176734
rect 180168 156058 180196 189042
rect 181444 171148 181496 171154
rect 181444 171090 181496 171096
rect 180248 163532 180300 163538
rect 180248 163474 180300 163480
rect 180156 156052 180208 156058
rect 180156 155994 180208 156000
rect 180260 141574 180288 163474
rect 180248 141568 180300 141574
rect 180248 141510 180300 141516
rect 180064 132456 180116 132462
rect 180064 132398 180116 132404
rect 180156 128376 180208 128382
rect 180156 128318 180208 128324
rect 178684 127628 178736 127634
rect 178684 127570 178736 127576
rect 178040 127016 178092 127022
rect 178040 126958 178092 126964
rect 178052 123486 178080 126958
rect 180064 124364 180116 124370
rect 180064 124306 180116 124312
rect 178684 124296 178736 124302
rect 178684 124238 178736 124244
rect 178040 123480 178092 123486
rect 178040 123422 178092 123428
rect 177304 118652 177356 118658
rect 177304 118594 177356 118600
rect 178696 105602 178724 124238
rect 180076 106962 180104 124306
rect 180168 121446 180196 128318
rect 181456 126274 181484 171090
rect 181548 160818 181576 195978
rect 182916 179512 182968 179518
rect 182916 179454 182968 179460
rect 181628 165640 181680 165646
rect 181628 165582 181680 165588
rect 181536 160812 181588 160818
rect 181536 160754 181588 160760
rect 181640 143546 181668 165582
rect 182824 160132 182876 160138
rect 182824 160074 182876 160080
rect 181628 143540 181680 143546
rect 181628 143482 181680 143488
rect 181444 126268 181496 126274
rect 181444 126210 181496 126216
rect 181536 125724 181588 125730
rect 181536 125666 181588 125672
rect 180156 121440 180208 121446
rect 180156 121382 180208 121388
rect 181548 108322 181576 125666
rect 181536 108316 181588 108322
rect 181536 108258 181588 108264
rect 180064 106956 180116 106962
rect 180064 106898 180116 106904
rect 178684 105596 178736 105602
rect 178684 105538 178736 105544
rect 175924 102808 175976 102814
rect 175924 102750 175976 102756
rect 182836 102134 182864 160074
rect 182928 139330 182956 179454
rect 183020 160886 183048 198698
rect 198002 198248 198058 198257
rect 198002 198183 198058 198192
rect 198016 197402 198044 198183
rect 198004 197396 198056 197402
rect 198004 197338 198056 197344
rect 198646 197160 198702 197169
rect 198646 197095 198702 197104
rect 198002 196072 198058 196081
rect 198002 196007 198004 196016
rect 198056 196007 198058 196016
rect 198004 195978 198056 195984
rect 198094 194984 198150 194993
rect 198094 194919 198150 194928
rect 198108 194614 198136 194919
rect 198096 194608 198148 194614
rect 198096 194550 198148 194556
rect 197726 193896 197782 193905
rect 197726 193831 197782 193840
rect 197740 193254 197768 193831
rect 197728 193248 197780 193254
rect 197728 193190 197780 193196
rect 197634 192808 197690 192817
rect 197634 192743 197690 192752
rect 197648 191894 197676 192743
rect 197636 191888 197688 191894
rect 197636 191830 197688 191836
rect 198094 191720 198150 191729
rect 198094 191655 198150 191664
rect 198108 191078 198136 191655
rect 191196 191072 191248 191078
rect 191196 191014 191248 191020
rect 198096 191072 198148 191078
rect 198096 191014 198148 191020
rect 188436 189168 188488 189174
rect 188436 189110 188488 189116
rect 184388 186448 184440 186454
rect 184388 186390 184440 186396
rect 184296 178152 184348 178158
rect 184296 178094 184348 178100
rect 184204 176724 184256 176730
rect 184204 176666 184256 176672
rect 183008 160880 183060 160886
rect 183008 160822 183060 160828
rect 182916 139324 182968 139330
rect 182916 139266 182968 139272
rect 184216 135182 184244 176666
rect 184308 141438 184336 178094
rect 184400 177342 184428 186390
rect 186964 185632 187016 185638
rect 186964 185574 187016 185580
rect 185584 182300 185636 182306
rect 185584 182242 185636 182248
rect 184388 177336 184440 177342
rect 184388 177278 184440 177284
rect 185596 143546 185624 182242
rect 186976 154562 187004 185574
rect 187056 173256 187108 173262
rect 187056 173198 187108 173204
rect 186964 154556 187016 154562
rect 186964 154498 187016 154504
rect 186964 150476 187016 150482
rect 186964 150418 187016 150424
rect 186320 143608 186372 143614
rect 186320 143550 186372 143556
rect 185584 143540 185636 143546
rect 185584 143482 185636 143488
rect 186332 142866 186360 143550
rect 186320 142860 186372 142866
rect 186320 142802 186372 142808
rect 184296 141432 184348 141438
rect 184296 141374 184348 141380
rect 186976 136610 187004 150418
rect 187068 150414 187096 173198
rect 188344 165708 188396 165714
rect 188344 165650 188396 165656
rect 187148 157412 187200 157418
rect 187148 157354 187200 157360
rect 187056 150408 187108 150414
rect 187056 150350 187108 150356
rect 187160 144226 187188 157354
rect 187148 144220 187200 144226
rect 187148 144162 187200 144168
rect 187056 142180 187108 142186
rect 187056 142122 187108 142128
rect 186964 136604 187016 136610
rect 186964 136546 187016 136552
rect 187068 135250 187096 142122
rect 187056 135244 187108 135250
rect 187056 135186 187108 135192
rect 184204 135176 184256 135182
rect 184204 135118 184256 135124
rect 186320 129804 186372 129810
rect 186320 129746 186372 129752
rect 184204 125656 184256 125662
rect 184204 125598 184256 125604
rect 184216 110430 184244 125598
rect 186332 125594 186360 129746
rect 186320 125588 186372 125594
rect 186320 125530 186372 125536
rect 186964 124908 187016 124914
rect 186964 124850 187016 124856
rect 186976 111790 187004 124850
rect 188356 113150 188384 165650
rect 188448 158030 188476 189110
rect 188528 177404 188580 177410
rect 188528 177346 188580 177352
rect 188436 158024 188488 158030
rect 188436 157966 188488 157972
rect 188540 148986 188568 177346
rect 189724 174548 189776 174554
rect 189724 174490 189776 174496
rect 188528 148980 188580 148986
rect 188528 148922 188580 148928
rect 189736 147626 189764 174490
rect 191104 169788 191156 169794
rect 191104 169730 191156 169736
rect 189724 147620 189776 147626
rect 189724 147562 189776 147568
rect 191116 121378 191144 169730
rect 191208 160750 191236 191014
rect 197358 190632 197414 190641
rect 197358 190567 197414 190576
rect 197372 190534 197400 190567
rect 197360 190528 197412 190534
rect 197360 190470 197412 190476
rect 197910 189544 197966 189553
rect 197910 189479 197966 189488
rect 197924 189106 197952 189479
rect 197912 189100 197964 189106
rect 197912 189042 197964 189048
rect 197358 188456 197414 188465
rect 197358 188391 197414 188400
rect 197372 187746 197400 188391
rect 197360 187740 197412 187746
rect 197360 187682 197412 187688
rect 197542 187368 197598 187377
rect 197542 187303 197598 187312
rect 197556 186386 197584 187303
rect 197544 186380 197596 186386
rect 197544 186322 197596 186328
rect 197634 186280 197690 186289
rect 195336 186244 195388 186250
rect 197634 186215 197636 186224
rect 195336 186186 195388 186192
rect 197688 186215 197690 186224
rect 197636 186186 197688 186192
rect 192484 181484 192536 181490
rect 192484 181426 192536 181432
rect 191288 176384 191340 176390
rect 191288 176326 191340 176332
rect 191196 160744 191248 160750
rect 191196 160686 191248 160692
rect 191300 149054 191328 176326
rect 192496 166326 192524 181426
rect 193864 180872 193916 180878
rect 193864 180814 193916 180820
rect 192576 169788 192628 169794
rect 192576 169730 192628 169736
rect 192484 166320 192536 166326
rect 192484 166262 192536 166268
rect 192484 164348 192536 164354
rect 192484 164290 192536 164296
rect 191380 160132 191432 160138
rect 191380 160074 191432 160080
rect 191288 149048 191340 149054
rect 191288 148990 191340 148996
rect 191392 140758 191420 160074
rect 191380 140752 191432 140758
rect 191380 140694 191432 140700
rect 191104 121372 191156 121378
rect 191104 121314 191156 121320
rect 191748 120760 191800 120766
rect 191748 120702 191800 120708
rect 191760 120018 191788 120702
rect 191748 120012 191800 120018
rect 191748 119954 191800 119960
rect 188344 113144 188396 113150
rect 188344 113086 188396 113092
rect 186964 111784 187016 111790
rect 186964 111726 187016 111732
rect 184204 110424 184256 110430
rect 184204 110366 184256 110372
rect 192496 110362 192524 164290
rect 192588 149734 192616 169730
rect 192668 153264 192720 153270
rect 192668 153206 192720 153212
rect 192576 149728 192628 149734
rect 192576 149670 192628 149676
rect 192680 137970 192708 153206
rect 193876 147762 193904 180814
rect 193956 168564 194008 168570
rect 193956 168506 194008 168512
rect 193864 147756 193916 147762
rect 193864 147698 193916 147704
rect 193968 144906 193996 168506
rect 195244 167136 195296 167142
rect 195244 167078 195296 167084
rect 193956 144900 194008 144906
rect 193956 144842 194008 144848
rect 192668 137964 192720 137970
rect 192668 137906 192720 137912
rect 195256 114918 195284 167078
rect 195348 153202 195376 186186
rect 197358 185056 197414 185065
rect 197358 184991 197414 185000
rect 197372 184210 197400 184991
rect 197360 184204 197412 184210
rect 197360 184146 197412 184152
rect 198370 183968 198426 183977
rect 198370 183903 198426 183912
rect 198384 183802 198412 183903
rect 196716 183796 196768 183802
rect 196716 183738 196768 183744
rect 198372 183796 198424 183802
rect 198372 183738 198424 183744
rect 195428 175296 195480 175302
rect 195428 175238 195480 175244
rect 195440 156942 195468 175238
rect 196624 168428 196676 168434
rect 196624 168370 196676 168376
rect 195428 156936 195480 156942
rect 195428 156878 195480 156884
rect 195520 156052 195572 156058
rect 195520 155994 195572 156000
rect 195336 153196 195388 153202
rect 195336 153138 195388 153144
rect 195532 139398 195560 155994
rect 195520 139392 195572 139398
rect 195520 139334 195572 139340
rect 196636 117230 196664 168370
rect 196728 151638 196756 183738
rect 197726 182880 197782 182889
rect 197726 182815 197782 182824
rect 197740 182238 197768 182815
rect 197728 182232 197780 182238
rect 197728 182174 197780 182180
rect 197358 181792 197414 181801
rect 197358 181727 197414 181736
rect 197372 181490 197400 181727
rect 197360 181484 197412 181490
rect 197360 181426 197412 181432
rect 198660 180794 198688 197095
rect 199396 189038 199424 199514
rect 199856 198830 199884 199543
rect 199948 198966 199976 199718
rect 203536 199714 203564 199838
rect 206744 199786 206796 199792
rect 200028 199708 200080 199714
rect 200028 199650 200080 199656
rect 203524 199708 203576 199714
rect 203524 199650 203576 199656
rect 203708 199708 203760 199714
rect 203708 199650 203760 199656
rect 199936 198960 199988 198966
rect 199936 198902 199988 198908
rect 199844 198824 199896 198830
rect 199844 198766 199896 198772
rect 200040 197826 200068 199650
rect 203720 199510 203748 199650
rect 204074 199608 204130 199617
rect 204074 199543 204130 199552
rect 207662 199608 207718 199617
rect 207662 199543 207718 199552
rect 204088 199510 204116 199543
rect 207676 199510 207704 199543
rect 210344 199510 210372 199974
rect 210424 199844 210476 199850
rect 210424 199786 210476 199792
rect 210436 199510 210464 199786
rect 210528 199510 210556 199974
rect 287612 199912 287664 199918
rect 287612 199854 287664 199860
rect 294788 199912 294840 199918
rect 294840 199860 295182 199866
rect 294788 199854 295182 199860
rect 213184 199776 213236 199782
rect 213184 199718 213236 199724
rect 244188 199776 244240 199782
rect 244188 199718 244240 199724
rect 249248 199776 249300 199782
rect 249248 199718 249300 199724
rect 211250 199608 211306 199617
rect 211250 199543 211306 199552
rect 211264 199510 211292 199543
rect 213196 199510 213224 199718
rect 213276 199708 213328 199714
rect 213276 199650 213328 199656
rect 213288 199510 213316 199650
rect 215024 199640 215076 199646
rect 215024 199582 215076 199588
rect 215036 199510 215064 199582
rect 244200 199510 244228 199718
rect 246304 199708 246356 199714
rect 246304 199650 246356 199656
rect 246210 199608 246266 199617
rect 246210 199543 246266 199552
rect 246224 199510 246252 199543
rect 246316 199510 246344 199650
rect 246486 199608 246542 199617
rect 246486 199543 246542 199552
rect 246500 199510 246528 199543
rect 249260 199510 249288 199718
rect 287072 199578 287362 199594
rect 287060 199572 287362 199578
rect 287112 199566 287362 199572
rect 287060 199514 287112 199520
rect 287624 199510 287652 199854
rect 294800 199838 295182 199854
rect 289636 199776 289688 199782
rect 293224 199776 293276 199782
rect 289688 199724 289938 199730
rect 289636 199718 289938 199724
rect 293224 199718 293276 199724
rect 287704 199708 287756 199714
rect 289648 199702 289938 199718
rect 287704 199650 287756 199656
rect 287716 199510 287744 199650
rect 291292 199640 291344 199646
rect 291344 199588 291686 199594
rect 291292 199582 291686 199588
rect 291304 199566 291686 199582
rect 293236 199510 293264 199718
rect 296628 199708 296680 199714
rect 296628 199650 296680 199656
rect 296640 199594 296668 199650
rect 296640 199566 296930 199594
rect 203708 199504 203760 199510
rect 203708 199446 203760 199452
rect 204076 199504 204128 199510
rect 204076 199446 204128 199452
rect 207664 199504 207716 199510
rect 207664 199446 207716 199452
rect 210332 199504 210384 199510
rect 210332 199446 210384 199452
rect 210424 199504 210476 199510
rect 210424 199446 210476 199452
rect 210516 199504 210568 199510
rect 211160 199504 211212 199510
rect 210516 199446 210568 199452
rect 210818 199452 211160 199458
rect 210818 199446 211212 199452
rect 211252 199504 211304 199510
rect 211252 199446 211304 199452
rect 213184 199504 213236 199510
rect 213184 199446 213236 199452
rect 213276 199504 213328 199510
rect 213276 199446 213328 199452
rect 215024 199504 215076 199510
rect 238024 199504 238076 199510
rect 215024 199446 215076 199452
rect 237774 199452 238024 199458
rect 237774 199446 238076 199452
rect 244188 199504 244240 199510
rect 244188 199446 244240 199452
rect 246212 199504 246264 199510
rect 246212 199446 246264 199452
rect 246304 199504 246356 199510
rect 246304 199446 246356 199452
rect 246488 199504 246540 199510
rect 246488 199446 246540 199452
rect 249248 199504 249300 199510
rect 249248 199446 249300 199452
rect 287612 199504 287664 199510
rect 287612 199446 287664 199452
rect 287704 199504 287756 199510
rect 287704 199446 287756 199452
rect 293224 199504 293276 199510
rect 293224 199446 293276 199452
rect 294144 199504 294196 199510
rect 294196 199452 294262 199458
rect 294144 199446 294262 199452
rect 210818 199430 211200 199446
rect 237774 199430 238064 199446
rect 294156 199430 294262 199446
rect 199948 197810 200068 197826
rect 199936 197804 200068 197810
rect 199988 197798 200068 197804
rect 199936 197746 199988 197752
rect 304276 193186 304304 200398
rect 304264 193180 304316 193186
rect 304264 193122 304316 193128
rect 580172 193180 580224 193186
rect 580172 193122 580224 193128
rect 580184 192545 580212 193122
rect 580170 192536 580226 192545
rect 580170 192471 580226 192480
rect 199384 189032 199436 189038
rect 199384 188974 199436 188980
rect 198660 180766 198872 180794
rect 197358 180704 197414 180713
rect 197358 180639 197414 180648
rect 197372 179450 197400 180639
rect 198094 179616 198150 179625
rect 198094 179551 198150 179560
rect 197360 179444 197412 179450
rect 197360 179386 197412 179392
rect 197910 178528 197966 178537
rect 197910 178463 197966 178472
rect 197924 178090 197952 178463
rect 197912 178084 197964 178090
rect 197912 178026 197964 178032
rect 197818 177440 197874 177449
rect 198108 177410 198136 179551
rect 197818 177375 197874 177384
rect 198096 177404 198148 177410
rect 197832 176390 197860 177375
rect 198096 177346 198148 177352
rect 198188 177336 198240 177342
rect 198188 177278 198240 177284
rect 197820 176384 197872 176390
rect 197358 176352 197414 176361
rect 197820 176326 197872 176332
rect 197358 176287 197414 176296
rect 197372 174554 197400 176287
rect 197360 174548 197412 174554
rect 197360 174490 197412 174496
rect 197358 174176 197414 174185
rect 197358 174111 197414 174120
rect 196808 173052 196860 173058
rect 196808 172994 196860 173000
rect 196716 151632 196768 151638
rect 196716 151574 196768 151580
rect 196820 146198 196848 172994
rect 197372 171834 197400 174111
rect 198096 173188 198148 173194
rect 198096 173130 198148 173136
rect 197360 171828 197412 171834
rect 197360 171770 197412 171776
rect 197726 170776 197782 170785
rect 197726 170711 197782 170720
rect 197740 169794 197768 170711
rect 197728 169788 197780 169794
rect 197728 169730 197780 169736
rect 197450 169688 197506 169697
rect 197450 169623 197506 169632
rect 197358 166424 197414 166433
rect 197358 166359 197414 166368
rect 197372 165646 197400 166359
rect 197360 165640 197412 165646
rect 197360 165582 197412 165588
rect 197358 164248 197414 164257
rect 197358 164183 197414 164192
rect 197372 163538 197400 164183
rect 197360 163532 197412 163538
rect 197360 163474 197412 163480
rect 197464 162178 197492 169623
rect 197726 168600 197782 168609
rect 197726 168535 197728 168544
rect 197780 168535 197782 168544
rect 197728 168506 197780 168512
rect 197910 167512 197966 167521
rect 197910 167447 197966 167456
rect 197924 167074 197952 167447
rect 197912 167068 197964 167074
rect 197912 167010 197964 167016
rect 197634 165336 197690 165345
rect 197634 165271 197690 165280
rect 197648 164286 197676 165271
rect 197636 164280 197688 164286
rect 197636 164222 197688 164228
rect 197634 163160 197690 163169
rect 197634 163095 197690 163104
rect 197648 162246 197676 163095
rect 197636 162240 197688 162246
rect 197636 162182 197688 162188
rect 197452 162172 197504 162178
rect 197452 162114 197504 162120
rect 197358 162072 197414 162081
rect 197358 162007 197414 162016
rect 197372 160138 197400 162007
rect 197360 160132 197412 160138
rect 197360 160074 197412 160080
rect 197542 159896 197598 159905
rect 197542 159831 197598 159840
rect 197556 158778 197584 159831
rect 197910 158808 197966 158817
rect 197544 158772 197596 158778
rect 197910 158743 197966 158752
rect 197544 158714 197596 158720
rect 197358 157720 197414 157729
rect 197358 157655 197414 157664
rect 197372 157418 197400 157655
rect 197360 157412 197412 157418
rect 197360 157354 197412 157360
rect 197924 156058 197952 158743
rect 198004 156936 198056 156942
rect 198004 156878 198056 156884
rect 197912 156052 197964 156058
rect 197912 155994 197964 156000
rect 197726 155408 197782 155417
rect 197726 155343 197782 155352
rect 197740 154630 197768 155343
rect 197728 154624 197780 154630
rect 197728 154566 197780 154572
rect 197360 154556 197412 154562
rect 197360 154498 197412 154504
rect 197372 154329 197400 154498
rect 197358 154320 197414 154329
rect 197358 154255 197414 154264
rect 197360 153264 197412 153270
rect 197358 153232 197360 153241
rect 197412 153232 197414 153241
rect 197358 153167 197414 153176
rect 197450 151056 197506 151065
rect 197450 150991 197506 151000
rect 197464 150482 197492 150991
rect 197452 150476 197504 150482
rect 197452 150418 197504 150424
rect 197360 150408 197412 150414
rect 197360 150350 197412 150356
rect 197372 149977 197400 150350
rect 197358 149968 197414 149977
rect 197358 149903 197414 149912
rect 197542 148880 197598 148889
rect 197542 148815 197598 148824
rect 197556 147694 197584 148815
rect 197544 147688 197596 147694
rect 197544 147630 197596 147636
rect 197360 146940 197412 146946
rect 197360 146882 197412 146888
rect 196808 146192 196860 146198
rect 196808 146134 196860 146140
rect 197372 145625 197400 146882
rect 197358 145616 197414 145625
rect 197358 145551 197414 145560
rect 197450 144528 197506 144537
rect 197450 144463 197506 144472
rect 197464 143614 197492 144463
rect 197452 143608 197504 143614
rect 197452 143550 197504 143556
rect 197360 143540 197412 143546
rect 197360 143482 197412 143488
rect 197372 143449 197400 143482
rect 197358 143440 197414 143449
rect 197358 143375 197414 143384
rect 197358 142216 197414 142225
rect 197358 142151 197360 142160
rect 197412 142151 197414 142160
rect 197360 142122 197412 142128
rect 197358 140040 197414 140049
rect 197358 139975 197414 139984
rect 197372 139466 197400 139975
rect 197360 139460 197412 139466
rect 197360 139402 197412 139408
rect 197542 137864 197598 137873
rect 197542 137799 197598 137808
rect 197556 136678 197584 137799
rect 197544 136672 197596 136678
rect 197544 136614 197596 136620
rect 197360 135176 197412 135182
rect 197360 135118 197412 135124
rect 197372 134609 197400 135118
rect 197358 134600 197414 134609
rect 197358 134535 197414 134544
rect 197450 133512 197506 133521
rect 197450 133447 197506 133456
rect 197464 132530 197492 133447
rect 197452 132524 197504 132530
rect 197452 132466 197504 132472
rect 197360 132456 197412 132462
rect 197358 132424 197360 132433
rect 197412 132424 197414 132433
rect 197358 132359 197414 132368
rect 197912 131776 197964 131782
rect 197912 131718 197964 131724
rect 197924 131345 197952 131718
rect 197910 131336 197966 131345
rect 197910 131271 197966 131280
rect 197452 130416 197504 130422
rect 197452 130358 197504 130364
rect 197360 129736 197412 129742
rect 197360 129678 197412 129684
rect 197372 129169 197400 129678
rect 197358 129160 197414 129169
rect 197358 129095 197414 129104
rect 197360 126948 197412 126954
rect 197360 126890 197412 126896
rect 197372 126857 197400 126890
rect 197358 126848 197414 126857
rect 197358 126783 197414 126792
rect 197464 125769 197492 130358
rect 198016 130257 198044 156878
rect 198108 147801 198136 173130
rect 198200 152153 198228 177278
rect 198554 175264 198610 175273
rect 198554 175199 198610 175208
rect 198568 173942 198596 175199
rect 198556 173936 198608 173942
rect 198556 173878 198608 173884
rect 198462 173088 198518 173097
rect 198462 173023 198464 173032
rect 198516 173023 198518 173032
rect 198464 172994 198516 173000
rect 198738 172000 198794 172009
rect 198738 171935 198794 171944
rect 198462 160984 198518 160993
rect 198462 160919 198518 160928
rect 198476 159390 198504 160919
rect 198464 159384 198516 159390
rect 198464 159326 198516 159332
rect 198464 158024 198516 158030
rect 198464 157966 198516 157972
rect 198476 156505 198504 157966
rect 198462 156496 198518 156505
rect 198462 156431 198518 156440
rect 198186 152144 198242 152153
rect 198186 152079 198242 152088
rect 198094 147792 198150 147801
rect 198094 147727 198150 147736
rect 198096 147688 198148 147694
rect 198096 147630 198148 147636
rect 198108 142154 198136 147630
rect 198186 146704 198242 146713
rect 198186 146639 198242 146648
rect 198200 146334 198228 146639
rect 198188 146328 198240 146334
rect 198188 146270 198240 146276
rect 198752 146266 198780 171935
rect 198740 146260 198792 146266
rect 198740 146202 198792 146208
rect 198108 142126 198228 142154
rect 198200 141137 198228 142126
rect 198464 141432 198516 141438
rect 198464 141374 198516 141380
rect 198186 141128 198242 141137
rect 198186 141063 198242 141072
rect 198188 139324 198240 139330
rect 198188 139266 198240 139272
rect 198200 138961 198228 139266
rect 198186 138952 198242 138961
rect 198186 138887 198242 138896
rect 198476 136785 198504 141374
rect 198462 136776 198518 136785
rect 198462 136711 198518 136720
rect 198186 135688 198242 135697
rect 198186 135623 198242 135632
rect 198200 135318 198228 135623
rect 198188 135312 198240 135318
rect 198188 135254 198240 135260
rect 198002 130248 198058 130257
rect 198002 130183 198058 130192
rect 198096 128308 198148 128314
rect 198096 128250 198148 128256
rect 198108 127945 198136 128250
rect 198094 127936 198150 127945
rect 198094 127871 198150 127880
rect 198004 127628 198056 127634
rect 198004 127570 198056 127576
rect 197912 126268 197964 126274
rect 197912 126210 197964 126216
rect 197450 125760 197506 125769
rect 197450 125695 197506 125704
rect 197636 125588 197688 125594
rect 197636 125530 197688 125536
rect 197648 124681 197676 125530
rect 197634 124672 197690 124681
rect 197634 124607 197690 124616
rect 197924 123593 197952 126210
rect 197910 123584 197966 123593
rect 197910 123519 197966 123528
rect 197636 123480 197688 123486
rect 197636 123422 197688 123428
rect 197360 122732 197412 122738
rect 197360 122674 197412 122680
rect 197372 122505 197400 122674
rect 197358 122496 197414 122505
rect 197358 122431 197414 122440
rect 197544 121440 197596 121446
rect 197358 121408 197414 121417
rect 197544 121382 197596 121388
rect 197358 121343 197360 121352
rect 197412 121343 197414 121352
rect 197360 121314 197412 121320
rect 197556 120329 197584 121382
rect 197542 120320 197598 120329
rect 197542 120255 197598 120264
rect 197360 118652 197412 118658
rect 197360 118594 197412 118600
rect 197372 118153 197400 118594
rect 197358 118144 197414 118153
rect 197358 118079 197414 118088
rect 196624 117224 196676 117230
rect 196624 117166 196676 117172
rect 197648 115977 197676 123422
rect 197634 115968 197690 115977
rect 197634 115903 197690 115912
rect 195244 114912 195296 114918
rect 197912 114912 197964 114918
rect 195244 114854 195296 114860
rect 197910 114880 197912 114889
rect 197964 114880 197966 114889
rect 197910 114815 197966 114824
rect 197360 114504 197412 114510
rect 197360 114446 197412 114452
rect 197372 113665 197400 114446
rect 197358 113656 197414 113665
rect 197358 113591 197414 113600
rect 197360 113144 197412 113150
rect 197360 113086 197412 113092
rect 197372 112577 197400 113086
rect 197358 112568 197414 112577
rect 197358 112503 197414 112512
rect 197360 111784 197412 111790
rect 197360 111726 197412 111732
rect 197372 111489 197400 111726
rect 197358 111480 197414 111489
rect 197358 111415 197414 111424
rect 197544 110424 197596 110430
rect 197358 110392 197414 110401
rect 192484 110356 192536 110362
rect 197544 110366 197596 110372
rect 197358 110327 197360 110336
rect 192484 110298 192536 110304
rect 197412 110327 197414 110336
rect 197360 110298 197412 110304
rect 197556 109313 197584 110366
rect 197542 109304 197598 109313
rect 197542 109239 197598 109248
rect 197544 108316 197596 108322
rect 197544 108258 197596 108264
rect 197556 107137 197584 108258
rect 198016 108225 198044 127570
rect 198844 122806 198872 180766
rect 580276 179217 580304 200738
rect 582380 198756 582432 198762
rect 582380 198698 582432 198704
rect 580262 179208 580318 179217
rect 580262 179143 580318 179152
rect 582392 165889 582420 198698
rect 582378 165880 582434 165889
rect 582378 165815 582434 165824
rect 198832 122800 198884 122806
rect 198832 122742 198884 122748
rect 198280 120012 198332 120018
rect 198280 119954 198332 119960
rect 198292 119241 198320 119954
rect 198278 119232 198334 119241
rect 198278 119167 198334 119176
rect 198464 117224 198516 117230
rect 198464 117166 198516 117172
rect 198476 117065 198504 117166
rect 198462 117056 198518 117065
rect 198462 116991 198518 117000
rect 198002 108216 198058 108225
rect 198002 108151 198058 108160
rect 197542 107128 197598 107137
rect 197542 107063 197598 107072
rect 198096 106956 198148 106962
rect 198096 106898 198148 106904
rect 197452 105596 197504 105602
rect 197452 105538 197504 105544
rect 197464 102785 197492 105538
rect 198108 104961 198136 106898
rect 198556 106276 198608 106282
rect 198556 106218 198608 106224
rect 198568 106049 198596 106218
rect 198554 106040 198610 106049
rect 198554 105975 198610 105984
rect 198094 104952 198150 104961
rect 198094 104887 198150 104896
rect 197544 104848 197596 104854
rect 197544 104790 197596 104796
rect 197556 103873 197584 104790
rect 197542 103864 197598 103873
rect 197542 103799 197598 103808
rect 198096 102808 198148 102814
rect 197450 102776 197506 102785
rect 198096 102750 198148 102756
rect 197450 102711 197506 102720
rect 182824 102128 182876 102134
rect 182824 102070 182876 102076
rect 197912 102128 197964 102134
rect 197912 102070 197964 102076
rect 197924 101697 197952 102070
rect 197910 101688 197966 101697
rect 197910 101623 197966 101632
rect 198108 100609 198136 102750
rect 199934 101008 199990 101017
rect 199934 100943 199990 100952
rect 199948 100706 199976 100943
rect 568580 100768 568632 100774
rect 298558 100736 298614 100745
rect 200592 100706 200698 100722
rect 202248 100706 202354 100722
rect 199936 100700 199988 100706
rect 199936 100642 199988 100648
rect 200580 100700 200698 100706
rect 200632 100694 200698 100700
rect 202236 100700 202354 100706
rect 200580 100642 200632 100648
rect 202288 100694 202354 100700
rect 295458 100706 295564 100722
rect 295458 100700 295576 100706
rect 295458 100694 295524 100700
rect 202236 100642 202288 100648
rect 298494 100694 298558 100722
rect 568580 100710 568632 100716
rect 298558 100671 298614 100680
rect 295524 100642 295576 100648
rect 198094 100600 198150 100609
rect 198094 100535 198150 100544
rect 297914 100464 297970 100473
rect 297850 100422 297914 100450
rect 297914 100399 297970 100408
rect 297914 100328 297970 100337
rect 297970 100286 298034 100314
rect 297914 100263 297970 100272
rect 211724 100162 211830 100178
rect 211528 100156 211580 100162
rect 211528 100098 211580 100104
rect 211712 100156 211830 100162
rect 211764 100150 211830 100156
rect 211712 100098 211764 100104
rect 147588 99816 147640 99822
rect 147588 99758 147640 99764
rect 144828 98048 144880 98054
rect 144828 97990 144880 97996
rect 143448 94648 143500 94654
rect 143448 94590 143500 94596
rect 142068 93288 142120 93294
rect 142068 93230 142120 93236
rect 140044 59356 140096 59362
rect 140044 59298 140096 59304
rect 142080 3602 142108 93230
rect 138848 3596 138900 3602
rect 138848 3538 138900 3544
rect 139308 3596 139360 3602
rect 139308 3538 139360 3544
rect 141240 3596 141292 3602
rect 141240 3538 141292 3544
rect 142068 3596 142120 3602
rect 142068 3538 142120 3544
rect 138860 480 138888 3538
rect 140044 2236 140096 2242
rect 140044 2178 140096 2184
rect 140056 480 140084 2178
rect 141252 480 141280 3538
rect 143460 2922 143488 94590
rect 144736 76832 144788 76838
rect 144736 76774 144788 76780
rect 143540 3596 143592 3602
rect 143540 3538 143592 3544
rect 142436 2916 142488 2922
rect 142436 2858 142488 2864
rect 143448 2916 143500 2922
rect 143448 2858 143500 2864
rect 142448 480 142476 2858
rect 143552 480 143580 3538
rect 144748 480 144776 76774
rect 144840 3602 144868 97990
rect 145932 3664 145984 3670
rect 145932 3606 145984 3612
rect 144828 3596 144880 3602
rect 144828 3538 144880 3544
rect 145944 480 145972 3606
rect 147600 3194 147628 99758
rect 156604 99680 156656 99686
rect 156604 99622 156656 99628
rect 155868 99612 155920 99618
rect 155868 99554 155920 99560
rect 153106 94480 153162 94489
rect 153106 94415 153162 94424
rect 148968 93356 149020 93362
rect 148968 93298 149020 93304
rect 148980 3602 149008 93298
rect 153016 76900 153068 76906
rect 153016 76842 153068 76848
rect 149520 3664 149572 3670
rect 149520 3606 149572 3612
rect 148324 3596 148376 3602
rect 148324 3538 148376 3544
rect 148968 3596 149020 3602
rect 148968 3538 149020 3544
rect 147128 3188 147180 3194
rect 147128 3130 147180 3136
rect 147588 3188 147640 3194
rect 147588 3130 147640 3136
rect 147140 480 147168 3130
rect 148336 480 148364 3538
rect 149532 480 149560 3606
rect 151820 3324 151872 3330
rect 151820 3266 151872 3272
rect 150624 2304 150676 2310
rect 150624 2246 150676 2252
rect 150636 480 150664 2246
rect 151832 480 151860 3266
rect 153028 480 153056 76842
rect 153120 3398 153148 94415
rect 155880 3398 155908 99554
rect 153108 3392 153160 3398
rect 153108 3334 153160 3340
rect 154212 3392 154264 3398
rect 154212 3334 154264 3340
rect 155408 3392 155460 3398
rect 155408 3334 155460 3340
rect 155868 3392 155920 3398
rect 155868 3334 155920 3340
rect 154224 480 154252 3334
rect 155420 480 155448 3334
rect 156616 3330 156644 99622
rect 197268 98932 197320 98938
rect 197268 98874 197320 98880
rect 180064 98864 180116 98870
rect 180064 98806 180116 98812
rect 173164 98796 173216 98802
rect 173164 98738 173216 98744
rect 162124 98728 162176 98734
rect 162124 98670 162176 98676
rect 159364 96008 159416 96014
rect 159364 95950 159416 95956
rect 158628 94716 158680 94722
rect 158628 94658 158680 94664
rect 158640 3398 158668 94658
rect 158904 3800 158956 3806
rect 158904 3742 158956 3748
rect 157800 3392 157852 3398
rect 157800 3334 157852 3340
rect 158628 3392 158680 3398
rect 158628 3334 158680 3340
rect 156604 3324 156656 3330
rect 156604 3266 156656 3272
rect 156696 3324 156748 3330
rect 156696 3266 156748 3272
rect 156708 1714 156736 3266
rect 156616 1686 156736 1714
rect 156616 480 156644 1686
rect 157812 480 157840 3334
rect 158916 480 158944 3742
rect 159376 3738 159404 95950
rect 161388 80844 161440 80850
rect 161388 80786 161440 80792
rect 161296 4140 161348 4146
rect 161296 4082 161348 4088
rect 159364 3732 159416 3738
rect 159364 3674 159416 3680
rect 160100 3188 160152 3194
rect 160100 3130 160152 3136
rect 160112 480 160140 3130
rect 161308 480 161336 4082
rect 161400 3194 161428 80786
rect 162136 4146 162164 98670
rect 165528 98116 165580 98122
rect 165528 98058 165580 98064
rect 162216 90704 162268 90710
rect 162216 90646 162268 90652
rect 162124 4140 162176 4146
rect 162124 4082 162176 4088
rect 162228 3330 162256 90646
rect 164148 80912 164200 80918
rect 164148 80854 164200 80860
rect 162492 3732 162544 3738
rect 162492 3674 162544 3680
rect 162216 3324 162268 3330
rect 162216 3266 162268 3272
rect 161388 3188 161440 3194
rect 161388 3130 161440 3136
rect 162504 480 162532 3674
rect 164160 3398 164188 80854
rect 165540 3398 165568 98058
rect 166908 94784 166960 94790
rect 166908 94726 166960 94732
rect 166920 3398 166948 94726
rect 169666 94616 169722 94625
rect 169666 94551 169722 94560
rect 168288 82408 168340 82414
rect 168288 82350 168340 82356
rect 168300 3398 168328 82350
rect 169680 6914 169708 94551
rect 171048 92132 171100 92138
rect 171048 92074 171100 92080
rect 170404 82340 170456 82346
rect 170404 82282 170456 82288
rect 169588 6886 169708 6914
rect 168380 4140 168432 4146
rect 168380 4082 168432 4088
rect 163688 3392 163740 3398
rect 163688 3334 163740 3340
rect 164148 3392 164200 3398
rect 164148 3334 164200 3340
rect 164884 3392 164936 3398
rect 164884 3334 164936 3340
rect 165528 3392 165580 3398
rect 165528 3334 165580 3340
rect 166080 3392 166132 3398
rect 166080 3334 166132 3340
rect 166908 3392 166960 3398
rect 166908 3334 166960 3340
rect 167184 3392 167236 3398
rect 167184 3334 167236 3340
rect 168288 3392 168340 3398
rect 168288 3334 168340 3340
rect 163700 480 163728 3334
rect 164896 480 164924 3334
rect 166092 480 166120 3334
rect 167196 480 167224 3334
rect 168392 480 168420 4082
rect 169588 480 169616 6886
rect 170416 3806 170444 82282
rect 171060 6914 171088 92074
rect 172428 76968 172480 76974
rect 172428 76910 172480 76916
rect 170784 6886 171088 6914
rect 170404 3800 170456 3806
rect 170404 3742 170456 3748
rect 170784 480 170812 6886
rect 171784 4004 171836 4010
rect 171784 3946 171836 3952
rect 171796 3670 171824 3946
rect 171876 3936 171928 3942
rect 171876 3878 171928 3884
rect 171784 3664 171836 3670
rect 171784 3606 171836 3612
rect 171888 3602 171916 3878
rect 172440 3602 172468 76910
rect 173176 4146 173204 98738
rect 178684 96144 178736 96150
rect 178684 96086 178736 96092
rect 177946 91896 178002 91905
rect 177946 91831 178002 91840
rect 177304 89344 177356 89350
rect 177304 89286 177356 89292
rect 175188 82476 175240 82482
rect 175188 82418 175240 82424
rect 173164 4140 173216 4146
rect 173164 4082 173216 4088
rect 173164 3800 173216 3806
rect 173164 3742 173216 3748
rect 171876 3596 171928 3602
rect 171876 3538 171928 3544
rect 171968 3596 172020 3602
rect 171968 3538 172020 3544
rect 172428 3596 172480 3602
rect 172428 3538 172480 3544
rect 171980 480 172008 3538
rect 173176 480 173204 3742
rect 175200 3534 175228 82418
rect 174268 3528 174320 3534
rect 174268 3470 174320 3476
rect 175188 3528 175240 3534
rect 175188 3470 175240 3476
rect 174280 480 174308 3470
rect 176660 3052 176712 3058
rect 176660 2994 176712 3000
rect 175464 2984 175516 2990
rect 175464 2926 175516 2932
rect 175476 480 175504 2926
rect 176672 480 176700 2994
rect 177316 2990 177344 89286
rect 177960 6914 177988 91831
rect 177868 6886 177988 6914
rect 177304 2984 177356 2990
rect 177304 2926 177356 2932
rect 177868 480 177896 6886
rect 178696 3602 178724 96086
rect 178776 89412 178828 89418
rect 178776 89354 178828 89360
rect 178684 3596 178736 3602
rect 178684 3538 178736 3544
rect 178788 3058 178816 89354
rect 180076 3534 180104 98806
rect 195336 97912 195388 97918
rect 195336 97854 195388 97860
rect 188342 97336 188398 97345
rect 188342 97271 188398 97280
rect 186962 96112 187018 96121
rect 183468 96076 183520 96082
rect 186962 96047 187018 96056
rect 183468 96018 183520 96024
rect 181444 94852 181496 94858
rect 181444 94794 181496 94800
rect 181456 3738 181484 94794
rect 181536 90772 181588 90778
rect 181536 90714 181588 90720
rect 181548 4010 181576 90714
rect 182824 83768 182876 83774
rect 182824 83710 182876 83716
rect 181536 4004 181588 4010
rect 181536 3946 181588 3952
rect 182836 3942 182864 83710
rect 182824 3936 182876 3942
rect 182824 3878 182876 3884
rect 181444 3732 181496 3738
rect 181444 3674 181496 3680
rect 183480 3534 183508 96018
rect 184848 93424 184900 93430
rect 184848 93366 184900 93372
rect 184204 85128 184256 85134
rect 184204 85070 184256 85076
rect 179052 3528 179104 3534
rect 179052 3470 179104 3476
rect 180064 3528 180116 3534
rect 180064 3470 180116 3476
rect 180248 3528 180300 3534
rect 180248 3470 180300 3476
rect 182548 3528 182600 3534
rect 182548 3470 182600 3476
rect 183468 3528 183520 3534
rect 183468 3470 183520 3476
rect 183744 3528 183796 3534
rect 183744 3470 183796 3476
rect 178776 3052 178828 3058
rect 178776 2994 178828 3000
rect 179064 480 179092 3470
rect 180260 480 180288 3470
rect 181444 3392 181496 3398
rect 181444 3334 181496 3340
rect 181456 480 181484 3334
rect 182560 480 182588 3470
rect 183756 480 183784 3470
rect 184216 3398 184244 85070
rect 184860 3534 184888 93366
rect 186228 92200 186280 92206
rect 186228 92142 186280 92148
rect 186240 3534 186268 92142
rect 184848 3528 184900 3534
rect 184848 3470 184900 3476
rect 184940 3528 184992 3534
rect 184940 3470 184992 3476
rect 186228 3528 186280 3534
rect 186228 3470 186280 3476
rect 184204 3392 184256 3398
rect 184204 3334 184256 3340
rect 184952 480 184980 3470
rect 186976 2922 187004 96047
rect 188356 91798 188384 97271
rect 192484 96212 192536 96218
rect 192484 96154 192536 96160
rect 191748 93492 191800 93498
rect 191748 93434 191800 93440
rect 188344 91792 188396 91798
rect 188344 91734 188396 91740
rect 188988 91792 189040 91798
rect 188988 91734 189040 91740
rect 188342 86184 188398 86193
rect 188342 86119 188398 86128
rect 187056 85196 187108 85202
rect 187056 85138 187108 85144
rect 187068 3806 187096 85138
rect 187056 3800 187108 3806
rect 187056 3742 187108 3748
rect 188356 3534 188384 86119
rect 189000 3534 189028 91734
rect 191656 83836 191708 83842
rect 191656 83778 191708 83784
rect 190368 82544 190420 82550
rect 190368 82486 190420 82492
rect 189724 3868 189776 3874
rect 189724 3810 189776 3816
rect 187332 3528 187384 3534
rect 187332 3470 187384 3476
rect 188344 3528 188396 3534
rect 188344 3470 188396 3476
rect 188528 3528 188580 3534
rect 188528 3470 188580 3476
rect 188988 3528 189040 3534
rect 188988 3470 189040 3476
rect 186136 2916 186188 2922
rect 186136 2858 186188 2864
rect 186964 2916 187016 2922
rect 186964 2858 187016 2864
rect 186148 480 186176 2858
rect 187344 480 187372 3470
rect 188540 480 188568 3470
rect 189736 480 189764 3810
rect 190380 3806 190408 82486
rect 191668 16574 191696 83778
rect 191576 16546 191696 16574
rect 190368 3800 190420 3806
rect 190368 3742 190420 3748
rect 190828 3528 190880 3534
rect 190828 3470 190880 3476
rect 190840 480 190868 3470
rect 191576 3058 191604 16546
rect 191760 6914 191788 93434
rect 191668 6886 191788 6914
rect 191668 3534 191696 6886
rect 192496 3874 192524 96154
rect 195242 94752 195298 94761
rect 195242 94687 195298 94696
rect 194506 90400 194562 90409
rect 194506 90335 194562 90344
rect 193128 87984 193180 87990
rect 193128 87926 193180 87932
rect 192484 3868 192536 3874
rect 192484 3810 192536 3816
rect 193140 3670 193168 87926
rect 194520 6914 194548 90335
rect 194428 6886 194548 6914
rect 193220 4004 193272 4010
rect 193220 3946 193272 3952
rect 193128 3664 193180 3670
rect 193128 3606 193180 3612
rect 191656 3528 191708 3534
rect 191656 3470 191708 3476
rect 191564 3052 191616 3058
rect 191564 2994 191616 3000
rect 192024 3052 192076 3058
rect 192024 2994 192076 3000
rect 192036 480 192064 2994
rect 193232 480 193260 3946
rect 194428 480 194456 6886
rect 195256 3602 195284 94687
rect 195348 91866 195376 97854
rect 195336 91860 195388 91866
rect 195336 91802 195388 91808
rect 195888 91860 195940 91866
rect 195888 91802 195940 91808
rect 195900 6914 195928 91802
rect 197176 88052 197228 88058
rect 197176 87994 197228 88000
rect 195624 6886 195928 6914
rect 195244 3596 195296 3602
rect 195244 3538 195296 3544
rect 195624 480 195652 6886
rect 196820 598 197032 626
rect 196820 480 196848 598
rect 197004 490 197032 598
rect 197188 490 197216 87994
rect 197280 3670 197308 98874
rect 200132 97345 200160 100028
rect 200316 98666 200344 100028
rect 200304 98660 200356 98666
rect 200304 98602 200356 98608
rect 200118 97336 200174 97345
rect 200118 97271 200174 97280
rect 199384 96688 199436 96694
rect 199384 96630 199436 96636
rect 198648 93560 198700 93566
rect 198648 93502 198700 93508
rect 197268 3664 197320 3670
rect 197268 3606 197320 3612
rect 198660 3534 198688 93502
rect 199396 24138 199424 96630
rect 200028 96280 200080 96286
rect 200028 96222 200080 96228
rect 199384 24132 199436 24138
rect 199384 24074 199436 24080
rect 200040 3806 200068 96222
rect 200500 95946 200528 100028
rect 200868 97209 200896 100028
rect 201052 100014 201158 100042
rect 201236 100014 201342 100042
rect 200854 97200 200910 97209
rect 200854 97135 200910 97144
rect 200762 96792 200818 96801
rect 200762 96727 200818 96736
rect 200488 95940 200540 95946
rect 200488 95882 200540 95888
rect 200396 94512 200448 94518
rect 200396 94454 200448 94460
rect 199108 3800 199160 3806
rect 199108 3742 199160 3748
rect 200028 3800 200080 3806
rect 200028 3742 200080 3748
rect 197912 3528 197964 3534
rect 197912 3470 197964 3476
rect 198648 3528 198700 3534
rect 198648 3470 198700 3476
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197004 462 197216 490
rect 197924 480 197952 3470
rect 199120 480 199148 3742
rect 200304 3528 200356 3534
rect 200304 3470 200356 3476
rect 200316 480 200344 3470
rect 200408 2106 200436 94454
rect 200776 51746 200804 96727
rect 200946 96656 201002 96665
rect 200946 96591 201002 96600
rect 200960 76566 200988 96591
rect 200948 76560 201000 76566
rect 200948 76502 201000 76508
rect 201052 68338 201080 100014
rect 201236 94518 201264 100014
rect 201408 98660 201460 98666
rect 201408 98602 201460 98608
rect 201224 94512 201276 94518
rect 201224 94454 201276 94460
rect 201040 68332 201092 68338
rect 201040 68274 201092 68280
rect 200764 51740 200816 51746
rect 200764 51682 200816 51688
rect 201420 3534 201448 98602
rect 201512 95849 201540 100028
rect 201498 95840 201554 95849
rect 201498 95775 201554 95784
rect 201592 94920 201644 94926
rect 201592 94862 201644 94868
rect 201604 84862 201632 94862
rect 201696 86290 201724 100028
rect 201880 96694 201908 100028
rect 202156 97918 202184 100028
rect 202432 100014 202538 100042
rect 202616 100014 202722 100042
rect 202144 97912 202196 97918
rect 202144 97854 202196 97860
rect 202144 97640 202196 97646
rect 202144 97582 202196 97588
rect 201960 96960 202012 96966
rect 201960 96902 202012 96908
rect 201868 96688 201920 96694
rect 201868 96630 201920 96636
rect 201684 86284 201736 86290
rect 201684 86226 201736 86232
rect 201592 84856 201644 84862
rect 201592 84798 201644 84804
rect 201408 3528 201460 3534
rect 201408 3470 201460 3476
rect 201500 3528 201552 3534
rect 201972 3505 202000 96902
rect 201500 3470 201552 3476
rect 201958 3496 202014 3505
rect 200396 2100 200448 2106
rect 200396 2042 200448 2048
rect 201512 480 201540 3470
rect 201958 3431 202014 3440
rect 202156 2242 202184 97582
rect 202432 94926 202460 100014
rect 202616 96966 202644 100014
rect 202604 96960 202656 96966
rect 202604 96902 202656 96908
rect 202604 96824 202656 96830
rect 202604 96766 202656 96772
rect 202420 94920 202472 94926
rect 202420 94862 202472 94868
rect 202616 89714 202644 96766
rect 202892 96665 202920 100028
rect 203168 96937 203196 100028
rect 203154 96928 203210 96937
rect 203154 96863 203210 96872
rect 202878 96656 202934 96665
rect 202878 96591 202934 96600
rect 203352 94926 203380 100028
rect 203444 100014 203550 100042
rect 203628 100014 203734 100042
rect 203812 100014 203918 100042
rect 203340 94920 203392 94926
rect 203340 94862 203392 94868
rect 203444 91746 203472 100014
rect 203524 94920 203576 94926
rect 203524 94862 203576 94868
rect 202340 89686 202644 89714
rect 203260 91718 203472 91746
rect 202236 84856 202288 84862
rect 202236 84798 202288 84804
rect 202248 4010 202276 84798
rect 202340 73914 202368 89686
rect 202328 73908 202380 73914
rect 202328 73850 202380 73856
rect 202236 4004 202288 4010
rect 202236 3946 202288 3952
rect 203260 3466 203288 91718
rect 203536 86954 203564 94862
rect 203628 93158 203656 100014
rect 203616 93152 203668 93158
rect 203616 93094 203668 93100
rect 203812 91934 203840 100014
rect 204180 94450 204208 100028
rect 204260 96892 204312 96898
rect 204260 96834 204312 96840
rect 204168 94444 204220 94450
rect 204168 94386 204220 94392
rect 203800 91928 203852 91934
rect 203800 91870 203852 91876
rect 204272 90438 204300 96834
rect 204364 96665 204392 100028
rect 204350 96656 204406 96665
rect 204350 96591 204406 96600
rect 204444 94512 204496 94518
rect 204444 94454 204496 94460
rect 204260 90432 204312 90438
rect 204260 90374 204312 90380
rect 203352 86926 203564 86954
rect 203352 68406 203380 86926
rect 204456 82113 204484 94454
rect 204548 87553 204576 100028
rect 204640 100014 204746 100042
rect 204640 94518 204668 100014
rect 204916 97306 204944 100028
rect 205192 98705 205220 100028
rect 205284 100014 205390 100042
rect 205468 100014 205574 100042
rect 205178 98696 205234 98705
rect 205178 98631 205234 98640
rect 204904 97300 204956 97306
rect 204904 97242 204956 97248
rect 204628 94512 204680 94518
rect 204628 94454 204680 94460
rect 204628 94376 204680 94382
rect 204628 94318 204680 94324
rect 204534 87544 204590 87553
rect 204534 87479 204590 87488
rect 204442 82104 204498 82113
rect 204442 82039 204498 82048
rect 203340 68400 203392 68406
rect 203340 68342 203392 68348
rect 204640 18630 204668 94318
rect 205284 84194 205312 100014
rect 205468 94382 205496 100014
rect 205744 96665 205772 100028
rect 205928 96937 205956 100028
rect 206204 97578 206232 100028
rect 206296 100014 206402 100042
rect 206480 100014 206586 100042
rect 206664 100014 206770 100042
rect 206848 100014 206954 100042
rect 207124 100014 207230 100042
rect 206192 97572 206244 97578
rect 206192 97514 206244 97520
rect 205914 96928 205970 96937
rect 205914 96863 205970 96872
rect 205730 96656 205786 96665
rect 205730 96591 205786 96600
rect 206296 94738 206324 100014
rect 206480 99374 206508 100014
rect 205928 94710 206324 94738
rect 206388 99346 206508 99374
rect 205456 94376 205508 94382
rect 205456 94318 205508 94324
rect 205928 93226 205956 94710
rect 206388 94602 206416 99346
rect 206468 97572 206520 97578
rect 206468 97514 206520 97520
rect 206020 94574 206416 94602
rect 205916 93220 205968 93226
rect 205916 93162 205968 93168
rect 205100 84166 205312 84194
rect 205100 73846 205128 84166
rect 205088 73840 205140 73846
rect 205088 73782 205140 73788
rect 206020 71058 206048 94574
rect 206480 89714 206508 97514
rect 206664 97374 206692 100014
rect 206652 97368 206704 97374
rect 206652 97310 206704 97316
rect 206296 89686 206508 89714
rect 206296 89010 206324 89686
rect 206284 89004 206336 89010
rect 206284 88946 206336 88952
rect 206848 84194 206876 100014
rect 206928 96688 206980 96694
rect 206928 96630 206980 96636
rect 206940 90506 206968 96630
rect 206928 90500 206980 90506
rect 206928 90442 206980 90448
rect 206664 84166 206876 84194
rect 206664 82142 206692 84166
rect 206652 82136 206704 82142
rect 206652 82078 206704 82084
rect 207124 77994 207152 100014
rect 207400 96801 207428 100028
rect 207492 100014 207598 100042
rect 207492 97492 207520 100014
rect 207492 97464 207612 97492
rect 207480 97300 207532 97306
rect 207480 97242 207532 97248
rect 207386 96792 207442 96801
rect 207386 96727 207442 96736
rect 207492 84194 207520 97242
rect 207584 87650 207612 97464
rect 207664 97368 207716 97374
rect 207664 97310 207716 97316
rect 207572 87644 207624 87650
rect 207572 87586 207624 87592
rect 207308 84166 207520 84194
rect 207112 77988 207164 77994
rect 207112 77930 207164 77936
rect 207308 71126 207336 84166
rect 207296 71120 207348 71126
rect 207296 71062 207348 71068
rect 206008 71052 206060 71058
rect 206008 70994 206060 71000
rect 204628 18624 204680 18630
rect 204628 18566 204680 18572
rect 203892 3800 203944 3806
rect 203892 3742 203944 3748
rect 203248 3460 203300 3466
rect 203248 3402 203300 3408
rect 202694 3360 202750 3369
rect 202694 3295 202750 3304
rect 202144 2236 202196 2242
rect 202144 2178 202196 2184
rect 202708 480 202736 3295
rect 203904 480 203932 3742
rect 207388 3664 207440 3670
rect 207388 3606 207440 3612
rect 205088 3596 205140 3602
rect 205088 3538 205140 3544
rect 205100 480 205128 3538
rect 206192 2100 206244 2106
rect 206192 2042 206244 2048
rect 206204 480 206232 2042
rect 207400 480 207428 3606
rect 207676 2310 207704 97310
rect 207768 97306 207796 100028
rect 207952 97442 207980 100028
rect 207940 97436 207992 97442
rect 207940 97378 207992 97384
rect 207756 97300 207808 97306
rect 207756 97242 207808 97248
rect 207756 96960 207808 96966
rect 207756 96902 207808 96908
rect 207768 89049 207796 96902
rect 208228 96830 208256 100028
rect 208216 96824 208268 96830
rect 208216 96766 208268 96772
rect 208412 96665 208440 100028
rect 208398 96656 208454 96665
rect 208398 96591 208454 96600
rect 208492 94512 208544 94518
rect 208492 94454 208544 94460
rect 207754 89040 207810 89049
rect 207754 88975 207810 88984
rect 208504 79422 208532 94454
rect 208596 84930 208624 100028
rect 208780 98841 208808 100028
rect 208872 100014 209070 100042
rect 209148 100014 209254 100042
rect 208766 98832 208822 98841
rect 208766 98767 208822 98776
rect 208872 94602 208900 100014
rect 208688 94574 208900 94602
rect 208688 87718 208716 94574
rect 209148 89714 209176 100014
rect 209424 96898 209452 100028
rect 209516 100014 209622 100042
rect 209412 96892 209464 96898
rect 209412 96834 209464 96840
rect 209228 96824 209280 96830
rect 209228 96766 209280 96772
rect 208872 89686 209176 89714
rect 208676 87712 208728 87718
rect 208676 87654 208728 87660
rect 208584 84924 208636 84930
rect 208584 84866 208636 84872
rect 208492 79416 208544 79422
rect 208492 79358 208544 79364
rect 208872 71194 208900 89686
rect 209240 84194 209268 96766
rect 209516 94518 209544 100014
rect 209792 96665 209820 100028
rect 209884 100014 210082 100042
rect 209778 96656 209834 96665
rect 209778 96591 209834 96600
rect 209884 94602 209912 100014
rect 210252 97510 210280 100028
rect 210344 100014 210450 100042
rect 210240 97504 210292 97510
rect 210240 97446 210292 97452
rect 210344 94602 210372 100014
rect 210620 96694 210648 100028
rect 210712 100014 210818 100042
rect 210896 100014 211094 100042
rect 210608 96688 210660 96694
rect 210608 96630 210660 96636
rect 209792 94574 209912 94602
rect 209976 94574 210372 94602
rect 209504 94512 209556 94518
rect 209504 94454 209556 94460
rect 209792 90370 209820 94574
rect 209872 94512 209924 94518
rect 209872 94454 209924 94460
rect 209780 90364 209832 90370
rect 209780 90306 209832 90312
rect 209056 84166 209268 84194
rect 208860 71188 208912 71194
rect 208860 71130 208912 71136
rect 209056 4826 209084 84166
rect 209884 71330 209912 94454
rect 209872 71324 209924 71330
rect 209872 71266 209924 71272
rect 209976 71262 210004 94574
rect 210712 94466 210740 100014
rect 210792 96688 210844 96694
rect 210792 96630 210844 96636
rect 210160 94438 210740 94466
rect 209964 71256 210016 71262
rect 209964 71198 210016 71204
rect 209044 4820 209096 4826
rect 209044 4762 209096 4768
rect 208584 4004 208636 4010
rect 208584 3946 208636 3952
rect 207664 2304 207716 2310
rect 207664 2246 207716 2252
rect 208596 480 208624 3946
rect 209780 3256 209832 3262
rect 209780 3198 209832 3204
rect 209792 480 209820 3198
rect 210160 2174 210188 94438
rect 210804 89714 210832 96630
rect 210896 94518 210924 100014
rect 211264 99414 211292 100028
rect 211252 99408 211304 99414
rect 211252 99350 211304 99356
rect 211448 96665 211476 100028
rect 211434 96656 211490 96665
rect 211434 96591 211490 96600
rect 211540 94602 211568 100098
rect 211646 100014 211752 100042
rect 211724 98274 211752 100014
rect 211724 98246 211936 98274
rect 211804 96756 211856 96762
rect 211804 96698 211856 96704
rect 211448 94574 211568 94602
rect 210884 94512 210936 94518
rect 210884 94454 210936 94460
rect 211448 92002 211476 94574
rect 211528 94512 211580 94518
rect 211528 94454 211580 94460
rect 211436 91996 211488 92002
rect 211436 91938 211488 91944
rect 210436 89686 210832 89714
rect 210436 87786 210464 89686
rect 210424 87780 210476 87786
rect 210424 87722 210476 87728
rect 211540 47598 211568 94454
rect 211816 86358 211844 96698
rect 211804 86352 211856 86358
rect 211804 86294 211856 86300
rect 211908 84998 211936 98246
rect 212092 96694 212120 100028
rect 212184 100014 212290 100042
rect 212368 100014 212474 100042
rect 212080 96688 212132 96694
rect 212080 96630 212132 96636
rect 212184 94518 212212 100014
rect 212172 94512 212224 94518
rect 212172 94454 212224 94460
rect 212368 90574 212396 100014
rect 212644 96665 212672 100028
rect 212630 96656 212686 96665
rect 212630 96591 212686 96600
rect 212724 94920 212776 94926
rect 212724 94862 212776 94868
rect 212356 90568 212408 90574
rect 212356 90510 212408 90516
rect 212736 87854 212764 94862
rect 212724 87848 212776 87854
rect 212724 87790 212776 87796
rect 211896 84992 211948 84998
rect 211896 84934 211948 84940
rect 212828 79354 212856 100028
rect 213104 99482 213132 100028
rect 213196 100014 213302 100042
rect 213380 100014 213486 100042
rect 213092 99476 213144 99482
rect 213092 99418 213144 99424
rect 213196 94926 213224 100014
rect 213380 99374 213408 100014
rect 213288 99346 213408 99374
rect 213184 94920 213236 94926
rect 213184 94862 213236 94868
rect 213288 94602 213316 99346
rect 213656 96966 213684 100028
rect 213736 97300 213788 97306
rect 213736 97242 213788 97248
rect 213644 96960 213696 96966
rect 213644 96902 213696 96908
rect 213368 96688 213420 96694
rect 213368 96630 213420 96636
rect 212920 94574 213316 94602
rect 212816 79348 212868 79354
rect 212816 79290 212868 79296
rect 211528 47592 211580 47598
rect 211528 47534 211580 47540
rect 212920 43450 212948 94574
rect 213380 89714 213408 96630
rect 213196 89686 213408 89714
rect 213748 89714 213776 97242
rect 213840 96830 213868 100028
rect 213828 96824 213880 96830
rect 213828 96766 213880 96772
rect 214116 96665 214144 100028
rect 214102 96656 214158 96665
rect 214102 96591 214158 96600
rect 214012 94512 214064 94518
rect 214012 94454 214064 94460
rect 213748 89686 213868 89714
rect 213196 83502 213224 89686
rect 213184 83496 213236 83502
rect 213184 83438 213236 83444
rect 212908 43444 212960 43450
rect 212908 43386 212960 43392
rect 213184 43444 213236 43450
rect 213184 43386 213236 43392
rect 211804 35216 211856 35222
rect 211804 35158 211856 35164
rect 210976 8968 211028 8974
rect 210976 8910 211028 8916
rect 210148 2168 210200 2174
rect 210148 2110 210200 2116
rect 210988 480 211016 8910
rect 211816 4010 211844 35158
rect 211804 4004 211856 4010
rect 211804 3946 211856 3952
rect 212172 3392 212224 3398
rect 212172 3334 212224 3340
rect 212184 480 212212 3334
rect 213196 3262 213224 43386
rect 213840 11778 213868 89686
rect 214024 73982 214052 94454
rect 214196 94444 214248 94450
rect 214196 94386 214248 94392
rect 214208 89214 214236 94386
rect 214300 89282 214328 100028
rect 214392 100014 214498 100042
rect 214682 100014 214788 100042
rect 214392 94518 214420 100014
rect 214564 97028 214616 97034
rect 214564 96970 214616 96976
rect 214380 94512 214432 94518
rect 214380 94454 214432 94460
rect 214288 89276 214340 89282
rect 214288 89218 214340 89224
rect 214196 89208 214248 89214
rect 214196 89150 214248 89156
rect 214576 82210 214604 96970
rect 214564 82204 214616 82210
rect 214564 82146 214616 82152
rect 214012 73976 214064 73982
rect 214012 73918 214064 73924
rect 214760 15910 214788 100014
rect 214852 94450 214880 100028
rect 215128 96762 215156 100028
rect 215326 100014 215432 100042
rect 215300 98116 215352 98122
rect 215300 98058 215352 98064
rect 215312 97850 215340 98058
rect 215300 97844 215352 97850
rect 215300 97786 215352 97792
rect 215404 97050 215432 100014
rect 215496 97578 215524 100028
rect 215484 97572 215536 97578
rect 215484 97514 215536 97520
rect 215312 97022 215432 97050
rect 215312 96830 215340 97022
rect 215392 96960 215444 96966
rect 215680 96937 215708 100028
rect 215772 100014 215878 100042
rect 215956 100014 216154 100042
rect 216232 100014 216338 100042
rect 216416 100014 216522 100042
rect 215392 96902 215444 96908
rect 215666 96928 215722 96937
rect 215300 96824 215352 96830
rect 215300 96766 215352 96772
rect 215116 96756 215168 96762
rect 215116 96698 215168 96704
rect 214840 94444 214892 94450
rect 214840 94386 214892 94392
rect 215404 80714 215432 96902
rect 215666 96863 215722 96872
rect 215576 95464 215628 95470
rect 215576 95406 215628 95412
rect 215588 87922 215616 95406
rect 215576 87916 215628 87922
rect 215576 87858 215628 87864
rect 215392 80708 215444 80714
rect 215392 80650 215444 80656
rect 214748 15904 214800 15910
rect 214748 15846 214800 15852
rect 215772 13122 215800 100014
rect 215956 96966 215984 100014
rect 215944 96960 215996 96966
rect 215944 96902 215996 96908
rect 215944 96824 215996 96830
rect 215944 96766 215996 96772
rect 215956 74050 215984 96766
rect 216232 95470 216260 100014
rect 216220 95464 216272 95470
rect 216220 95406 216272 95412
rect 216416 83570 216444 100014
rect 216692 96937 216720 100028
rect 216864 96960 216916 96966
rect 216678 96928 216734 96937
rect 216864 96902 216916 96908
rect 216678 96863 216734 96872
rect 216772 96892 216824 96898
rect 216772 96834 216824 96840
rect 216784 83638 216812 96834
rect 216876 86426 216904 96902
rect 216968 96830 216996 100028
rect 217060 100014 217166 100042
rect 217350 100014 217456 100042
rect 216956 96824 217008 96830
rect 216956 96766 217008 96772
rect 216864 86420 216916 86426
rect 216864 86362 216916 86368
rect 216772 83632 216824 83638
rect 216772 83574 216824 83580
rect 216404 83564 216456 83570
rect 216404 83506 216456 83512
rect 215944 74044 215996 74050
rect 215944 73986 215996 73992
rect 217060 17270 217088 100014
rect 217324 97776 217376 97782
rect 217324 97718 217376 97724
rect 217336 80782 217364 97718
rect 217428 90642 217456 100014
rect 217520 96966 217548 100028
rect 217612 100014 217718 100042
rect 217508 96960 217560 96966
rect 217508 96902 217560 96908
rect 217612 96898 217640 100014
rect 217980 99550 218008 100028
rect 217968 99544 218020 99550
rect 217968 99486 218020 99492
rect 218164 97034 218192 100028
rect 218152 97028 218204 97034
rect 218152 96970 218204 96976
rect 218244 96960 218296 96966
rect 218348 96937 218376 100028
rect 218244 96902 218296 96908
rect 218334 96928 218390 96937
rect 217600 96892 217652 96898
rect 217600 96834 217652 96840
rect 217416 90636 217468 90642
rect 217416 90578 217468 90584
rect 218256 86494 218284 96902
rect 218334 96863 218390 96872
rect 218428 96892 218480 96898
rect 218428 96834 218480 96840
rect 218244 86488 218296 86494
rect 218244 86430 218296 86436
rect 217324 80776 217376 80782
rect 217324 80718 217376 80724
rect 218440 79490 218468 96834
rect 218532 89078 218560 100028
rect 218624 100014 218730 100042
rect 218808 100014 219006 100042
rect 219084 100014 219190 100042
rect 219268 100014 219374 100042
rect 218624 96966 218652 100014
rect 218612 96960 218664 96966
rect 218612 96902 218664 96908
rect 218520 89072 218572 89078
rect 218520 89014 218572 89020
rect 218808 83706 218836 100014
rect 219084 89146 219112 100014
rect 219268 96898 219296 100014
rect 219544 97617 219572 100028
rect 219728 97782 219756 100028
rect 219716 97776 219768 97782
rect 219716 97718 219768 97724
rect 219530 97608 219586 97617
rect 219530 97543 219586 97552
rect 219808 97028 219860 97034
rect 219808 96970 219860 96976
rect 219256 96892 219308 96898
rect 219256 96834 219308 96840
rect 219624 96892 219676 96898
rect 219624 96834 219676 96840
rect 219072 89140 219124 89146
rect 219072 89082 219124 89088
rect 219636 85066 219664 96834
rect 219624 85060 219676 85066
rect 219624 85002 219676 85008
rect 218796 83700 218848 83706
rect 218796 83642 218848 83648
rect 218428 79484 218480 79490
rect 218428 79426 218480 79432
rect 219820 71398 219848 96970
rect 219900 96960 219952 96966
rect 219900 96902 219952 96908
rect 219912 79558 219940 96902
rect 220004 86562 220032 100028
rect 220096 100014 220202 100042
rect 220280 100014 220386 100042
rect 220464 100014 220570 100042
rect 220648 100014 220754 100042
rect 220096 96898 220124 100014
rect 220280 96966 220308 100014
rect 220268 96960 220320 96966
rect 220268 96902 220320 96908
rect 220084 96892 220136 96898
rect 220084 96834 220136 96840
rect 220464 86630 220492 100014
rect 220648 97034 220676 100014
rect 220636 97028 220688 97034
rect 220636 96970 220688 96976
rect 221016 96937 221044 100028
rect 221002 96928 221058 96937
rect 221002 96863 221058 96872
rect 221200 86698 221228 100028
rect 221292 100014 221398 100042
rect 221476 100014 221582 100042
rect 221188 86692 221240 86698
rect 221188 86634 221240 86640
rect 220452 86624 220504 86630
rect 220452 86566 220504 86572
rect 219992 86556 220044 86562
rect 219992 86498 220044 86504
rect 219900 79552 219952 79558
rect 219900 79494 219952 79500
rect 220728 77988 220780 77994
rect 220728 77930 220780 77936
rect 219808 71392 219860 71398
rect 219808 71334 219860 71340
rect 219348 42084 219400 42090
rect 219348 42026 219400 42032
rect 217048 17264 217100 17270
rect 217048 17206 217100 17212
rect 215760 13116 215812 13122
rect 215760 13058 215812 13064
rect 217968 13116 218020 13122
rect 217968 13058 218020 13064
rect 213840 11750 213960 11778
rect 213368 3664 213420 3670
rect 213368 3606 213420 3612
rect 213184 3256 213236 3262
rect 213184 3198 213236 3204
rect 213380 480 213408 3606
rect 213932 3466 213960 11750
rect 216588 10328 216640 10334
rect 216588 10270 216640 10276
rect 213920 3460 213972 3466
rect 213920 3402 213972 3408
rect 214472 3460 214524 3466
rect 214472 3402 214524 3408
rect 214484 480 214512 3402
rect 216600 3262 216628 10270
rect 217980 3466 218008 13058
rect 219360 3738 219388 42026
rect 220452 3800 220504 3806
rect 220452 3742 220504 3748
rect 218060 3732 218112 3738
rect 218060 3674 218112 3680
rect 219348 3732 219400 3738
rect 219348 3674 219400 3680
rect 216864 3460 216916 3466
rect 216864 3402 216916 3408
rect 217968 3460 218020 3466
rect 217968 3402 218020 3408
rect 215668 3256 215720 3262
rect 215668 3198 215720 3204
rect 216588 3256 216640 3262
rect 216588 3198 216640 3204
rect 215680 480 215708 3198
rect 216876 480 216904 3402
rect 218072 480 218100 3674
rect 219256 3596 219308 3602
rect 219256 3538 219308 3544
rect 219268 480 219296 3538
rect 220464 480 220492 3742
rect 220740 3466 220768 77930
rect 221292 68474 221320 100014
rect 221476 76634 221504 100014
rect 221752 94586 221780 100028
rect 222028 96150 222056 100028
rect 222016 96144 222068 96150
rect 222016 96086 222068 96092
rect 222212 95985 222240 100028
rect 222292 97028 222344 97034
rect 222292 96970 222344 96976
rect 222198 95976 222254 95985
rect 222198 95911 222254 95920
rect 221740 94580 221792 94586
rect 221740 94522 221792 94528
rect 222304 82278 222332 96970
rect 222396 96937 222424 100028
rect 222382 96928 222438 96937
rect 222382 96863 222438 96872
rect 222580 92070 222608 100028
rect 222660 96960 222712 96966
rect 222660 96902 222712 96908
rect 222568 92064 222620 92070
rect 222568 92006 222620 92012
rect 222292 82272 222344 82278
rect 222292 82214 222344 82220
rect 222672 76702 222700 96902
rect 222764 96014 222792 100028
rect 222856 100014 223054 100042
rect 223132 100014 223238 100042
rect 223316 100014 223422 100042
rect 222856 99754 222884 100014
rect 222844 99748 222896 99754
rect 222844 99690 222896 99696
rect 223132 97034 223160 100014
rect 223120 97028 223172 97034
rect 223120 96970 223172 96976
rect 223316 96966 223344 100014
rect 223488 97436 223540 97442
rect 223488 97378 223540 97384
rect 223304 96960 223356 96966
rect 223304 96902 223356 96908
rect 223500 96694 223528 97378
rect 223592 96937 223620 100028
rect 223790 100014 223896 100042
rect 223672 96960 223724 96966
rect 223578 96928 223634 96937
rect 223672 96902 223724 96908
rect 223578 96863 223634 96872
rect 222844 96688 222896 96694
rect 222844 96630 222896 96636
rect 223488 96688 223540 96694
rect 223488 96630 223540 96636
rect 222752 96008 222804 96014
rect 222752 95950 222804 95956
rect 222660 76696 222712 76702
rect 222660 76638 222712 76644
rect 221464 76628 221516 76634
rect 221464 76570 221516 76576
rect 221280 68468 221332 68474
rect 221280 68410 221332 68416
rect 222856 10334 222884 96630
rect 222936 95260 222988 95266
rect 222936 95202 222988 95208
rect 222948 76974 222976 95202
rect 223488 81456 223540 81462
rect 223488 81398 223540 81404
rect 222936 76968 222988 76974
rect 222936 76910 222988 76916
rect 222844 10328 222896 10334
rect 222844 10270 222896 10276
rect 223500 3466 223528 81398
rect 223684 76838 223712 96902
rect 223672 76832 223724 76838
rect 223672 76774 223724 76780
rect 223868 76770 223896 100014
rect 224052 97646 224080 100028
rect 224144 100014 224250 100042
rect 224040 97640 224092 97646
rect 224040 97582 224092 97588
rect 224144 93294 224172 100014
rect 224224 96892 224276 96898
rect 224224 96834 224276 96840
rect 224132 93288 224184 93294
rect 224132 93230 224184 93236
rect 224236 82414 224264 96834
rect 224420 94654 224448 100028
rect 224604 97986 224632 100028
rect 224696 100014 224802 100042
rect 224592 97980 224644 97986
rect 224592 97922 224644 97928
rect 224696 96966 224724 100014
rect 224684 96960 224736 96966
rect 224684 96902 224736 96908
rect 224408 94648 224460 94654
rect 224408 94590 224460 94596
rect 224868 93152 224920 93158
rect 224868 93094 224920 93100
rect 224224 82408 224276 82414
rect 224224 82350 224276 82356
rect 223856 76764 223908 76770
rect 223856 76706 223908 76712
rect 224880 3466 224908 93094
rect 225064 83774 225092 100028
rect 225156 100014 225262 100042
rect 225156 99822 225184 100014
rect 225144 99816 225196 99822
rect 225144 99758 225196 99764
rect 225432 99374 225460 100028
rect 225248 99346 225460 99374
rect 225524 100014 225630 100042
rect 225248 93362 225276 99346
rect 225236 93356 225288 93362
rect 225236 93298 225288 93304
rect 225524 90778 225552 100014
rect 225892 97510 225920 100028
rect 226076 99686 226104 100028
rect 226168 100014 226274 100042
rect 226064 99680 226116 99686
rect 226064 99622 226116 99628
rect 226168 99374 226196 100014
rect 225984 99346 226196 99374
rect 225880 97504 225932 97510
rect 225880 97446 225932 97452
rect 225512 90772 225564 90778
rect 225512 90714 225564 90720
rect 225984 90658 226012 99346
rect 226064 97368 226116 97374
rect 226064 97310 226116 97316
rect 225340 90630 226012 90658
rect 225052 83768 225104 83774
rect 225052 83710 225104 83716
rect 225340 76906 225368 90630
rect 226076 89714 226104 97310
rect 226444 96665 226472 100028
rect 226628 99618 226656 100028
rect 226720 100014 226918 100042
rect 226616 99612 226668 99618
rect 226616 99554 226668 99560
rect 226720 99374 226748 100014
rect 226628 99346 226748 99374
rect 226430 96656 226486 96665
rect 226430 96591 226486 96600
rect 226628 90710 226656 99346
rect 226984 96756 227036 96762
rect 226984 96698 227036 96704
rect 226708 94580 226760 94586
rect 226708 94522 226760 94528
rect 226616 90704 226668 90710
rect 226616 90646 226668 90652
rect 225616 89686 226104 89714
rect 225328 76900 225380 76906
rect 225328 76842 225380 76848
rect 225616 8974 225644 89686
rect 226720 80850 226748 94522
rect 226996 92138 227024 96698
rect 227088 94722 227116 100028
rect 227180 100014 227286 100042
rect 227364 100014 227470 100042
rect 227076 94716 227128 94722
rect 227076 94658 227128 94664
rect 226984 92132 227036 92138
rect 226984 92074 227036 92080
rect 227180 89714 227208 100014
rect 227364 94586 227392 100014
rect 227640 98734 227668 100028
rect 227628 98728 227680 98734
rect 227628 98670 227680 98676
rect 227916 94858 227944 100028
rect 228008 100014 228114 100042
rect 227904 94852 227956 94858
rect 227904 94794 227956 94800
rect 227352 94580 227404 94586
rect 227352 94522 227404 94528
rect 227628 94444 227680 94450
rect 227628 94386 227680 94392
rect 226812 89686 227208 89714
rect 226812 82346 226840 89686
rect 226984 83496 227036 83502
rect 226984 83438 227036 83444
rect 226800 82340 226852 82346
rect 226800 82282 226852 82288
rect 226708 80844 226760 80850
rect 226708 80786 226760 80792
rect 225604 8968 225656 8974
rect 225604 8910 225656 8916
rect 225144 3936 225196 3942
rect 225144 3878 225196 3884
rect 220728 3460 220780 3466
rect 220728 3402 220780 3408
rect 221556 3460 221608 3466
rect 221556 3402 221608 3408
rect 222752 3460 222804 3466
rect 222752 3402 222804 3408
rect 223488 3460 223540 3466
rect 223488 3402 223540 3408
rect 223948 3460 224000 3466
rect 223948 3402 224000 3408
rect 224868 3460 224920 3466
rect 224868 3402 224920 3408
rect 221568 480 221596 3402
rect 222764 480 222792 3402
rect 223960 480 223988 3402
rect 225156 480 225184 3878
rect 226340 3868 226392 3874
rect 226340 3810 226392 3816
rect 226352 480 226380 3810
rect 226996 3670 227024 83438
rect 227640 6914 227668 94386
rect 228008 80918 228036 100014
rect 228284 97850 228312 100028
rect 228376 100014 228482 100042
rect 228272 97844 228324 97850
rect 228272 97786 228324 97792
rect 228376 94858 228404 100014
rect 228456 97504 228508 97510
rect 228456 97446 228508 97452
rect 228364 94852 228416 94858
rect 228364 94794 228416 94800
rect 228364 94716 228416 94722
rect 228364 94658 228416 94664
rect 227996 80912 228048 80918
rect 227996 80854 228048 80860
rect 227548 6886 227668 6914
rect 226984 3664 227036 3670
rect 226984 3606 227036 3612
rect 227548 480 227576 6886
rect 228376 3398 228404 94658
rect 228468 81462 228496 97446
rect 228652 96898 228680 100028
rect 228928 98802 228956 100028
rect 228916 98796 228968 98802
rect 228916 98738 228968 98744
rect 228640 96892 228692 96898
rect 228640 96834 228692 96840
rect 228548 96688 228600 96694
rect 228548 96630 228600 96636
rect 228560 88058 228588 96630
rect 229112 94625 229140 100028
rect 229296 96762 229324 100028
rect 229388 100014 229494 100042
rect 229572 100014 229678 100042
rect 229756 100014 229954 100042
rect 230032 100014 230138 100042
rect 230216 100014 230322 100042
rect 229284 96756 229336 96762
rect 229284 96698 229336 96704
rect 229388 95266 229416 100014
rect 229572 99374 229600 100014
rect 229480 99346 229600 99374
rect 229376 95260 229428 95266
rect 229376 95202 229428 95208
rect 229098 94616 229154 94625
rect 229008 94580 229060 94586
rect 229480 94602 229508 99346
rect 229098 94551 229154 94560
rect 229204 94574 229508 94602
rect 229008 94522 229060 94528
rect 228548 88052 228600 88058
rect 228548 87994 228600 88000
rect 228456 81456 228508 81462
rect 228456 81398 228508 81404
rect 229020 6914 229048 94522
rect 229204 85202 229232 94574
rect 229376 94512 229428 94518
rect 229376 94454 229428 94460
rect 229388 89418 229416 94454
rect 229376 89412 229428 89418
rect 229376 89354 229428 89360
rect 229192 85196 229244 85202
rect 229192 85138 229244 85144
rect 229756 84194 229784 100014
rect 230032 89350 230060 100014
rect 230216 94518 230244 100014
rect 230492 96801 230520 100028
rect 230676 98870 230704 100028
rect 230664 98864 230716 98870
rect 230664 98806 230716 98812
rect 230478 96792 230534 96801
rect 230478 96727 230534 96736
rect 230952 96665 230980 100028
rect 231044 100014 231150 100042
rect 230938 96656 230994 96665
rect 230938 96591 230994 96600
rect 230204 94512 230256 94518
rect 230204 94454 230256 94460
rect 230020 89344 230072 89350
rect 230020 89286 230072 89292
rect 230388 87644 230440 87650
rect 230388 87586 230440 87592
rect 229572 84166 229784 84194
rect 229572 82482 229600 84166
rect 229560 82476 229612 82482
rect 229560 82418 229612 82424
rect 228744 6886 229048 6914
rect 228364 3392 228416 3398
rect 228364 3334 228416 3340
rect 228744 480 228772 6886
rect 229836 3460 229888 3466
rect 229836 3402 229888 3408
rect 229848 480 229876 3402
rect 230400 3194 230428 87586
rect 231044 85134 231072 100014
rect 231216 97980 231268 97986
rect 231216 97922 231268 97928
rect 231122 96520 231178 96529
rect 231122 96455 231178 96464
rect 231032 85128 231084 85134
rect 231032 85070 231084 85076
rect 231136 3806 231164 96455
rect 231228 42090 231256 97922
rect 231320 96082 231348 100028
rect 231412 100014 231518 100042
rect 231596 100014 231702 100042
rect 231308 96076 231360 96082
rect 231308 96018 231360 96024
rect 231412 93430 231440 100014
rect 231400 93424 231452 93430
rect 231400 93366 231452 93372
rect 231596 92206 231624 100014
rect 231964 96121 231992 100028
rect 232148 96665 232176 100028
rect 232240 100014 232346 100042
rect 232134 96656 232190 96665
rect 232134 96591 232190 96600
rect 231950 96112 232006 96121
rect 231950 96047 232006 96056
rect 231584 92200 231636 92206
rect 231584 92142 231636 92148
rect 232240 91798 232268 100014
rect 232516 96218 232544 100028
rect 232608 100014 232714 100042
rect 232792 100014 232990 100042
rect 233068 100014 233174 100042
rect 232504 96212 232556 96218
rect 232504 96154 232556 96160
rect 232608 93498 232636 100014
rect 232596 93492 232648 93498
rect 232596 93434 232648 93440
rect 232228 91792 232280 91798
rect 232228 91734 232280 91740
rect 231768 91112 231820 91118
rect 231768 91054 231820 91060
rect 231216 42084 231268 42090
rect 231216 42026 231268 42032
rect 231124 3800 231176 3806
rect 231124 3742 231176 3748
rect 231780 3534 231808 91054
rect 232792 89714 232820 100014
rect 232240 89686 232820 89714
rect 232240 83842 232268 89686
rect 232504 85604 232556 85610
rect 232504 85546 232556 85552
rect 232228 83836 232280 83842
rect 232228 83778 232280 83784
rect 232516 3874 232544 85546
rect 233068 84862 233096 100014
rect 233344 96665 233372 100028
rect 233436 100014 233542 100042
rect 233330 96656 233386 96665
rect 233330 96591 233386 96600
rect 233436 91866 233464 100014
rect 233804 96694 233832 100028
rect 233896 100014 234002 100042
rect 234080 100014 234186 100042
rect 233792 96688 233844 96694
rect 233792 96630 233844 96636
rect 233896 93566 233924 100014
rect 233884 93560 233936 93566
rect 233884 93502 233936 93508
rect 233424 91860 233476 91866
rect 233424 91802 233476 91808
rect 233148 91384 233200 91390
rect 233148 91326 233200 91332
rect 233056 84856 233108 84862
rect 233056 84798 233108 84804
rect 232504 3868 232556 3874
rect 232504 3810 232556 3816
rect 233160 3534 233188 91326
rect 233608 89956 233660 89962
rect 233608 89898 233660 89904
rect 233424 4480 233476 4486
rect 233424 4422 233476 4428
rect 231032 3528 231084 3534
rect 231032 3470 231084 3476
rect 231768 3528 231820 3534
rect 231768 3470 231820 3476
rect 232228 3528 232280 3534
rect 232228 3470 232280 3476
rect 233148 3528 233200 3534
rect 233148 3470 233200 3476
rect 230388 3188 230440 3194
rect 230388 3130 230440 3136
rect 231044 480 231072 3470
rect 232240 480 232268 3470
rect 233436 480 233464 4422
rect 233620 3602 233648 89898
rect 234080 84194 234108 100014
rect 234356 98666 234384 100028
rect 234448 100014 234554 100042
rect 234344 98660 234396 98666
rect 234344 98602 234396 98608
rect 234448 89962 234476 100014
rect 234528 97708 234580 97714
rect 234528 97650 234580 97656
rect 234436 89956 234488 89962
rect 234436 89898 234488 89904
rect 233896 84166 234108 84194
rect 233896 82550 233924 84166
rect 233884 82544 233936 82550
rect 233884 82486 233936 82492
rect 233882 81560 233938 81569
rect 233882 81495 233938 81504
rect 233896 3670 233924 81495
rect 234540 6914 234568 97650
rect 234712 96960 234764 96966
rect 234712 96902 234764 96908
rect 234724 35222 234752 96902
rect 234816 96694 234844 100028
rect 235000 99482 235028 100028
rect 234988 99476 235040 99482
rect 234988 99418 235040 99424
rect 234988 99272 235040 99278
rect 234988 99214 235040 99220
rect 234896 97164 234948 97170
rect 234896 97106 234948 97112
rect 234804 96688 234856 96694
rect 234804 96630 234856 96636
rect 234908 87990 234936 97106
rect 235000 96286 235028 99214
rect 235184 97170 235212 100028
rect 235276 100014 235382 100042
rect 235172 97164 235224 97170
rect 235172 97106 235224 97112
rect 235276 96778 235304 100014
rect 235552 98938 235580 100028
rect 235644 100014 235842 100042
rect 236026 100014 236132 100042
rect 235540 98932 235592 98938
rect 235540 98874 235592 98880
rect 235644 96966 235672 100014
rect 235632 96960 235684 96966
rect 235632 96902 235684 96908
rect 235092 96750 235304 96778
rect 234988 96280 235040 96286
rect 234988 96222 235040 96228
rect 234896 87984 234948 87990
rect 234896 87926 234948 87932
rect 234712 35216 234764 35222
rect 234712 35158 234764 35164
rect 234540 6886 234660 6914
rect 233884 3664 233936 3670
rect 233884 3606 233936 3612
rect 233608 3596 233660 3602
rect 233608 3538 233660 3544
rect 234632 480 234660 6886
rect 235092 2106 235120 96750
rect 236104 96694 236132 100014
rect 236196 97374 236224 100028
rect 236184 97368 236236 97374
rect 236184 97310 236236 97316
rect 236276 96960 236328 96966
rect 236276 96902 236328 96908
rect 235264 96688 235316 96694
rect 235264 96630 235316 96636
rect 236092 96688 236144 96694
rect 236092 96630 236144 96636
rect 235276 3369 235304 96630
rect 236288 13122 236316 96902
rect 236380 94654 236408 100028
rect 236368 94648 236420 94654
rect 236368 94590 236420 94596
rect 236564 83502 236592 100028
rect 236840 97306 236868 100028
rect 237024 97442 237052 100028
rect 237116 100014 237222 100042
rect 237012 97436 237064 97442
rect 237012 97378 237064 97384
rect 236828 97300 236880 97306
rect 236828 97242 236880 97248
rect 236644 97164 236696 97170
rect 236644 97106 236696 97112
rect 236656 91118 236684 97106
rect 237116 96966 237144 100014
rect 237392 97986 237420 100028
rect 237380 97980 237432 97986
rect 237380 97922 237432 97928
rect 237380 97844 237432 97850
rect 237380 97786 237432 97792
rect 237104 96960 237156 96966
rect 237104 96902 237156 96908
rect 236736 96688 236788 96694
rect 236736 96630 236788 96636
rect 236644 91112 236696 91118
rect 236644 91054 236696 91060
rect 236552 83496 236604 83502
rect 236552 83438 236604 83444
rect 236748 43450 236776 96630
rect 237392 94518 237420 97786
rect 237576 96937 237604 100028
rect 237852 96937 237880 100028
rect 237944 100014 238050 100042
rect 237562 96928 237618 96937
rect 237562 96863 237618 96872
rect 237838 96928 237894 96937
rect 237838 96863 237894 96872
rect 237944 96778 237972 100014
rect 238220 97510 238248 100028
rect 238312 100014 238418 100042
rect 238496 100014 238602 100042
rect 238208 97504 238260 97510
rect 238208 97446 238260 97452
rect 237484 96750 237972 96778
rect 237380 94512 237432 94518
rect 237380 94454 237432 94460
rect 237484 77994 237512 96750
rect 237656 96688 237708 96694
rect 237656 96630 237708 96636
rect 237472 77988 237524 77994
rect 237472 77930 237524 77936
rect 236736 43444 236788 43450
rect 236736 43386 236788 43392
rect 236276 13116 236328 13122
rect 236276 13058 236328 13064
rect 237668 3942 237696 96630
rect 238312 93158 238340 100014
rect 238496 96694 238524 100014
rect 238668 97980 238720 97986
rect 238668 97922 238720 97928
rect 238484 96688 238536 96694
rect 238484 96630 238536 96636
rect 238300 93152 238352 93158
rect 238300 93094 238352 93100
rect 238680 22778 238708 97922
rect 238864 85610 238892 100028
rect 238944 98320 238996 98326
rect 238944 98262 238996 98268
rect 238852 85604 238904 85610
rect 238852 85546 238904 85552
rect 238956 23594 238984 98262
rect 239048 97850 239076 100028
rect 239232 99482 239260 100028
rect 239220 99476 239272 99482
rect 239220 99418 239272 99424
rect 239220 99272 239272 99278
rect 239220 99214 239272 99220
rect 239036 97844 239088 97850
rect 239036 97786 239088 97792
rect 239128 96824 239180 96830
rect 239128 96766 239180 96772
rect 238944 23588 238996 23594
rect 238944 23530 238996 23536
rect 238668 22772 238720 22778
rect 238668 22714 238720 22720
rect 238024 22092 238076 22098
rect 238024 22034 238076 22040
rect 237656 3936 237708 3942
rect 237656 3878 237708 3884
rect 238036 3534 238064 22034
rect 239140 4486 239168 96766
rect 239232 94586 239260 99214
rect 239416 98326 239444 100028
rect 239404 98320 239456 98326
rect 239404 98262 239456 98268
rect 239600 97170 239628 100028
rect 239692 100014 239890 100042
rect 239968 100014 240074 100042
rect 239588 97164 239640 97170
rect 239588 97106 239640 97112
rect 239220 94580 239272 94586
rect 239220 94522 239272 94528
rect 239692 91390 239720 100014
rect 239968 96830 239996 100014
rect 240244 97714 240272 100028
rect 240232 97708 240284 97714
rect 240232 97650 240284 97656
rect 239956 96824 240008 96830
rect 239956 96766 240008 96772
rect 240140 96688 240192 96694
rect 240140 96630 240192 96636
rect 239680 91384 239732 91390
rect 239680 91326 239732 91332
rect 239128 4480 239180 4486
rect 239128 4422 239180 4428
rect 238116 3732 238168 3738
rect 238116 3674 238168 3680
rect 237012 3528 237064 3534
rect 237012 3470 237064 3476
rect 238024 3528 238076 3534
rect 238024 3470 238076 3476
rect 235262 3360 235318 3369
rect 235262 3295 235318 3304
rect 235816 3188 235868 3194
rect 235816 3130 235868 3136
rect 235080 2100 235132 2106
rect 235080 2042 235132 2048
rect 235828 480 235856 3130
rect 237024 480 237052 3470
rect 238128 480 238156 3674
rect 239312 3664 239364 3670
rect 239312 3606 239364 3612
rect 239324 480 239352 3606
rect 240152 490 240180 96630
rect 240324 96212 240376 96218
rect 240324 96154 240376 96160
rect 240336 68338 240364 96154
rect 240428 87650 240456 100028
rect 240508 96960 240560 96966
rect 240508 96902 240560 96908
rect 240416 87644 240468 87650
rect 240416 87586 240468 87592
rect 240520 80850 240548 96902
rect 240508 80844 240560 80850
rect 240508 80786 240560 80792
rect 240324 68332 240376 68338
rect 240324 68274 240376 68280
rect 240232 23588 240284 23594
rect 240232 23530 240284 23536
rect 240244 3466 240272 23530
rect 240612 22098 240640 100028
rect 240704 100014 240902 100042
rect 240980 100014 241086 100042
rect 240704 96218 240732 100014
rect 240980 96966 241008 100014
rect 240968 96960 241020 96966
rect 240968 96902 241020 96908
rect 241256 96694 241284 100028
rect 241440 97986 241468 100028
rect 241428 97980 241480 97986
rect 241428 97922 241480 97928
rect 241624 96762 241652 100028
rect 241900 96830 241928 100028
rect 242084 96966 242112 100028
rect 242282 100014 242388 100042
rect 242466 100014 242664 100042
rect 242072 96960 242124 96966
rect 242072 96902 242124 96908
rect 241888 96824 241940 96830
rect 241888 96766 241940 96772
rect 241612 96756 241664 96762
rect 241612 96698 241664 96704
rect 241244 96688 241296 96694
rect 241244 96630 241296 96636
rect 240692 96212 240744 96218
rect 240692 96154 240744 96160
rect 242360 93854 242388 100014
rect 242532 96960 242584 96966
rect 242532 96902 242584 96908
rect 242636 96914 242664 100014
rect 242728 97578 242756 100028
rect 242716 97572 242768 97578
rect 242716 97514 242768 97520
rect 242360 93826 242480 93854
rect 241520 22772 241572 22778
rect 241520 22714 241572 22720
rect 240600 22092 240652 22098
rect 240600 22034 240652 22040
rect 241532 16574 241560 22714
rect 241532 16546 241744 16574
rect 240232 3460 240284 3466
rect 240232 3402 240284 3408
rect 240336 598 240548 626
rect 240336 490 240364 598
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240152 462 240364 490
rect 240520 480 240548 598
rect 241716 480 241744 16546
rect 242452 4214 242480 93826
rect 242544 75886 242572 96902
rect 242636 96886 242848 96914
rect 242624 96824 242676 96830
rect 242624 96766 242676 96772
rect 242532 75880 242584 75886
rect 242532 75822 242584 75828
rect 242636 41478 242664 96766
rect 242716 96756 242768 96762
rect 242716 96698 242768 96704
rect 242624 41472 242676 41478
rect 242624 41414 242676 41420
rect 242728 28966 242756 96698
rect 242820 91798 242848 96886
rect 242912 96830 242940 100028
rect 242900 96824 242952 96830
rect 242900 96766 242952 96772
rect 243096 96762 243124 100028
rect 243280 97170 243308 100028
rect 243268 97164 243320 97170
rect 243268 97106 243320 97112
rect 243464 97102 243492 100028
rect 243754 100014 243860 100042
rect 243452 97096 243504 97102
rect 243452 97038 243504 97044
rect 243832 96914 243860 100014
rect 243924 97034 243952 100028
rect 243912 97028 243964 97034
rect 243912 96970 243964 96976
rect 243832 96886 244044 96914
rect 243820 96824 243872 96830
rect 243820 96766 243872 96772
rect 243084 96756 243136 96762
rect 243084 96698 243136 96704
rect 242808 91792 242860 91798
rect 242808 91734 242860 91740
rect 243832 42770 243860 96766
rect 243912 96756 243964 96762
rect 243912 96698 243964 96704
rect 243924 84862 243952 96698
rect 243912 84856 243964 84862
rect 243912 84798 243964 84804
rect 244016 77994 244044 96886
rect 244004 77988 244056 77994
rect 244004 77930 244056 77936
rect 244108 47598 244136 100028
rect 244188 97028 244240 97034
rect 244188 96970 244240 96976
rect 244200 93158 244228 96970
rect 244292 96898 244320 100028
rect 244476 97442 244504 100028
rect 244766 100014 244872 100042
rect 244464 97436 244516 97442
rect 244464 97378 244516 97384
rect 244280 96892 244332 96898
rect 244280 96834 244332 96840
rect 244844 93854 244872 100014
rect 244936 96966 244964 100028
rect 245120 97306 245148 100028
rect 245108 97300 245160 97306
rect 245108 97242 245160 97248
rect 244924 96960 244976 96966
rect 244924 96902 244976 96908
rect 244844 93826 245240 93854
rect 244188 93152 244240 93158
rect 244188 93094 244240 93100
rect 245212 79354 245240 93826
rect 245200 79348 245252 79354
rect 245200 79290 245252 79296
rect 245304 76566 245332 100028
rect 245502 100014 245608 100042
rect 245476 96960 245528 96966
rect 245476 96902 245528 96908
rect 245384 96892 245436 96898
rect 245384 96834 245436 96840
rect 245292 76560 245344 76566
rect 245292 76502 245344 76508
rect 244280 75880 244332 75886
rect 244280 75822 244332 75828
rect 244096 47592 244148 47598
rect 244096 47534 244148 47540
rect 243820 42764 243872 42770
rect 243820 42706 243872 42712
rect 242900 41472 242952 41478
rect 242900 41414 242952 41420
rect 242716 28960 242768 28966
rect 242716 28902 242768 28908
rect 242912 11762 242940 41414
rect 244292 16574 244320 75822
rect 245396 75206 245424 96834
rect 245384 75200 245436 75206
rect 245384 75142 245436 75148
rect 244292 16546 245240 16574
rect 242900 11756 242952 11762
rect 242900 11698 242952 11704
rect 244096 11756 244148 11762
rect 244096 11698 244148 11704
rect 242440 4208 242492 4214
rect 242440 4150 242492 4156
rect 242900 3460 242952 3466
rect 242900 3402 242952 3408
rect 242912 480 242940 3402
rect 244108 480 244136 11698
rect 245212 480 245240 16546
rect 245488 6322 245516 96902
rect 245476 6316 245528 6322
rect 245476 6258 245528 6264
rect 245580 3602 245608 100014
rect 245764 97510 245792 100028
rect 245752 97504 245804 97510
rect 245752 97446 245804 97452
rect 245948 96762 245976 100028
rect 246132 97238 246160 100028
rect 246316 97374 246344 100028
rect 246514 100014 246712 100042
rect 246304 97368 246356 97374
rect 246304 97310 246356 97316
rect 246120 97232 246172 97238
rect 246120 97174 246172 97180
rect 246304 97164 246356 97170
rect 246304 97106 246356 97112
rect 245936 96756 245988 96762
rect 245936 96698 245988 96704
rect 246316 76634 246344 97106
rect 246396 97096 246448 97102
rect 246396 97038 246448 97044
rect 246408 86290 246436 97038
rect 246684 96914 246712 100014
rect 246776 97034 246804 100028
rect 246764 97028 246816 97034
rect 246764 96970 246816 96976
rect 246960 96937 246988 100028
rect 247144 97034 247172 100028
rect 247328 97646 247356 100028
rect 247316 97640 247368 97646
rect 247316 97582 247368 97588
rect 247132 97028 247184 97034
rect 247132 96970 247184 96976
rect 246946 96928 247002 96937
rect 246684 96886 246896 96914
rect 246764 96756 246816 96762
rect 246764 96698 246816 96704
rect 246396 86284 246448 86290
rect 246396 86226 246448 86232
rect 246304 76628 246356 76634
rect 246304 76570 246356 76576
rect 246776 51746 246804 96698
rect 246764 51740 246816 51746
rect 246764 51682 246816 51688
rect 245660 28960 245712 28966
rect 245660 28902 245712 28908
rect 245568 3596 245620 3602
rect 245568 3538 245620 3544
rect 245672 3466 245700 28902
rect 246868 28286 246896 96886
rect 246946 96863 247002 96872
rect 247512 96830 247540 100028
rect 247684 97572 247736 97578
rect 247684 97514 247736 97520
rect 246948 96824 247000 96830
rect 246948 96766 247000 96772
rect 247500 96824 247552 96830
rect 247500 96766 247552 96772
rect 246856 28280 246908 28286
rect 246856 28222 246908 28228
rect 246396 4208 246448 4214
rect 246396 4150 246448 4156
rect 245660 3460 245712 3466
rect 245660 3402 245712 3408
rect 246408 480 246436 4150
rect 246960 3534 246988 96766
rect 247696 45830 247724 97514
rect 247788 96966 247816 100028
rect 247986 100014 248092 100042
rect 248170 100014 248276 100042
rect 247776 96960 247828 96966
rect 247776 96902 247828 96908
rect 248064 89010 248092 100014
rect 248144 96960 248196 96966
rect 248144 96902 248196 96908
rect 248248 96914 248276 100014
rect 248340 99006 248368 100028
rect 248328 99000 248380 99006
rect 248328 98942 248380 98948
rect 248052 89004 248104 89010
rect 248052 88946 248104 88952
rect 248156 82142 248184 96902
rect 248248 96886 248368 96914
rect 248236 96824 248288 96830
rect 248236 96766 248288 96772
rect 248144 82136 248196 82142
rect 248144 82078 248196 82084
rect 248248 71058 248276 96766
rect 248236 71052 248288 71058
rect 248236 70994 248288 71000
rect 247684 45824 247736 45830
rect 247684 45766 247736 45772
rect 248340 6254 248368 96886
rect 248524 96694 248552 100028
rect 248800 96898 248828 100028
rect 248984 97102 249012 100028
rect 248972 97096 249024 97102
rect 248972 97038 249024 97044
rect 249168 96966 249196 100028
rect 249366 100014 249472 100042
rect 249064 96960 249116 96966
rect 249064 96902 249116 96908
rect 249156 96960 249208 96966
rect 249156 96902 249208 96908
rect 248788 96892 248840 96898
rect 248788 96834 248840 96840
rect 248512 96688 248564 96694
rect 248512 96630 248564 96636
rect 248420 45824 248472 45830
rect 248420 45766 248472 45772
rect 248328 6248 248380 6254
rect 248328 6190 248380 6196
rect 247592 3868 247644 3874
rect 247592 3810 247644 3816
rect 246948 3528 247000 3534
rect 246948 3470 247000 3476
rect 247604 480 247632 3810
rect 248432 490 248460 45766
rect 249076 3466 249104 96902
rect 249444 96778 249472 100014
rect 249536 96937 249564 100028
rect 249708 96960 249760 96966
rect 249522 96928 249578 96937
rect 249708 96902 249760 96908
rect 249522 96863 249578 96872
rect 249616 96892 249668 96898
rect 249616 96834 249668 96840
rect 249444 96750 249564 96778
rect 249432 96688 249484 96694
rect 249432 96630 249484 96636
rect 249444 87718 249472 96630
rect 249432 87712 249484 87718
rect 249432 87654 249484 87660
rect 249536 87650 249564 96750
rect 249524 87644 249576 87650
rect 249524 87586 249576 87592
rect 249628 46238 249656 96834
rect 249616 46232 249668 46238
rect 249616 46174 249668 46180
rect 249720 6186 249748 96902
rect 249812 96762 249840 100028
rect 249996 96966 250024 100028
rect 249984 96960 250036 96966
rect 249984 96902 250036 96908
rect 250180 96830 250208 100028
rect 250168 96824 250220 96830
rect 250168 96766 250220 96772
rect 249800 96756 249852 96762
rect 249800 96698 249852 96704
rect 250364 94518 250392 100028
rect 250654 100014 250760 100042
rect 250444 97232 250496 97238
rect 250444 97174 250496 97180
rect 250352 94512 250404 94518
rect 250352 94454 250404 94460
rect 249892 68332 249944 68338
rect 249892 68274 249944 68280
rect 249800 42764 249852 42770
rect 249800 42706 249852 42712
rect 249708 6180 249760 6186
rect 249708 6122 249760 6128
rect 249812 3482 249840 42706
rect 249904 3738 249932 68274
rect 250456 42090 250484 97174
rect 250732 96914 250760 100014
rect 250824 97034 250852 100028
rect 250812 97028 250864 97034
rect 250812 96970 250864 96976
rect 251008 96937 251036 100028
rect 251088 97028 251140 97034
rect 251088 96970 251140 96976
rect 250994 96928 251050 96937
rect 250732 96886 250944 96914
rect 250812 96824 250864 96830
rect 250812 96766 250864 96772
rect 250444 42084 250496 42090
rect 250444 42026 250496 42032
rect 250824 7750 250852 96766
rect 250916 80782 250944 96886
rect 250994 96863 251050 96872
rect 250996 96756 251048 96762
rect 250996 96698 251048 96704
rect 250904 80776 250956 80782
rect 250904 80718 250956 80724
rect 251008 73846 251036 96698
rect 251100 96121 251128 96970
rect 251192 96830 251220 100028
rect 251180 96824 251232 96830
rect 251180 96766 251232 96772
rect 251376 96354 251404 100028
rect 251652 96762 251680 100028
rect 251850 100014 251956 100042
rect 251824 97300 251876 97306
rect 251824 97242 251876 97248
rect 251640 96756 251692 96762
rect 251640 96698 251692 96704
rect 251364 96348 251416 96354
rect 251364 96290 251416 96296
rect 251086 96112 251142 96121
rect 251086 96047 251142 96056
rect 251836 78062 251864 97242
rect 251928 96914 251956 100014
rect 252020 97073 252048 100028
rect 252006 97064 252062 97073
rect 252204 97034 252232 100028
rect 252006 96999 252062 97008
rect 252192 97028 252244 97034
rect 252192 96970 252244 96976
rect 252388 96937 252416 100028
rect 252664 97714 252692 100028
rect 252652 97708 252704 97714
rect 252652 97650 252704 97656
rect 252374 96928 252430 96937
rect 251928 96886 252324 96914
rect 252192 96824 252244 96830
rect 252192 96766 252244 96772
rect 252204 80714 252232 96766
rect 252296 89418 252324 96886
rect 252374 96863 252430 96872
rect 252376 96756 252428 96762
rect 252376 96698 252428 96704
rect 252284 89412 252336 89418
rect 252284 89354 252336 89360
rect 252388 88058 252416 96698
rect 252848 96694 252876 100028
rect 253032 96762 253060 100028
rect 253216 99822 253244 100028
rect 253414 100014 253612 100042
rect 253204 99816 253256 99822
rect 253204 99758 253256 99764
rect 253204 97640 253256 97646
rect 253204 97582 253256 97588
rect 253020 96756 253072 96762
rect 253020 96698 253072 96704
rect 252836 96688 252888 96694
rect 252836 96630 252888 96636
rect 252376 88052 252428 88058
rect 252376 87994 252428 88000
rect 252560 86284 252612 86290
rect 252560 86226 252612 86232
rect 252192 80708 252244 80714
rect 252192 80650 252244 80656
rect 251824 78056 251876 78062
rect 251824 77998 251876 78004
rect 251180 76628 251232 76634
rect 251180 76570 251232 76576
rect 250996 73840 251048 73846
rect 250996 73782 251048 73788
rect 251192 11762 251220 76570
rect 251180 11756 251232 11762
rect 251180 11698 251232 11704
rect 252376 11756 252428 11762
rect 252376 11698 252428 11704
rect 250812 7744 250864 7750
rect 250812 7686 250864 7692
rect 249892 3732 249944 3738
rect 249892 3674 249944 3680
rect 249064 3460 249116 3466
rect 249812 3454 250024 3482
rect 249064 3402 249116 3408
rect 248616 598 248828 626
rect 248616 490 248644 598
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248432 462 248644 490
rect 248800 480 248828 598
rect 249996 480 250024 3454
rect 251180 3188 251232 3194
rect 251180 3130 251232 3136
rect 251192 480 251220 3130
rect 252388 480 252416 11698
rect 252572 3482 252600 86226
rect 252652 80844 252704 80850
rect 252652 80786 252704 80792
rect 252664 3670 252692 80786
rect 253216 69698 253244 97582
rect 253296 97028 253348 97034
rect 253296 96970 253348 96976
rect 253308 89350 253336 96970
rect 253584 96778 253612 100014
rect 253676 96937 253704 100028
rect 253860 97306 253888 100028
rect 253848 97300 253900 97306
rect 253848 97242 253900 97248
rect 253662 96928 253718 96937
rect 254044 96898 254072 100028
rect 253662 96863 253718 96872
rect 254032 96892 254084 96898
rect 254032 96834 254084 96840
rect 253584 96750 253796 96778
rect 253664 96688 253716 96694
rect 253664 96630 253716 96636
rect 253676 90778 253704 96630
rect 253664 90772 253716 90778
rect 253664 90714 253716 90720
rect 253296 89344 253348 89350
rect 253296 89286 253348 89292
rect 253768 86562 253796 96750
rect 253848 96756 253900 96762
rect 253848 96698 253900 96704
rect 253756 86556 253808 86562
rect 253756 86498 253808 86504
rect 253860 81122 253888 96698
rect 254228 94858 254256 100028
rect 254412 96762 254440 100028
rect 254688 96966 254716 100028
rect 254584 96960 254636 96966
rect 254584 96902 254636 96908
rect 254676 96960 254728 96966
rect 254676 96902 254728 96908
rect 254400 96756 254452 96762
rect 254400 96698 254452 96704
rect 254216 94852 254268 94858
rect 254216 94794 254268 94800
rect 253848 81116 253900 81122
rect 253848 81058 253900 81064
rect 254596 80850 254624 96902
rect 254584 80844 254636 80850
rect 254584 80786 254636 80792
rect 253204 69692 253256 69698
rect 253204 69634 253256 69640
rect 254872 9382 254900 100028
rect 255056 98870 255084 100028
rect 255044 98864 255096 98870
rect 255044 98806 255096 98812
rect 255044 96960 255096 96966
rect 255240 96937 255268 100028
rect 255044 96902 255096 96908
rect 255226 96928 255282 96937
rect 255056 87990 255084 96902
rect 255136 96892 255188 96898
rect 255424 96898 255452 100028
rect 255700 99754 255728 100028
rect 255688 99748 255740 99754
rect 255688 99690 255740 99696
rect 255780 97096 255832 97102
rect 255780 97038 255832 97044
rect 255226 96863 255282 96872
rect 255412 96892 255464 96898
rect 255136 96834 255188 96840
rect 255412 96834 255464 96840
rect 255044 87984 255096 87990
rect 255044 87926 255096 87932
rect 255148 86698 255176 96834
rect 255792 93854 255820 97038
rect 255884 96966 255912 100028
rect 255964 97436 256016 97442
rect 255964 97378 256016 97384
rect 255872 96960 255924 96966
rect 255872 96902 255924 96908
rect 255976 96778 256004 97378
rect 256068 96937 256096 100028
rect 256266 100014 256372 100042
rect 256054 96928 256110 96937
rect 256054 96863 256110 96872
rect 255976 96750 256096 96778
rect 255792 93826 256004 93854
rect 255320 93152 255372 93158
rect 255320 93094 255372 93100
rect 255136 86692 255188 86698
rect 255136 86634 255188 86640
rect 255332 16574 255360 93094
rect 255332 16546 255912 16574
rect 254860 9376 254912 9382
rect 254860 9318 254912 9324
rect 252652 3664 252704 3670
rect 252652 3606 252704 3612
rect 254676 3664 254728 3670
rect 254676 3606 254728 3612
rect 252572 3454 253520 3482
rect 253492 480 253520 3454
rect 254688 480 254716 3606
rect 255884 480 255912 16546
rect 255976 3369 256004 93826
rect 256068 72622 256096 96750
rect 256344 93498 256372 100014
rect 256436 97850 256464 100028
rect 256424 97844 256476 97850
rect 256424 97786 256476 97792
rect 256516 96960 256568 96966
rect 256516 96902 256568 96908
rect 256332 93492 256384 93498
rect 256332 93434 256384 93440
rect 256528 86630 256556 96902
rect 256608 96892 256660 96898
rect 256608 96834 256660 96840
rect 256516 86624 256568 86630
rect 256516 86566 256568 86572
rect 256620 81054 256648 96834
rect 256712 96286 256740 100028
rect 256896 97782 256924 100028
rect 256884 97776 256936 97782
rect 256884 97718 256936 97724
rect 256700 96280 256752 96286
rect 256700 96222 256752 96228
rect 257080 94926 257108 100028
rect 257264 96694 257292 100028
rect 257462 100014 257660 100042
rect 257344 97504 257396 97510
rect 257344 97446 257396 97452
rect 257252 96688 257304 96694
rect 257252 96630 257304 96636
rect 257068 94920 257120 94926
rect 257068 94862 257120 94868
rect 256608 81048 256660 81054
rect 256608 80990 256660 80996
rect 257356 78130 257384 97446
rect 257632 96778 257660 100014
rect 257724 96937 257752 100028
rect 257908 97374 257936 100028
rect 257896 97368 257948 97374
rect 257896 97310 257948 97316
rect 257710 96928 257766 96937
rect 257710 96863 257766 96872
rect 257632 96750 257936 96778
rect 257804 96688 257856 96694
rect 257804 96630 257856 96636
rect 257344 78124 257396 78130
rect 257344 78066 257396 78072
rect 256056 72616 256108 72622
rect 256056 72558 256108 72564
rect 257816 47598 257844 96630
rect 257908 93430 257936 96750
rect 258092 96150 258120 100028
rect 258276 97034 258304 100028
rect 258264 97028 258316 97034
rect 258264 96970 258316 96976
rect 258552 96966 258580 100028
rect 258540 96960 258592 96966
rect 258540 96902 258592 96908
rect 258736 96898 258764 100028
rect 258920 96937 258948 100028
rect 259104 97073 259132 100028
rect 259288 99618 259316 100028
rect 259276 99612 259328 99618
rect 259276 99554 259328 99560
rect 259564 97102 259592 100028
rect 259552 97096 259604 97102
rect 259090 97064 259146 97073
rect 259552 97038 259604 97044
rect 259090 96999 259146 97008
rect 259276 97028 259328 97034
rect 259276 96970 259328 96976
rect 259092 96960 259144 96966
rect 258906 96928 258962 96937
rect 258724 96892 258776 96898
rect 259092 96902 259144 96908
rect 258906 96863 258962 96872
rect 258724 96834 258776 96840
rect 258724 96756 258776 96762
rect 258724 96698 258776 96704
rect 258080 96144 258132 96150
rect 258080 96086 258132 96092
rect 257896 93424 257948 93430
rect 257896 93366 257948 93372
rect 258080 91792 258132 91798
rect 258080 91734 258132 91740
rect 256700 47592 256752 47598
rect 256700 47534 256752 47540
rect 257804 47592 257856 47598
rect 257804 47534 257856 47540
rect 255962 3360 256018 3369
rect 255962 3295 256018 3304
rect 256712 490 256740 47534
rect 258092 3874 258120 91734
rect 258172 84856 258224 84862
rect 258172 84798 258224 84804
rect 258080 3868 258132 3874
rect 258080 3810 258132 3816
rect 258184 3194 258212 84798
rect 258736 6526 258764 96698
rect 259104 70038 259132 96902
rect 259184 96892 259236 96898
rect 259184 96834 259236 96840
rect 259196 93362 259224 96834
rect 259184 93356 259236 93362
rect 259184 93298 259236 93304
rect 259288 87922 259316 96970
rect 259748 96966 259776 100028
rect 259932 99686 259960 100028
rect 259920 99680 259972 99686
rect 259920 99622 259972 99628
rect 260012 97232 260064 97238
rect 260012 97174 260064 97180
rect 259736 96960 259788 96966
rect 259736 96902 259788 96908
rect 260024 93854 260052 97174
rect 260116 96898 260144 100028
rect 260196 97776 260248 97782
rect 260196 97718 260248 97724
rect 260104 96892 260156 96898
rect 260104 96834 260156 96840
rect 260024 93826 260144 93854
rect 259276 87916 259328 87922
rect 259276 87858 259328 87864
rect 259460 72616 259512 72622
rect 259460 72558 259512 72564
rect 259092 70032 259144 70038
rect 259092 69974 259144 69980
rect 258724 6520 258776 6526
rect 258724 6462 258776 6468
rect 258264 3732 258316 3738
rect 258264 3674 258316 3680
rect 258172 3188 258224 3194
rect 258172 3130 258224 3136
rect 256896 598 257108 626
rect 256896 490 256924 598
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 256712 462 256924 490
rect 257080 480 257108 598
rect 258276 480 258304 3674
rect 259472 480 259500 72558
rect 260116 7614 260144 93826
rect 260208 7682 260236 97718
rect 260300 97510 260328 100028
rect 260288 97504 260340 97510
rect 260288 97446 260340 97452
rect 260288 97368 260340 97374
rect 260288 97310 260340 97316
rect 260300 75478 260328 97310
rect 260576 96937 260604 100028
rect 260760 97073 260788 100028
rect 260746 97064 260802 97073
rect 260746 96999 260802 97008
rect 260748 96960 260800 96966
rect 260562 96928 260618 96937
rect 260748 96902 260800 96908
rect 260562 96863 260618 96872
rect 260656 96892 260708 96898
rect 260656 96834 260708 96840
rect 260668 90710 260696 96834
rect 260656 90704 260708 90710
rect 260656 90646 260708 90652
rect 260288 75472 260340 75478
rect 260288 75414 260340 75420
rect 260760 11898 260788 96902
rect 260944 96898 260972 100028
rect 261128 97374 261156 100028
rect 261116 97368 261168 97374
rect 261116 97310 261168 97316
rect 261312 97034 261340 100028
rect 261300 97028 261352 97034
rect 261300 96970 261352 96976
rect 260932 96892 260984 96898
rect 260932 96834 260984 96840
rect 261588 96830 261616 100028
rect 261668 96960 261720 96966
rect 261668 96902 261720 96908
rect 261576 96824 261628 96830
rect 261576 96766 261628 96772
rect 261680 93854 261708 96902
rect 261772 96694 261800 100028
rect 261864 100014 261970 100042
rect 261760 96688 261812 96694
rect 261760 96630 261812 96636
rect 261680 93826 261800 93854
rect 260840 79348 260892 79354
rect 260840 79290 260892 79296
rect 260748 11892 260800 11898
rect 260748 11834 260800 11840
rect 260196 7676 260248 7682
rect 260196 7618 260248 7624
rect 260104 7608 260156 7614
rect 260104 7550 260156 7556
rect 259828 6316 259880 6322
rect 259828 6258 259880 6264
rect 259840 3262 259868 6258
rect 260852 3482 260880 79290
rect 261772 72758 261800 93826
rect 261864 85202 261892 100014
rect 262140 96966 262168 100028
rect 262128 96960 262180 96966
rect 262128 96902 262180 96908
rect 262036 96892 262088 96898
rect 262036 96834 262088 96840
rect 261944 96824 261996 96830
rect 261944 96766 261996 96772
rect 261852 85196 261904 85202
rect 261852 85138 261904 85144
rect 261956 79490 261984 96766
rect 262048 79558 262076 96834
rect 262324 96694 262352 100028
rect 262600 96966 262628 100028
rect 262588 96960 262640 96966
rect 262784 96937 262812 100028
rect 262982 100014 263088 100042
rect 262864 98184 262916 98190
rect 262864 98126 262916 98132
rect 262876 97714 262904 98126
rect 262864 97708 262916 97714
rect 262864 97650 262916 97656
rect 262864 97504 262916 97510
rect 262864 97446 262916 97452
rect 262588 96902 262640 96908
rect 262770 96928 262826 96937
rect 262770 96863 262826 96872
rect 262128 96688 262180 96694
rect 262128 96630 262180 96636
rect 262312 96688 262364 96694
rect 262312 96630 262364 96636
rect 262140 92070 262168 96630
rect 262128 92064 262180 92070
rect 262128 92006 262180 92012
rect 262876 79626 262904 97446
rect 262956 97028 263008 97034
rect 262956 96970 263008 96976
rect 262968 85270 262996 96970
rect 263060 96778 263088 100014
rect 263152 96898 263180 100028
rect 263336 96937 263364 100028
rect 263508 96960 263560 96966
rect 263322 96928 263378 96937
rect 263140 96892 263192 96898
rect 263508 96902 263560 96908
rect 263322 96863 263378 96872
rect 263140 96834 263192 96840
rect 263060 96750 263456 96778
rect 263324 96688 263376 96694
rect 263324 96630 263376 96636
rect 263336 93294 263364 96630
rect 263324 93288 263376 93294
rect 263324 93230 263376 93236
rect 263428 92002 263456 96750
rect 263416 91996 263468 92002
rect 263416 91938 263468 91944
rect 262956 85264 263008 85270
rect 262956 85206 263008 85212
rect 262864 79620 262916 79626
rect 262864 79562 262916 79568
rect 262036 79552 262088 79558
rect 262036 79494 262088 79500
rect 261944 79484 261996 79490
rect 261944 79426 261996 79432
rect 262220 78056 262272 78062
rect 262220 77998 262272 78004
rect 261760 72752 261812 72758
rect 261760 72694 261812 72700
rect 262232 16574 262260 77998
rect 263520 72690 263548 96902
rect 263612 94586 263640 100028
rect 263796 97510 263824 100028
rect 263784 97504 263836 97510
rect 263784 97446 263836 97452
rect 263980 96898 264008 100028
rect 264164 96966 264192 100028
rect 264244 97096 264296 97102
rect 264244 97038 264296 97044
rect 264152 96960 264204 96966
rect 264152 96902 264204 96908
rect 263968 96892 264020 96898
rect 263968 96834 264020 96840
rect 263600 94580 263652 94586
rect 263600 94522 263652 94528
rect 263600 76560 263652 76566
rect 263600 76502 263652 76508
rect 263508 72684 263560 72690
rect 263508 72626 263560 72632
rect 262864 28280 262916 28286
rect 262864 28222 262916 28228
rect 262232 16546 262536 16574
rect 260668 3454 260880 3482
rect 259828 3256 259880 3262
rect 259828 3198 259880 3204
rect 260668 480 260696 3454
rect 261760 3256 261812 3262
rect 261760 3198 261812 3204
rect 261772 480 261800 3198
rect 262508 490 262536 16546
rect 262876 3806 262904 28222
rect 263612 16574 263640 76502
rect 264256 75410 264284 97038
rect 264348 96937 264376 100028
rect 264624 97102 264652 100028
rect 264612 97096 264664 97102
rect 264808 97073 264836 100028
rect 264992 97782 265020 100028
rect 264980 97776 265032 97782
rect 264980 97718 265032 97724
rect 264612 97038 264664 97044
rect 264794 97064 264850 97073
rect 264794 96999 264850 97008
rect 264704 96960 264756 96966
rect 264334 96928 264390 96937
rect 264704 96902 264756 96908
rect 264334 96863 264390 96872
rect 264336 96824 264388 96830
rect 264336 96766 264388 96772
rect 264348 85134 264376 96766
rect 264336 85128 264388 85134
rect 264336 85070 264388 85076
rect 264244 75404 264296 75410
rect 264244 75346 264296 75352
rect 263612 16546 264192 16574
rect 262864 3800 262916 3806
rect 262864 3742 262916 3748
rect 262784 598 262996 626
rect 262784 490 262812 598
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262508 462 262812 490
rect 262968 480 262996 598
rect 264164 480 264192 16546
rect 264716 9314 264744 96902
rect 264796 96892 264848 96898
rect 264796 96834 264848 96840
rect 264808 11830 264836 96834
rect 265176 96830 265204 100028
rect 265360 97578 265388 100028
rect 265348 97572 265400 97578
rect 265348 97514 265400 97520
rect 265636 96966 265664 100028
rect 265624 96960 265676 96966
rect 265624 96902 265676 96908
rect 265820 96898 265848 100028
rect 265900 97096 265952 97102
rect 265900 97038 265952 97044
rect 265808 96892 265860 96898
rect 265808 96834 265860 96840
rect 265164 96824 265216 96830
rect 265164 96766 265216 96772
rect 265912 94790 265940 97038
rect 265900 94784 265952 94790
rect 265900 94726 265952 94732
rect 266004 91934 266032 100028
rect 266084 96960 266136 96966
rect 266188 96937 266216 100028
rect 266084 96902 266136 96908
rect 266174 96928 266230 96937
rect 265992 91928 266044 91934
rect 265992 91870 266044 91876
rect 266096 85066 266124 96902
rect 266174 96863 266230 96872
rect 266268 96892 266320 96898
rect 266268 96834 266320 96840
rect 266176 96824 266228 96830
rect 266176 96766 266228 96772
rect 266084 85060 266136 85066
rect 266084 85002 266136 85008
rect 266188 69970 266216 96766
rect 266176 69964 266228 69970
rect 266176 69906 266228 69912
rect 266280 14550 266308 96834
rect 266372 96762 266400 100028
rect 266648 96966 266676 100028
rect 266636 96960 266688 96966
rect 266636 96902 266688 96908
rect 266832 96898 266860 100028
rect 267030 100014 267136 100042
rect 266820 96892 266872 96898
rect 266820 96834 266872 96840
rect 266360 96756 266412 96762
rect 266360 96698 266412 96704
rect 267108 93854 267136 100014
rect 267200 96830 267228 100028
rect 267476 97073 267504 100028
rect 267462 97064 267518 97073
rect 267462 96999 267518 97008
rect 267372 96960 267424 96966
rect 267660 96937 267688 100028
rect 267844 98802 267872 100028
rect 267832 98796 267884 98802
rect 267832 98738 267884 98744
rect 268028 97170 268056 100028
rect 268016 97164 268068 97170
rect 268016 97106 268068 97112
rect 267372 96902 267424 96908
rect 267646 96928 267702 96937
rect 267188 96824 267240 96830
rect 267188 96766 267240 96772
rect 267108 93826 267320 93854
rect 266360 78124 266412 78130
rect 266360 78066 266412 78072
rect 266372 16574 266400 78066
rect 267004 71052 267056 71058
rect 267004 70994 267056 71000
rect 266372 16546 266584 16574
rect 266268 14544 266320 14550
rect 266268 14486 266320 14492
rect 264796 11824 264848 11830
rect 264796 11766 264848 11772
rect 264704 9308 264756 9314
rect 264704 9250 264756 9256
rect 265348 3596 265400 3602
rect 265348 3538 265400 3544
rect 265360 480 265388 3538
rect 266556 480 266584 16546
rect 267016 3602 267044 70994
rect 267292 68406 267320 93826
rect 267384 86494 267412 96902
rect 267556 96892 267608 96898
rect 267646 96863 267702 96872
rect 267556 96834 267608 96840
rect 267464 96756 267516 96762
rect 267464 96698 267516 96704
rect 267372 86488 267424 86494
rect 267372 86430 267424 86436
rect 267476 78198 267504 96698
rect 267464 78192 267516 78198
rect 267464 78134 267516 78140
rect 267568 71262 267596 96834
rect 268212 96830 268240 100028
rect 268502 100014 268608 100042
rect 268686 100014 268792 100042
rect 268870 100014 268976 100042
rect 268384 97504 268436 97510
rect 268384 97446 268436 97452
rect 267648 96824 267700 96830
rect 267648 96766 267700 96772
rect 268200 96824 268252 96830
rect 268200 96766 268252 96772
rect 267660 91798 267688 96766
rect 267648 91792 267700 91798
rect 267648 91734 267700 91740
rect 267832 77988 267884 77994
rect 267832 77930 267884 77936
rect 267556 71256 267608 71262
rect 267556 71198 267608 71204
rect 267280 68400 267332 68406
rect 267280 68342 267332 68348
rect 267740 42084 267792 42090
rect 267740 42026 267792 42032
rect 267004 3596 267056 3602
rect 267004 3538 267056 3544
rect 267752 3482 267780 42026
rect 267844 3670 267872 77930
rect 268396 16574 268424 97446
rect 268580 87854 268608 100014
rect 268764 96914 268792 100014
rect 268764 96886 268884 96914
rect 268568 87848 268620 87854
rect 268568 87790 268620 87796
rect 268856 83842 268884 96886
rect 268844 83836 268896 83842
rect 268844 83778 268896 83784
rect 268948 78130 268976 100014
rect 269040 96937 269068 100028
rect 269026 96928 269082 96937
rect 269026 96863 269082 96872
rect 269224 96830 269252 100028
rect 269500 96966 269528 100028
rect 269488 96960 269540 96966
rect 269488 96902 269540 96908
rect 269684 96898 269712 100028
rect 269882 100014 269988 100042
rect 269764 97572 269816 97578
rect 269764 97514 269816 97520
rect 269672 96892 269724 96898
rect 269672 96834 269724 96840
rect 269028 96824 269080 96830
rect 269028 96766 269080 96772
rect 269212 96824 269264 96830
rect 269212 96766 269264 96772
rect 268936 78124 268988 78130
rect 268936 78066 268988 78072
rect 269040 42090 269068 96766
rect 269776 91866 269804 97514
rect 269960 93854 269988 100014
rect 270052 96762 270080 100028
rect 270236 96937 270264 100028
rect 270408 96960 270460 96966
rect 270222 96928 270278 96937
rect 270408 96902 270460 96908
rect 270222 96863 270278 96872
rect 270316 96892 270368 96898
rect 270316 96834 270368 96840
rect 270224 96824 270276 96830
rect 270224 96766 270276 96772
rect 270040 96756 270092 96762
rect 270040 96698 270092 96704
rect 269960 93826 270172 93854
rect 269764 91860 269816 91866
rect 269764 91802 269816 91808
rect 270144 83774 270172 93826
rect 270132 83768 270184 83774
rect 270132 83710 270184 83716
rect 269212 75200 269264 75206
rect 269212 75142 269264 75148
rect 269028 42084 269080 42090
rect 269028 42026 269080 42032
rect 268396 16546 268516 16574
rect 268488 3670 268516 16546
rect 269224 3738 269252 75142
rect 270236 71194 270264 96766
rect 270224 71188 270276 71194
rect 270224 71130 270276 71136
rect 270328 9246 270356 96834
rect 270316 9240 270368 9246
rect 270316 9182 270368 9188
rect 270420 7614 270448 96902
rect 270512 96830 270540 100028
rect 270696 96966 270724 100028
rect 270880 97034 270908 100028
rect 270868 97028 270920 97034
rect 270868 96970 270920 96976
rect 270684 96960 270736 96966
rect 270684 96902 270736 96908
rect 271064 96898 271092 100028
rect 271248 96937 271276 100028
rect 271538 100014 271644 100042
rect 271616 97050 271644 100014
rect 271708 97209 271736 100028
rect 271694 97200 271750 97209
rect 271694 97135 271750 97144
rect 271512 97028 271564 97034
rect 271616 97022 271828 97050
rect 271512 96970 271564 96976
rect 271420 96960 271472 96966
rect 271234 96928 271290 96937
rect 271052 96892 271104 96898
rect 271420 96902 271472 96908
rect 271234 96863 271290 96872
rect 271052 96834 271104 96840
rect 270500 96824 270552 96830
rect 270500 96766 270552 96772
rect 271432 10334 271460 96902
rect 271524 90642 271552 96970
rect 271604 96892 271656 96898
rect 271604 96834 271656 96840
rect 271512 90636 271564 90642
rect 271512 90578 271564 90584
rect 271616 83706 271644 96834
rect 271696 96824 271748 96830
rect 271696 96766 271748 96772
rect 271604 83700 271656 83706
rect 271604 83642 271656 83648
rect 271708 71126 271736 96766
rect 271800 90574 271828 97022
rect 271892 96898 271920 100028
rect 271880 96892 271932 96898
rect 271880 96834 271932 96840
rect 272076 94722 272104 100028
rect 272260 96966 272288 100028
rect 272550 100014 272656 100042
rect 272734 100014 272840 100042
rect 272248 96960 272300 96966
rect 272248 96902 272300 96908
rect 272064 94716 272116 94722
rect 272064 94658 272116 94664
rect 272628 93854 272656 100014
rect 272812 96914 272840 100014
rect 272904 97073 272932 100028
rect 273088 97646 273116 100028
rect 273076 97640 273128 97646
rect 273076 97582 273128 97588
rect 272890 97064 272946 97073
rect 272890 96999 272946 97008
rect 273076 96960 273128 96966
rect 272812 96886 272932 96914
rect 273076 96902 273128 96908
rect 272628 93826 272840 93854
rect 271788 90568 271840 90574
rect 271788 90510 271840 90516
rect 271696 71120 271748 71126
rect 271696 71062 271748 71068
rect 272812 66910 272840 93826
rect 272904 80986 272932 96886
rect 272984 96892 273036 96898
rect 272984 96834 273036 96840
rect 272892 80980 272944 80986
rect 272892 80922 272944 80928
rect 272996 77994 273024 96834
rect 272984 77988 273036 77994
rect 272984 77930 273036 77936
rect 273088 74186 273116 96902
rect 273272 96898 273300 100028
rect 273260 96892 273312 96898
rect 273260 96834 273312 96840
rect 273548 96694 273576 100028
rect 273746 100014 273852 100042
rect 273536 96688 273588 96694
rect 273536 96630 273588 96636
rect 273824 93854 273852 100014
rect 273916 96966 273944 100028
rect 274114 100014 274220 100042
rect 273904 96960 273956 96966
rect 273904 96902 273956 96908
rect 274088 96892 274140 96898
rect 274088 96834 274140 96840
rect 274100 96642 274128 96834
rect 274192 96778 274220 100014
rect 274284 96937 274312 100028
rect 274560 97073 274588 100028
rect 274744 97238 274772 100028
rect 274732 97232 274784 97238
rect 274732 97174 274784 97180
rect 274546 97064 274602 97073
rect 274546 96999 274602 97008
rect 274548 96960 274600 96966
rect 274270 96928 274326 96937
rect 274548 96902 274600 96908
rect 274270 96863 274326 96872
rect 274192 96750 274496 96778
rect 274364 96688 274416 96694
rect 274100 96614 274312 96642
rect 274364 96630 274416 96636
rect 273824 93826 274220 93854
rect 273076 74180 273128 74186
rect 273076 74122 273128 74128
rect 272800 66904 272852 66910
rect 272800 66846 272852 66852
rect 274192 53106 274220 93826
rect 274284 90506 274312 96614
rect 274272 90500 274324 90506
rect 274272 90442 274324 90448
rect 274376 72554 274404 96630
rect 274364 72548 274416 72554
rect 274364 72490 274416 72496
rect 274468 69902 274496 96750
rect 274560 90438 274588 96902
rect 274928 96762 274956 100028
rect 275112 96830 275140 100028
rect 275284 97368 275336 97374
rect 275284 97310 275336 97316
rect 275296 96914 275324 97310
rect 275388 97102 275416 100028
rect 275586 100014 275692 100042
rect 275376 97096 275428 97102
rect 275376 97038 275428 97044
rect 275664 96914 275692 100014
rect 275756 97918 275784 100028
rect 275744 97912 275796 97918
rect 275744 97854 275796 97860
rect 275940 97073 275968 100028
rect 275926 97064 275982 97073
rect 276124 97034 276152 100028
rect 275926 96999 275982 97008
rect 276112 97028 276164 97034
rect 276112 96970 276164 96976
rect 275296 96886 275416 96914
rect 275664 96886 275968 96914
rect 276400 96898 276428 100028
rect 276584 96966 276612 100028
rect 276768 97510 276796 100028
rect 276756 97504 276808 97510
rect 276756 97446 276808 97452
rect 276756 97164 276808 97170
rect 276756 97106 276808 97112
rect 276664 97096 276716 97102
rect 276664 97038 276716 97044
rect 276572 96960 276624 96966
rect 276572 96902 276624 96908
rect 275100 96824 275152 96830
rect 275100 96766 275152 96772
rect 274916 96756 274968 96762
rect 274916 96698 274968 96704
rect 275284 96688 275336 96694
rect 275284 96630 275336 96636
rect 274548 90432 274600 90438
rect 274548 90374 274600 90380
rect 275296 78062 275324 96630
rect 275388 92138 275416 96886
rect 275744 96824 275796 96830
rect 275744 96766 275796 96772
rect 275376 92132 275428 92138
rect 275376 92074 275428 92080
rect 275756 90370 275784 96766
rect 275836 96756 275888 96762
rect 275836 96698 275888 96704
rect 275744 90364 275796 90370
rect 275744 90306 275796 90312
rect 275284 78056 275336 78062
rect 275284 77998 275336 78004
rect 274456 69896 274508 69902
rect 274456 69838 274508 69844
rect 275848 68338 275876 96698
rect 275836 68332 275888 68338
rect 275836 68274 275888 68280
rect 275940 62830 275968 96886
rect 276388 96892 276440 96898
rect 276388 96834 276440 96840
rect 276676 69834 276704 97038
rect 276768 72622 276796 97106
rect 276952 96937 276980 100028
rect 277136 97578 277164 100028
rect 277124 97572 277176 97578
rect 277124 97514 277176 97520
rect 277412 97209 277440 100028
rect 277398 97200 277454 97209
rect 277398 97135 277454 97144
rect 277308 97028 277360 97034
rect 277308 96970 277360 96976
rect 277124 96960 277176 96966
rect 276938 96928 276994 96937
rect 277124 96902 277176 96908
rect 276938 96863 276994 96872
rect 277136 83570 277164 96902
rect 277216 96892 277268 96898
rect 277216 96834 277268 96840
rect 277124 83564 277176 83570
rect 277124 83506 277176 83512
rect 277228 76702 277256 96834
rect 277216 76696 277268 76702
rect 277216 76638 277268 76644
rect 276756 72616 276808 72622
rect 276756 72558 276808 72564
rect 276664 69828 276716 69834
rect 276664 69770 276716 69776
rect 276112 69692 276164 69698
rect 276112 69634 276164 69640
rect 275928 62824 275980 62830
rect 275282 62792 275338 62801
rect 275928 62766 275980 62772
rect 275282 62727 275338 62736
rect 274180 53100 274232 53106
rect 274180 53042 274232 53048
rect 273260 51740 273312 51746
rect 273260 51682 273312 51688
rect 271420 10328 271472 10334
rect 271420 10270 271472 10276
rect 270040 7608 270092 7614
rect 270040 7550 270092 7556
rect 270408 7608 270460 7614
rect 270408 7550 270460 7556
rect 269212 3732 269264 3738
rect 269212 3674 269264 3680
rect 267832 3664 267884 3670
rect 267832 3606 267884 3612
rect 268476 3664 268528 3670
rect 268476 3606 268528 3612
rect 267752 3454 268424 3482
rect 267832 3392 267884 3398
rect 267832 3334 267884 3340
rect 267844 626 267872 3334
rect 267752 598 267872 626
rect 267752 480 267780 598
rect 268396 490 268424 3454
rect 268672 598 268884 626
rect 268672 490 268700 598
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268396 462 268700 490
rect 268856 480 268884 598
rect 270052 480 270080 7550
rect 271236 3800 271288 3806
rect 271236 3742 271288 3748
rect 271248 480 271276 3742
rect 272432 3528 272484 3534
rect 272432 3470 272484 3476
rect 272444 480 272472 3470
rect 273272 3398 273300 51682
rect 273626 6216 273682 6225
rect 273626 6151 273682 6160
rect 273260 3392 273312 3398
rect 273260 3334 273312 3340
rect 273640 480 273668 6151
rect 275296 3466 275324 62727
rect 276124 6914 276152 69634
rect 277320 17270 277348 96970
rect 277596 96694 277624 100028
rect 277780 96966 277808 100028
rect 277768 96960 277820 96966
rect 277768 96902 277820 96908
rect 277964 96898 277992 100028
rect 278162 100014 278360 100042
rect 278438 100014 278544 100042
rect 277952 96892 278004 96898
rect 277952 96834 278004 96840
rect 277584 96688 277636 96694
rect 277584 96630 277636 96636
rect 278332 89214 278360 100014
rect 278412 96960 278464 96966
rect 278412 96902 278464 96908
rect 278320 89208 278372 89214
rect 278320 89150 278372 89156
rect 278424 84998 278452 96902
rect 278516 96778 278544 100014
rect 278608 96937 278636 100028
rect 278792 98054 278820 100028
rect 278780 98048 278832 98054
rect 278780 97990 278832 97996
rect 278594 96928 278650 96937
rect 278976 96898 279004 100028
rect 279174 100014 279372 100042
rect 279450 100014 279556 100042
rect 279634 100014 279740 100042
rect 279344 97730 279372 100014
rect 279344 97702 279464 97730
rect 279436 97646 279464 97702
rect 279332 97640 279384 97646
rect 279332 97582 279384 97588
rect 279424 97640 279476 97646
rect 279424 97582 279476 97588
rect 278594 96863 278650 96872
rect 278688 96892 278740 96898
rect 278688 96834 278740 96840
rect 278964 96892 279016 96898
rect 278964 96834 279016 96840
rect 278516 96750 278636 96778
rect 278504 96688 278556 96694
rect 278504 96630 278556 96636
rect 278412 84992 278464 84998
rect 278412 84934 278464 84940
rect 278516 76770 278544 96630
rect 278504 76764 278556 76770
rect 278504 76706 278556 76712
rect 278608 69766 278636 96750
rect 278596 69760 278648 69766
rect 278596 69702 278648 69708
rect 278700 19990 278728 96834
rect 279344 93854 279372 97582
rect 279424 97232 279476 97238
rect 279424 97174 279476 97180
rect 279436 96642 279464 97174
rect 279528 96778 279556 100014
rect 279712 96948 279740 100014
rect 279804 97510 279832 100028
rect 279792 97504 279844 97510
rect 279792 97446 279844 97452
rect 279988 97073 280016 100028
rect 279974 97064 280030 97073
rect 279974 96999 280030 97008
rect 280172 96966 280200 100028
rect 280160 96960 280212 96966
rect 279712 96920 280016 96948
rect 279528 96750 279924 96778
rect 279436 96614 279556 96642
rect 279344 93826 279464 93854
rect 278780 82136 278832 82142
rect 278780 82078 278832 82084
rect 278688 19984 278740 19990
rect 278688 19926 278740 19932
rect 277308 17264 277360 17270
rect 277308 17206 277360 17212
rect 276032 6886 276152 6914
rect 274824 3460 274876 3466
rect 274824 3402 274876 3408
rect 275284 3460 275336 3466
rect 275284 3402 275336 3408
rect 274836 480 274864 3402
rect 276032 480 276060 6886
rect 277124 3596 277176 3602
rect 277124 3538 277176 3544
rect 277136 480 277164 3538
rect 278792 3534 278820 82078
rect 279436 76634 279464 93826
rect 279528 83638 279556 96614
rect 279896 89146 279924 96750
rect 279884 89140 279936 89146
rect 279884 89082 279936 89088
rect 279516 83632 279568 83638
rect 279516 83574 279568 83580
rect 279988 82414 280016 96920
rect 280160 96902 280212 96908
rect 280068 96892 280120 96898
rect 280068 96834 280120 96840
rect 279976 82408 280028 82414
rect 279976 82350 280028 82356
rect 279424 76628 279476 76634
rect 279424 76570 279476 76576
rect 280080 69698 280108 96834
rect 280448 96762 280476 100028
rect 280632 96830 280660 100028
rect 280712 97912 280764 97918
rect 280712 97854 280764 97860
rect 280620 96824 280672 96830
rect 280620 96766 280672 96772
rect 280436 96756 280488 96762
rect 280436 96698 280488 96704
rect 280724 90409 280752 97854
rect 280816 96898 280844 100028
rect 281000 97850 281028 100028
rect 280988 97844 281040 97850
rect 280988 97786 281040 97792
rect 281184 96937 281212 100028
rect 281356 96960 281408 96966
rect 281170 96928 281226 96937
rect 280804 96892 280856 96898
rect 281460 96937 281488 100028
rect 281356 96902 281408 96908
rect 281446 96928 281502 96937
rect 281170 96863 281226 96872
rect 281264 96892 281316 96898
rect 280804 96834 280856 96840
rect 281264 96834 281316 96840
rect 281172 96824 281224 96830
rect 281172 96766 281224 96772
rect 280710 90400 280766 90409
rect 280710 90335 280766 90344
rect 281184 89282 281212 96766
rect 281172 89276 281224 89282
rect 281172 89218 281224 89224
rect 281276 82346 281304 96834
rect 281264 82340 281316 82346
rect 281264 82282 281316 82288
rect 281368 71058 281396 96902
rect 281446 96863 281502 96872
rect 281644 96830 281672 100028
rect 281828 96966 281856 100028
rect 281816 96960 281868 96966
rect 281816 96902 281868 96908
rect 282012 96898 282040 100028
rect 282210 100014 282408 100042
rect 282380 97374 282408 100014
rect 282472 98666 282500 100028
rect 282670 100014 282776 100042
rect 282460 98660 282512 98666
rect 282460 98602 282512 98608
rect 282368 97368 282420 97374
rect 282368 97310 282420 97316
rect 282184 97300 282236 97306
rect 282184 97242 282236 97248
rect 282000 96892 282052 96898
rect 282000 96834 282052 96840
rect 281632 96824 281684 96830
rect 281632 96766 281684 96772
rect 281448 96756 281500 96762
rect 281448 96698 281500 96704
rect 281356 71052 281408 71058
rect 281356 70994 281408 71000
rect 280068 69692 280120 69698
rect 280068 69634 280120 69640
rect 281460 51746 281488 96698
rect 282196 92206 282224 97242
rect 282460 96960 282512 96966
rect 282460 96902 282512 96908
rect 282184 92200 282236 92206
rect 282184 92142 282236 92148
rect 282472 89078 282500 96902
rect 282644 96892 282696 96898
rect 282644 96834 282696 96840
rect 282550 91216 282606 91225
rect 282550 91151 282606 91160
rect 282460 89072 282512 89078
rect 282460 89014 282512 89020
rect 281540 89004 281592 89010
rect 281540 88946 281592 88952
rect 281448 51740 281500 51746
rect 281448 51682 281500 51688
rect 280712 6248 280764 6254
rect 280712 6190 280764 6196
rect 278320 3528 278372 3534
rect 278320 3470 278372 3476
rect 278780 3528 278832 3534
rect 278780 3470 278832 3476
rect 279516 3528 279568 3534
rect 279516 3470 279568 3476
rect 278332 480 278360 3470
rect 279528 480 279556 3470
rect 280724 480 280752 6190
rect 281552 3534 281580 88946
rect 282564 79422 282592 91151
rect 282656 82482 282684 96834
rect 282644 82476 282696 82482
rect 282644 82418 282696 82424
rect 282552 79416 282604 79422
rect 282552 79358 282604 79364
rect 282748 75342 282776 100014
rect 282840 96937 282868 100028
rect 283024 97889 283052 100028
rect 283010 97880 283066 97889
rect 283010 97815 283066 97824
rect 283208 96966 283236 100028
rect 283380 99000 283432 99006
rect 283380 98942 283432 98948
rect 283196 96960 283248 96966
rect 282826 96928 282882 96937
rect 283196 96902 283248 96908
rect 282826 96863 282882 96872
rect 282828 96824 282880 96830
rect 282828 96766 282880 96772
rect 282736 75336 282788 75342
rect 282736 75278 282788 75284
rect 282840 21418 282868 96766
rect 283392 93854 283420 98942
rect 283484 96694 283512 100028
rect 283668 98734 283696 100028
rect 283866 100014 283972 100042
rect 283656 98728 283708 98734
rect 283656 98670 283708 98676
rect 283564 98048 283616 98054
rect 283564 97990 283616 97996
rect 283472 96688 283524 96694
rect 283472 96630 283524 96636
rect 283392 93826 283512 93854
rect 282828 21412 282880 21418
rect 282828 21354 282880 21360
rect 283484 5574 283512 93826
rect 283576 93158 283604 97990
rect 283840 96960 283892 96966
rect 283840 96902 283892 96908
rect 283564 93152 283616 93158
rect 283564 93094 283616 93100
rect 283852 89010 283880 96902
rect 283944 96778 283972 100014
rect 284036 96937 284064 100028
rect 284312 98841 284340 100028
rect 284298 98832 284354 98841
rect 284298 98767 284354 98776
rect 284022 96928 284078 96937
rect 284022 96863 284078 96872
rect 284496 96830 284524 100028
rect 284484 96824 284536 96830
rect 283944 96750 284248 96778
rect 284484 96766 284536 96772
rect 284680 96762 284708 100028
rect 284864 98977 284892 100028
rect 285062 100014 285260 100042
rect 285338 100014 285444 100042
rect 285522 100014 285628 100042
rect 284850 98968 284906 98977
rect 284850 98903 284906 98912
rect 285232 96948 285260 100014
rect 285416 96948 285444 100014
rect 285232 96920 285352 96948
rect 285416 96920 285536 96948
rect 285220 96824 285272 96830
rect 285220 96766 285272 96772
rect 284116 96688 284168 96694
rect 284116 96630 284168 96636
rect 283840 89004 283892 89010
rect 283840 88946 283892 88952
rect 284128 82278 284156 96630
rect 284116 82272 284168 82278
rect 284116 82214 284168 82220
rect 284220 75274 284248 96750
rect 284668 96756 284720 96762
rect 284668 96698 284720 96704
rect 284208 75268 284260 75274
rect 284208 75210 284260 75216
rect 285232 75206 285260 96766
rect 285220 75200 285272 75206
rect 285220 75142 285272 75148
rect 285324 74118 285352 96920
rect 285404 96756 285456 96762
rect 285404 96698 285456 96704
rect 285312 74112 285364 74118
rect 285312 74054 285364 74060
rect 285416 65550 285444 96698
rect 285404 65544 285456 65550
rect 285404 65486 285456 65492
rect 285508 13122 285536 96920
rect 285496 13116 285548 13122
rect 285496 13058 285548 13064
rect 285600 6390 285628 100014
rect 285692 96898 285720 100028
rect 285772 98048 285824 98054
rect 285772 97990 285824 97996
rect 285784 97889 285812 97990
rect 285770 97880 285826 97889
rect 285770 97815 285826 97824
rect 285680 96892 285732 96898
rect 285680 96834 285732 96840
rect 285876 96830 285904 100028
rect 285864 96824 285916 96830
rect 285864 96766 285916 96772
rect 286060 96082 286088 100028
rect 286336 96966 286364 100028
rect 286534 100014 286640 100042
rect 286324 96960 286376 96966
rect 286324 96902 286376 96908
rect 286048 96076 286100 96082
rect 286048 96018 286100 96024
rect 285680 87712 285732 87718
rect 285680 87654 285732 87660
rect 285588 6384 285640 6390
rect 285588 6326 285640 6332
rect 281908 5568 281960 5574
rect 281908 5510 281960 5516
rect 283472 5568 283524 5574
rect 283472 5510 283524 5516
rect 281540 3528 281592 3534
rect 281540 3470 281592 3476
rect 281920 480 281948 5510
rect 284300 3528 284352 3534
rect 284300 3470 284352 3476
rect 283104 2984 283156 2990
rect 283104 2926 283156 2932
rect 283116 480 283144 2926
rect 284312 480 284340 3470
rect 285402 3360 285458 3369
rect 285402 3295 285458 3304
rect 285416 480 285444 3295
rect 285692 2990 285720 87654
rect 286612 46238 286640 100014
rect 286704 99550 286732 100028
rect 286692 99544 286744 99550
rect 286692 99486 286744 99492
rect 286692 96960 286744 96966
rect 286888 96937 286916 100028
rect 286692 96902 286744 96908
rect 286874 96928 286930 96937
rect 286704 87718 286732 96902
rect 286784 96892 286836 96898
rect 287072 96898 287100 100028
rect 286874 96863 286930 96872
rect 287060 96892 287112 96898
rect 286784 96834 286836 96840
rect 287060 96834 287112 96840
rect 286692 87712 286744 87718
rect 286692 87654 286744 87660
rect 286796 84862 286824 96834
rect 286876 96824 286928 96830
rect 286876 96766 286928 96772
rect 286784 84856 286836 84862
rect 286784 84798 286836 84804
rect 286888 82210 286916 96766
rect 287348 96014 287376 100028
rect 287532 96966 287560 100028
rect 287730 100014 287836 100042
rect 287520 96960 287572 96966
rect 287520 96902 287572 96908
rect 287336 96008 287388 96014
rect 287336 95950 287388 95956
rect 287808 93854 287836 100014
rect 287900 99482 287928 100028
rect 288098 100014 288296 100042
rect 287888 99476 287940 99482
rect 287888 99418 287940 99424
rect 288072 96960 288124 96966
rect 288072 96902 288124 96908
rect 287978 95840 288034 95849
rect 287978 95775 288034 95784
rect 287992 95130 288020 95775
rect 287980 95124 288032 95130
rect 287980 95066 288032 95072
rect 287808 93826 288020 93854
rect 287060 87644 287112 87650
rect 287060 87586 287112 87592
rect 286876 82204 286928 82210
rect 286876 82146 286928 82152
rect 285772 46232 285824 46238
rect 285772 46174 285824 46180
rect 286600 46232 286652 46238
rect 286600 46174 286652 46180
rect 285784 3534 285812 46174
rect 287072 16574 287100 87586
rect 287072 16546 287376 16574
rect 286600 6180 286652 6186
rect 286600 6122 286652 6128
rect 285772 3528 285824 3534
rect 285772 3470 285824 3476
rect 285680 2984 285732 2990
rect 285680 2926 285732 2932
rect 286612 480 286640 6122
rect 287348 490 287376 16546
rect 287992 9110 288020 93826
rect 288084 87786 288112 96902
rect 288164 96892 288216 96898
rect 288164 96834 288216 96840
rect 288072 87780 288124 87786
rect 288072 87722 288124 87728
rect 288176 84930 288204 96834
rect 288164 84924 288216 84930
rect 288164 84866 288216 84872
rect 288268 74050 288296 100014
rect 288360 96937 288388 100028
rect 288346 96928 288402 96937
rect 288346 96863 288402 96872
rect 288544 95946 288572 100028
rect 288728 96966 288756 100028
rect 288716 96960 288768 96966
rect 288716 96902 288768 96908
rect 288912 96830 288940 100028
rect 289096 99414 289124 100028
rect 289084 99408 289136 99414
rect 289084 99350 289136 99356
rect 288900 96824 288952 96830
rect 288900 96766 288952 96772
rect 288532 95940 288584 95946
rect 288532 95882 288584 95888
rect 289084 94512 289136 94518
rect 289084 94454 289136 94460
rect 288256 74044 288308 74050
rect 288256 73986 288308 73992
rect 287980 9104 288032 9110
rect 287980 9046 288032 9052
rect 288992 3460 289044 3466
rect 288992 3402 289044 3408
rect 287624 598 287836 626
rect 287624 490 287652 598
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287348 462 287652 490
rect 287808 480 287836 598
rect 289004 480 289032 3402
rect 289096 2922 289124 94454
rect 289372 9042 289400 100028
rect 289452 96960 289504 96966
rect 289452 96902 289504 96908
rect 289464 87650 289492 96902
rect 289452 87644 289504 87650
rect 289452 87586 289504 87592
rect 289556 73982 289584 100028
rect 289636 96824 289688 96830
rect 289636 96766 289688 96772
rect 289544 73976 289596 73982
rect 289544 73918 289596 73924
rect 289648 14482 289676 96766
rect 289740 95985 289768 100028
rect 289924 96898 289952 100028
rect 290108 96966 290136 100028
rect 290096 96960 290148 96966
rect 290096 96902 290148 96908
rect 289912 96892 289964 96898
rect 289912 96834 289964 96840
rect 290384 96694 290412 100028
rect 290568 96830 290596 100028
rect 290752 97034 290780 100028
rect 290936 99657 290964 100028
rect 291028 100014 291134 100042
rect 290922 99648 290978 99657
rect 290922 99583 290978 99592
rect 290740 97028 290792 97034
rect 290740 96970 290792 96976
rect 290832 96960 290884 96966
rect 291028 96948 291056 100014
rect 291108 97028 291160 97034
rect 291108 96970 291160 96976
rect 290832 96902 290884 96908
rect 290936 96920 291056 96948
rect 290740 96892 290792 96898
rect 290740 96834 290792 96840
rect 290556 96824 290608 96830
rect 290556 96766 290608 96772
rect 290372 96688 290424 96694
rect 290372 96630 290424 96636
rect 289726 95976 289782 95985
rect 289726 95911 289782 95920
rect 290752 87689 290780 96834
rect 290738 87680 290794 87689
rect 290738 87615 290794 87624
rect 290844 86426 290872 96902
rect 290832 86420 290884 86426
rect 290832 86362 290884 86368
rect 290936 82142 290964 96920
rect 291016 96824 291068 96830
rect 291016 96766 291068 96772
rect 290924 82136 290976 82142
rect 290924 82078 290976 82084
rect 291028 73914 291056 96766
rect 291016 73908 291068 73914
rect 291016 73850 291068 73856
rect 291120 24138 291148 96970
rect 291396 96694 291424 100028
rect 291580 98705 291608 100028
rect 291566 98696 291622 98705
rect 291566 98631 291622 98640
rect 291660 97844 291712 97850
rect 291660 97786 291712 97792
rect 291672 97442 291700 97786
rect 291660 97436 291712 97442
rect 291660 97378 291712 97384
rect 291764 96966 291792 100028
rect 291752 96960 291804 96966
rect 291752 96902 291804 96908
rect 291948 96898 291976 100028
rect 291936 96892 291988 96898
rect 291936 96834 291988 96840
rect 291200 96688 291252 96694
rect 291200 96630 291252 96636
rect 291384 96688 291436 96694
rect 291384 96630 291436 96636
rect 291212 95849 291240 96630
rect 291198 95840 291254 95849
rect 291198 95775 291254 95784
rect 291200 80844 291252 80850
rect 291200 80786 291252 80792
rect 291108 24132 291160 24138
rect 291108 24074 291160 24080
rect 291212 16574 291240 80786
rect 292224 39370 292252 100028
rect 292408 96937 292436 100028
rect 292592 97481 292620 100028
rect 292578 97472 292634 97481
rect 292578 97407 292634 97416
rect 292776 96966 292804 100028
rect 292488 96960 292540 96966
rect 292394 96928 292450 96937
rect 292304 96892 292356 96898
rect 292488 96902 292540 96908
rect 292764 96960 292816 96966
rect 292764 96902 292816 96908
rect 292394 96863 292450 96872
rect 292304 96834 292356 96840
rect 292316 80918 292344 96834
rect 292396 96688 292448 96694
rect 292396 96630 292448 96636
rect 292304 80912 292356 80918
rect 292304 80854 292356 80860
rect 292408 72486 292436 96630
rect 292500 93226 292528 96902
rect 292960 96898 292988 100028
rect 293250 100014 293356 100042
rect 293328 97050 293356 100014
rect 293420 97170 293448 100028
rect 293604 97345 293632 100028
rect 293590 97336 293646 97345
rect 293590 97271 293646 97280
rect 293408 97164 293460 97170
rect 293408 97106 293460 97112
rect 293328 97022 293724 97050
rect 293500 96960 293552 96966
rect 293500 96902 293552 96908
rect 292948 96892 293000 96898
rect 292948 96834 293000 96840
rect 292488 93220 292540 93226
rect 292488 93162 292540 93168
rect 292396 72480 292448 72486
rect 292396 72422 292448 72428
rect 292212 39364 292264 39370
rect 292212 39306 292264 39312
rect 291212 16546 291424 16574
rect 289636 14476 289688 14482
rect 289636 14418 289688 14424
rect 289360 9036 289412 9042
rect 289360 8978 289412 8984
rect 290188 4140 290240 4146
rect 290188 4082 290240 4088
rect 289084 2916 289136 2922
rect 289084 2858 289136 2864
rect 290200 480 290228 4082
rect 291396 480 291424 16546
rect 292580 7744 292632 7750
rect 292580 7686 292632 7692
rect 292592 480 292620 7686
rect 293512 6322 293540 96902
rect 293592 96892 293644 96898
rect 293592 96834 293644 96840
rect 293604 87553 293632 96834
rect 293590 87544 293646 87553
rect 293590 87479 293646 87488
rect 293696 80850 293724 97022
rect 293684 80844 293736 80850
rect 293684 80786 293736 80792
rect 293788 15910 293816 100028
rect 293972 99521 294000 100028
rect 293958 99512 294014 99521
rect 293958 99447 294014 99456
rect 293868 97164 293920 97170
rect 293868 97106 293920 97112
rect 293880 93906 293908 97106
rect 294248 96898 294276 100028
rect 294236 96892 294288 96898
rect 294236 96834 294288 96840
rect 294432 96830 294460 100028
rect 294616 96966 294644 100028
rect 294604 96960 294656 96966
rect 294604 96902 294656 96908
rect 294420 96824 294472 96830
rect 294420 96766 294472 96772
rect 294800 96762 294828 100028
rect 294984 96937 295012 100028
rect 295064 96960 295116 96966
rect 294970 96928 295026 96937
rect 295260 96937 295288 100028
rect 295064 96902 295116 96908
rect 295246 96928 295302 96937
rect 294970 96863 295026 96872
rect 294972 96824 295024 96830
rect 294972 96766 295024 96772
rect 294788 96756 294840 96762
rect 294788 96698 294840 96704
rect 294604 94580 294656 94586
rect 294604 94522 294656 94528
rect 293868 93900 293920 93906
rect 293868 93842 293920 93848
rect 293776 15904 293828 15910
rect 293776 15846 293828 15852
rect 294616 6458 294644 94522
rect 294696 93152 294748 93158
rect 294696 93094 294748 93100
rect 294708 9178 294736 93094
rect 294984 80889 295012 96766
rect 295076 90681 295104 96902
rect 295156 96892 295208 96898
rect 295246 96863 295302 96872
rect 295156 96834 295208 96840
rect 295062 90672 295118 90681
rect 295062 90607 295118 90616
rect 295168 86358 295196 96834
rect 295628 96830 295656 100028
rect 295812 97481 295840 100028
rect 296010 100014 296208 100042
rect 295798 97472 295854 97481
rect 295798 97407 295854 97416
rect 296076 97164 296128 97170
rect 296076 97106 296128 97112
rect 295616 96824 295668 96830
rect 295616 96766 295668 96772
rect 295248 96756 295300 96762
rect 295248 96698 295300 96704
rect 295260 93158 295288 96698
rect 295984 95124 296036 95130
rect 295984 95066 296036 95072
rect 295248 93152 295300 93158
rect 295248 93094 295300 93100
rect 295156 86352 295208 86358
rect 295156 86294 295208 86300
rect 294970 80880 295026 80889
rect 294970 80815 295026 80824
rect 295340 80776 295392 80782
rect 295340 80718 295392 80724
rect 294696 9172 294748 9178
rect 294696 9114 294748 9120
rect 294604 6452 294656 6458
rect 294604 6394 294656 6400
rect 293500 6316 293552 6322
rect 293500 6258 293552 6264
rect 295352 3534 295380 80718
rect 295996 11762 296024 95066
rect 296088 94586 296116 97106
rect 296180 96948 296208 100014
rect 296272 97102 296300 100028
rect 296456 97170 296484 100028
rect 296548 100014 296654 100042
rect 296444 97164 296496 97170
rect 296444 97106 296496 97112
rect 296260 97096 296312 97102
rect 296260 97038 296312 97044
rect 296548 96948 296576 100014
rect 296628 97096 296680 97102
rect 296628 97038 296680 97044
rect 296180 96920 296392 96948
rect 296260 96824 296312 96830
rect 296260 96766 296312 96772
rect 296076 94580 296128 94586
rect 296076 94522 296128 94528
rect 296074 80744 296130 80753
rect 296074 80679 296130 80688
rect 296088 16574 296116 80679
rect 296272 76566 296300 96766
rect 296364 86290 296392 96920
rect 296456 96920 296576 96948
rect 296352 86284 296404 86290
rect 296352 86226 296404 86232
rect 296456 86193 296484 96920
rect 296442 86184 296498 86193
rect 296442 86119 296498 86128
rect 296640 84194 296668 97038
rect 296824 96762 296852 100028
rect 296812 96756 296864 96762
rect 296812 96698 296864 96704
rect 297008 94518 297036 100028
rect 297284 96830 297312 100028
rect 297482 100014 297588 100042
rect 297666 100014 297772 100042
rect 297560 96948 297588 100014
rect 297744 97050 297772 100014
rect 297744 97022 298048 97050
rect 297560 96920 297956 96948
rect 297272 96824 297324 96830
rect 297272 96766 297324 96772
rect 297824 96824 297876 96830
rect 297824 96766 297876 96772
rect 297732 96756 297784 96762
rect 297732 96698 297784 96704
rect 296996 94512 297048 94518
rect 296996 94454 297048 94460
rect 297364 93900 297416 93906
rect 297364 93842 297416 93848
rect 296548 84166 296668 84194
rect 296548 80782 296576 84166
rect 296536 80776 296588 80782
rect 296536 80718 296588 80724
rect 296260 76560 296312 76566
rect 296260 76502 296312 76508
rect 296088 16546 296208 16574
rect 295984 11756 296036 11762
rect 295984 11698 296036 11704
rect 296076 3596 296128 3602
rect 296076 3538 296128 3544
rect 294880 3528 294932 3534
rect 294880 3470 294932 3476
rect 295340 3528 295392 3534
rect 295340 3470 295392 3476
rect 293684 2916 293736 2922
rect 293684 2858 293736 2864
rect 293696 480 293724 2858
rect 294892 480 294920 3470
rect 296088 480 296116 3538
rect 296180 3262 296208 16546
rect 297376 6254 297404 93842
rect 297744 80714 297772 96698
rect 297836 83502 297864 96766
rect 297824 83496 297876 83502
rect 297824 83438 297876 83444
rect 297928 80753 297956 96920
rect 298020 96626 298048 97022
rect 298008 96620 298060 96626
rect 298008 96562 298060 96568
rect 298296 94489 298324 100028
rect 298664 96694 298692 100028
rect 298848 96966 298876 100028
rect 299046 100014 299244 100042
rect 298836 96960 298888 96966
rect 298836 96902 298888 96908
rect 299216 96812 299244 100014
rect 299308 96937 299336 100028
rect 299388 96960 299440 96966
rect 299294 96928 299350 96937
rect 299388 96902 299440 96908
rect 299294 96863 299350 96872
rect 299216 96784 299336 96812
rect 298652 96688 298704 96694
rect 298652 96630 298704 96636
rect 299204 96688 299256 96694
rect 299204 96630 299256 96636
rect 298744 96620 298796 96626
rect 298744 96562 298796 96568
rect 298282 94480 298338 94489
rect 298282 94415 298338 94424
rect 297914 80744 297970 80753
rect 297456 80708 297508 80714
rect 297456 80650 297508 80656
rect 297732 80708 297784 80714
rect 297914 80679 297970 80688
rect 297732 80650 297784 80656
rect 297364 6248 297416 6254
rect 297364 6190 297416 6196
rect 297468 3534 297496 80650
rect 298100 73840 298152 73846
rect 298100 73782 298152 73788
rect 298112 4146 298140 73782
rect 298756 6186 298784 96562
rect 299216 79354 299244 96630
rect 299204 79348 299256 79354
rect 299204 79290 299256 79296
rect 299308 73846 299336 96784
rect 299296 73840 299348 73846
rect 299296 73782 299348 73788
rect 299400 8974 299428 96902
rect 299492 96898 299520 100028
rect 299676 97306 299704 100028
rect 299664 97300 299716 97306
rect 299664 97242 299716 97248
rect 299860 96966 299888 100028
rect 320180 99816 320232 99822
rect 320180 99758 320232 99764
rect 306380 98184 306432 98190
rect 306380 98126 306432 98132
rect 300584 97776 300636 97782
rect 300584 97718 300636 97724
rect 299848 96960 299900 96966
rect 299848 96902 299900 96908
rect 299480 96892 299532 96898
rect 299480 96834 299532 96840
rect 300596 96218 300624 97718
rect 304998 97472 305054 97481
rect 304998 97407 305054 97416
rect 300768 96960 300820 96966
rect 300768 96902 300820 96908
rect 300676 96892 300728 96898
rect 300676 96834 300728 96840
rect 300584 96212 300636 96218
rect 300584 96154 300636 96160
rect 300688 64190 300716 96834
rect 300676 64184 300728 64190
rect 300676 64126 300728 64132
rect 300124 39364 300176 39370
rect 300124 39306 300176 39312
rect 299388 8968 299440 8974
rect 299388 8910 299440 8916
rect 298744 6180 298796 6186
rect 298744 6122 298796 6128
rect 298100 4140 298152 4146
rect 298100 4082 298152 4088
rect 297456 3528 297508 3534
rect 297456 3470 297508 3476
rect 298468 3528 298520 3534
rect 298468 3470 298520 3476
rect 296168 3256 296220 3262
rect 296168 3198 296220 3204
rect 297272 3256 297324 3262
rect 297272 3198 297324 3204
rect 297284 480 297312 3198
rect 298480 480 298508 3470
rect 300136 3466 300164 39306
rect 300780 35222 300808 96902
rect 302332 96348 302384 96354
rect 302332 96290 302384 96296
rect 302238 94616 302294 94625
rect 302238 94551 302294 94560
rect 300860 89412 300912 89418
rect 300860 89354 300912 89360
rect 300768 35216 300820 35222
rect 300768 35158 300820 35164
rect 300872 16574 300900 89354
rect 300872 16546 301544 16574
rect 300768 3528 300820 3534
rect 300768 3470 300820 3476
rect 300124 3460 300176 3466
rect 300124 3402 300176 3408
rect 299664 3392 299716 3398
rect 299664 3334 299716 3340
rect 299676 480 299704 3334
rect 300780 480 300808 3470
rect 301516 490 301544 16546
rect 302252 3210 302280 94551
rect 302344 3398 302372 96290
rect 303710 96112 303766 96121
rect 303710 96047 303766 96056
rect 303620 89344 303672 89350
rect 303620 89286 303672 89292
rect 302332 3392 302384 3398
rect 302332 3334 302384 3340
rect 302252 3182 303200 3210
rect 301792 598 302004 626
rect 301792 490 301820 598
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301516 462 301820 490
rect 301976 480 302004 598
rect 303172 480 303200 3182
rect 303632 626 303660 89286
rect 303724 3602 303752 96047
rect 305012 94654 305040 97407
rect 305000 94648 305052 94654
rect 305000 94590 305052 94596
rect 303712 3596 303764 3602
rect 303712 3538 303764 3544
rect 305550 2000 305606 2009
rect 305550 1935 305606 1944
rect 303632 598 303936 626
rect 303908 490 303936 598
rect 304184 598 304396 626
rect 304184 490 304212 598
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 303908 462 304212 490
rect 304368 480 304396 598
rect 305564 480 305592 1935
rect 306392 490 306420 98126
rect 309876 97708 309928 97714
rect 309876 97650 309928 97656
rect 307024 90772 307076 90778
rect 307024 90714 307076 90720
rect 307036 2922 307064 90714
rect 309140 88052 309192 88058
rect 309140 87994 309192 88000
rect 307852 81116 307904 81122
rect 307852 81058 307904 81064
rect 307864 11694 307892 81058
rect 307852 11688 307904 11694
rect 307852 11630 307904 11636
rect 309048 11688 309100 11694
rect 309048 11630 309100 11636
rect 307024 2916 307076 2922
rect 307024 2858 307076 2864
rect 307944 2916 307996 2922
rect 307944 2858 307996 2864
rect 306576 598 306788 626
rect 306576 490 306604 598
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306392 462 306604 490
rect 306760 480 306788 598
rect 307956 480 307984 2858
rect 309060 480 309088 11630
rect 309152 3534 309180 87994
rect 309888 86562 309916 97650
rect 312542 97336 312598 97345
rect 312542 97271 312598 97280
rect 312556 93294 312584 97271
rect 318064 94920 318116 94926
rect 318064 94862 318116 94868
rect 316040 94852 316092 94858
rect 316040 94794 316092 94800
rect 311164 93288 311216 93294
rect 311164 93230 311216 93236
rect 312544 93288 312596 93294
rect 312544 93230 312596 93236
rect 309784 86556 309836 86562
rect 309784 86498 309836 86504
rect 309876 86556 309928 86562
rect 309876 86498 309928 86504
rect 309796 3534 309824 86498
rect 310244 3732 310296 3738
rect 310244 3674 310296 3680
rect 309140 3528 309192 3534
rect 309140 3470 309192 3476
rect 309784 3528 309836 3534
rect 309784 3470 309836 3476
rect 310256 480 310284 3674
rect 311176 3602 311204 93230
rect 313280 92200 313332 92206
rect 313280 92142 313332 92148
rect 311256 86692 311308 86698
rect 311256 86634 311308 86640
rect 311164 3596 311216 3602
rect 311164 3538 311216 3544
rect 311268 3194 311296 86634
rect 311898 82104 311954 82113
rect 311898 82039 311954 82048
rect 311912 16574 311940 82039
rect 313292 16574 313320 92142
rect 316052 16574 316080 94794
rect 317420 87984 317472 87990
rect 317420 87926 317472 87932
rect 316682 76800 316738 76809
rect 316682 76735 316738 76744
rect 311912 16546 312216 16574
rect 313292 16546 313872 16574
rect 316052 16546 316264 16574
rect 311440 3528 311492 3534
rect 311440 3470 311492 3476
rect 311256 3188 311308 3194
rect 311256 3130 311308 3136
rect 311452 480 311480 3470
rect 312188 490 312216 16546
rect 312464 598 312676 626
rect 312464 490 312492 598
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312188 462 312492 490
rect 312648 480 312676 598
rect 313844 480 313872 16546
rect 315028 3188 315080 3194
rect 315028 3130 315080 3136
rect 315040 480 315068 3130
rect 316236 480 316264 16546
rect 316696 2990 316724 76735
rect 317432 12434 317460 87926
rect 318076 16574 318104 94862
rect 318076 16546 318196 16574
rect 317432 12406 318104 12434
rect 317328 6520 317380 6526
rect 317328 6462 317380 6468
rect 316684 2984 316736 2990
rect 316684 2926 316736 2932
rect 317340 480 317368 6462
rect 318076 490 318104 12406
rect 318168 3806 318196 16546
rect 319720 9376 319772 9382
rect 319720 9318 319772 9324
rect 318156 3800 318208 3806
rect 318156 3742 318208 3748
rect 318352 598 318564 626
rect 318352 490 318380 598
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318076 462 318380 490
rect 318536 480 318564 598
rect 319732 480 319760 9318
rect 320192 3942 320220 99758
rect 323584 99748 323636 99754
rect 323584 99690 323636 99696
rect 322940 81048 322992 81054
rect 322940 80990 322992 80996
rect 320180 3936 320232 3942
rect 320180 3878 320232 3884
rect 320916 3120 320968 3126
rect 320916 3062 320968 3068
rect 320928 480 320956 3062
rect 322112 2984 322164 2990
rect 322112 2926 322164 2932
rect 322124 480 322152 2926
rect 322952 490 322980 80990
rect 323596 4146 323624 99690
rect 331864 99680 331916 99686
rect 331864 99622 331916 99628
rect 529938 99648 529994 99657
rect 324412 98864 324464 98870
rect 324412 98806 324464 98812
rect 324424 12434 324452 98806
rect 328460 98116 328512 98122
rect 328460 98058 328512 98064
rect 327080 93492 327132 93498
rect 327080 93434 327132 93440
rect 324504 86624 324556 86630
rect 324504 86566 324556 86572
rect 324516 16574 324544 86566
rect 326342 73808 326398 73817
rect 326342 73743 326398 73752
rect 326356 16574 326384 73743
rect 327092 16574 327120 93434
rect 327722 79656 327778 79665
rect 327722 79591 327778 79600
rect 324516 16546 325648 16574
rect 326356 16546 326476 16574
rect 327092 16546 327672 16574
rect 324332 12406 324452 12434
rect 323584 4140 323636 4146
rect 323584 4082 323636 4088
rect 324332 3126 324360 12406
rect 324412 4140 324464 4146
rect 324412 4082 324464 4088
rect 324320 3120 324372 3126
rect 324320 3062 324372 3068
rect 323136 598 323348 626
rect 323136 490 323164 598
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 322952 462 323164 490
rect 323320 480 323348 598
rect 324424 480 324452 4082
rect 325620 480 325648 16546
rect 326342 11928 326398 11937
rect 326342 11863 326398 11872
rect 326356 490 326384 11863
rect 326448 3942 326476 16546
rect 326436 3936 326488 3942
rect 326436 3878 326488 3884
rect 327644 2774 327672 16546
rect 327736 3874 327764 79591
rect 328472 16574 328500 98058
rect 329840 96280 329892 96286
rect 329840 96222 329892 96228
rect 329852 16574 329880 96222
rect 328472 16546 328776 16574
rect 329852 16546 330432 16574
rect 327724 3868 327776 3874
rect 327724 3810 327776 3816
rect 327644 2746 328040 2774
rect 326632 598 326844 626
rect 326632 490 326660 598
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326356 462 326660 490
rect 326816 480 326844 598
rect 328012 480 328040 2746
rect 328748 490 328776 16546
rect 329024 598 329236 626
rect 329024 490 329052 598
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 328748 462 329052 490
rect 329208 480 329236 598
rect 330404 480 330432 16546
rect 331588 7676 331640 7682
rect 331588 7618 331640 7624
rect 331600 480 331628 7618
rect 331876 3942 331904 99622
rect 345020 99612 345072 99618
rect 529938 99583 529994 99592
rect 345020 99554 345072 99560
rect 338120 96144 338172 96150
rect 338120 96086 338172 96092
rect 333980 93424 334032 93430
rect 333980 93366 334032 93372
rect 332692 47592 332744 47598
rect 332692 47534 332744 47540
rect 332704 11694 332732 47534
rect 333992 16574 334020 93366
rect 336004 93356 336056 93362
rect 336004 93298 336056 93304
rect 333992 16546 334664 16574
rect 332692 11688 332744 11694
rect 332692 11630 332744 11636
rect 333888 11688 333940 11694
rect 333888 11630 333940 11636
rect 331864 3936 331916 3942
rect 331864 3878 331916 3884
rect 332692 3596 332744 3602
rect 332692 3538 332744 3544
rect 332704 480 332732 3538
rect 333900 480 333928 11630
rect 334636 490 334664 16546
rect 336016 3330 336044 93298
rect 336740 75472 336792 75478
rect 336740 75414 336792 75420
rect 336096 72752 336148 72758
rect 336096 72694 336148 72700
rect 336108 3806 336136 72694
rect 336752 16574 336780 75414
rect 338132 16574 338160 96086
rect 341524 89276 341576 89282
rect 341524 89218 341576 89224
rect 339500 87916 339552 87922
rect 339500 87858 339552 87864
rect 336752 16546 337056 16574
rect 338132 16546 338712 16574
rect 336096 3800 336148 3806
rect 336096 3742 336148 3748
rect 336280 3732 336332 3738
rect 336280 3674 336332 3680
rect 336004 3324 336056 3330
rect 336004 3266 336056 3272
rect 334912 598 335124 626
rect 334912 490 334940 598
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 334636 462 334940 490
rect 335096 480 335124 598
rect 336292 480 336320 3674
rect 337028 490 337056 16546
rect 337304 598 337516 626
rect 337304 490 337332 598
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337028 462 337332 490
rect 337488 480 337516 598
rect 338684 480 338712 16546
rect 339512 490 339540 87858
rect 340972 70032 341024 70038
rect 340972 69974 341024 69980
rect 339696 598 339908 626
rect 339696 490 339724 598
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339512 462 339724 490
rect 339880 480 339908 598
rect 340984 480 341012 69974
rect 341536 3602 341564 89218
rect 342258 84960 342314 84969
rect 342258 84895 342314 84904
rect 342272 16574 342300 84895
rect 345032 16574 345060 99554
rect 504364 99544 504416 99550
rect 504364 99486 504416 99492
rect 493322 98968 493378 98977
rect 493322 98903 493378 98912
rect 394700 98796 394752 98802
rect 394700 98738 394752 98744
rect 353944 97640 353996 97646
rect 353944 97582 353996 97588
rect 351918 93392 351974 93401
rect 351918 93327 351974 93336
rect 347044 90704 347096 90710
rect 347044 90646 347096 90652
rect 346400 75404 346452 75410
rect 346400 75346 346452 75352
rect 346412 16574 346440 75346
rect 342272 16546 342944 16574
rect 345032 16546 345336 16574
rect 346412 16546 346992 16574
rect 341524 3596 341576 3602
rect 341524 3538 341576 3544
rect 342168 3324 342220 3330
rect 342168 3266 342220 3272
rect 342180 480 342208 3266
rect 342916 490 342944 16546
rect 344560 3868 344612 3874
rect 344560 3810 344612 3816
rect 343192 598 343404 626
rect 343192 490 343220 598
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 342916 462 343220 490
rect 343376 480 343404 598
rect 344572 480 344600 3810
rect 345308 490 345336 16546
rect 345584 598 345796 626
rect 345584 490 345612 598
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345308 462 345612 490
rect 345768 480 345796 598
rect 346964 480 346992 16546
rect 347056 3126 347084 90646
rect 350540 79620 350592 79626
rect 350540 79562 350592 79568
rect 350552 16574 350580 79562
rect 351932 16574 351960 93327
rect 353298 72448 353354 72457
rect 353298 72383 353354 72392
rect 353312 16574 353340 72383
rect 353956 22778 353984 97582
rect 378140 96212 378192 96218
rect 378140 96154 378192 96160
rect 375380 94784 375432 94790
rect 375380 94726 375432 94732
rect 356060 92132 356112 92138
rect 356060 92074 356112 92080
rect 354680 79552 354732 79558
rect 354680 79494 354732 79500
rect 353944 22772 353996 22778
rect 353944 22714 353996 22720
rect 354692 16574 354720 79494
rect 356072 16574 356100 92074
rect 358820 92064 358872 92070
rect 358820 92006 358872 92012
rect 357440 85264 357492 85270
rect 357440 85206 357492 85212
rect 350552 16546 351224 16574
rect 351932 16546 352880 16574
rect 353312 16546 353616 16574
rect 354692 16546 355272 16574
rect 356072 16546 356376 16574
rect 348056 11892 348108 11898
rect 348056 11834 348108 11840
rect 347044 3120 347096 3126
rect 347044 3062 347096 3068
rect 348068 480 348096 11834
rect 349252 3800 349304 3806
rect 349252 3742 349304 3748
rect 349264 480 349292 3742
rect 350448 3120 350500 3126
rect 350448 3062 350500 3068
rect 350460 480 350488 3062
rect 351196 490 351224 16546
rect 351472 598 351684 626
rect 351472 490 351500 598
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351196 462 351500 490
rect 351656 480 351684 598
rect 352852 480 352880 16546
rect 353588 490 353616 16546
rect 353864 598 354076 626
rect 353864 490 353892 598
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 353588 462 353892 490
rect 354048 480 354076 598
rect 355244 480 355272 16546
rect 356348 480 356376 16546
rect 357452 6914 357480 85206
rect 357532 79484 357584 79490
rect 357532 79426 357584 79432
rect 357544 11694 357572 79426
rect 358832 16574 358860 92006
rect 364984 91996 365036 92002
rect 364984 91938 365036 91944
rect 360200 85196 360252 85202
rect 360200 85138 360252 85144
rect 360212 16574 360240 85138
rect 363602 79520 363658 79529
rect 363602 79455 363658 79464
rect 358832 16546 359504 16574
rect 360212 16546 361160 16574
rect 357532 11688 357584 11694
rect 357532 11630 357584 11636
rect 358728 11688 358780 11694
rect 358728 11630 358780 11636
rect 357452 6886 357572 6914
rect 357544 480 357572 6886
rect 358740 480 358768 11630
rect 359476 490 359504 16546
rect 359752 598 359964 626
rect 359752 490 359780 598
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359476 462 359780 490
rect 359936 480 359964 598
rect 361132 480 361160 16546
rect 363616 4078 363644 79455
rect 364340 72684 364392 72690
rect 364340 72626 364392 72632
rect 364352 16574 364380 72626
rect 364352 16546 364656 16574
rect 363604 4072 363656 4078
rect 363604 4014 363656 4020
rect 362316 3732 362368 3738
rect 362316 3674 362368 3680
rect 362328 480 362356 3674
rect 363512 3528 363564 3534
rect 363512 3470 363564 3476
rect 363524 480 363552 3470
rect 364628 480 364656 16546
rect 364996 3534 365024 91938
rect 374644 91928 374696 91934
rect 374644 91870 374696 91876
rect 370502 90672 370558 90681
rect 370502 90607 370558 90616
rect 367100 85128 367152 85134
rect 367100 85070 367152 85076
rect 367112 6914 367140 85070
rect 367742 30968 367798 30977
rect 367742 30903 367798 30912
rect 367756 16574 367784 30903
rect 367756 16546 367876 16574
rect 367112 6886 367784 6914
rect 365812 4072 365864 4078
rect 365812 4014 365864 4020
rect 364984 3528 365036 3534
rect 364984 3470 365036 3476
rect 365824 480 365852 4014
rect 367008 3528 367060 3534
rect 367008 3470 367060 3476
rect 367020 480 367048 3470
rect 367756 490 367784 6886
rect 367848 3330 367876 16546
rect 370516 3534 370544 90607
rect 373998 71224 374054 71233
rect 373998 71159 374054 71168
rect 372896 11824 372948 11830
rect 372896 11766 372948 11772
rect 370596 6452 370648 6458
rect 370596 6394 370648 6400
rect 370504 3528 370556 3534
rect 370504 3470 370556 3476
rect 367836 3324 367888 3330
rect 367836 3266 367888 3272
rect 369400 3324 369452 3330
rect 369400 3266 369452 3272
rect 368032 598 368244 626
rect 368032 490 368060 598
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 367756 462 368060 490
rect 368216 480 368244 598
rect 369412 480 369440 3266
rect 370608 480 370636 6394
rect 371700 3664 371752 3670
rect 371700 3606 371752 3612
rect 371712 480 371740 3606
rect 372908 480 372936 11766
rect 374012 3398 374040 71159
rect 374092 9308 374144 9314
rect 374092 9250 374144 9256
rect 374000 3392 374052 3398
rect 374000 3334 374052 3340
rect 374104 480 374132 9250
rect 374656 3670 374684 91870
rect 375392 16574 375420 94726
rect 376758 91760 376814 91769
rect 376758 91695 376814 91704
rect 376772 16574 376800 91695
rect 378152 16574 378180 96154
rect 380900 91860 380952 91866
rect 380900 91802 380952 91808
rect 378784 69964 378836 69970
rect 378784 69906 378836 69912
rect 375392 16546 376064 16574
rect 376772 16546 377720 16574
rect 378152 16546 378456 16574
rect 374644 3664 374696 3670
rect 374644 3606 374696 3612
rect 375288 3392 375340 3398
rect 375288 3334 375340 3340
rect 375300 480 375328 3334
rect 376036 490 376064 16546
rect 376312 598 376524 626
rect 376312 490 376340 598
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376036 462 376340 490
rect 376496 480 376524 598
rect 377692 480 377720 16546
rect 378428 490 378456 16546
rect 378796 3398 378824 69906
rect 380912 16574 380940 91802
rect 389824 91792 389876 91798
rect 389824 91734 389876 91740
rect 385684 89208 385736 89214
rect 385684 89150 385736 89156
rect 382280 85060 382332 85066
rect 382280 85002 382332 85008
rect 382292 16574 382320 85002
rect 385038 75304 385094 75313
rect 385038 75239 385094 75248
rect 385052 16574 385080 75239
rect 380912 16546 381216 16574
rect 382292 16546 382412 16574
rect 385052 16546 385632 16574
rect 378784 3392 378836 3398
rect 378784 3334 378836 3340
rect 379980 3392 380032 3398
rect 379980 3334 380032 3340
rect 378704 598 378916 626
rect 378704 490 378732 598
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378428 462 378732 490
rect 378888 480 378916 598
rect 379992 480 380020 3334
rect 381188 480 381216 16546
rect 382384 480 382412 16546
rect 383568 14544 383620 14550
rect 383568 14486 383620 14492
rect 383580 480 383608 14486
rect 384764 3664 384816 3670
rect 384764 3606 384816 3612
rect 384776 480 384804 3606
rect 385604 3482 385632 16546
rect 385696 3670 385724 89150
rect 387800 86488 387852 86494
rect 387800 86430 387852 86436
rect 386420 78192 386472 78198
rect 386420 78134 386472 78140
rect 386432 16574 386460 78134
rect 386432 16546 386736 16574
rect 385684 3664 385736 3670
rect 385684 3606 385736 3612
rect 385604 3454 386000 3482
rect 385972 480 386000 3454
rect 386708 490 386736 16546
rect 386984 598 387196 626
rect 386984 490 387012 598
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 386708 462 387012 490
rect 387168 480 387196 598
rect 387812 490 387840 86430
rect 389180 71256 389232 71262
rect 389180 71198 389232 71204
rect 389192 16574 389220 71198
rect 389192 16546 389496 16574
rect 388088 598 388300 626
rect 388088 490 388116 598
rect 387126 -960 387238 480
rect 387812 462 388116 490
rect 388272 480 388300 598
rect 389468 480 389496 16546
rect 389836 3058 389864 91734
rect 391938 84824 391994 84833
rect 391938 84759 391994 84768
rect 390652 68400 390704 68406
rect 390652 68342 390704 68348
rect 389824 3052 389876 3058
rect 389824 2994 389876 3000
rect 390664 480 390692 68342
rect 391952 16574 391980 84759
rect 393318 78160 393374 78169
rect 393318 78095 393374 78104
rect 393332 16574 393360 78095
rect 394712 16574 394740 98738
rect 475384 98728 475436 98734
rect 475384 98670 475436 98676
rect 443644 97572 443696 97578
rect 443644 97514 443696 97520
rect 403622 97200 403678 97209
rect 403622 97135 403678 97144
rect 396724 87848 396776 87854
rect 396724 87790 396776 87796
rect 396080 72616 396132 72622
rect 396080 72558 396132 72564
rect 391952 16546 392624 16574
rect 393332 16546 394280 16574
rect 394712 16546 395384 16574
rect 391848 3052 391900 3058
rect 391848 2994 391900 3000
rect 391860 480 391888 2994
rect 392596 490 392624 16546
rect 392872 598 393084 626
rect 392872 490 392900 598
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 392596 462 392900 490
rect 393056 480 393084 598
rect 394252 480 394280 16546
rect 395356 480 395384 16546
rect 396092 490 396120 72558
rect 396736 3398 396764 87790
rect 398932 83836 398984 83842
rect 398932 83778 398984 83784
rect 397460 42084 397512 42090
rect 397460 42026 397512 42032
rect 397472 16574 397500 42026
rect 397472 16546 397776 16574
rect 396724 3392 396776 3398
rect 396724 3334 396776 3340
rect 396368 598 396580 626
rect 396368 490 396396 598
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396092 462 396396 490
rect 396552 480 396580 598
rect 397748 480 397776 16546
rect 398944 11830 398972 83778
rect 400220 78124 400272 78130
rect 400220 78066 400272 78072
rect 400232 16574 400260 78066
rect 403070 76664 403126 76673
rect 403070 76599 403126 76608
rect 402980 71188 403032 71194
rect 402980 71130 403032 71136
rect 400232 16546 400904 16574
rect 398932 11824 398984 11830
rect 398932 11766 398984 11772
rect 400128 11824 400180 11830
rect 400128 11766 400180 11772
rect 398932 3392 398984 3398
rect 398932 3334 398984 3340
rect 398944 480 398972 3334
rect 400140 480 400168 11766
rect 400876 490 400904 16546
rect 402520 4140 402572 4146
rect 402520 4082 402572 4088
rect 401152 598 401364 626
rect 401152 490 401180 598
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 400876 462 401180 490
rect 401336 480 401364 598
rect 402532 480 402560 4082
rect 402992 3482 403020 71130
rect 403084 4146 403112 76599
rect 403636 72622 403664 97135
rect 421012 94716 421064 94722
rect 421012 94658 421064 94664
rect 412640 90636 412692 90642
rect 412640 90578 412692 90584
rect 406384 83768 406436 83774
rect 406384 83710 406436 83716
rect 403624 72616 403676 72622
rect 403624 72558 403676 72564
rect 406016 9240 406068 9246
rect 406016 9182 406068 9188
rect 404820 7608 404872 7614
rect 404820 7550 404872 7556
rect 403072 4140 403124 4146
rect 403072 4082 403124 4088
rect 402992 3454 403664 3482
rect 403636 480 403664 3454
rect 404832 480 404860 7550
rect 406028 480 406056 9182
rect 406396 3398 406424 83710
rect 411904 80980 411956 80986
rect 411904 80922 411956 80928
rect 407212 78056 407264 78062
rect 407212 77998 407264 78004
rect 407224 11830 407252 77998
rect 409970 76528 410026 76537
rect 409970 76463 410026 76472
rect 409880 71120 409932 71126
rect 409880 71062 409932 71068
rect 407212 11824 407264 11830
rect 407212 11766 407264 11772
rect 408408 11824 408460 11830
rect 408408 11766 408460 11772
rect 406384 3392 406436 3398
rect 406384 3334 406436 3340
rect 407212 3392 407264 3398
rect 407212 3334 407264 3340
rect 407224 480 407252 3334
rect 408420 480 408448 11766
rect 409892 3738 409920 71062
rect 409880 3732 409932 3738
rect 409880 3674 409932 3680
rect 409984 3482 410012 76463
rect 411812 10328 411864 10334
rect 411812 10270 411864 10276
rect 410800 3732 410852 3738
rect 410800 3674 410852 3680
rect 409616 3454 410012 3482
rect 409616 480 409644 3454
rect 410812 480 410840 3674
rect 411824 3482 411852 10270
rect 411916 3738 411944 80922
rect 411904 3732 411956 3738
rect 411904 3674 411956 3680
rect 411824 3454 411944 3482
rect 411916 480 411944 3454
rect 412652 490 412680 90578
rect 416872 90568 416924 90574
rect 416872 90510 416924 90516
rect 414020 83700 414072 83706
rect 414020 83642 414072 83648
rect 414032 16574 414060 83642
rect 415398 78024 415454 78033
rect 415398 77959 415454 77968
rect 415412 16574 415440 77959
rect 414032 16546 414336 16574
rect 415412 16546 415532 16574
rect 412928 598 413140 626
rect 412928 490 412956 598
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 412652 462 412956 490
rect 413112 480 413140 598
rect 414308 480 414336 16546
rect 415504 480 415532 16546
rect 416780 11756 416832 11762
rect 416780 11698 416832 11704
rect 416792 3806 416820 11698
rect 416780 3800 416832 3806
rect 416780 3742 416832 3748
rect 416884 3482 416912 90510
rect 418160 77988 418212 77994
rect 418160 77930 418212 77936
rect 418172 16574 418200 77930
rect 420920 74180 420972 74186
rect 420920 74122 420972 74128
rect 418172 16546 418568 16574
rect 417884 3800 417936 3806
rect 417884 3742 417936 3748
rect 416700 3454 416912 3482
rect 416700 480 416728 3454
rect 417896 480 417924 3742
rect 418540 490 418568 16546
rect 420184 3392 420236 3398
rect 420184 3334 420236 3340
rect 418816 598 419028 626
rect 418816 490 418844 598
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418540 462 418844 490
rect 419000 480 419028 598
rect 420196 480 420224 3334
rect 420932 490 420960 74122
rect 421024 3398 421052 94658
rect 429842 90536 429898 90545
rect 427912 90500 427964 90506
rect 429842 90471 429898 90480
rect 427912 90442 427964 90448
rect 425060 86556 425112 86562
rect 425060 86498 425112 86504
rect 423770 83600 423826 83609
rect 423770 83535 423826 83544
rect 422300 66904 422352 66910
rect 422300 66846 422352 66852
rect 422312 16574 422340 66846
rect 422312 16546 422616 16574
rect 421012 3392 421064 3398
rect 421012 3334 421064 3340
rect 421208 598 421420 626
rect 421208 490 421236 598
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 420932 462 421236 490
rect 421392 480 421420 598
rect 422588 480 422616 16546
rect 423784 11762 423812 83535
rect 425072 16574 425100 86498
rect 427820 72548 427872 72554
rect 427820 72490 427872 72496
rect 425072 16546 425744 16574
rect 423772 11756 423824 11762
rect 423772 11698 423824 11704
rect 424968 11756 425020 11762
rect 424968 11698 425020 11704
rect 423772 3732 423824 3738
rect 423772 3674 423824 3680
rect 423784 480 423812 3674
rect 424980 480 425008 11698
rect 425716 490 425744 16546
rect 427268 3392 427320 3398
rect 427268 3334 427320 3340
rect 425992 598 426204 626
rect 425992 490 426020 598
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 425716 462 426020 490
rect 426176 480 426204 598
rect 427280 480 427308 3334
rect 427832 3210 427860 72490
rect 427924 3398 427952 90442
rect 429200 53100 429252 53106
rect 429200 53042 429252 53048
rect 427912 3392 427964 3398
rect 427912 3334 427964 3340
rect 427832 3182 428504 3210
rect 428476 480 428504 3182
rect 429212 490 429240 53042
rect 429856 2922 429884 90471
rect 430580 90432 430632 90438
rect 430580 90374 430632 90380
rect 440238 90400 440294 90409
rect 430592 16574 430620 90374
rect 438952 90364 439004 90370
rect 440238 90335 440294 90344
rect 438952 90306 439004 90312
rect 434720 83632 434772 83638
rect 434720 83574 434772 83580
rect 432604 76764 432656 76770
rect 432604 76706 432656 76712
rect 431224 69896 431276 69902
rect 431224 69838 431276 69844
rect 430592 16546 430896 16574
rect 429844 2916 429896 2922
rect 429844 2858 429896 2864
rect 429488 598 429700 626
rect 429488 490 429516 598
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429212 462 429516 490
rect 429672 480 429700 598
rect 430868 480 430896 16546
rect 431236 4146 431264 69838
rect 432510 11792 432566 11801
rect 432510 11727 432566 11736
rect 431224 4140 431276 4146
rect 431224 4082 431276 4088
rect 432052 4140 432104 4146
rect 432052 4082 432104 4088
rect 432064 480 432092 4082
rect 432524 3482 432552 11727
rect 432616 3738 432644 76706
rect 434732 16574 434760 83574
rect 436744 76696 436796 76702
rect 436744 76638 436796 76644
rect 436100 68332 436152 68338
rect 436100 68274 436152 68280
rect 436112 16574 436140 68274
rect 434732 16546 435128 16574
rect 436112 16546 436692 16574
rect 432604 3732 432656 3738
rect 432604 3674 432656 3680
rect 432524 3454 433288 3482
rect 433260 480 433288 3454
rect 434444 2916 434496 2922
rect 434444 2858 434496 2864
rect 434456 480 434484 2858
rect 435100 490 435128 16546
rect 436664 3482 436692 16546
rect 436756 3806 436784 76638
rect 438860 69828 438912 69834
rect 438860 69770 438912 69776
rect 436744 3800 436796 3806
rect 436744 3742 436796 3748
rect 436664 3454 436784 3482
rect 435376 598 435588 626
rect 435376 490 435404 598
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435100 462 435404 490
rect 435560 480 435588 598
rect 436756 480 436784 3454
rect 437940 3052 437992 3058
rect 437940 2994 437992 3000
rect 437952 480 437980 2994
rect 438872 2938 438900 69770
rect 438964 3058 438992 90306
rect 440252 3398 440280 90335
rect 441618 83464 441674 83473
rect 441618 83399 441674 83408
rect 440332 62824 440384 62830
rect 440332 62766 440384 62772
rect 440240 3392 440292 3398
rect 440240 3334 440292 3340
rect 438952 3052 439004 3058
rect 438952 2994 439004 3000
rect 438872 2910 439176 2938
rect 439148 480 439176 2910
rect 440344 480 440372 62766
rect 441632 16574 441660 83399
rect 443000 17264 443052 17270
rect 443000 17206 443052 17212
rect 443012 16574 443040 17206
rect 441632 16546 442672 16574
rect 443012 16546 443408 16574
rect 441528 3392 441580 3398
rect 441528 3334 441580 3340
rect 441540 480 441568 3334
rect 442644 480 442672 16546
rect 443380 490 443408 16546
rect 443656 5574 443684 97514
rect 454684 97504 454736 97510
rect 454684 97446 454736 97452
rect 449164 84992 449216 84998
rect 449164 84934 449216 84940
rect 445760 83564 445812 83570
rect 445760 83506 445812 83512
rect 443644 5568 443696 5574
rect 443644 5510 443696 5516
rect 445024 3800 445076 3806
rect 445024 3742 445076 3748
rect 443656 598 443868 626
rect 443656 490 443684 598
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443380 462 443684 490
rect 443840 480 443868 598
rect 445036 480 445064 3742
rect 445772 490 445800 83506
rect 447782 77888 447838 77897
rect 447782 77823 447838 77832
rect 447416 5568 447468 5574
rect 447416 5510 447468 5516
rect 446048 598 446260 626
rect 446048 490 446076 598
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 445772 462 446076 490
rect 446232 480 446260 598
rect 447428 480 447456 5510
rect 447796 3058 447824 77823
rect 448612 76628 448664 76634
rect 448612 76570 448664 76576
rect 448624 16574 448652 76570
rect 448624 16546 449112 16574
rect 449084 3482 449112 16546
rect 449176 3874 449204 84934
rect 453304 82476 453356 82482
rect 453304 82418 453356 82424
rect 450542 79384 450598 79393
rect 450542 79319 450598 79328
rect 449900 72616 449952 72622
rect 449900 72558 449952 72564
rect 449912 6914 449940 72558
rect 450556 16574 450584 79319
rect 453316 16574 453344 82418
rect 454040 19984 454092 19990
rect 454040 19926 454092 19932
rect 450556 16546 450676 16574
rect 453316 16546 453436 16574
rect 449912 6886 450584 6914
rect 449164 3868 449216 3874
rect 449164 3810 449216 3816
rect 450556 3482 450584 6886
rect 450648 3806 450676 16546
rect 453304 3868 453356 3874
rect 453304 3810 453356 3816
rect 450636 3800 450688 3806
rect 450636 3742 450688 3748
rect 452108 3732 452160 3738
rect 452108 3674 452160 3680
rect 449084 3454 449848 3482
rect 450556 3454 450952 3482
rect 447784 3052 447836 3058
rect 447784 2994 447836 3000
rect 448612 3052 448664 3058
rect 448612 2994 448664 3000
rect 448624 480 448652 2994
rect 449820 480 449848 3454
rect 450924 480 450952 3454
rect 452120 480 452148 3674
rect 453316 480 453344 3810
rect 453408 3738 453436 16546
rect 453396 3732 453448 3738
rect 453396 3674 453448 3680
rect 454052 490 454080 19926
rect 454696 7614 454724 97446
rect 461584 97436 461636 97442
rect 461584 97378 461636 97384
rect 457444 89140 457496 89146
rect 457444 89082 457496 89088
rect 456892 69760 456944 69766
rect 456892 69702 456944 69708
rect 454684 7608 454736 7614
rect 454684 7550 454736 7556
rect 455696 3664 455748 3670
rect 455696 3606 455748 3612
rect 454328 598 454540 626
rect 454328 490 454356 598
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454052 462 454356 490
rect 454512 480 454540 598
rect 455708 480 455736 3606
rect 456904 480 456932 69702
rect 457456 3126 457484 89082
rect 459560 69692 459612 69698
rect 459560 69634 459612 69640
rect 459572 16574 459600 69634
rect 460940 22772 460992 22778
rect 460940 22714 460992 22720
rect 459572 16546 459968 16574
rect 459192 9172 459244 9178
rect 459192 9114 459244 9120
rect 458088 3800 458140 3806
rect 458088 3742 458140 3748
rect 457444 3120 457496 3126
rect 457444 3062 457496 3068
rect 458100 480 458128 3742
rect 459204 480 459232 9114
rect 459940 490 459968 16546
rect 460952 6914 460980 22714
rect 461596 10334 461624 97378
rect 468484 97368 468536 97374
rect 468484 97310 468536 97316
rect 465078 89176 465134 89185
rect 465078 89111 465134 89120
rect 463700 82408 463752 82414
rect 463700 82350 463752 82356
rect 463712 16574 463740 82350
rect 465092 16574 465120 89111
rect 466460 71052 466512 71058
rect 466460 70994 466512 71000
rect 466472 16574 466500 70994
rect 467840 51740 467892 51746
rect 467840 51682 467892 51688
rect 467852 16574 467880 51682
rect 463712 16546 464016 16574
rect 465092 16546 465856 16574
rect 466472 16546 467512 16574
rect 467852 16546 468248 16574
rect 461584 10328 461636 10334
rect 461584 10270 461636 10276
rect 460952 6886 461624 6914
rect 460216 598 460428 626
rect 460216 490 460244 598
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 459940 462 460244 490
rect 460400 480 460428 598
rect 461596 480 461624 6886
rect 462780 3120 462832 3126
rect 462780 3062 462832 3068
rect 462792 480 462820 3062
rect 463988 480 464016 16546
rect 465172 7608 465224 7614
rect 465172 7550 465224 7556
rect 465184 480 465212 7550
rect 465828 490 465856 16546
rect 466104 598 466316 626
rect 466104 490 466132 598
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 465828 462 466132 490
rect 466288 480 466316 598
rect 467484 480 467512 16546
rect 468220 490 468248 16546
rect 468496 7614 468524 97310
rect 472622 86320 472678 86329
rect 472622 86255 472678 86264
rect 470600 82340 470652 82346
rect 470600 82282 470652 82288
rect 468484 7608 468536 7614
rect 468484 7550 468536 7556
rect 469864 3596 469916 3602
rect 469864 3538 469916 3544
rect 468496 598 468708 626
rect 468496 490 468524 598
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468220 462 468524 490
rect 468680 480 468708 598
rect 469876 480 469904 3538
rect 470612 490 470640 82282
rect 472256 10328 472308 10334
rect 472256 10270 472308 10276
rect 470888 598 471100 626
rect 470888 490 470916 598
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 470612 462 470916 490
rect 471072 480 471100 598
rect 472268 480 472296 10270
rect 472636 3602 472664 86255
rect 474740 21412 474792 21418
rect 474740 21354 474792 21360
rect 474752 6914 474780 21354
rect 475396 16574 475424 98670
rect 479524 98660 479576 98666
rect 479524 98602 479576 98608
rect 476120 89072 476172 89078
rect 476120 89014 476172 89020
rect 476132 16574 476160 89014
rect 475396 16546 475516 16574
rect 476132 16546 476528 16574
rect 474752 6886 475424 6914
rect 474554 4856 474610 4865
rect 474554 4791 474610 4800
rect 472624 3596 472676 3602
rect 472624 3538 472676 3544
rect 473452 3596 473504 3602
rect 473452 3538 473504 3544
rect 473464 480 473492 3538
rect 474568 480 474596 4791
rect 475396 3482 475424 6886
rect 475488 3670 475516 16546
rect 475476 3664 475528 3670
rect 475476 3606 475528 3612
rect 475396 3454 475792 3482
rect 475764 480 475792 3454
rect 476500 490 476528 16546
rect 479340 7608 479392 7614
rect 479340 7550 479392 7556
rect 478144 3732 478196 3738
rect 478144 3674 478196 3680
rect 476776 598 476988 626
rect 476776 490 476804 598
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476500 462 476804 490
rect 476960 480 476988 598
rect 478156 480 478184 3674
rect 479352 480 479380 7550
rect 479536 3058 479564 98602
rect 483020 98048 483072 98054
rect 483020 97990 483072 97996
rect 481640 79416 481692 79422
rect 481640 79358 481692 79364
rect 481652 3602 481680 79358
rect 481732 75336 481784 75342
rect 481732 75278 481784 75284
rect 481640 3596 481692 3602
rect 481640 3538 481692 3544
rect 479524 3052 479576 3058
rect 479524 2994 479576 3000
rect 480536 3052 480588 3058
rect 480536 2994 480588 3000
rect 480548 480 480576 2994
rect 481744 480 481772 75278
rect 483032 16574 483060 97990
rect 489918 93256 489974 93265
rect 489918 93191 489974 93200
rect 484400 89004 484452 89010
rect 484400 88946 484452 88952
rect 484412 16574 484440 88946
rect 489184 87780 489236 87786
rect 489184 87722 489236 87728
rect 485780 82272 485832 82278
rect 485780 82214 485832 82220
rect 485792 16574 485820 82214
rect 488540 75268 488592 75274
rect 488540 75210 488592 75216
rect 488552 16574 488580 75210
rect 483032 16546 484072 16574
rect 484412 16546 484808 16574
rect 485792 16546 486464 16574
rect 488552 16546 488856 16574
rect 482836 3596 482888 3602
rect 482836 3538 482888 3544
rect 482848 480 482876 3538
rect 484044 480 484072 16546
rect 484780 490 484808 16546
rect 485056 598 485268 626
rect 485056 490 485084 598
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 484780 462 485084 490
rect 485240 480 485268 598
rect 486436 480 486464 16546
rect 487620 3664 487672 3670
rect 487620 3606 487672 3612
rect 487632 480 487660 3606
rect 488828 480 488856 16546
rect 489196 3602 489224 87722
rect 489184 3596 489236 3602
rect 489184 3538 489236 3544
rect 489932 480 489960 93191
rect 491300 75200 491352 75206
rect 491300 75142 491352 75148
rect 491312 16574 491340 75142
rect 492680 65544 492732 65550
rect 492680 65486 492732 65492
rect 492692 16574 492720 65486
rect 491312 16546 492352 16574
rect 492692 16546 493088 16574
rect 491116 3664 491168 3670
rect 491116 3606 491168 3612
rect 491128 480 491156 3606
rect 492324 480 492352 16546
rect 493060 490 493088 16546
rect 493336 3398 493364 98903
rect 494058 98832 494114 98841
rect 494058 98767 494114 98776
rect 494072 3670 494100 98767
rect 500960 96076 501012 96082
rect 500960 96018 501012 96024
rect 497462 95976 497518 95985
rect 497462 95911 497518 95920
rect 495440 74112 495492 74118
rect 495440 74054 495492 74060
rect 494060 3664 494112 3670
rect 494060 3606 494112 3612
rect 493324 3392 493376 3398
rect 493324 3334 493376 3340
rect 494704 3392 494756 3398
rect 494704 3334 494756 3340
rect 493336 598 493548 626
rect 493336 490 493364 598
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493060 462 493364 490
rect 493520 480 493548 598
rect 494716 480 494744 3334
rect 495452 490 495480 74054
rect 497096 13116 497148 13122
rect 497096 13058 497148 13064
rect 495728 598 495940 626
rect 495728 490 495756 598
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495452 462 495756 490
rect 495912 480 495940 598
rect 497108 480 497136 13058
rect 497476 3670 497504 95911
rect 499580 82204 499632 82210
rect 499580 82146 499632 82152
rect 499592 16574 499620 82146
rect 500972 16574 501000 96018
rect 502340 87712 502392 87718
rect 502340 87654 502392 87660
rect 502352 16574 502380 87654
rect 503720 46232 503772 46238
rect 503720 46174 503772 46180
rect 499592 16546 500632 16574
rect 500972 16546 501368 16574
rect 502352 16546 503024 16574
rect 498200 6384 498252 6390
rect 498200 6326 498252 6332
rect 497464 3664 497516 3670
rect 497464 3606 497516 3612
rect 498212 480 498240 6326
rect 499396 3732 499448 3738
rect 499396 3674 499448 3680
rect 499408 480 499436 3674
rect 500604 480 500632 16546
rect 501340 490 501368 16546
rect 501616 598 501828 626
rect 501616 490 501644 598
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501340 462 501644 490
rect 501800 480 501828 598
rect 502996 480 503024 16546
rect 503732 490 503760 46174
rect 504376 3398 504404 99486
rect 512000 99476 512052 99482
rect 512000 99418 512052 99424
rect 507860 96008 507912 96014
rect 507860 95950 507912 95956
rect 506480 84924 506532 84930
rect 506480 84866 506532 84872
rect 506492 16574 506520 84866
rect 507872 16574 507900 95950
rect 510712 84856 510764 84862
rect 510712 84798 510764 84804
rect 506492 16546 507256 16574
rect 507872 16546 508912 16574
rect 506480 3800 506532 3806
rect 506480 3742 506532 3748
rect 504364 3392 504416 3398
rect 504364 3334 504416 3340
rect 505376 3392 505428 3398
rect 505376 3334 505428 3340
rect 504008 598 504220 626
rect 504008 490 504036 598
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 503732 462 504036 490
rect 504192 480 504220 598
rect 505388 480 505416 3334
rect 506492 480 506520 3742
rect 507228 490 507256 16546
rect 507504 598 507716 626
rect 507504 490 507532 598
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507228 462 507532 490
rect 507688 480 507716 598
rect 508884 480 508912 16546
rect 510724 3738 510752 84798
rect 511264 9104 511316 9110
rect 511264 9046 511316 9052
rect 510712 3732 510764 3738
rect 510712 3674 510764 3680
rect 510068 3596 510120 3602
rect 510068 3538 510120 3544
rect 510080 480 510108 3538
rect 511276 480 511304 9046
rect 512012 490 512040 99418
rect 520372 99408 520424 99414
rect 520372 99350 520424 99356
rect 518900 95940 518952 95946
rect 518900 95882 518952 95888
rect 515404 86420 515456 86426
rect 515404 86362 515456 86368
rect 513380 74044 513432 74050
rect 513380 73986 513432 73992
rect 513392 16574 513420 73986
rect 514758 71088 514814 71097
rect 514758 71023 514814 71032
rect 513392 16546 513604 16574
rect 512288 598 512500 626
rect 512288 490 512316 598
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512012 462 512316 490
rect 512472 480 512500 598
rect 513576 480 513604 16546
rect 514772 480 514800 71023
rect 515416 3874 515444 86362
rect 517610 75168 517666 75177
rect 517610 75103 517666 75112
rect 517520 14476 517572 14482
rect 517520 14418 517572 14424
rect 515404 3868 515456 3874
rect 515404 3810 515456 3816
rect 517152 3800 517204 3806
rect 517152 3742 517204 3748
rect 515956 3732 516008 3738
rect 515956 3674 516008 3680
rect 515968 480 515996 3674
rect 517164 480 517192 3742
rect 517532 626 517560 14418
rect 517624 3942 517652 75103
rect 517612 3936 517664 3942
rect 517612 3878 517664 3884
rect 518912 3738 518940 95882
rect 518900 3732 518952 3738
rect 518900 3674 518952 3680
rect 520384 3602 520412 99350
rect 525798 95840 525854 95849
rect 525798 95775 525854 95784
rect 525064 82136 525116 82142
rect 525064 82078 525116 82084
rect 522302 80880 522358 80889
rect 522302 80815 522358 80824
rect 521660 73976 521712 73982
rect 521660 73918 521712 73924
rect 521672 16574 521700 73918
rect 521672 16546 521884 16574
rect 520740 9036 520792 9042
rect 520740 8978 520792 8984
rect 519544 3596 519596 3602
rect 519544 3538 519596 3544
rect 520372 3596 520424 3602
rect 520372 3538 520424 3544
rect 517532 598 517928 626
rect 517900 490 517928 598
rect 518176 598 518388 626
rect 518176 490 518204 598
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 517900 462 518204 490
rect 518360 480 518388 598
rect 519556 480 519584 3538
rect 520752 480 520780 8978
rect 521856 480 521884 16546
rect 522316 3602 522344 80815
rect 525076 3806 525104 82078
rect 525812 16574 525840 95775
rect 528652 87644 528704 87650
rect 528652 87586 528704 87592
rect 527180 73908 527232 73914
rect 527180 73850 527232 73856
rect 527192 16574 527220 73850
rect 528560 24132 528612 24138
rect 528560 24074 528612 24080
rect 525812 16546 526208 16574
rect 527192 16546 527864 16574
rect 525432 3868 525484 3874
rect 525432 3810 525484 3816
rect 525064 3800 525116 3806
rect 525064 3742 525116 3748
rect 523040 3664 523092 3670
rect 523040 3606 523092 3612
rect 524236 3664 524288 3670
rect 524236 3606 524288 3612
rect 522304 3596 522356 3602
rect 522304 3538 522356 3544
rect 523052 480 523080 3606
rect 524248 480 524276 3606
rect 525444 480 525472 3810
rect 526180 490 526208 16546
rect 526456 598 526668 626
rect 526456 490 526484 598
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526180 462 526484 490
rect 526640 480 526668 598
rect 527836 480 527864 16546
rect 528572 490 528600 24074
rect 528664 3738 528692 87586
rect 529952 16574 529980 99583
rect 550638 99512 550694 99521
rect 550638 99447 550694 99456
rect 532698 98696 532754 98705
rect 532698 98631 532754 98640
rect 531412 72480 531464 72486
rect 531412 72422 531464 72428
rect 531424 16574 531452 72422
rect 532712 16574 532740 98631
rect 539600 93288 539652 93294
rect 539600 93230 539652 93236
rect 538218 87816 538274 87825
rect 538218 87751 538274 87760
rect 536838 87680 536894 87689
rect 536838 87615 536894 87624
rect 535460 80912 535512 80918
rect 535460 80854 535512 80860
rect 535472 16574 535500 80854
rect 529952 16546 530164 16574
rect 531424 16546 532096 16574
rect 532712 16546 533752 16574
rect 535472 16546 536144 16574
rect 528652 3732 528704 3738
rect 528652 3674 528704 3680
rect 528848 598 529060 626
rect 528848 490 528876 598
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528572 462 528876 490
rect 529032 480 529060 598
rect 530136 480 530164 16546
rect 531320 3800 531372 3806
rect 531320 3742 531372 3748
rect 531332 480 531360 3742
rect 532068 490 532096 16546
rect 532344 598 532556 626
rect 532344 490 532372 598
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532068 462 532372 490
rect 532528 480 532556 598
rect 533724 480 533752 16546
rect 534908 3732 534960 3738
rect 534908 3674 534960 3680
rect 534920 480 534948 3674
rect 536116 480 536144 16546
rect 536852 3670 536880 87615
rect 538232 16574 538260 87751
rect 538232 16546 538444 16574
rect 536840 3664 536892 3670
rect 536840 3606 536892 3612
rect 537208 3460 537260 3466
rect 537208 3402 537260 3408
rect 537220 480 537248 3402
rect 538416 480 538444 16546
rect 539612 480 539640 93230
rect 546592 93220 546644 93226
rect 546592 93162 546644 93168
rect 542360 80844 542412 80850
rect 542360 80786 542412 80792
rect 542372 16574 542400 80786
rect 542372 16546 542768 16574
rect 540796 6316 540848 6322
rect 540796 6258 540848 6264
rect 540808 480 540836 6258
rect 541992 3664 542044 3670
rect 541992 3606 542044 3612
rect 542004 480 542032 3606
rect 542740 490 542768 16546
rect 546500 15904 546552 15910
rect 546500 15846 546552 15852
rect 545486 11656 545542 11665
rect 545486 11591 545542 11600
rect 544384 6248 544436 6254
rect 544384 6190 544436 6196
rect 543016 598 543228 626
rect 543016 490 543044 598
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 542740 462 543044 490
rect 543200 480 543228 598
rect 544396 480 544424 6190
rect 545500 480 545528 11591
rect 546512 3482 546540 15846
rect 546604 3738 546632 93162
rect 547880 86352 547932 86358
rect 547880 86294 547932 86300
rect 547892 16574 547920 86294
rect 547892 16546 548656 16574
rect 546592 3732 546644 3738
rect 546592 3674 546644 3680
rect 546512 3454 546724 3482
rect 546696 480 546724 3454
rect 547880 3120 547932 3126
rect 547880 3062 547932 3068
rect 547892 480 547920 3062
rect 548628 490 548656 16546
rect 550272 3596 550324 3602
rect 550272 3538 550324 3544
rect 548904 598 549116 626
rect 548904 490 548932 598
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 548628 462 548932 490
rect 549088 480 549116 598
rect 550284 480 550312 3538
rect 550652 3126 550680 99447
rect 557540 94648 557592 94654
rect 557540 94590 557592 94596
rect 553398 93120 553454 93129
rect 553398 93055 553454 93064
rect 553412 16574 553440 93055
rect 554778 87544 554834 87553
rect 554778 87479 554834 87488
rect 553412 16546 553808 16574
rect 552664 3596 552716 3602
rect 552664 3538 552716 3544
rect 551468 3528 551520 3534
rect 551468 3470 551520 3476
rect 550640 3120 550692 3126
rect 550640 3062 550692 3068
rect 551480 480 551508 3470
rect 552676 480 552704 3538
rect 553780 480 553808 16546
rect 554792 3670 554820 87479
rect 557552 16574 557580 94590
rect 561680 94580 561732 94586
rect 561680 94522 561732 94528
rect 560300 80776 560352 80782
rect 560300 80718 560352 80724
rect 560312 16574 560340 80718
rect 561692 16574 561720 94522
rect 565820 94512 565872 94518
rect 565820 94454 565872 94460
rect 564440 93152 564492 93158
rect 564440 93094 564492 93100
rect 557552 16546 558592 16574
rect 560312 16546 560432 16574
rect 561692 16546 562088 16574
rect 556160 3800 556212 3806
rect 556160 3742 556212 3748
rect 554780 3664 554832 3670
rect 554780 3606 554832 3612
rect 554964 3460 555016 3466
rect 554964 3402 555016 3408
rect 554976 480 555004 3402
rect 556172 480 556200 3742
rect 557356 3664 557408 3670
rect 557356 3606 557408 3612
rect 557368 480 557396 3606
rect 558564 480 558592 16546
rect 559748 3528 559800 3534
rect 559748 3470 559800 3476
rect 559760 480 559788 3470
rect 560404 490 560432 16546
rect 560680 598 560892 626
rect 560680 490 560708 598
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560404 462 560708 490
rect 560864 480 560892 598
rect 562060 480 562088 16546
rect 564452 3754 564480 93094
rect 563244 3732 563296 3738
rect 563244 3674 563296 3680
rect 564360 3726 564480 3754
rect 563256 480 563284 3674
rect 564360 3602 564388 3726
rect 564348 3596 564400 3602
rect 564348 3538 564400 3544
rect 564440 3596 564492 3602
rect 564440 3538 564492 3544
rect 564452 480 564480 3538
rect 565832 3482 565860 94454
rect 566832 3868 566884 3874
rect 566832 3810 566884 3816
rect 565648 3454 565860 3482
rect 565648 480 565676 3454
rect 566844 480 566872 3810
rect 568592 3806 568620 100710
rect 574098 89040 574154 89049
rect 574098 88975 574154 88984
rect 572720 86284 572772 86290
rect 572720 86226 572772 86232
rect 571340 83496 571392 83502
rect 571340 83438 571392 83444
rect 569960 76560 570012 76566
rect 569960 76502 570012 76508
rect 569132 6180 569184 6186
rect 569132 6122 569184 6128
rect 568580 3800 568632 3806
rect 568580 3742 568632 3748
rect 568026 3360 568082 3369
rect 568026 3295 568082 3304
rect 568040 480 568068 3295
rect 569144 480 569172 6122
rect 569972 3670 570000 76502
rect 571352 3874 571380 83438
rect 572732 16574 572760 86226
rect 572732 16546 572852 16574
rect 571340 3868 571392 3874
rect 571340 3810 571392 3816
rect 572720 3868 572772 3874
rect 572720 3810 572772 3816
rect 570328 3800 570380 3806
rect 570328 3742 570380 3748
rect 569960 3664 570012 3670
rect 569960 3606 570012 3612
rect 570340 480 570368 3742
rect 571524 3664 571576 3670
rect 571524 3606 571576 3612
rect 571536 480 571564 3606
rect 572732 480 572760 3810
rect 572824 3534 572852 16546
rect 574112 3534 574140 88975
rect 575570 86184 575626 86193
rect 575570 86119 575626 86128
rect 575112 3936 575164 3942
rect 575112 3878 575164 3884
rect 572812 3528 572864 3534
rect 572812 3470 572864 3476
rect 574100 3528 574152 3534
rect 574100 3470 574152 3476
rect 573916 3460 573968 3466
rect 573916 3402 573968 3408
rect 573928 480 573956 3402
rect 575124 480 575152 3878
rect 575584 3738 575612 86119
rect 579618 80744 579674 80753
rect 578240 80708 578292 80714
rect 579618 80679 579674 80688
rect 578240 80650 578292 80656
rect 576308 8968 576360 8974
rect 576308 8910 576360 8916
rect 575572 3732 575624 3738
rect 575572 3674 575624 3680
rect 576320 480 576348 8910
rect 578252 3602 578280 80650
rect 578240 3596 578292 3602
rect 578240 3538 578292 3544
rect 577412 3528 577464 3534
rect 577412 3470 577464 3476
rect 577424 480 577452 3470
rect 579632 3369 579660 80679
rect 582378 50280 582434 50289
rect 582378 50215 582434 50224
rect 582194 3632 582250 3641
rect 582194 3567 582250 3576
rect 580998 3496 581054 3505
rect 580998 3431 581054 3440
rect 579618 3360 579674 3369
rect 579618 3295 579674 3304
rect 578608 3052 578660 3058
rect 578608 2994 578660 3000
rect 578620 480 578648 2994
rect 581012 480 581040 3431
rect 582208 480 582236 3567
rect 582392 3058 582420 50215
rect 582484 19825 582512 204274
rect 583128 203561 583156 537775
rect 583206 511320 583262 511329
rect 583206 511255 583262 511264
rect 583220 204950 583248 511255
rect 583298 484664 583354 484673
rect 583298 484599 583354 484608
rect 583312 209098 583340 484599
rect 583404 458862 583432 683839
rect 583482 577280 583538 577289
rect 583482 577215 583538 577224
rect 583392 458856 583444 458862
rect 583392 458798 583444 458804
rect 583390 404968 583446 404977
rect 583390 404903 583446 404912
rect 583300 209092 583352 209098
rect 583300 209034 583352 209040
rect 583404 207738 583432 404903
rect 583496 403646 583524 577215
rect 583666 524784 583722 524793
rect 583666 524719 583722 524728
rect 583574 471064 583630 471073
rect 583574 470999 583630 471008
rect 583484 403640 583536 403646
rect 583484 403582 583536 403588
rect 583484 343256 583536 343262
rect 583484 343198 583536 343204
rect 583392 207732 583444 207738
rect 583392 207674 583444 207680
rect 583208 204944 583260 204950
rect 583208 204886 583260 204892
rect 583392 204400 583444 204406
rect 583392 204342 583444 204348
rect 583114 203552 583170 203561
rect 583114 203487 583170 203496
rect 583024 203108 583076 203114
rect 583024 203050 583076 203056
rect 582656 203040 582708 203046
rect 582656 202982 582708 202988
rect 582668 86193 582696 202982
rect 583036 99521 583064 203050
rect 583208 201952 583260 201958
rect 583208 201894 583260 201900
rect 583116 198076 583168 198082
rect 583116 198018 583168 198024
rect 583128 112849 583156 198018
rect 583220 126041 583248 201894
rect 583300 201612 583352 201618
rect 583300 201554 583352 201560
rect 583312 139369 583340 201554
rect 583404 152697 583432 204342
rect 583496 202201 583524 343198
rect 583588 300150 583616 470999
rect 583680 354006 583708 524719
rect 583668 354000 583720 354006
rect 583668 353942 583720 353948
rect 583576 300144 583628 300150
rect 583576 300086 583628 300092
rect 583576 202972 583628 202978
rect 583576 202914 583628 202920
rect 583482 202192 583538 202201
rect 583482 202127 583538 202136
rect 583482 200152 583538 200161
rect 583482 200087 583538 200096
rect 583390 152688 583446 152697
rect 583390 152623 583446 152632
rect 583298 139360 583354 139369
rect 583298 139295 583354 139304
rect 583206 126032 583262 126041
rect 583206 125967 583262 125976
rect 583114 112840 583170 112849
rect 583114 112775 583170 112784
rect 583390 102232 583446 102241
rect 583390 102167 583446 102176
rect 583114 101008 583170 101017
rect 583114 100943 583170 100952
rect 583022 99512 583078 99521
rect 583022 99447 583078 99456
rect 582932 97300 582984 97306
rect 582932 97242 582984 97248
rect 582654 86184 582710 86193
rect 582654 86119 582710 86128
rect 582840 79348 582892 79354
rect 582840 79290 582892 79296
rect 582748 73840 582800 73846
rect 582748 73782 582800 73788
rect 582656 64184 582708 64190
rect 582656 64126 582708 64132
rect 582564 35216 582616 35222
rect 582564 35158 582616 35164
rect 582470 19816 582526 19825
rect 582470 19751 582526 19760
rect 582576 3346 582604 35158
rect 582668 3505 582696 64126
rect 582760 3534 582788 73782
rect 582852 3942 582880 79290
rect 582840 3936 582892 3942
rect 582840 3878 582892 3884
rect 582944 3641 582972 97242
rect 582930 3632 582986 3641
rect 582930 3567 582986 3576
rect 582748 3528 582800 3534
rect 582654 3496 582710 3505
rect 582748 3470 582800 3476
rect 583128 3466 583156 100943
rect 583206 100872 583262 100881
rect 583206 100807 583262 100816
rect 583220 3806 583248 100807
rect 583298 94480 583354 94489
rect 583298 94415 583354 94424
rect 583312 3874 583340 94415
rect 583404 6914 583432 102167
rect 583496 16574 583524 200087
rect 583588 46889 583616 202914
rect 583668 200184 583720 200190
rect 583668 200126 583720 200132
rect 583680 60217 583708 200126
rect 583772 198898 583800 696895
rect 583852 202904 583904 202910
rect 583852 202846 583904 202852
rect 583760 198892 583812 198898
rect 583760 198834 583812 198840
rect 583760 198008 583812 198014
rect 583760 197950 583812 197956
rect 583772 73273 583800 197950
rect 583758 73264 583814 73273
rect 583758 73199 583814 73208
rect 583666 60208 583722 60217
rect 583666 60143 583722 60152
rect 583574 46880 583630 46889
rect 583574 46815 583630 46824
rect 583864 32881 583892 202846
rect 583850 32872 583906 32881
rect 583850 32807 583906 32816
rect 583496 16546 583616 16574
rect 583404 6886 583524 6914
rect 583588 6905 583616 16546
rect 583300 3868 583352 3874
rect 583300 3810 583352 3816
rect 583208 3800 583260 3806
rect 583208 3742 583260 3748
rect 583496 3670 583524 6886
rect 583574 6896 583630 6905
rect 583574 6831 583630 6840
rect 583484 3664 583536 3670
rect 583484 3606 583536 3612
rect 582654 3431 582710 3440
rect 583116 3460 583168 3466
rect 583116 3402 583168 3408
rect 582576 3318 583432 3346
rect 582380 3052 582432 3058
rect 582380 2994 582432 3000
rect 583404 480 583432 3318
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 3514 671200 3570 671256
rect 3422 658144 3478 658200
rect 3422 632068 3424 632088
rect 3424 632068 3476 632088
rect 3476 632068 3478 632088
rect 3422 632032 3478 632068
rect 3146 619112 3202 619168
rect 3238 606056 3294 606112
rect 3330 579944 3386 580000
rect 3422 566888 3478 566944
rect 3422 553832 3478 553888
rect 3422 527856 3478 527912
rect 3422 514820 3478 514856
rect 3422 514800 3424 514820
rect 3424 514800 3476 514820
rect 3476 514800 3478 514820
rect 3422 501744 3478 501800
rect 3054 475632 3110 475688
rect 3146 449520 3202 449576
rect 2870 410488 2926 410544
rect 3146 358400 3202 358456
rect 3330 345344 3386 345400
rect 3330 319232 3386 319288
rect 3054 267144 3110 267200
rect 3054 241032 3110 241088
rect 3514 462576 3570 462632
rect 3514 423544 3570 423600
rect 3514 397468 3516 397488
rect 3516 397468 3568 397488
rect 3568 397468 3570 397488
rect 3514 397432 3570 397468
rect 3514 371320 3570 371376
rect 3514 306176 3570 306232
rect 3514 293120 3570 293176
rect 3514 254088 3570 254144
rect 3146 214920 3202 214976
rect 73066 205128 73122 205184
rect 106186 203632 106242 203688
rect 3238 201864 3294 201920
rect 3238 162832 3294 162888
rect 3514 188808 3570 188864
rect 3422 149776 3478 149832
rect 3238 136720 3294 136776
rect 3422 110608 3478 110664
rect 3422 97552 3478 97608
rect 3146 84632 3202 84688
rect 3422 71576 3478 71632
rect 3054 58520 3110 58576
rect 3422 45500 3424 45520
rect 3424 45500 3476 45520
rect 3476 45500 3478 45520
rect 3422 45464 3478 45500
rect 2870 32408 2926 32464
rect 3422 19352 3478 19408
rect 3422 6432 3478 6488
rect 15842 100952 15898 101008
rect 30286 98640 30342 98696
rect 18602 95784 18658 95840
rect 15934 3440 15990 3496
rect 26146 93064 26202 93120
rect 28262 91704 28318 91760
rect 27526 87488 27582 87544
rect 34426 93200 34482 93256
rect 35254 82048 35310 82104
rect 35806 73752 35862 73808
rect 46202 97144 46258 97200
rect 49606 80688 49662 80744
rect 57886 84768 57942 84824
rect 75182 87624 75238 87680
rect 80702 98776 80758 98832
rect 79966 88984 80022 89040
rect 83462 84904 83518 84960
rect 92386 73888 92442 73944
rect 97906 89120 97962 89176
rect 101494 79328 101550 79384
rect 130382 95920 130438 95976
rect 125506 93336 125562 93392
rect 107566 44784 107622 44840
rect 114466 77832 114522 77888
rect 122746 79464 122802 79520
rect 133234 83408 133290 83464
rect 200394 200096 200450 200152
rect 222382 202136 222438 202192
rect 231674 204856 231730 204912
rect 230386 203496 230442 203552
rect 237194 206216 237250 206272
rect 235998 204992 236054 205048
rect 242530 207576 242586 207632
rect 242990 202816 243046 202872
rect 244922 202816 244978 202872
rect 244738 202680 244794 202736
rect 246026 202680 246082 202736
rect 250626 202544 250682 202600
rect 252650 202816 252706 202872
rect 253386 202544 253442 202600
rect 255318 203632 255374 203688
rect 255134 202816 255190 202872
rect 255318 201864 255374 201920
rect 255962 203768 256018 203824
rect 258630 205128 258686 205184
rect 257710 201864 257766 201920
rect 259182 202816 259238 202872
rect 260378 202816 260434 202872
rect 268198 203768 268254 203824
rect 305642 207576 305698 207632
rect 582470 670656 582526 670712
rect 580170 458088 580226 458144
rect 580170 431568 580226 431624
rect 580170 418240 580226 418296
rect 580906 378392 580962 378448
rect 580170 365064 580226 365120
rect 579894 351908 579896 351928
rect 579896 351908 579948 351928
rect 579948 351908 579950 351928
rect 579894 351872 579950 351908
rect 580170 325216 580226 325272
rect 580170 312024 580226 312080
rect 580906 298696 580962 298752
rect 580170 272176 580226 272232
rect 580170 258848 580226 258904
rect 580170 232328 580226 232384
rect 580170 219000 580226 219056
rect 580170 205692 580226 205728
rect 580170 205672 580172 205692
rect 580172 205672 580224 205692
rect 580224 205672 580226 205692
rect 582562 644000 582618 644056
rect 582654 630808 582710 630864
rect 582470 206216 582526 206272
rect 582746 617480 582802 617536
rect 582838 590960 582894 591016
rect 583758 696904 583814 696960
rect 583390 683848 583446 683904
rect 583022 564304 583078 564360
rect 582930 245520 582986 245576
rect 582654 204992 582710 205048
rect 583114 537784 583170 537840
rect 583022 204856 583078 204912
rect 199842 199552 199898 199608
rect 198002 199280 198058 199336
rect 170402 173236 170458 173292
rect 169298 161492 169354 161528
rect 169298 161472 169300 161492
rect 169300 161472 169352 161492
rect 169352 161472 169354 161492
rect 169390 144200 169446 144256
rect 172426 189216 172482 189272
rect 171782 187720 171838 187776
rect 172426 186768 172482 186824
rect 171782 185408 171838 185464
rect 171690 184184 171746 184240
rect 172426 183660 172482 183696
rect 172426 183640 172428 183660
rect 172428 183640 172480 183660
rect 172480 183640 172482 183660
rect 172426 182416 172482 182472
rect 172426 181056 172482 181112
rect 172058 179832 172114 179888
rect 172150 178608 172206 178664
rect 172242 177248 172298 177304
rect 172426 176740 172428 176760
rect 172428 176740 172480 176760
rect 172480 176740 172482 176760
rect 172426 176704 172482 176740
rect 172426 175344 172482 175400
rect 171966 174120 172022 174176
rect 171782 169768 171838 169824
rect 171138 164736 171194 164792
rect 171690 163376 171746 163432
rect 171690 153176 171746 153232
rect 171506 152632 171562 152688
rect 171322 150456 171378 150512
rect 171506 149368 171562 149424
rect 171322 148316 171324 148336
rect 171324 148316 171376 148336
rect 171376 148316 171378 148336
rect 171322 148280 171378 148316
rect 171690 147736 171746 147792
rect 171322 143520 171378 143576
rect 171690 142976 171746 143032
rect 171506 141888 171562 141944
rect 171506 140800 171562 140856
rect 171690 139712 171746 139768
rect 171322 138624 171378 138680
rect 170494 137536 170550 137592
rect 171506 136992 171562 137048
rect 171690 135904 171746 135960
rect 171506 135360 171562 135416
rect 171506 134272 171562 134328
rect 171690 132776 171746 132832
rect 171690 132232 171746 132288
rect 171690 130600 171746 130656
rect 170402 129512 170458 129568
rect 171598 128968 171654 129024
rect 171690 127880 171746 127936
rect 171690 124616 171746 124672
rect 171874 162988 171930 163024
rect 171874 162968 171876 162988
rect 171876 162968 171928 162988
rect 171928 162968 171930 162988
rect 171874 160384 171930 160440
rect 172242 171672 172298 171728
rect 172242 170312 172298 170368
rect 172426 168544 172482 168600
rect 172426 167320 172482 167376
rect 172426 165960 172482 166016
rect 171874 149912 171930 149968
rect 172242 153720 172298 153776
rect 172334 152088 172390 152144
rect 172334 151544 172390 151600
rect 172426 151000 172482 151056
rect 171966 146648 172022 146704
rect 172150 146124 172206 146160
rect 172150 146104 172152 146124
rect 172152 146104 172204 146124
rect 172204 146104 172206 146124
rect 172426 148824 172482 148880
rect 172426 147192 172482 147248
rect 172426 145560 172482 145616
rect 172334 145016 172390 145072
rect 172242 144472 172298 144528
rect 172426 142432 172482 142488
rect 172426 141344 172482 141400
rect 172426 140256 172482 140312
rect 172426 139204 172428 139224
rect 172428 139204 172480 139224
rect 172480 139204 172482 139224
rect 172426 139168 172482 139204
rect 171966 138080 172022 138136
rect 172426 136448 172482 136504
rect 171874 134816 171930 134872
rect 171874 133864 171930 133920
rect 172426 133356 172428 133376
rect 172428 133356 172480 133376
rect 172480 133356 172482 133376
rect 172426 133320 172482 133356
rect 172426 131724 172428 131744
rect 172428 131724 172480 131744
rect 172480 131724 172482 131744
rect 172426 131688 172482 131724
rect 172426 131164 172482 131200
rect 172426 131144 172428 131164
rect 172428 131144 172480 131164
rect 172480 131144 172482 131164
rect 172058 130056 172114 130112
rect 172426 128444 172482 128480
rect 172426 128424 172428 128444
rect 172428 128424 172480 128444
rect 172480 128424 172482 128444
rect 172058 127336 172114 127392
rect 172334 126792 172390 126848
rect 172150 126248 172206 126304
rect 171874 125160 171930 125216
rect 172426 125724 172482 125760
rect 172426 125704 172428 125724
rect 172428 125704 172480 125724
rect 172480 125704 172482 125724
rect 172426 124228 172482 124264
rect 172426 124208 172428 124228
rect 172428 124208 172480 124228
rect 172480 124208 172482 124228
rect 198002 198192 198058 198248
rect 198646 197104 198702 197160
rect 198002 196036 198058 196072
rect 198002 196016 198004 196036
rect 198004 196016 198056 196036
rect 198056 196016 198058 196036
rect 198094 194928 198150 194984
rect 197726 193840 197782 193896
rect 197634 192752 197690 192808
rect 198094 191664 198150 191720
rect 197358 190576 197414 190632
rect 197910 189488 197966 189544
rect 197358 188400 197414 188456
rect 197542 187312 197598 187368
rect 197634 186244 197690 186280
rect 197634 186224 197636 186244
rect 197636 186224 197688 186244
rect 197688 186224 197690 186244
rect 197358 185000 197414 185056
rect 198370 183912 198426 183968
rect 197726 182824 197782 182880
rect 197358 181736 197414 181792
rect 204074 199552 204130 199608
rect 207662 199552 207718 199608
rect 211250 199552 211306 199608
rect 246210 199552 246266 199608
rect 246486 199552 246542 199608
rect 580170 192480 580226 192536
rect 197358 180648 197414 180704
rect 198094 179560 198150 179616
rect 197910 178472 197966 178528
rect 197818 177384 197874 177440
rect 197358 176296 197414 176352
rect 197358 174120 197414 174176
rect 197726 170720 197782 170776
rect 197450 169632 197506 169688
rect 197358 166368 197414 166424
rect 197358 164192 197414 164248
rect 197726 168564 197782 168600
rect 197726 168544 197728 168564
rect 197728 168544 197780 168564
rect 197780 168544 197782 168564
rect 197910 167456 197966 167512
rect 197634 165280 197690 165336
rect 197634 163104 197690 163160
rect 197358 162016 197414 162072
rect 197542 159840 197598 159896
rect 197910 158752 197966 158808
rect 197358 157664 197414 157720
rect 197726 155352 197782 155408
rect 197358 154264 197414 154320
rect 197358 153212 197360 153232
rect 197360 153212 197412 153232
rect 197412 153212 197414 153232
rect 197358 153176 197414 153212
rect 197450 151000 197506 151056
rect 197358 149912 197414 149968
rect 197542 148824 197598 148880
rect 197358 145560 197414 145616
rect 197450 144472 197506 144528
rect 197358 143384 197414 143440
rect 197358 142180 197414 142216
rect 197358 142160 197360 142180
rect 197360 142160 197412 142180
rect 197412 142160 197414 142180
rect 197358 139984 197414 140040
rect 197542 137808 197598 137864
rect 197358 134544 197414 134600
rect 197450 133456 197506 133512
rect 197358 132404 197360 132424
rect 197360 132404 197412 132424
rect 197412 132404 197414 132424
rect 197358 132368 197414 132404
rect 197910 131280 197966 131336
rect 197358 129104 197414 129160
rect 197358 126792 197414 126848
rect 198554 175208 198610 175264
rect 198462 173052 198518 173088
rect 198462 173032 198464 173052
rect 198464 173032 198516 173052
rect 198516 173032 198518 173052
rect 198738 171944 198794 172000
rect 198462 160928 198518 160984
rect 198462 156440 198518 156496
rect 198186 152088 198242 152144
rect 198094 147736 198150 147792
rect 198186 146648 198242 146704
rect 198186 141072 198242 141128
rect 198186 138896 198242 138952
rect 198462 136720 198518 136776
rect 198186 135632 198242 135688
rect 198002 130192 198058 130248
rect 198094 127880 198150 127936
rect 197450 125704 197506 125760
rect 197634 124616 197690 124672
rect 197910 123528 197966 123584
rect 197358 122440 197414 122496
rect 197358 121372 197414 121408
rect 197358 121352 197360 121372
rect 197360 121352 197412 121372
rect 197412 121352 197414 121372
rect 197542 120264 197598 120320
rect 197358 118088 197414 118144
rect 197634 115912 197690 115968
rect 197910 114860 197912 114880
rect 197912 114860 197964 114880
rect 197964 114860 197966 114880
rect 197910 114824 197966 114860
rect 197358 113600 197414 113656
rect 197358 112512 197414 112568
rect 197358 111424 197414 111480
rect 197358 110356 197414 110392
rect 197358 110336 197360 110356
rect 197360 110336 197412 110356
rect 197412 110336 197414 110356
rect 197542 109248 197598 109304
rect 580262 179152 580318 179208
rect 582378 165824 582434 165880
rect 198278 119176 198334 119232
rect 198462 117000 198518 117056
rect 198002 108160 198058 108216
rect 197542 107072 197598 107128
rect 198554 105984 198610 106040
rect 198094 104896 198150 104952
rect 197542 103808 197598 103864
rect 197450 102720 197506 102776
rect 197910 101632 197966 101688
rect 199934 100952 199990 101008
rect 298558 100680 298614 100736
rect 198094 100544 198150 100600
rect 297914 100408 297970 100464
rect 297914 100272 297970 100328
rect 153106 94424 153162 94480
rect 169666 94560 169722 94616
rect 177946 91840 178002 91896
rect 188342 97280 188398 97336
rect 186962 96056 187018 96112
rect 188342 86128 188398 86184
rect 195242 94696 195298 94752
rect 194506 90344 194562 90400
rect 200118 97280 200174 97336
rect 200854 97144 200910 97200
rect 200762 96736 200818 96792
rect 200946 96600 201002 96656
rect 201498 95784 201554 95840
rect 201958 3440 202014 3496
rect 203154 96872 203210 96928
rect 202878 96600 202934 96656
rect 204350 96600 204406 96656
rect 205178 98640 205234 98696
rect 204534 87488 204590 87544
rect 204442 82048 204498 82104
rect 205914 96872 205970 96928
rect 205730 96600 205786 96656
rect 207386 96736 207442 96792
rect 202694 3304 202750 3360
rect 208398 96600 208454 96656
rect 207754 88984 207810 89040
rect 208766 98776 208822 98832
rect 209778 96600 209834 96656
rect 211434 96600 211490 96656
rect 212630 96600 212686 96656
rect 214102 96600 214158 96656
rect 215666 96872 215722 96928
rect 216678 96872 216734 96928
rect 218334 96872 218390 96928
rect 219530 97552 219586 97608
rect 221002 96872 221058 96928
rect 222198 95920 222254 95976
rect 222382 96872 222438 96928
rect 223578 96872 223634 96928
rect 226430 96600 226486 96656
rect 229098 94560 229154 94616
rect 230478 96736 230534 96792
rect 230938 96600 230994 96656
rect 231122 96464 231178 96520
rect 232134 96600 232190 96656
rect 231950 96056 232006 96112
rect 233330 96600 233386 96656
rect 233882 81504 233938 81560
rect 237562 96872 237618 96928
rect 237838 96872 237894 96928
rect 235262 3304 235318 3360
rect 246946 96872 247002 96928
rect 249522 96872 249578 96928
rect 250994 96872 251050 96928
rect 251086 96056 251142 96112
rect 252006 97008 252062 97064
rect 252374 96872 252430 96928
rect 253662 96872 253718 96928
rect 255226 96872 255282 96928
rect 256054 96872 256110 96928
rect 257710 96872 257766 96928
rect 259090 97008 259146 97064
rect 258906 96872 258962 96928
rect 255962 3304 256018 3360
rect 260746 97008 260802 97064
rect 260562 96872 260618 96928
rect 262770 96872 262826 96928
rect 263322 96872 263378 96928
rect 264794 97008 264850 97064
rect 264334 96872 264390 96928
rect 266174 96872 266230 96928
rect 267462 97008 267518 97064
rect 267646 96872 267702 96928
rect 269026 96872 269082 96928
rect 270222 96872 270278 96928
rect 271694 97144 271750 97200
rect 271234 96872 271290 96928
rect 272890 97008 272946 97064
rect 274546 97008 274602 97064
rect 274270 96872 274326 96928
rect 275926 97008 275982 97064
rect 277398 97144 277454 97200
rect 276938 96872 276994 96928
rect 275282 62736 275338 62792
rect 273626 6160 273682 6216
rect 278594 96872 278650 96928
rect 279974 97008 280030 97064
rect 281170 96872 281226 96928
rect 280710 90344 280766 90400
rect 281446 96872 281502 96928
rect 282550 91160 282606 91216
rect 283010 97824 283066 97880
rect 282826 96872 282882 96928
rect 284298 98776 284354 98832
rect 284022 96872 284078 96928
rect 284850 98912 284906 98968
rect 285770 97824 285826 97880
rect 285402 3304 285458 3360
rect 286874 96872 286930 96928
rect 287978 95784 288034 95840
rect 288346 96872 288402 96928
rect 290922 99592 290978 99648
rect 289726 95920 289782 95976
rect 290738 87624 290794 87680
rect 291566 98640 291622 98696
rect 291198 95784 291254 95840
rect 292578 97416 292634 97472
rect 292394 96872 292450 96928
rect 293590 97280 293646 97336
rect 293590 87488 293646 87544
rect 293958 99456 294014 99512
rect 294970 96872 295026 96928
rect 295246 96872 295302 96928
rect 295062 90616 295118 90672
rect 295798 97416 295854 97472
rect 294970 80824 295026 80880
rect 296074 80688 296130 80744
rect 296442 86128 296498 86184
rect 299294 96872 299350 96928
rect 298282 94424 298338 94480
rect 297914 80688 297970 80744
rect 304998 97416 305054 97472
rect 302238 94560 302294 94616
rect 303710 96056 303766 96112
rect 305550 1944 305606 2000
rect 312542 97280 312598 97336
rect 311898 82048 311954 82104
rect 316682 76744 316738 76800
rect 326342 73752 326398 73808
rect 327722 79600 327778 79656
rect 326342 11872 326398 11928
rect 529938 99592 529994 99648
rect 342258 84904 342314 84960
rect 493322 98912 493378 98968
rect 351918 93336 351974 93392
rect 353298 72392 353354 72448
rect 363602 79464 363658 79520
rect 370502 90616 370558 90672
rect 367742 30912 367798 30968
rect 373998 71168 374054 71224
rect 376758 91704 376814 91760
rect 385038 75248 385094 75304
rect 391938 84768 391994 84824
rect 393318 78104 393374 78160
rect 403622 97144 403678 97200
rect 403070 76608 403126 76664
rect 409970 76472 410026 76528
rect 415398 77968 415454 78024
rect 429842 90480 429898 90536
rect 423770 83544 423826 83600
rect 440238 90344 440294 90400
rect 432510 11736 432566 11792
rect 441618 83408 441674 83464
rect 447782 77832 447838 77888
rect 450542 79328 450598 79384
rect 465078 89120 465134 89176
rect 472622 86264 472678 86320
rect 474554 4800 474610 4856
rect 489918 93200 489974 93256
rect 494058 98776 494114 98832
rect 497462 95920 497518 95976
rect 514758 71032 514814 71088
rect 517610 75112 517666 75168
rect 525798 95784 525854 95840
rect 522302 80824 522358 80880
rect 550638 99456 550694 99512
rect 532698 98640 532754 98696
rect 538218 87760 538274 87816
rect 536838 87624 536894 87680
rect 545486 11600 545542 11656
rect 553398 93064 553454 93120
rect 554778 87488 554834 87544
rect 574098 88984 574154 89040
rect 568026 3304 568082 3360
rect 575570 86128 575626 86184
rect 579618 80688 579674 80744
rect 582378 50224 582434 50280
rect 582194 3576 582250 3632
rect 580998 3440 581054 3496
rect 579618 3304 579674 3360
rect 583206 511264 583262 511320
rect 583298 484608 583354 484664
rect 583482 577224 583538 577280
rect 583390 404912 583446 404968
rect 583666 524728 583722 524784
rect 583574 471008 583630 471064
rect 583114 203496 583170 203552
rect 583482 202136 583538 202192
rect 583482 200096 583538 200152
rect 583390 152632 583446 152688
rect 583298 139304 583354 139360
rect 583206 125976 583262 126032
rect 583114 112784 583170 112840
rect 583390 102176 583446 102232
rect 583114 100952 583170 101008
rect 583022 99456 583078 99512
rect 582654 86128 582710 86184
rect 582470 19760 582526 19816
rect 582930 3576 582986 3632
rect 582654 3440 582710 3496
rect 583206 100816 583262 100872
rect 583298 94424 583354 94480
rect 583758 73208 583814 73264
rect 583666 60152 583722 60208
rect 583574 46824 583630 46880
rect 583850 32816 583906 32872
rect 583574 6840 583630 6896
<< metal3 >>
rect -960 697220 480 697460
rect 583520 697234 584960 697324
rect 583342 697174 584960 697234
rect 583342 697098 583402 697174
rect 583520 697098 584960 697174
rect 583342 697084 584960 697098
rect 583342 697038 583770 697084
rect 583710 696965 583770 697038
rect 583710 696960 583819 696965
rect 583710 696904 583758 696960
rect 583814 696904 583819 696960
rect 583710 696902 583819 696904
rect 583753 696899 583819 696902
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 583385 683906 583451 683909
rect 583520 683906 584960 683996
rect 583385 683904 584960 683906
rect 583385 683848 583390 683904
rect 583446 683848 584960 683904
rect 583385 683846 584960 683848
rect 583385 683843 583451 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3509 671258 3575 671261
rect -960 671256 3575 671258
rect -960 671200 3514 671256
rect 3570 671200 3575 671256
rect -960 671198 3575 671200
rect -960 671108 480 671198
rect 3509 671195 3575 671198
rect 582465 670714 582531 670717
rect 583520 670714 584960 670804
rect 582465 670712 584960 670714
rect 582465 670656 582470 670712
rect 582526 670656 584960 670712
rect 582465 670654 584960 670656
rect 582465 670651 582531 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3417 658202 3483 658205
rect -960 658200 3483 658202
rect -960 658144 3422 658200
rect 3478 658144 3483 658200
rect -960 658142 3483 658144
rect -960 658052 480 658142
rect 3417 658139 3483 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 582557 644058 582623 644061
rect 583520 644058 584960 644148
rect 582557 644056 584960 644058
rect 582557 644000 582562 644056
rect 582618 644000 584960 644056
rect 582557 643998 584960 644000
rect 582557 643995 582623 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 3417 632090 3483 632093
rect -960 632088 3483 632090
rect -960 632032 3422 632088
rect 3478 632032 3483 632088
rect -960 632030 3483 632032
rect -960 631940 480 632030
rect 3417 632027 3483 632030
rect 582649 630866 582715 630869
rect 583520 630866 584960 630956
rect 582649 630864 584960 630866
rect 582649 630808 582654 630864
rect 582710 630808 584960 630864
rect 582649 630806 584960 630808
rect 582649 630803 582715 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3141 619170 3207 619173
rect -960 619168 3207 619170
rect -960 619112 3146 619168
rect 3202 619112 3207 619168
rect -960 619110 3207 619112
rect -960 619020 480 619110
rect 3141 619107 3207 619110
rect 582741 617538 582807 617541
rect 583520 617538 584960 617628
rect 582741 617536 584960 617538
rect 582741 617480 582746 617536
rect 582802 617480 584960 617536
rect 582741 617478 584960 617480
rect 582741 617475 582807 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3233 606114 3299 606117
rect -960 606112 3299 606114
rect -960 606056 3238 606112
rect 3294 606056 3299 606112
rect -960 606054 3299 606056
rect -960 605964 480 606054
rect 3233 606051 3299 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 582833 591018 582899 591021
rect 583520 591018 584960 591108
rect 582833 591016 584960 591018
rect 582833 590960 582838 591016
rect 582894 590960 584960 591016
rect 582833 590958 584960 590960
rect 582833 590955 582899 590958
rect 583520 590868 584960 590958
rect -960 580002 480 580092
rect 3325 580002 3391 580005
rect -960 580000 3391 580002
rect -960 579944 3330 580000
rect 3386 579944 3391 580000
rect -960 579942 3391 579944
rect -960 579852 480 579942
rect 3325 579939 3391 579942
rect 583520 577690 584960 577780
rect 583342 577630 584960 577690
rect 583342 577554 583402 577630
rect 583520 577554 584960 577630
rect 583342 577540 584960 577554
rect 583342 577494 583586 577540
rect 583526 577285 583586 577494
rect 583477 577280 583586 577285
rect 583477 577224 583482 577280
rect 583538 577224 583586 577280
rect 583477 577222 583586 577224
rect 583477 577219 583543 577222
rect -960 566946 480 567036
rect 3417 566946 3483 566949
rect -960 566944 3483 566946
rect -960 566888 3422 566944
rect 3478 566888 3483 566944
rect -960 566886 3483 566888
rect -960 566796 480 566886
rect 3417 566883 3483 566886
rect 583017 564362 583083 564365
rect 583520 564362 584960 564452
rect 583017 564360 584960 564362
rect 583017 564304 583022 564360
rect 583078 564304 584960 564360
rect 583017 564302 584960 564304
rect 583017 564299 583083 564302
rect 583520 564212 584960 564302
rect -960 553890 480 553980
rect 3417 553890 3483 553893
rect -960 553888 3483 553890
rect -960 553832 3422 553888
rect 3478 553832 3483 553888
rect -960 553830 3483 553832
rect -960 553740 480 553830
rect 3417 553827 3483 553830
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 583109 537842 583175 537845
rect 583520 537842 584960 537932
rect 583109 537840 584960 537842
rect 583109 537784 583114 537840
rect 583170 537784 584960 537840
rect 583109 537782 584960 537784
rect 583109 537779 583175 537782
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect 3417 527914 3483 527917
rect -960 527912 3483 527914
rect -960 527856 3422 527912
rect 3478 527856 3483 527912
rect -960 527854 3483 527856
rect -960 527764 480 527854
rect 3417 527851 3483 527854
rect 583661 524786 583727 524789
rect 583526 524784 583727 524786
rect 583526 524728 583666 524784
rect 583722 524728 583727 524784
rect 583526 524726 583727 524728
rect 583526 524650 583586 524726
rect 583661 524723 583727 524726
rect 583342 524604 583586 524650
rect 583342 524590 584960 524604
rect 583342 524514 583402 524590
rect 583520 524514 584960 524590
rect 583342 524454 584960 524514
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 3417 514858 3483 514861
rect -960 514856 3483 514858
rect -960 514800 3422 514856
rect 3478 514800 3483 514856
rect -960 514798 3483 514800
rect -960 514708 480 514798
rect 3417 514795 3483 514798
rect 583201 511322 583267 511325
rect 583520 511322 584960 511412
rect 583201 511320 584960 511322
rect 583201 511264 583206 511320
rect 583262 511264 584960 511320
rect 583201 511262 584960 511264
rect 583201 511259 583267 511262
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect 3417 501802 3483 501805
rect -960 501800 3483 501802
rect -960 501744 3422 501800
rect 3478 501744 3483 501800
rect -960 501742 3483 501744
rect -960 501652 480 501742
rect 3417 501739 3483 501742
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 583293 484666 583359 484669
rect 583520 484666 584960 484756
rect 583293 484664 584960 484666
rect 583293 484608 583298 484664
rect 583354 484608 584960 484664
rect 583293 484606 584960 484608
rect 583293 484603 583359 484606
rect 583520 484516 584960 484606
rect -960 475690 480 475780
rect 3049 475690 3115 475693
rect -960 475688 3115 475690
rect -960 475632 3054 475688
rect 3110 475632 3115 475688
rect -960 475630 3115 475632
rect -960 475540 480 475630
rect 3049 475627 3115 475630
rect 583520 471474 584960 471564
rect 583342 471414 584960 471474
rect 583342 471338 583402 471414
rect 583520 471338 584960 471414
rect 583342 471324 584960 471338
rect 583342 471278 583586 471324
rect 583526 471069 583586 471278
rect 583526 471064 583635 471069
rect 583526 471008 583574 471064
rect 583630 471008 583635 471064
rect 583526 471006 583635 471008
rect 583569 471003 583635 471006
rect -960 462634 480 462724
rect 3509 462634 3575 462637
rect -960 462632 3575 462634
rect -960 462576 3514 462632
rect 3570 462576 3575 462632
rect -960 462574 3575 462576
rect -960 462484 480 462574
rect 3509 462571 3575 462574
rect 580165 458146 580231 458149
rect 583520 458146 584960 458236
rect 580165 458144 584960 458146
rect 580165 458088 580170 458144
rect 580226 458088 584960 458144
rect 580165 458086 584960 458088
rect 580165 458083 580231 458086
rect 583520 457996 584960 458086
rect -960 449578 480 449668
rect 3141 449578 3207 449581
rect -960 449576 3207 449578
rect -960 449520 3146 449576
rect 3202 449520 3207 449576
rect -960 449518 3207 449520
rect -960 449428 480 449518
rect 3141 449515 3207 449518
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 580165 431626 580231 431629
rect 583520 431626 584960 431716
rect 580165 431624 584960 431626
rect 580165 431568 580170 431624
rect 580226 431568 584960 431624
rect 580165 431566 584960 431568
rect 580165 431563 580231 431566
rect 583520 431476 584960 431566
rect -960 423602 480 423692
rect 3509 423602 3575 423605
rect -960 423600 3575 423602
rect -960 423544 3514 423600
rect 3570 423544 3575 423600
rect -960 423542 3575 423544
rect -960 423452 480 423542
rect 3509 423539 3575 423542
rect 580165 418298 580231 418301
rect 583520 418298 584960 418388
rect 580165 418296 584960 418298
rect 580165 418240 580170 418296
rect 580226 418240 584960 418296
rect 580165 418238 584960 418240
rect 580165 418235 580231 418238
rect 583520 418148 584960 418238
rect -960 410546 480 410636
rect 2865 410546 2931 410549
rect -960 410544 2931 410546
rect -960 410488 2870 410544
rect 2926 410488 2931 410544
rect -960 410486 2931 410488
rect -960 410396 480 410486
rect 2865 410483 2931 410486
rect 583385 404970 583451 404973
rect 583520 404970 584960 405060
rect 583385 404968 584960 404970
rect 583385 404912 583390 404968
rect 583446 404912 584960 404968
rect 583385 404910 584960 404912
rect 583385 404907 583451 404910
rect 583520 404820 584960 404910
rect -960 397490 480 397580
rect 3509 397490 3575 397493
rect -960 397488 3575 397490
rect -960 397432 3514 397488
rect 3570 397432 3575 397488
rect -960 397430 3575 397432
rect -960 397340 480 397430
rect 3509 397427 3575 397430
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 580901 378450 580967 378453
rect 583520 378450 584960 378540
rect 580901 378448 584960 378450
rect 580901 378392 580906 378448
rect 580962 378392 584960 378448
rect 580901 378390 584960 378392
rect 580901 378387 580967 378390
rect 583520 378300 584960 378390
rect -960 371378 480 371468
rect 3509 371378 3575 371381
rect -960 371376 3575 371378
rect -960 371320 3514 371376
rect 3570 371320 3575 371376
rect -960 371318 3575 371320
rect -960 371228 480 371318
rect 3509 371315 3575 371318
rect 580165 365122 580231 365125
rect 583520 365122 584960 365212
rect 580165 365120 584960 365122
rect 580165 365064 580170 365120
rect 580226 365064 584960 365120
rect 580165 365062 584960 365064
rect 580165 365059 580231 365062
rect 583520 364972 584960 365062
rect -960 358458 480 358548
rect 3141 358458 3207 358461
rect -960 358456 3207 358458
rect -960 358400 3146 358456
rect 3202 358400 3207 358456
rect -960 358398 3207 358400
rect -960 358308 480 358398
rect 3141 358395 3207 358398
rect 579889 351930 579955 351933
rect 583520 351930 584960 352020
rect 579889 351928 584960 351930
rect 579889 351872 579894 351928
rect 579950 351872 584960 351928
rect 579889 351870 584960 351872
rect 579889 351867 579955 351870
rect 583520 351780 584960 351870
rect -960 345402 480 345492
rect 3325 345402 3391 345405
rect -960 345400 3391 345402
rect -960 345344 3330 345400
rect 3386 345344 3391 345400
rect -960 345342 3391 345344
rect -960 345252 480 345342
rect 3325 345339 3391 345342
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 580165 325274 580231 325277
rect 583520 325274 584960 325364
rect 580165 325272 584960 325274
rect 580165 325216 580170 325272
rect 580226 325216 584960 325272
rect 580165 325214 584960 325216
rect 580165 325211 580231 325214
rect 583520 325124 584960 325214
rect -960 319290 480 319380
rect 3325 319290 3391 319293
rect -960 319288 3391 319290
rect -960 319232 3330 319288
rect 3386 319232 3391 319288
rect -960 319230 3391 319232
rect -960 319140 480 319230
rect 3325 319227 3391 319230
rect 580165 312082 580231 312085
rect 583520 312082 584960 312172
rect 580165 312080 584960 312082
rect 580165 312024 580170 312080
rect 580226 312024 584960 312080
rect 580165 312022 584960 312024
rect 580165 312019 580231 312022
rect 583520 311932 584960 312022
rect -960 306234 480 306324
rect 3509 306234 3575 306237
rect -960 306232 3575 306234
rect -960 306176 3514 306232
rect 3570 306176 3575 306232
rect -960 306174 3575 306176
rect -960 306084 480 306174
rect 3509 306171 3575 306174
rect 580901 298754 580967 298757
rect 583520 298754 584960 298844
rect 580901 298752 584960 298754
rect 580901 298696 580906 298752
rect 580962 298696 584960 298752
rect 580901 298694 584960 298696
rect 580901 298691 580967 298694
rect 583520 298604 584960 298694
rect -960 293178 480 293268
rect 3509 293178 3575 293181
rect -960 293176 3575 293178
rect -960 293120 3514 293176
rect 3570 293120 3575 293176
rect -960 293118 3575 293120
rect -960 293028 480 293118
rect 3509 293115 3575 293118
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 580165 272234 580231 272237
rect 583520 272234 584960 272324
rect 580165 272232 584960 272234
rect 580165 272176 580170 272232
rect 580226 272176 584960 272232
rect 580165 272174 584960 272176
rect 580165 272171 580231 272174
rect 583520 272084 584960 272174
rect -960 267202 480 267292
rect 3049 267202 3115 267205
rect -960 267200 3115 267202
rect -960 267144 3054 267200
rect 3110 267144 3115 267200
rect -960 267142 3115 267144
rect -960 267052 480 267142
rect 3049 267139 3115 267142
rect 580165 258906 580231 258909
rect 583520 258906 584960 258996
rect 580165 258904 584960 258906
rect 580165 258848 580170 258904
rect 580226 258848 584960 258904
rect 580165 258846 584960 258848
rect 580165 258843 580231 258846
rect 583520 258756 584960 258846
rect -960 254146 480 254236
rect 3509 254146 3575 254149
rect -960 254144 3575 254146
rect -960 254088 3514 254144
rect 3570 254088 3575 254144
rect -960 254086 3575 254088
rect -960 253996 480 254086
rect 3509 254083 3575 254086
rect 582925 245578 582991 245581
rect 583520 245578 584960 245668
rect 582925 245576 584960 245578
rect 582925 245520 582930 245576
rect 582986 245520 584960 245576
rect 582925 245518 584960 245520
rect 582925 245515 582991 245518
rect 583520 245428 584960 245518
rect -960 241090 480 241180
rect 3049 241090 3115 241093
rect -960 241088 3115 241090
rect -960 241032 3054 241088
rect 3110 241032 3115 241088
rect -960 241030 3115 241032
rect -960 240940 480 241030
rect 3049 241027 3115 241030
rect 580165 232386 580231 232389
rect 583520 232386 584960 232476
rect 580165 232384 584960 232386
rect 580165 232328 580170 232384
rect 580226 232328 584960 232384
rect 580165 232326 584960 232328
rect 580165 232323 580231 232326
rect 583520 232236 584960 232326
rect -960 227884 480 228124
rect 580165 219058 580231 219061
rect 583520 219058 584960 219148
rect 580165 219056 584960 219058
rect 580165 219000 580170 219056
rect 580226 219000 584960 219056
rect 580165 218998 584960 219000
rect 580165 218995 580231 218998
rect 583520 218908 584960 218998
rect -960 214978 480 215068
rect 3141 214978 3207 214981
rect -960 214976 3207 214978
rect -960 214920 3146 214976
rect 3202 214920 3207 214976
rect -960 214918 3207 214920
rect -960 214828 480 214918
rect 3141 214915 3207 214918
rect 242525 207634 242591 207637
rect 305637 207634 305703 207637
rect 242525 207632 305703 207634
rect 242525 207576 242530 207632
rect 242586 207576 305642 207632
rect 305698 207576 305703 207632
rect 242525 207574 305703 207576
rect 242525 207571 242591 207574
rect 305637 207571 305703 207574
rect 237189 206274 237255 206277
rect 582465 206274 582531 206277
rect 237189 206272 582531 206274
rect 237189 206216 237194 206272
rect 237250 206216 582470 206272
rect 582526 206216 582531 206272
rect 237189 206214 582531 206216
rect 237189 206211 237255 206214
rect 582465 206211 582531 206214
rect 580165 205730 580231 205733
rect 583520 205730 584960 205820
rect 580165 205728 584960 205730
rect 580165 205672 580170 205728
rect 580226 205672 584960 205728
rect 580165 205670 584960 205672
rect 580165 205667 580231 205670
rect 583520 205580 584960 205670
rect 73061 205186 73127 205189
rect 258625 205186 258691 205189
rect 73061 205184 258691 205186
rect 73061 205128 73066 205184
rect 73122 205128 258630 205184
rect 258686 205128 258691 205184
rect 73061 205126 258691 205128
rect 73061 205123 73127 205126
rect 258625 205123 258691 205126
rect 235993 205050 236059 205053
rect 582649 205050 582715 205053
rect 235993 205048 582715 205050
rect 235993 204992 235998 205048
rect 236054 204992 582654 205048
rect 582710 204992 582715 205048
rect 235993 204990 582715 204992
rect 235993 204987 236059 204990
rect 582649 204987 582715 204990
rect 231669 204914 231735 204917
rect 583017 204914 583083 204917
rect 231669 204912 583083 204914
rect 231669 204856 231674 204912
rect 231730 204856 583022 204912
rect 583078 204856 583083 204912
rect 231669 204854 583083 204856
rect 231669 204851 231735 204854
rect 583017 204851 583083 204854
rect 255957 203826 256023 203829
rect 268193 203826 268259 203829
rect 255957 203824 268259 203826
rect 255957 203768 255962 203824
rect 256018 203768 268198 203824
rect 268254 203768 268259 203824
rect 255957 203766 268259 203768
rect 255957 203763 256023 203766
rect 268193 203763 268259 203766
rect 106181 203690 106247 203693
rect 255313 203690 255379 203693
rect 106181 203688 255379 203690
rect 106181 203632 106186 203688
rect 106242 203632 255318 203688
rect 255374 203632 255379 203688
rect 106181 203630 255379 203632
rect 106181 203627 106247 203630
rect 255313 203627 255379 203630
rect 230381 203554 230447 203557
rect 583109 203554 583175 203557
rect 230381 203552 583175 203554
rect 230381 203496 230386 203552
rect 230442 203496 583114 203552
rect 583170 203496 583175 203552
rect 230381 203494 583175 203496
rect 230381 203491 230447 203494
rect 583109 203491 583175 203494
rect 242985 202874 243051 202877
rect 244917 202874 244983 202877
rect 242985 202872 244983 202874
rect 242985 202816 242990 202872
rect 243046 202816 244922 202872
rect 244978 202816 244983 202872
rect 242985 202814 244983 202816
rect 242985 202811 243051 202814
rect 244917 202811 244983 202814
rect 252645 202874 252711 202877
rect 255129 202874 255195 202877
rect 252645 202872 255195 202874
rect 252645 202816 252650 202872
rect 252706 202816 255134 202872
rect 255190 202816 255195 202872
rect 252645 202814 255195 202816
rect 252645 202811 252711 202814
rect 255129 202811 255195 202814
rect 259177 202874 259243 202877
rect 260373 202874 260439 202877
rect 259177 202872 260439 202874
rect 259177 202816 259182 202872
rect 259238 202816 260378 202872
rect 260434 202816 260439 202872
rect 259177 202814 260439 202816
rect 259177 202811 259243 202814
rect 260373 202811 260439 202814
rect 244733 202738 244799 202741
rect 246021 202738 246087 202741
rect 244733 202736 246087 202738
rect 244733 202680 244738 202736
rect 244794 202680 246026 202736
rect 246082 202680 246087 202736
rect 244733 202678 246087 202680
rect 244733 202675 244799 202678
rect 246021 202675 246087 202678
rect 250621 202602 250687 202605
rect 253381 202602 253447 202605
rect 250621 202600 253447 202602
rect 250621 202544 250626 202600
rect 250682 202544 253386 202600
rect 253442 202544 253447 202600
rect 250621 202542 253447 202544
rect 250621 202539 250687 202542
rect 253381 202539 253447 202542
rect 222377 202194 222443 202197
rect 583477 202194 583543 202197
rect 222377 202192 583543 202194
rect 222377 202136 222382 202192
rect 222438 202136 583482 202192
rect 583538 202136 583543 202192
rect 222377 202134 583543 202136
rect 222377 202131 222443 202134
rect 583477 202131 583543 202134
rect -960 201922 480 202012
rect 3233 201922 3299 201925
rect -960 201920 3299 201922
rect -960 201864 3238 201920
rect 3294 201864 3299 201920
rect -960 201862 3299 201864
rect -960 201772 480 201862
rect 3233 201859 3299 201862
rect 255313 201922 255379 201925
rect 257705 201922 257771 201925
rect 255313 201920 257771 201922
rect 255313 201864 255318 201920
rect 255374 201864 257710 201920
rect 257766 201864 257771 201920
rect 255313 201862 257771 201864
rect 255313 201859 255379 201862
rect 257705 201859 257771 201862
rect 200389 200154 200455 200157
rect 583477 200154 583543 200157
rect 200389 200152 583543 200154
rect 200389 200096 200394 200152
rect 200450 200096 583482 200152
rect 583538 200096 583543 200152
rect 200389 200094 583543 200096
rect 200389 200091 200455 200094
rect 583477 200091 583543 200094
rect 199837 199610 199903 199613
rect 204069 199610 204135 199613
rect 199837 199608 204135 199610
rect 199837 199552 199842 199608
rect 199898 199552 204074 199608
rect 204130 199552 204135 199608
rect 199837 199550 204135 199552
rect 199837 199547 199903 199550
rect 204069 199547 204135 199550
rect 207657 199610 207723 199613
rect 211245 199610 211311 199613
rect 207657 199608 211311 199610
rect 207657 199552 207662 199608
rect 207718 199552 211250 199608
rect 211306 199552 211311 199608
rect 207657 199550 211311 199552
rect 207657 199547 207723 199550
rect 211245 199547 211311 199550
rect 246205 199610 246271 199613
rect 246481 199610 246547 199613
rect 246205 199608 246547 199610
rect 246205 199552 246210 199608
rect 246266 199552 246486 199608
rect 246542 199552 246547 199608
rect 246205 199550 246547 199552
rect 246205 199547 246271 199550
rect 246481 199547 246547 199550
rect 197997 199338 198063 199341
rect 197997 199336 200100 199338
rect 197997 199280 198002 199336
rect 198058 199280 200100 199336
rect 197997 199278 200100 199280
rect 197997 199275 198063 199278
rect 197997 198250 198063 198253
rect 197997 198248 200100 198250
rect 197997 198192 198002 198248
rect 198058 198192 200100 198248
rect 197997 198190 200100 198192
rect 197997 198187 198063 198190
rect 198641 197162 198707 197165
rect 198641 197160 200100 197162
rect 198641 197104 198646 197160
rect 198702 197104 200100 197160
rect 198641 197102 200100 197104
rect 198641 197099 198707 197102
rect 197997 196074 198063 196077
rect 197997 196072 200100 196074
rect 197997 196016 198002 196072
rect 198058 196016 200100 196072
rect 197997 196014 200100 196016
rect 197997 196011 198063 196014
rect 198089 194986 198155 194989
rect 198089 194984 200100 194986
rect 198089 194928 198094 194984
rect 198150 194928 200100 194984
rect 198089 194926 200100 194928
rect 198089 194923 198155 194926
rect 197721 193898 197787 193901
rect 197721 193896 200100 193898
rect 197721 193840 197726 193896
rect 197782 193840 200100 193896
rect 197721 193838 200100 193840
rect 197721 193835 197787 193838
rect 197629 192810 197695 192813
rect 197629 192808 200100 192810
rect 197629 192752 197634 192808
rect 197690 192752 200100 192808
rect 197629 192750 200100 192752
rect 197629 192747 197695 192750
rect 580165 192538 580231 192541
rect 583520 192538 584960 192628
rect 580165 192536 584960 192538
rect 580165 192480 580170 192536
rect 580226 192480 584960 192536
rect 580165 192478 584960 192480
rect 580165 192475 580231 192478
rect 583520 192388 584960 192478
rect 198089 191722 198155 191725
rect 198089 191720 200100 191722
rect 198089 191664 198094 191720
rect 198150 191664 200100 191720
rect 198089 191662 200100 191664
rect 198089 191659 198155 191662
rect 197353 190634 197419 190637
rect 197353 190632 200100 190634
rect 197353 190576 197358 190632
rect 197414 190576 200100 190632
rect 197353 190574 200100 190576
rect 197353 190571 197419 190574
rect 197905 189546 197971 189549
rect 197905 189544 200100 189546
rect 197905 189488 197910 189544
rect 197966 189488 200100 189544
rect 197905 189486 200100 189488
rect 197905 189483 197971 189486
rect 169894 189274 169954 189448
rect 172421 189274 172487 189277
rect 169894 189272 172487 189274
rect 169894 189216 172426 189272
rect 172482 189216 172487 189272
rect 169894 189214 172487 189216
rect 172421 189211 172487 189214
rect -960 188866 480 188956
rect 3509 188866 3575 188869
rect -960 188864 3575 188866
rect -960 188808 3514 188864
rect 3570 188808 3575 188864
rect -960 188806 3575 188808
rect -960 188716 480 188806
rect 3509 188803 3575 188806
rect 197353 188458 197419 188461
rect 197353 188456 200100 188458
rect 197353 188400 197358 188456
rect 197414 188400 200100 188456
rect 197353 188398 200100 188400
rect 197353 188395 197419 188398
rect 169894 187778 169954 188360
rect 171777 187778 171843 187781
rect 169894 187776 171843 187778
rect 169894 187720 171782 187776
rect 171838 187720 171843 187776
rect 169894 187718 171843 187720
rect 171777 187715 171843 187718
rect 197537 187370 197603 187373
rect 197537 187368 200100 187370
rect 197537 187312 197542 187368
rect 197598 187312 200100 187368
rect 197537 187310 200100 187312
rect 197537 187307 197603 187310
rect 169894 186826 169954 187136
rect 172421 186826 172487 186829
rect 169894 186824 172487 186826
rect 169894 186768 172426 186824
rect 172482 186768 172487 186824
rect 169894 186766 172487 186768
rect 172421 186763 172487 186766
rect 197629 186282 197695 186285
rect 197629 186280 200100 186282
rect 197629 186224 197634 186280
rect 197690 186224 200100 186280
rect 197629 186222 200100 186224
rect 197629 186219 197695 186222
rect 169894 185466 169954 186048
rect 171777 185466 171843 185469
rect 169894 185464 171843 185466
rect 169894 185408 171782 185464
rect 171838 185408 171843 185464
rect 169894 185406 171843 185408
rect 171777 185403 171843 185406
rect 197353 185058 197419 185061
rect 197353 185056 200100 185058
rect 197353 185000 197358 185056
rect 197414 185000 200100 185056
rect 197353 184998 200100 185000
rect 197353 184995 197419 184998
rect 169894 184242 169954 184824
rect 171685 184242 171751 184245
rect 169894 184240 171751 184242
rect 169894 184184 171690 184240
rect 171746 184184 171751 184240
rect 169894 184182 171751 184184
rect 171685 184179 171751 184182
rect 198365 183970 198431 183973
rect 198365 183968 200100 183970
rect 198365 183912 198370 183968
rect 198426 183912 200100 183968
rect 198365 183910 200100 183912
rect 198365 183907 198431 183910
rect 169894 183698 169954 183736
rect 172421 183698 172487 183701
rect 169894 183696 172487 183698
rect 169894 183640 172426 183696
rect 172482 183640 172487 183696
rect 169894 183638 172487 183640
rect 172421 183635 172487 183638
rect 197721 182882 197787 182885
rect 197721 182880 200100 182882
rect 197721 182824 197726 182880
rect 197782 182824 200100 182880
rect 197721 182822 200100 182824
rect 197721 182819 197787 182822
rect 169894 182474 169954 182512
rect 172421 182474 172487 182477
rect 169894 182472 172487 182474
rect 169894 182416 172426 182472
rect 172482 182416 172487 182472
rect 169894 182414 172487 182416
rect 172421 182411 172487 182414
rect 197353 181794 197419 181797
rect 197353 181792 200100 181794
rect 197353 181736 197358 181792
rect 197414 181736 200100 181792
rect 197353 181734 200100 181736
rect 197353 181731 197419 181734
rect 169894 181114 169954 181424
rect 172421 181114 172487 181117
rect 169894 181112 172487 181114
rect 169894 181056 172426 181112
rect 172482 181056 172487 181112
rect 169894 181054 172487 181056
rect 172421 181051 172487 181054
rect 197353 180706 197419 180709
rect 197353 180704 200100 180706
rect 197353 180648 197358 180704
rect 197414 180648 200100 180704
rect 197353 180646 200100 180648
rect 197353 180643 197419 180646
rect 169894 179890 169954 180200
rect 172053 179890 172119 179893
rect 169894 179888 172119 179890
rect 169894 179832 172058 179888
rect 172114 179832 172119 179888
rect 169894 179830 172119 179832
rect 172053 179827 172119 179830
rect 198089 179618 198155 179621
rect 198089 179616 200100 179618
rect 198089 179560 198094 179616
rect 198150 179560 200100 179616
rect 198089 179558 200100 179560
rect 198089 179555 198155 179558
rect 580257 179210 580323 179213
rect 583520 179210 584960 179300
rect 580257 179208 584960 179210
rect 580257 179152 580262 179208
rect 580318 179152 584960 179208
rect 580257 179150 584960 179152
rect 580257 179147 580323 179150
rect 169894 178666 169954 179112
rect 583520 179060 584960 179150
rect 172145 178666 172211 178669
rect 169894 178664 172211 178666
rect 169894 178608 172150 178664
rect 172206 178608 172211 178664
rect 169894 178606 172211 178608
rect 172145 178603 172211 178606
rect 197905 178530 197971 178533
rect 197905 178528 200100 178530
rect 197905 178472 197910 178528
rect 197966 178472 200100 178528
rect 197905 178470 200100 178472
rect 197905 178467 197971 178470
rect 169894 177306 169954 177888
rect 197813 177442 197879 177445
rect 197813 177440 200100 177442
rect 197813 177384 197818 177440
rect 197874 177384 200100 177440
rect 197813 177382 200100 177384
rect 197813 177379 197879 177382
rect 172237 177306 172303 177309
rect 169894 177304 172303 177306
rect 169894 177248 172242 177304
rect 172298 177248 172303 177304
rect 169894 177246 172303 177248
rect 172237 177243 172303 177246
rect 169894 176762 169954 176800
rect 172421 176762 172487 176765
rect 169894 176760 172487 176762
rect 169894 176704 172426 176760
rect 172482 176704 172487 176760
rect 169894 176702 172487 176704
rect 172421 176699 172487 176702
rect 197353 176354 197419 176357
rect 197353 176352 200100 176354
rect 197353 176296 197358 176352
rect 197414 176296 200100 176352
rect 197353 176294 200100 176296
rect 197353 176291 197419 176294
rect -960 175796 480 176036
rect 169894 175402 169954 175576
rect 172421 175402 172487 175405
rect 169894 175400 172487 175402
rect 169894 175344 172426 175400
rect 172482 175344 172487 175400
rect 169894 175342 172487 175344
rect 172421 175339 172487 175342
rect 198549 175266 198615 175269
rect 198549 175264 200100 175266
rect 198549 175208 198554 175264
rect 198610 175208 200100 175264
rect 198549 175206 200100 175208
rect 198549 175203 198615 175206
rect 169894 174178 169954 174488
rect 171961 174178 172027 174181
rect 169894 174176 172027 174178
rect 169894 174120 171966 174176
rect 172022 174120 172027 174176
rect 169894 174118 172027 174120
rect 171961 174115 172027 174118
rect 197353 174178 197419 174181
rect 197353 174176 200100 174178
rect 197353 174120 197358 174176
rect 197414 174120 200100 174176
rect 197353 174118 200100 174120
rect 197353 174115 197419 174118
rect 170397 173294 170463 173297
rect 169924 173292 170463 173294
rect 169924 173236 170402 173292
rect 170458 173236 170463 173292
rect 169924 173234 170463 173236
rect 170397 173231 170463 173234
rect 198457 173090 198523 173093
rect 198457 173088 200100 173090
rect 198457 173032 198462 173088
rect 198518 173032 200100 173088
rect 198457 173030 200100 173032
rect 198457 173027 198523 173030
rect 169894 171730 169954 172176
rect 198733 172002 198799 172005
rect 198733 172000 200100 172002
rect 198733 171944 198738 172000
rect 198794 171944 200100 172000
rect 198733 171942 200100 171944
rect 198733 171939 198799 171942
rect 172237 171730 172303 171733
rect 169894 171728 172303 171730
rect 169894 171672 172242 171728
rect 172298 171672 172303 171728
rect 169894 171670 172303 171672
rect 172237 171667 172303 171670
rect 169894 170370 169954 170952
rect 197721 170778 197787 170781
rect 197721 170776 200100 170778
rect 197721 170720 197726 170776
rect 197782 170720 200100 170776
rect 197721 170718 200100 170720
rect 197721 170715 197787 170718
rect 172237 170370 172303 170373
rect 169894 170368 172303 170370
rect 169894 170312 172242 170368
rect 172298 170312 172303 170368
rect 169894 170310 172303 170312
rect 172237 170307 172303 170310
rect 169894 169826 169954 169864
rect 171777 169826 171843 169829
rect 169894 169824 171843 169826
rect 169894 169768 171782 169824
rect 171838 169768 171843 169824
rect 169894 169766 171843 169768
rect 171777 169763 171843 169766
rect 197445 169690 197511 169693
rect 197445 169688 200100 169690
rect 197445 169632 197450 169688
rect 197506 169632 200100 169688
rect 197445 169630 200100 169632
rect 197445 169627 197511 169630
rect 169894 168602 169954 168640
rect 172421 168602 172487 168605
rect 169894 168600 172487 168602
rect 169894 168544 172426 168600
rect 172482 168544 172487 168600
rect 169894 168542 172487 168544
rect 172421 168539 172487 168542
rect 197721 168602 197787 168605
rect 197721 168600 200100 168602
rect 197721 168544 197726 168600
rect 197782 168544 200100 168600
rect 197721 168542 200100 168544
rect 197721 168539 197787 168542
rect 169894 167378 169954 167552
rect 197905 167514 197971 167517
rect 197905 167512 200100 167514
rect 197905 167456 197910 167512
rect 197966 167456 200100 167512
rect 197905 167454 200100 167456
rect 197905 167451 197971 167454
rect 172421 167378 172487 167381
rect 169894 167376 172487 167378
rect 169894 167320 172426 167376
rect 172482 167320 172487 167376
rect 169894 167318 172487 167320
rect 172421 167315 172487 167318
rect 197353 166426 197419 166429
rect 197353 166424 200100 166426
rect 197353 166368 197358 166424
rect 197414 166368 200100 166424
rect 197353 166366 200100 166368
rect 197353 166363 197419 166366
rect 169894 166018 169954 166328
rect 172421 166018 172487 166021
rect 169894 166016 172487 166018
rect 169894 165960 172426 166016
rect 172482 165960 172487 166016
rect 169894 165958 172487 165960
rect 172421 165955 172487 165958
rect 582373 165882 582439 165885
rect 583520 165882 584960 165972
rect 582373 165880 584960 165882
rect 582373 165824 582378 165880
rect 582434 165824 584960 165880
rect 582373 165822 584960 165824
rect 582373 165819 582439 165822
rect 583520 165732 584960 165822
rect 197629 165338 197695 165341
rect 197629 165336 200100 165338
rect 197629 165280 197634 165336
rect 197690 165280 200100 165336
rect 197629 165278 200100 165280
rect 197629 165275 197695 165278
rect 169894 164794 169954 165240
rect 171133 164794 171199 164797
rect 169894 164792 171199 164794
rect 169894 164736 171138 164792
rect 171194 164736 171199 164792
rect 169894 164734 171199 164736
rect 171133 164731 171199 164734
rect 197353 164250 197419 164253
rect 197353 164248 200100 164250
rect 197353 164192 197358 164248
rect 197414 164192 200100 164248
rect 197353 164190 200100 164192
rect 197353 164187 197419 164190
rect 169894 163434 169954 164016
rect 171685 163434 171751 163437
rect 169894 163432 171751 163434
rect 169894 163376 171690 163432
rect 171746 163376 171751 163432
rect 169894 163374 171751 163376
rect 171685 163371 171751 163374
rect 197629 163162 197695 163165
rect 197629 163160 200100 163162
rect 197629 163104 197634 163160
rect 197690 163104 200100 163160
rect 197629 163102 200100 163104
rect 197629 163099 197695 163102
rect 171869 163026 171935 163029
rect 169894 163024 171935 163026
rect -960 162890 480 162980
rect 169894 162968 171874 163024
rect 171930 162968 171935 163024
rect 169894 162966 171935 162968
rect 169894 162928 169954 162966
rect 171869 162963 171935 162966
rect 3233 162890 3299 162893
rect -960 162888 3299 162890
rect -960 162832 3238 162888
rect 3294 162832 3299 162888
rect -960 162830 3299 162832
rect -960 162740 480 162830
rect 3233 162827 3299 162830
rect 197353 162074 197419 162077
rect 197353 162072 200100 162074
rect 197353 162016 197358 162072
rect 197414 162016 200100 162072
rect 197353 162014 200100 162016
rect 197353 162011 197419 162014
rect 169342 161533 169402 161704
rect 169293 161528 169402 161533
rect 169293 161472 169298 161528
rect 169354 161472 169402 161528
rect 169293 161470 169402 161472
rect 169293 161467 169359 161470
rect 198457 160986 198523 160989
rect 198457 160984 200100 160986
rect 198457 160928 198462 160984
rect 198518 160928 200100 160984
rect 198457 160926 200100 160928
rect 198457 160923 198523 160926
rect 169894 160442 169954 160616
rect 171869 160442 171935 160445
rect 169894 160440 171935 160442
rect 169894 160384 171874 160440
rect 171930 160384 171935 160440
rect 169894 160382 171935 160384
rect 171869 160379 171935 160382
rect 197537 159898 197603 159901
rect 197537 159896 200100 159898
rect 197537 159840 197542 159896
rect 197598 159840 200100 159896
rect 197537 159838 200100 159840
rect 197537 159835 197603 159838
rect 197905 158810 197971 158813
rect 197905 158808 200100 158810
rect 197905 158752 197910 158808
rect 197966 158752 200100 158808
rect 197905 158750 200100 158752
rect 197905 158747 197971 158750
rect 197353 157722 197419 157725
rect 197353 157720 200100 157722
rect 197353 157664 197358 157720
rect 197414 157664 200100 157720
rect 197353 157662 200100 157664
rect 197353 157659 197419 157662
rect 198457 156498 198523 156501
rect 198457 156496 200100 156498
rect 198457 156440 198462 156496
rect 198518 156440 200100 156496
rect 198457 156438 200100 156440
rect 198457 156435 198523 156438
rect 197721 155410 197787 155413
rect 197721 155408 200100 155410
rect 197721 155352 197726 155408
rect 197782 155352 200100 155408
rect 197721 155350 200100 155352
rect 197721 155347 197787 155350
rect 197353 154322 197419 154325
rect 197353 154320 200100 154322
rect 197353 154264 197358 154320
rect 197414 154264 200100 154320
rect 197353 154262 200100 154264
rect 197353 154259 197419 154262
rect 172237 153778 172303 153781
rect 169924 153776 172303 153778
rect 169924 153720 172242 153776
rect 172298 153720 172303 153776
rect 169924 153718 172303 153720
rect 172237 153715 172303 153718
rect 171685 153234 171751 153237
rect 169924 153232 171751 153234
rect 169924 153176 171690 153232
rect 171746 153176 171751 153232
rect 169924 153174 171751 153176
rect 171685 153171 171751 153174
rect 197353 153234 197419 153237
rect 197353 153232 200100 153234
rect 197353 153176 197358 153232
rect 197414 153176 200100 153232
rect 197353 153174 200100 153176
rect 197353 153171 197419 153174
rect 171501 152690 171567 152693
rect 169924 152688 171567 152690
rect 169924 152632 171506 152688
rect 171562 152632 171567 152688
rect 169924 152630 171567 152632
rect 171501 152627 171567 152630
rect 583385 152690 583451 152693
rect 583520 152690 584960 152780
rect 583385 152688 584960 152690
rect 583385 152632 583390 152688
rect 583446 152632 584960 152688
rect 583385 152630 584960 152632
rect 583385 152627 583451 152630
rect 583520 152540 584960 152630
rect 172329 152146 172395 152149
rect 169924 152144 172395 152146
rect 169924 152088 172334 152144
rect 172390 152088 172395 152144
rect 169924 152086 172395 152088
rect 172329 152083 172395 152086
rect 198181 152146 198247 152149
rect 198181 152144 200100 152146
rect 198181 152088 198186 152144
rect 198242 152088 200100 152144
rect 198181 152086 200100 152088
rect 198181 152083 198247 152086
rect 172329 151602 172395 151605
rect 169924 151600 172395 151602
rect 169924 151544 172334 151600
rect 172390 151544 172395 151600
rect 169924 151542 172395 151544
rect 172329 151539 172395 151542
rect 172421 151058 172487 151061
rect 169924 151056 172487 151058
rect 169924 151000 172426 151056
rect 172482 151000 172487 151056
rect 169924 150998 172487 151000
rect 172421 150995 172487 150998
rect 197445 151058 197511 151061
rect 197445 151056 200100 151058
rect 197445 151000 197450 151056
rect 197506 151000 200100 151056
rect 197445 150998 200100 151000
rect 197445 150995 197511 150998
rect 171317 150514 171383 150517
rect 169924 150512 171383 150514
rect 169924 150456 171322 150512
rect 171378 150456 171383 150512
rect 169924 150454 171383 150456
rect 171317 150451 171383 150454
rect 171869 149970 171935 149973
rect 169924 149968 171935 149970
rect -960 149834 480 149924
rect 169924 149912 171874 149968
rect 171930 149912 171935 149968
rect 169924 149910 171935 149912
rect 171869 149907 171935 149910
rect 197353 149970 197419 149973
rect 197353 149968 200100 149970
rect 197353 149912 197358 149968
rect 197414 149912 200100 149968
rect 197353 149910 200100 149912
rect 197353 149907 197419 149910
rect 3417 149834 3483 149837
rect -960 149832 3483 149834
rect -960 149776 3422 149832
rect 3478 149776 3483 149832
rect -960 149774 3483 149776
rect -960 149684 480 149774
rect 3417 149771 3483 149774
rect 171501 149426 171567 149429
rect 169924 149424 171567 149426
rect 169924 149368 171506 149424
rect 171562 149368 171567 149424
rect 169924 149366 171567 149368
rect 171501 149363 171567 149366
rect 172421 148882 172487 148885
rect 169924 148880 172487 148882
rect 169924 148824 172426 148880
rect 172482 148824 172487 148880
rect 169924 148822 172487 148824
rect 172421 148819 172487 148822
rect 197537 148882 197603 148885
rect 197537 148880 200100 148882
rect 197537 148824 197542 148880
rect 197598 148824 200100 148880
rect 197537 148822 200100 148824
rect 197537 148819 197603 148822
rect 171317 148338 171383 148341
rect 169924 148336 171383 148338
rect 169924 148280 171322 148336
rect 171378 148280 171383 148336
rect 169924 148278 171383 148280
rect 171317 148275 171383 148278
rect 171685 147794 171751 147797
rect 169924 147792 171751 147794
rect 169924 147736 171690 147792
rect 171746 147736 171751 147792
rect 169924 147734 171751 147736
rect 171685 147731 171751 147734
rect 198089 147794 198155 147797
rect 198089 147792 200100 147794
rect 198089 147736 198094 147792
rect 198150 147736 200100 147792
rect 198089 147734 200100 147736
rect 198089 147731 198155 147734
rect 172421 147250 172487 147253
rect 169924 147248 172487 147250
rect 169924 147192 172426 147248
rect 172482 147192 172487 147248
rect 169924 147190 172487 147192
rect 172421 147187 172487 147190
rect 171961 146706 172027 146709
rect 169924 146704 172027 146706
rect 169924 146648 171966 146704
rect 172022 146648 172027 146704
rect 169924 146646 172027 146648
rect 171961 146643 172027 146646
rect 198181 146706 198247 146709
rect 198181 146704 200100 146706
rect 198181 146648 198186 146704
rect 198242 146648 200100 146704
rect 198181 146646 200100 146648
rect 198181 146643 198247 146646
rect 172145 146162 172211 146165
rect 169924 146160 172211 146162
rect 169924 146104 172150 146160
rect 172206 146104 172211 146160
rect 169924 146102 172211 146104
rect 172145 146099 172211 146102
rect 172421 145618 172487 145621
rect 169924 145616 172487 145618
rect 169924 145560 172426 145616
rect 172482 145560 172487 145616
rect 169924 145558 172487 145560
rect 172421 145555 172487 145558
rect 197353 145618 197419 145621
rect 197353 145616 200100 145618
rect 197353 145560 197358 145616
rect 197414 145560 200100 145616
rect 197353 145558 200100 145560
rect 197353 145555 197419 145558
rect 172329 145074 172395 145077
rect 169924 145072 172395 145074
rect 169924 145016 172334 145072
rect 172390 145016 172395 145072
rect 169924 145014 172395 145016
rect 172329 145011 172395 145014
rect 172237 144530 172303 144533
rect 169924 144528 172303 144530
rect 169924 144472 172242 144528
rect 172298 144472 172303 144528
rect 169924 144470 172303 144472
rect 172237 144467 172303 144470
rect 197445 144530 197511 144533
rect 197445 144528 200100 144530
rect 197445 144472 197450 144528
rect 197506 144472 200100 144528
rect 197445 144470 200100 144472
rect 197445 144467 197511 144470
rect 169385 144258 169451 144261
rect 169342 144256 169451 144258
rect 169342 144200 169390 144256
rect 169446 144200 169451 144256
rect 169342 144195 169451 144200
rect 169342 144092 169402 144195
rect 171317 143578 171383 143581
rect 169924 143576 171383 143578
rect 169924 143520 171322 143576
rect 171378 143520 171383 143576
rect 169924 143518 171383 143520
rect 171317 143515 171383 143518
rect 197353 143442 197419 143445
rect 197353 143440 200100 143442
rect 197353 143384 197358 143440
rect 197414 143384 200100 143440
rect 197353 143382 200100 143384
rect 197353 143379 197419 143382
rect 171685 143034 171751 143037
rect 169924 143032 171751 143034
rect 169924 142976 171690 143032
rect 171746 142976 171751 143032
rect 169924 142974 171751 142976
rect 171685 142971 171751 142974
rect 172421 142490 172487 142493
rect 169924 142488 172487 142490
rect 169924 142432 172426 142488
rect 172482 142432 172487 142488
rect 169924 142430 172487 142432
rect 172421 142427 172487 142430
rect 197353 142218 197419 142221
rect 197353 142216 200100 142218
rect 197353 142160 197358 142216
rect 197414 142160 200100 142216
rect 197353 142158 200100 142160
rect 197353 142155 197419 142158
rect 171501 141946 171567 141949
rect 169924 141944 171567 141946
rect 169924 141888 171506 141944
rect 171562 141888 171567 141944
rect 169924 141886 171567 141888
rect 171501 141883 171567 141886
rect 172421 141402 172487 141405
rect 169924 141400 172487 141402
rect 169924 141344 172426 141400
rect 172482 141344 172487 141400
rect 169924 141342 172487 141344
rect 172421 141339 172487 141342
rect 198181 141130 198247 141133
rect 198181 141128 200100 141130
rect 198181 141072 198186 141128
rect 198242 141072 200100 141128
rect 198181 141070 200100 141072
rect 198181 141067 198247 141070
rect 171501 140858 171567 140861
rect 169924 140856 171567 140858
rect 169924 140800 171506 140856
rect 171562 140800 171567 140856
rect 169924 140798 171567 140800
rect 171501 140795 171567 140798
rect 172421 140314 172487 140317
rect 169924 140312 172487 140314
rect 169924 140256 172426 140312
rect 172482 140256 172487 140312
rect 169924 140254 172487 140256
rect 172421 140251 172487 140254
rect 197353 140042 197419 140045
rect 197353 140040 200100 140042
rect 197353 139984 197358 140040
rect 197414 139984 200100 140040
rect 197353 139982 200100 139984
rect 197353 139979 197419 139982
rect 171685 139770 171751 139773
rect 169924 139768 171751 139770
rect 169924 139712 171690 139768
rect 171746 139712 171751 139768
rect 169924 139710 171751 139712
rect 171685 139707 171751 139710
rect 583293 139362 583359 139365
rect 583520 139362 584960 139452
rect 583293 139360 584960 139362
rect 583293 139304 583298 139360
rect 583354 139304 584960 139360
rect 583293 139302 584960 139304
rect 583293 139299 583359 139302
rect 172421 139226 172487 139229
rect 169924 139224 172487 139226
rect 169924 139168 172426 139224
rect 172482 139168 172487 139224
rect 583520 139212 584960 139302
rect 169924 139166 172487 139168
rect 172421 139163 172487 139166
rect 198181 138954 198247 138957
rect 198181 138952 200100 138954
rect 198181 138896 198186 138952
rect 198242 138896 200100 138952
rect 198181 138894 200100 138896
rect 198181 138891 198247 138894
rect 171317 138682 171383 138685
rect 169924 138680 171383 138682
rect 169924 138624 171322 138680
rect 171378 138624 171383 138680
rect 169924 138622 171383 138624
rect 171317 138619 171383 138622
rect 171961 138138 172027 138141
rect 169924 138136 172027 138138
rect 169924 138080 171966 138136
rect 172022 138080 172027 138136
rect 169924 138078 172027 138080
rect 171961 138075 172027 138078
rect 197537 137866 197603 137869
rect 197537 137864 200100 137866
rect 197537 137808 197542 137864
rect 197598 137808 200100 137864
rect 197537 137806 200100 137808
rect 197537 137803 197603 137806
rect 170489 137594 170555 137597
rect 169924 137592 170555 137594
rect 169924 137536 170494 137592
rect 170550 137536 170555 137592
rect 169924 137534 170555 137536
rect 170489 137531 170555 137534
rect 171501 137050 171567 137053
rect 169924 137048 171567 137050
rect 169924 136992 171506 137048
rect 171562 136992 171567 137048
rect 169924 136990 171567 136992
rect 171501 136987 171567 136990
rect -960 136778 480 136868
rect 3233 136778 3299 136781
rect -960 136776 3299 136778
rect -960 136720 3238 136776
rect 3294 136720 3299 136776
rect -960 136718 3299 136720
rect -960 136628 480 136718
rect 3233 136715 3299 136718
rect 198457 136778 198523 136781
rect 198457 136776 200100 136778
rect 198457 136720 198462 136776
rect 198518 136720 200100 136776
rect 198457 136718 200100 136720
rect 198457 136715 198523 136718
rect 172421 136506 172487 136509
rect 169924 136504 172487 136506
rect 169924 136448 172426 136504
rect 172482 136448 172487 136504
rect 169924 136446 172487 136448
rect 172421 136443 172487 136446
rect 171685 135962 171751 135965
rect 169924 135960 171751 135962
rect 169924 135904 171690 135960
rect 171746 135904 171751 135960
rect 169924 135902 171751 135904
rect 171685 135899 171751 135902
rect 198181 135690 198247 135693
rect 198181 135688 200100 135690
rect 198181 135632 198186 135688
rect 198242 135632 200100 135688
rect 198181 135630 200100 135632
rect 198181 135627 198247 135630
rect 171501 135418 171567 135421
rect 169924 135416 171567 135418
rect 169924 135360 171506 135416
rect 171562 135360 171567 135416
rect 169924 135358 171567 135360
rect 171501 135355 171567 135358
rect 171869 134874 171935 134877
rect 169924 134872 171935 134874
rect 169924 134816 171874 134872
rect 171930 134816 171935 134872
rect 169924 134814 171935 134816
rect 171869 134811 171935 134814
rect 197353 134602 197419 134605
rect 197353 134600 200100 134602
rect 197353 134544 197358 134600
rect 197414 134544 200100 134600
rect 197353 134542 200100 134544
rect 197353 134539 197419 134542
rect 171501 134330 171567 134333
rect 169924 134328 171567 134330
rect 169924 134272 171506 134328
rect 171562 134272 171567 134328
rect 169924 134270 171567 134272
rect 171501 134267 171567 134270
rect 171869 133922 171935 133925
rect 169924 133920 171935 133922
rect 169924 133864 171874 133920
rect 171930 133864 171935 133920
rect 169924 133862 171935 133864
rect 171869 133859 171935 133862
rect 197445 133514 197511 133517
rect 197445 133512 200100 133514
rect 197445 133456 197450 133512
rect 197506 133456 200100 133512
rect 197445 133454 200100 133456
rect 197445 133451 197511 133454
rect 172421 133378 172487 133381
rect 169924 133376 172487 133378
rect 169924 133320 172426 133376
rect 172482 133320 172487 133376
rect 169924 133318 172487 133320
rect 172421 133315 172487 133318
rect 171685 132834 171751 132837
rect 169924 132832 171751 132834
rect 169924 132776 171690 132832
rect 171746 132776 171751 132832
rect 169924 132774 171751 132776
rect 171685 132771 171751 132774
rect 197353 132426 197419 132429
rect 197353 132424 200100 132426
rect 197353 132368 197358 132424
rect 197414 132368 200100 132424
rect 197353 132366 200100 132368
rect 197353 132363 197419 132366
rect 171685 132290 171751 132293
rect 169924 132288 171751 132290
rect 169924 132232 171690 132288
rect 171746 132232 171751 132288
rect 169924 132230 171751 132232
rect 171685 132227 171751 132230
rect 172421 131746 172487 131749
rect 169924 131744 172487 131746
rect 169924 131688 172426 131744
rect 172482 131688 172487 131744
rect 169924 131686 172487 131688
rect 172421 131683 172487 131686
rect 197905 131338 197971 131341
rect 197905 131336 200100 131338
rect 197905 131280 197910 131336
rect 197966 131280 200100 131336
rect 197905 131278 200100 131280
rect 197905 131275 197971 131278
rect 172421 131202 172487 131205
rect 169924 131200 172487 131202
rect 169924 131144 172426 131200
rect 172482 131144 172487 131200
rect 169924 131142 172487 131144
rect 172421 131139 172487 131142
rect 171685 130658 171751 130661
rect 169924 130656 171751 130658
rect 169924 130600 171690 130656
rect 171746 130600 171751 130656
rect 169924 130598 171751 130600
rect 171685 130595 171751 130598
rect 197997 130250 198063 130253
rect 197997 130248 200100 130250
rect 197997 130192 198002 130248
rect 198058 130192 200100 130248
rect 197997 130190 200100 130192
rect 197997 130187 198063 130190
rect 172053 130114 172119 130117
rect 169924 130112 172119 130114
rect 169924 130056 172058 130112
rect 172114 130056 172119 130112
rect 169924 130054 172119 130056
rect 172053 130051 172119 130054
rect 170397 129570 170463 129573
rect 169924 129568 170463 129570
rect 169924 129512 170402 129568
rect 170458 129512 170463 129568
rect 169924 129510 170463 129512
rect 170397 129507 170463 129510
rect 197353 129162 197419 129165
rect 197353 129160 200100 129162
rect 197353 129104 197358 129160
rect 197414 129104 200100 129160
rect 197353 129102 200100 129104
rect 197353 129099 197419 129102
rect 171593 129026 171659 129029
rect 169924 129024 171659 129026
rect 169924 128968 171598 129024
rect 171654 128968 171659 129024
rect 169924 128966 171659 128968
rect 171593 128963 171659 128966
rect 172421 128482 172487 128485
rect 169924 128480 172487 128482
rect 169924 128424 172426 128480
rect 172482 128424 172487 128480
rect 169924 128422 172487 128424
rect 172421 128419 172487 128422
rect 171685 127938 171751 127941
rect 169924 127936 171751 127938
rect 169924 127880 171690 127936
rect 171746 127880 171751 127936
rect 169924 127878 171751 127880
rect 171685 127875 171751 127878
rect 198089 127938 198155 127941
rect 198089 127936 200100 127938
rect 198089 127880 198094 127936
rect 198150 127880 200100 127936
rect 198089 127878 200100 127880
rect 198089 127875 198155 127878
rect 172053 127394 172119 127397
rect 169924 127392 172119 127394
rect 169924 127336 172058 127392
rect 172114 127336 172119 127392
rect 169924 127334 172119 127336
rect 172053 127331 172119 127334
rect 172329 126850 172395 126853
rect 169924 126848 172395 126850
rect 169924 126792 172334 126848
rect 172390 126792 172395 126848
rect 169924 126790 172395 126792
rect 172329 126787 172395 126790
rect 197353 126850 197419 126853
rect 197353 126848 200100 126850
rect 197353 126792 197358 126848
rect 197414 126792 200100 126848
rect 197353 126790 200100 126792
rect 197353 126787 197419 126790
rect 172145 126306 172211 126309
rect 169924 126304 172211 126306
rect 169924 126248 172150 126304
rect 172206 126248 172211 126304
rect 169924 126246 172211 126248
rect 172145 126243 172211 126246
rect 583201 126034 583267 126037
rect 583520 126034 584960 126124
rect 583201 126032 584960 126034
rect 583201 125976 583206 126032
rect 583262 125976 584960 126032
rect 583201 125974 584960 125976
rect 583201 125971 583267 125974
rect 583520 125884 584960 125974
rect 172421 125762 172487 125765
rect 169924 125760 172487 125762
rect 169924 125704 172426 125760
rect 172482 125704 172487 125760
rect 169924 125702 172487 125704
rect 172421 125699 172487 125702
rect 197445 125762 197511 125765
rect 197445 125760 200100 125762
rect 197445 125704 197450 125760
rect 197506 125704 200100 125760
rect 197445 125702 200100 125704
rect 197445 125699 197511 125702
rect 171869 125218 171935 125221
rect 169924 125216 171935 125218
rect 169924 125160 171874 125216
rect 171930 125160 171935 125216
rect 169924 125158 171935 125160
rect 171869 125155 171935 125158
rect 171685 124674 171751 124677
rect 169924 124672 171751 124674
rect 169924 124616 171690 124672
rect 171746 124616 171751 124672
rect 169924 124614 171751 124616
rect 171685 124611 171751 124614
rect 197629 124674 197695 124677
rect 197629 124672 200100 124674
rect 197629 124616 197634 124672
rect 197690 124616 200100 124672
rect 197629 124614 200100 124616
rect 197629 124611 197695 124614
rect 172421 124266 172487 124269
rect 169924 124264 172487 124266
rect 169924 124208 172426 124264
rect 172482 124208 172487 124264
rect 169924 124206 172487 124208
rect 172421 124203 172487 124206
rect -960 123572 480 123812
rect 197905 123586 197971 123589
rect 197905 123584 200100 123586
rect 197905 123528 197910 123584
rect 197966 123528 200100 123584
rect 197905 123526 200100 123528
rect 197905 123523 197971 123526
rect 197353 122498 197419 122501
rect 197353 122496 200100 122498
rect 197353 122440 197358 122496
rect 197414 122440 200100 122496
rect 197353 122438 200100 122440
rect 197353 122435 197419 122438
rect 197353 121410 197419 121413
rect 197353 121408 200100 121410
rect 197353 121352 197358 121408
rect 197414 121352 200100 121408
rect 197353 121350 200100 121352
rect 197353 121347 197419 121350
rect 197537 120322 197603 120325
rect 197537 120320 200100 120322
rect 197537 120264 197542 120320
rect 197598 120264 200100 120320
rect 197537 120262 200100 120264
rect 197537 120259 197603 120262
rect 198273 119234 198339 119237
rect 198273 119232 200100 119234
rect 198273 119176 198278 119232
rect 198334 119176 200100 119232
rect 198273 119174 200100 119176
rect 198273 119171 198339 119174
rect 197353 118146 197419 118149
rect 197353 118144 200100 118146
rect 197353 118088 197358 118144
rect 197414 118088 200100 118144
rect 197353 118086 200100 118088
rect 197353 118083 197419 118086
rect 198457 117058 198523 117061
rect 198457 117056 200100 117058
rect 198457 117000 198462 117056
rect 198518 117000 200100 117056
rect 198457 116998 200100 117000
rect 198457 116995 198523 116998
rect 197629 115970 197695 115973
rect 197629 115968 200100 115970
rect 197629 115912 197634 115968
rect 197690 115912 200100 115968
rect 197629 115910 200100 115912
rect 197629 115907 197695 115910
rect 197905 114882 197971 114885
rect 197905 114880 200100 114882
rect 197905 114824 197910 114880
rect 197966 114824 200100 114880
rect 197905 114822 200100 114824
rect 197905 114819 197971 114822
rect 197353 113658 197419 113661
rect 197353 113656 200100 113658
rect 197353 113600 197358 113656
rect 197414 113600 200100 113656
rect 197353 113598 200100 113600
rect 197353 113595 197419 113598
rect 583109 112842 583175 112845
rect 583520 112842 584960 112932
rect 583109 112840 584960 112842
rect 583109 112784 583114 112840
rect 583170 112784 584960 112840
rect 583109 112782 584960 112784
rect 583109 112779 583175 112782
rect 583520 112692 584960 112782
rect 197353 112570 197419 112573
rect 197353 112568 200100 112570
rect 197353 112512 197358 112568
rect 197414 112512 200100 112568
rect 197353 112510 200100 112512
rect 197353 112507 197419 112510
rect 197353 111482 197419 111485
rect 197353 111480 200100 111482
rect 197353 111424 197358 111480
rect 197414 111424 200100 111480
rect 197353 111422 200100 111424
rect 197353 111419 197419 111422
rect -960 110666 480 110756
rect 3417 110666 3483 110669
rect -960 110664 3483 110666
rect -960 110608 3422 110664
rect 3478 110608 3483 110664
rect -960 110606 3483 110608
rect -960 110516 480 110606
rect 3417 110603 3483 110606
rect 197353 110394 197419 110397
rect 197353 110392 200100 110394
rect 197353 110336 197358 110392
rect 197414 110336 200100 110392
rect 197353 110334 200100 110336
rect 197353 110331 197419 110334
rect 197537 109306 197603 109309
rect 197537 109304 200100 109306
rect 197537 109248 197542 109304
rect 197598 109248 200100 109304
rect 197537 109246 200100 109248
rect 197537 109243 197603 109246
rect 197997 108218 198063 108221
rect 197997 108216 200100 108218
rect 197997 108160 198002 108216
rect 198058 108160 200100 108216
rect 197997 108158 200100 108160
rect 197997 108155 198063 108158
rect 197537 107130 197603 107133
rect 197537 107128 200100 107130
rect 197537 107072 197542 107128
rect 197598 107072 200100 107128
rect 197537 107070 200100 107072
rect 197537 107067 197603 107070
rect 198549 106042 198615 106045
rect 198549 106040 200100 106042
rect 198549 105984 198554 106040
rect 198610 105984 200100 106040
rect 198549 105982 200100 105984
rect 198549 105979 198615 105982
rect 198089 104954 198155 104957
rect 198089 104952 200100 104954
rect 198089 104896 198094 104952
rect 198150 104896 200100 104952
rect 198089 104894 200100 104896
rect 198089 104891 198155 104894
rect 197537 103866 197603 103869
rect 197537 103864 200100 103866
rect 197537 103808 197542 103864
rect 197598 103808 200100 103864
rect 197537 103806 200100 103808
rect 197537 103803 197603 103806
rect 197445 102778 197511 102781
rect 197445 102776 200100 102778
rect 197445 102720 197450 102776
rect 197506 102720 200100 102776
rect 197445 102718 200100 102720
rect 197445 102715 197511 102718
rect 298134 102172 298140 102236
rect 298204 102234 298210 102236
rect 583385 102234 583451 102237
rect 298204 102232 583451 102234
rect 298204 102176 583390 102232
rect 583446 102176 583451 102232
rect 298204 102174 583451 102176
rect 298204 102172 298210 102174
rect 583385 102171 583451 102174
rect 197905 101690 197971 101693
rect 197905 101688 200100 101690
rect 197905 101632 197910 101688
rect 197966 101632 200100 101688
rect 197905 101630 200100 101632
rect 197905 101627 197971 101630
rect 15837 101010 15903 101013
rect 199929 101010 199995 101013
rect 583109 101010 583175 101013
rect 15837 101008 199995 101010
rect 15837 100952 15842 101008
rect 15898 100952 199934 101008
rect 199990 100952 199995 101008
rect 15837 100950 199995 100952
rect 15837 100947 15903 100950
rect 199929 100947 199995 100950
rect 298694 101008 583175 101010
rect 298694 100952 583114 101008
rect 583170 100952 583175 101008
rect 298694 100950 583175 100952
rect 298553 100738 298619 100741
rect 298694 100738 298754 100950
rect 583109 100947 583175 100950
rect 583201 100874 583267 100877
rect 298553 100736 298754 100738
rect 298553 100680 298558 100736
rect 298614 100680 298754 100736
rect 298553 100678 298754 100680
rect 298878 100872 583267 100874
rect 298878 100816 583206 100872
rect 583262 100816 583267 100872
rect 298878 100814 583267 100816
rect 298553 100675 298619 100678
rect 198089 100602 198155 100605
rect 198089 100600 200100 100602
rect 198089 100544 198094 100600
rect 198150 100544 200100 100600
rect 198089 100542 200100 100544
rect 198089 100539 198155 100542
rect 297909 100466 297975 100469
rect 298878 100466 298938 100814
rect 583201 100811 583267 100814
rect 297909 100464 298938 100466
rect 297909 100408 297914 100464
rect 297970 100408 298938 100464
rect 297909 100406 298938 100408
rect 297909 100403 297975 100406
rect 297909 100332 297975 100333
rect 297909 100330 297956 100332
rect 297864 100328 297956 100330
rect 297864 100272 297914 100328
rect 297864 100270 297956 100272
rect 297909 100268 297956 100270
rect 298020 100268 298026 100332
rect 297909 100267 297975 100268
rect 290917 99650 290983 99653
rect 529933 99650 529999 99653
rect 290917 99648 529999 99650
rect 290917 99592 290922 99648
rect 290978 99592 529938 99648
rect 529994 99592 529999 99648
rect 290917 99590 529999 99592
rect 290917 99587 290983 99590
rect 529933 99587 529999 99590
rect 293953 99514 294019 99517
rect 550633 99514 550699 99517
rect 293953 99512 550699 99514
rect 293953 99456 293958 99512
rect 294014 99456 550638 99512
rect 550694 99456 550699 99512
rect 293953 99454 550699 99456
rect 293953 99451 294019 99454
rect 550633 99451 550699 99454
rect 583017 99514 583083 99517
rect 583520 99514 584960 99604
rect 583017 99512 584960 99514
rect 583017 99456 583022 99512
rect 583078 99456 584960 99512
rect 583017 99454 584960 99456
rect 583017 99451 583083 99454
rect 583520 99364 584960 99454
rect 284845 98970 284911 98973
rect 493317 98970 493383 98973
rect 284845 98968 493383 98970
rect 284845 98912 284850 98968
rect 284906 98912 493322 98968
rect 493378 98912 493383 98968
rect 284845 98910 493383 98912
rect 284845 98907 284911 98910
rect 493317 98907 493383 98910
rect 80697 98834 80763 98837
rect 208761 98834 208827 98837
rect 80697 98832 208827 98834
rect 80697 98776 80702 98832
rect 80758 98776 208766 98832
rect 208822 98776 208827 98832
rect 80697 98774 208827 98776
rect 80697 98771 80763 98774
rect 208761 98771 208827 98774
rect 284293 98834 284359 98837
rect 494053 98834 494119 98837
rect 284293 98832 494119 98834
rect 284293 98776 284298 98832
rect 284354 98776 494058 98832
rect 494114 98776 494119 98832
rect 284293 98774 494119 98776
rect 284293 98771 284359 98774
rect 494053 98771 494119 98774
rect 30281 98698 30347 98701
rect 205173 98698 205239 98701
rect 30281 98696 205239 98698
rect 30281 98640 30286 98696
rect 30342 98640 205178 98696
rect 205234 98640 205239 98696
rect 30281 98638 205239 98640
rect 30281 98635 30347 98638
rect 205173 98635 205239 98638
rect 291561 98698 291627 98701
rect 532693 98698 532759 98701
rect 291561 98696 532759 98698
rect 291561 98640 291566 98696
rect 291622 98640 532698 98696
rect 532754 98640 532759 98696
rect 291561 98638 532759 98640
rect 291561 98635 291627 98638
rect 532693 98635 532759 98638
rect 283005 97882 283071 97885
rect 285765 97882 285831 97885
rect 283005 97880 285831 97882
rect 283005 97824 283010 97880
rect 283066 97824 285770 97880
rect 285826 97824 285831 97880
rect 283005 97822 285831 97824
rect 283005 97819 283071 97822
rect 285765 97819 285831 97822
rect -960 97610 480 97700
rect 3417 97610 3483 97613
rect -960 97608 3483 97610
rect -960 97552 3422 97608
rect 3478 97552 3483 97608
rect -960 97550 3483 97552
rect -960 97460 480 97550
rect 3417 97547 3483 97550
rect 219382 97548 219388 97612
rect 219452 97610 219458 97612
rect 219525 97610 219591 97613
rect 219452 97608 219591 97610
rect 219452 97552 219530 97608
rect 219586 97552 219591 97608
rect 219452 97550 219591 97552
rect 219452 97548 219458 97550
rect 219525 97547 219591 97550
rect 292573 97474 292639 97477
rect 295793 97474 295859 97477
rect 304993 97474 305059 97477
rect 292573 97472 294706 97474
rect 292573 97416 292578 97472
rect 292634 97416 294706 97472
rect 292573 97414 294706 97416
rect 292573 97411 292639 97414
rect 188337 97338 188403 97341
rect 200113 97338 200179 97341
rect 188337 97336 200179 97338
rect 188337 97280 188342 97336
rect 188398 97280 200118 97336
rect 200174 97280 200179 97336
rect 188337 97278 200179 97280
rect 188337 97275 188403 97278
rect 200113 97275 200179 97278
rect 292430 97276 292436 97340
rect 292500 97338 292506 97340
rect 293585 97338 293651 97341
rect 292500 97336 293651 97338
rect 292500 97280 293590 97336
rect 293646 97280 293651 97336
rect 292500 97278 293651 97280
rect 294646 97338 294706 97414
rect 295793 97472 305059 97474
rect 295793 97416 295798 97472
rect 295854 97416 304998 97472
rect 305054 97416 305059 97472
rect 295793 97414 305059 97416
rect 295793 97411 295859 97414
rect 304993 97411 305059 97414
rect 312537 97338 312603 97341
rect 294646 97336 312603 97338
rect 294646 97280 312542 97336
rect 312598 97280 312603 97336
rect 294646 97278 312603 97280
rect 292500 97276 292506 97278
rect 293585 97275 293651 97278
rect 312537 97275 312603 97278
rect 46197 97202 46263 97205
rect 200849 97202 200915 97205
rect 46197 97200 200915 97202
rect 46197 97144 46202 97200
rect 46258 97144 200854 97200
rect 200910 97144 200915 97200
rect 46197 97142 200915 97144
rect 46197 97139 46263 97142
rect 200849 97139 200915 97142
rect 271454 97140 271460 97204
rect 271524 97202 271530 97204
rect 271689 97202 271755 97205
rect 271524 97200 271755 97202
rect 271524 97144 271694 97200
rect 271750 97144 271755 97200
rect 271524 97142 271755 97144
rect 271524 97140 271530 97142
rect 271689 97139 271755 97142
rect 277393 97202 277459 97205
rect 403617 97202 403683 97205
rect 277393 97200 403683 97202
rect 277393 97144 277398 97200
rect 277454 97144 403622 97200
rect 403678 97144 403683 97200
rect 277393 97142 403683 97144
rect 277393 97139 277459 97142
rect 403617 97139 403683 97142
rect 252001 97066 252067 97069
rect 252502 97066 252508 97068
rect 252001 97064 252508 97066
rect 252001 97008 252006 97064
rect 252062 97008 252508 97064
rect 252001 97006 252508 97008
rect 252001 97003 252067 97006
rect 252502 97004 252508 97006
rect 252572 97004 252578 97068
rect 259085 97066 259151 97069
rect 259310 97066 259316 97068
rect 259085 97064 259316 97066
rect 259085 97008 259090 97064
rect 259146 97008 259316 97064
rect 259085 97006 259316 97008
rect 259085 97003 259151 97006
rect 259310 97004 259316 97006
rect 259380 97004 259386 97068
rect 260598 97004 260604 97068
rect 260668 97066 260674 97068
rect 260741 97066 260807 97069
rect 260668 97064 260807 97066
rect 260668 97008 260746 97064
rect 260802 97008 260807 97064
rect 260668 97006 260807 97008
rect 260668 97004 260674 97006
rect 260741 97003 260807 97006
rect 264462 97004 264468 97068
rect 264532 97066 264538 97068
rect 264789 97066 264855 97069
rect 267457 97068 267523 97069
rect 267406 97066 267412 97068
rect 264532 97064 264855 97066
rect 264532 97008 264794 97064
rect 264850 97008 264855 97064
rect 264532 97006 264855 97008
rect 267366 97006 267412 97066
rect 267476 97064 267523 97068
rect 267518 97008 267523 97064
rect 264532 97004 264538 97006
rect 264789 97003 264855 97006
rect 267406 97004 267412 97006
rect 267476 97004 267523 97008
rect 267457 97003 267523 97004
rect 272885 97066 272951 97069
rect 273110 97066 273116 97068
rect 272885 97064 273116 97066
rect 272885 97008 272890 97064
rect 272946 97008 273116 97064
rect 272885 97006 273116 97008
rect 272885 97003 272951 97006
rect 273110 97004 273116 97006
rect 273180 97004 273186 97068
rect 274214 97004 274220 97068
rect 274284 97066 274290 97068
rect 274541 97066 274607 97069
rect 274284 97064 274607 97066
rect 274284 97008 274546 97064
rect 274602 97008 274607 97064
rect 274284 97006 274607 97008
rect 274284 97004 274290 97006
rect 274541 97003 274607 97006
rect 275318 97004 275324 97068
rect 275388 97066 275394 97068
rect 275921 97066 275987 97069
rect 275388 97064 275987 97066
rect 275388 97008 275926 97064
rect 275982 97008 275987 97064
rect 275388 97006 275987 97008
rect 275388 97004 275394 97006
rect 275921 97003 275987 97006
rect 278998 97004 279004 97068
rect 279068 97066 279074 97068
rect 279969 97066 280035 97069
rect 279068 97064 280035 97066
rect 279068 97008 279974 97064
rect 280030 97008 280035 97064
rect 279068 97006 280035 97008
rect 279068 97004 279074 97006
rect 279969 97003 280035 97006
rect 202822 96868 202828 96932
rect 202892 96930 202898 96932
rect 203149 96930 203215 96933
rect 202892 96928 203215 96930
rect 202892 96872 203154 96928
rect 203210 96872 203215 96928
rect 202892 96870 203215 96872
rect 202892 96868 202898 96870
rect 203149 96867 203215 96870
rect 205909 96932 205975 96933
rect 205909 96928 205956 96932
rect 206020 96930 206026 96932
rect 205909 96872 205914 96928
rect 205909 96868 205956 96872
rect 206020 96870 206066 96930
rect 206020 96868 206026 96870
rect 215334 96868 215340 96932
rect 215404 96930 215410 96932
rect 215661 96930 215727 96933
rect 216673 96932 216739 96933
rect 216622 96930 216628 96932
rect 215404 96928 215727 96930
rect 215404 96872 215666 96928
rect 215722 96872 215727 96928
rect 215404 96870 215727 96872
rect 216582 96870 216628 96930
rect 216692 96928 216739 96932
rect 216734 96872 216739 96928
rect 215404 96868 215410 96870
rect 205909 96867 205975 96868
rect 215661 96867 215727 96870
rect 216622 96868 216628 96870
rect 216692 96868 216739 96872
rect 216673 96867 216739 96868
rect 218329 96930 218395 96933
rect 218646 96930 218652 96932
rect 218329 96928 218652 96930
rect 218329 96872 218334 96928
rect 218390 96872 218652 96928
rect 218329 96870 218652 96872
rect 218329 96867 218395 96870
rect 218646 96868 218652 96870
rect 218716 96868 218722 96932
rect 220854 96868 220860 96932
rect 220924 96930 220930 96932
rect 220997 96930 221063 96933
rect 222377 96932 222443 96933
rect 222326 96930 222332 96932
rect 220924 96928 221063 96930
rect 220924 96872 221002 96928
rect 221058 96872 221063 96928
rect 220924 96870 221063 96872
rect 222286 96870 222332 96930
rect 222396 96928 222443 96932
rect 222438 96872 222443 96928
rect 220924 96868 220930 96870
rect 220997 96867 221063 96870
rect 222326 96868 222332 96870
rect 222396 96868 222443 96872
rect 222377 96867 222443 96868
rect 223573 96932 223639 96933
rect 237557 96932 237623 96933
rect 223573 96928 223620 96932
rect 223684 96930 223690 96932
rect 223573 96872 223578 96928
rect 223573 96868 223620 96872
rect 223684 96870 223730 96930
rect 237557 96928 237604 96932
rect 237668 96930 237674 96932
rect 237833 96930 237899 96933
rect 237557 96872 237562 96928
rect 223684 96868 223690 96870
rect 237557 96868 237604 96872
rect 237668 96870 237714 96930
rect 237790 96928 237899 96930
rect 237790 96872 237838 96928
rect 237894 96872 237899 96928
rect 237668 96868 237674 96870
rect 223573 96867 223639 96868
rect 237557 96867 237623 96868
rect 237790 96867 237899 96872
rect 246798 96868 246804 96932
rect 246868 96930 246874 96932
rect 246941 96930 247007 96933
rect 246868 96928 247007 96930
rect 246868 96872 246946 96928
rect 247002 96872 247007 96928
rect 246868 96870 247007 96872
rect 246868 96868 246874 96870
rect 246941 96867 247007 96870
rect 249517 96932 249583 96933
rect 249517 96928 249564 96932
rect 249628 96930 249634 96932
rect 249517 96872 249522 96928
rect 249517 96868 249564 96872
rect 249628 96870 249674 96930
rect 249628 96868 249634 96870
rect 250846 96868 250852 96932
rect 250916 96930 250922 96932
rect 250989 96930 251055 96933
rect 252369 96932 252435 96933
rect 253657 96932 253723 96933
rect 252318 96930 252324 96932
rect 250916 96928 251055 96930
rect 250916 96872 250994 96928
rect 251050 96872 251055 96928
rect 250916 96870 251055 96872
rect 252278 96870 252324 96930
rect 252388 96928 252435 96932
rect 253606 96930 253612 96932
rect 252430 96872 252435 96928
rect 250916 96868 250922 96870
rect 249517 96867 249583 96868
rect 250989 96867 251055 96870
rect 252318 96868 252324 96870
rect 252388 96868 252435 96872
rect 253566 96870 253612 96930
rect 253676 96928 253723 96932
rect 253718 96872 253723 96928
rect 253606 96868 253612 96870
rect 253676 96868 253723 96872
rect 255078 96868 255084 96932
rect 255148 96930 255154 96932
rect 255221 96930 255287 96933
rect 255148 96928 255287 96930
rect 255148 96872 255226 96928
rect 255282 96872 255287 96928
rect 255148 96870 255287 96872
rect 255148 96868 255154 96870
rect 252369 96867 252435 96868
rect 253657 96867 253723 96868
rect 255221 96867 255287 96870
rect 256049 96930 256115 96933
rect 256550 96930 256556 96932
rect 256049 96928 256556 96930
rect 256049 96872 256054 96928
rect 256110 96872 256556 96928
rect 256049 96870 256556 96872
rect 256049 96867 256115 96870
rect 256550 96868 256556 96870
rect 256620 96868 256626 96932
rect 257286 96868 257292 96932
rect 257356 96930 257362 96932
rect 257705 96930 257771 96933
rect 257356 96928 257771 96930
rect 257356 96872 257710 96928
rect 257766 96872 257771 96928
rect 257356 96870 257771 96872
rect 257356 96868 257362 96870
rect 257705 96867 257771 96870
rect 258901 96930 258967 96933
rect 259126 96930 259132 96932
rect 258901 96928 259132 96930
rect 258901 96872 258906 96928
rect 258962 96872 259132 96928
rect 258901 96870 259132 96872
rect 258901 96867 258967 96870
rect 259126 96868 259132 96870
rect 259196 96868 259202 96932
rect 260414 96868 260420 96932
rect 260484 96930 260490 96932
rect 260557 96930 260623 96933
rect 260484 96928 260623 96930
rect 260484 96872 260562 96928
rect 260618 96872 260623 96928
rect 260484 96870 260623 96872
rect 260484 96868 260490 96870
rect 260557 96867 260623 96870
rect 262765 96930 262831 96933
rect 263317 96932 263383 96933
rect 263174 96930 263180 96932
rect 262765 96928 263180 96930
rect 262765 96872 262770 96928
rect 262826 96872 263180 96928
rect 262765 96870 263180 96872
rect 262765 96867 262831 96870
rect 263174 96868 263180 96870
rect 263244 96868 263250 96932
rect 263317 96928 263364 96932
rect 263428 96930 263434 96932
rect 264329 96930 264395 96933
rect 266169 96932 266235 96933
rect 267641 96932 267707 96933
rect 264646 96930 264652 96932
rect 263317 96872 263322 96928
rect 263317 96868 263364 96872
rect 263428 96870 263474 96930
rect 264329 96928 264652 96930
rect 264329 96872 264334 96928
rect 264390 96872 264652 96928
rect 264329 96870 264652 96872
rect 263428 96868 263434 96870
rect 263317 96867 263383 96868
rect 264329 96867 264395 96870
rect 264646 96868 264652 96870
rect 264716 96868 264722 96932
rect 266118 96930 266124 96932
rect 266078 96870 266124 96930
rect 266188 96928 266235 96932
rect 267590 96930 267596 96932
rect 266230 96872 266235 96928
rect 266118 96868 266124 96870
rect 266188 96868 266235 96872
rect 267550 96870 267596 96930
rect 267660 96928 267707 96932
rect 267702 96872 267707 96928
rect 267590 96868 267596 96870
rect 267660 96868 267707 96872
rect 268878 96868 268884 96932
rect 268948 96930 268954 96932
rect 269021 96930 269087 96933
rect 268948 96928 269087 96930
rect 268948 96872 269026 96928
rect 269082 96872 269087 96928
rect 268948 96870 269087 96872
rect 268948 96868 268954 96870
rect 266169 96867 266235 96868
rect 267641 96867 267707 96868
rect 269021 96867 269087 96870
rect 270217 96930 270283 96933
rect 270350 96930 270356 96932
rect 270217 96928 270356 96930
rect 270217 96872 270222 96928
rect 270278 96872 270356 96928
rect 270217 96870 270356 96872
rect 270217 96867 270283 96870
rect 270350 96868 270356 96870
rect 270420 96868 270426 96932
rect 271229 96930 271295 96933
rect 271638 96930 271644 96932
rect 271229 96928 271644 96930
rect 271229 96872 271234 96928
rect 271290 96872 271644 96928
rect 271229 96870 271644 96872
rect 271229 96867 271295 96870
rect 271638 96868 271644 96870
rect 271708 96868 271714 96932
rect 274265 96930 274331 96933
rect 274398 96930 274404 96932
rect 274265 96928 274404 96930
rect 274265 96872 274270 96928
rect 274326 96872 274404 96928
rect 274265 96870 274404 96872
rect 274265 96867 274331 96870
rect 274398 96868 274404 96870
rect 274468 96868 274474 96932
rect 276933 96930 276999 96933
rect 278589 96932 278655 96933
rect 281165 96932 281231 96933
rect 281441 96932 281507 96933
rect 277158 96930 277164 96932
rect 276933 96928 277164 96930
rect 276933 96872 276938 96928
rect 276994 96872 277164 96928
rect 276933 96870 277164 96872
rect 276933 96867 276999 96870
rect 277158 96868 277164 96870
rect 277228 96868 277234 96932
rect 278589 96928 278636 96932
rect 278700 96930 278706 96932
rect 278589 96872 278594 96928
rect 278589 96868 278636 96872
rect 278700 96870 278746 96930
rect 281165 96928 281212 96932
rect 281276 96930 281282 96932
rect 281165 96872 281170 96928
rect 278700 96868 278706 96870
rect 281165 96868 281212 96872
rect 281276 96870 281322 96930
rect 281276 96868 281282 96870
rect 281390 96868 281396 96932
rect 281460 96930 281507 96932
rect 281460 96928 281552 96930
rect 281502 96872 281552 96928
rect 281460 96870 281552 96872
rect 281460 96868 281507 96870
rect 282126 96868 282132 96932
rect 282196 96930 282202 96932
rect 282821 96930 282887 96933
rect 282196 96928 282887 96930
rect 282196 96872 282826 96928
rect 282882 96872 282887 96928
rect 282196 96870 282887 96872
rect 282196 96868 282202 96870
rect 278589 96867 278655 96868
rect 281165 96867 281231 96868
rect 281441 96867 281507 96868
rect 282821 96867 282887 96870
rect 284017 96930 284083 96933
rect 286869 96932 286935 96933
rect 284150 96930 284156 96932
rect 284017 96928 284156 96930
rect 284017 96872 284022 96928
rect 284078 96872 284156 96928
rect 284017 96870 284156 96872
rect 284017 96867 284083 96870
rect 284150 96868 284156 96870
rect 284220 96868 284226 96932
rect 286869 96928 286916 96932
rect 286980 96930 286986 96932
rect 286869 96872 286874 96928
rect 286869 96868 286916 96872
rect 286980 96870 287026 96930
rect 286980 96868 286986 96870
rect 288198 96868 288204 96932
rect 288268 96930 288274 96932
rect 288341 96930 288407 96933
rect 288268 96928 288407 96930
rect 288268 96872 288346 96928
rect 288402 96872 288407 96928
rect 288268 96870 288407 96872
rect 288268 96868 288274 96870
rect 286869 96867 286935 96868
rect 288341 96867 288407 96870
rect 292246 96868 292252 96932
rect 292316 96930 292322 96932
rect 292389 96930 292455 96933
rect 294965 96932 295031 96933
rect 295241 96932 295307 96933
rect 299289 96932 299355 96933
rect 294965 96930 295012 96932
rect 292316 96928 292455 96930
rect 292316 96872 292394 96928
rect 292450 96872 292455 96928
rect 292316 96870 292455 96872
rect 294920 96928 295012 96930
rect 294920 96872 294970 96928
rect 294920 96870 295012 96872
rect 292316 96868 292322 96870
rect 292389 96867 292455 96870
rect 294965 96868 295012 96870
rect 295076 96868 295082 96932
rect 295190 96930 295196 96932
rect 295150 96870 295196 96930
rect 295260 96928 295307 96932
rect 299238 96930 299244 96932
rect 295302 96872 295307 96928
rect 295190 96868 295196 96870
rect 295260 96868 295307 96872
rect 299198 96870 299244 96930
rect 299308 96928 299355 96932
rect 299350 96872 299355 96928
rect 299238 96868 299244 96870
rect 299308 96868 299355 96872
rect 294965 96867 295031 96868
rect 295241 96867 295307 96868
rect 299289 96867 299355 96868
rect 200757 96794 200823 96797
rect 207381 96794 207447 96797
rect 200757 96792 207447 96794
rect 200757 96736 200762 96792
rect 200818 96736 207386 96792
rect 207442 96736 207447 96792
rect 200757 96734 207447 96736
rect 200757 96731 200823 96734
rect 207381 96731 207447 96734
rect 230473 96794 230539 96797
rect 230606 96794 230612 96796
rect 230473 96792 230612 96794
rect 230473 96736 230478 96792
rect 230534 96736 230612 96792
rect 230473 96734 230612 96736
rect 230473 96731 230539 96734
rect 230606 96732 230612 96734
rect 230676 96732 230682 96796
rect 200941 96658 201007 96661
rect 202873 96658 202939 96661
rect 204345 96660 204411 96661
rect 204294 96658 204300 96660
rect 200941 96656 202939 96658
rect 200941 96600 200946 96656
rect 201002 96600 202878 96656
rect 202934 96600 202939 96656
rect 200941 96598 202939 96600
rect 204254 96598 204300 96658
rect 204364 96656 204411 96660
rect 204406 96600 204411 96656
rect 200941 96595 201007 96598
rect 202873 96595 202939 96598
rect 204294 96596 204300 96598
rect 204364 96596 204411 96600
rect 204345 96595 204411 96596
rect 205725 96660 205791 96661
rect 208393 96660 208459 96661
rect 205725 96656 205772 96660
rect 205836 96658 205842 96660
rect 208342 96658 208348 96660
rect 205725 96600 205730 96656
rect 205725 96596 205772 96600
rect 205836 96598 205882 96658
rect 208302 96598 208348 96658
rect 208412 96656 208459 96660
rect 209773 96660 209839 96661
rect 209773 96658 209820 96660
rect 208454 96600 208459 96656
rect 205836 96596 205842 96598
rect 208342 96596 208348 96598
rect 208412 96596 208459 96600
rect 209728 96656 209820 96658
rect 209728 96600 209778 96656
rect 209728 96598 209820 96600
rect 205725 96595 205791 96596
rect 208393 96595 208459 96596
rect 209773 96596 209820 96598
rect 209884 96596 209890 96660
rect 211429 96658 211495 96661
rect 212625 96660 212691 96661
rect 211654 96658 211660 96660
rect 211429 96656 211660 96658
rect 211429 96600 211434 96656
rect 211490 96600 211660 96656
rect 211429 96598 211660 96600
rect 209773 96595 209839 96596
rect 211429 96595 211495 96598
rect 211654 96596 211660 96598
rect 211724 96596 211730 96660
rect 212574 96658 212580 96660
rect 212534 96598 212580 96658
rect 212644 96656 212691 96660
rect 212686 96600 212691 96656
rect 212574 96596 212580 96598
rect 212644 96596 212691 96600
rect 213862 96596 213868 96660
rect 213932 96658 213938 96660
rect 214097 96658 214163 96661
rect 226425 96660 226491 96661
rect 226374 96658 226380 96660
rect 213932 96656 214163 96658
rect 213932 96600 214102 96656
rect 214158 96600 214163 96656
rect 213932 96598 214163 96600
rect 226334 96598 226380 96658
rect 226444 96656 226491 96660
rect 226486 96600 226491 96656
rect 213932 96596 213938 96598
rect 212625 96595 212691 96596
rect 214097 96595 214163 96598
rect 226374 96596 226380 96598
rect 226444 96596 226491 96600
rect 230422 96596 230428 96660
rect 230492 96658 230498 96660
rect 230933 96658 230999 96661
rect 230492 96656 230999 96658
rect 230492 96600 230938 96656
rect 230994 96600 230999 96656
rect 230492 96598 230999 96600
rect 230492 96596 230498 96598
rect 226425 96595 226491 96596
rect 230933 96595 230999 96598
rect 231894 96596 231900 96660
rect 231964 96658 231970 96660
rect 232129 96658 232195 96661
rect 231964 96656 232195 96658
rect 231964 96600 232134 96656
rect 232190 96600 232195 96656
rect 231964 96598 232195 96600
rect 231964 96596 231970 96598
rect 232129 96595 232195 96598
rect 233182 96596 233188 96660
rect 233252 96658 233258 96660
rect 233325 96658 233391 96661
rect 233252 96656 233391 96658
rect 233252 96600 233330 96656
rect 233386 96600 233391 96656
rect 233252 96598 233391 96600
rect 233252 96596 233258 96598
rect 233325 96595 233391 96598
rect 231117 96522 231183 96525
rect 237790 96522 237850 96867
rect 231117 96520 237850 96522
rect 231117 96464 231122 96520
rect 231178 96464 237850 96520
rect 231117 96462 237850 96464
rect 231117 96459 231183 96462
rect 186957 96114 187023 96117
rect 231945 96114 232011 96117
rect 186957 96112 232011 96114
rect 186957 96056 186962 96112
rect 187018 96056 231950 96112
rect 232006 96056 232011 96112
rect 186957 96054 232011 96056
rect 186957 96051 187023 96054
rect 231945 96051 232011 96054
rect 251081 96114 251147 96117
rect 303705 96114 303771 96117
rect 251081 96112 303771 96114
rect 251081 96056 251086 96112
rect 251142 96056 303710 96112
rect 303766 96056 303771 96112
rect 251081 96054 303771 96056
rect 251081 96051 251147 96054
rect 303705 96051 303771 96054
rect 130377 95978 130443 95981
rect 222193 95978 222259 95981
rect 130377 95976 222259 95978
rect 130377 95920 130382 95976
rect 130438 95920 222198 95976
rect 222254 95920 222259 95976
rect 130377 95918 222259 95920
rect 130377 95915 130443 95918
rect 222193 95915 222259 95918
rect 289721 95978 289787 95981
rect 497457 95978 497523 95981
rect 289721 95976 497523 95978
rect 289721 95920 289726 95976
rect 289782 95920 497462 95976
rect 497518 95920 497523 95976
rect 289721 95918 497523 95920
rect 289721 95915 289787 95918
rect 497457 95915 497523 95918
rect 18597 95842 18663 95845
rect 201493 95842 201559 95845
rect 18597 95840 201559 95842
rect 18597 95784 18602 95840
rect 18658 95784 201498 95840
rect 201554 95784 201559 95840
rect 18597 95782 201559 95784
rect 18597 95779 18663 95782
rect 201493 95779 201559 95782
rect 271454 95780 271460 95844
rect 271524 95842 271530 95844
rect 287973 95842 288039 95845
rect 271524 95840 288039 95842
rect 271524 95784 287978 95840
rect 288034 95784 288039 95840
rect 271524 95782 288039 95784
rect 271524 95780 271530 95782
rect 287973 95779 288039 95782
rect 291193 95842 291259 95845
rect 525793 95842 525859 95845
rect 291193 95840 525859 95842
rect 291193 95784 291198 95840
rect 291254 95784 525798 95840
rect 525854 95784 525859 95840
rect 291193 95782 525859 95784
rect 291193 95779 291259 95782
rect 525793 95779 525859 95782
rect 195237 94754 195303 94757
rect 230422 94754 230428 94756
rect 195237 94752 230428 94754
rect 195237 94696 195242 94752
rect 195298 94696 230428 94752
rect 195237 94694 230428 94696
rect 195237 94691 195303 94694
rect 230422 94692 230428 94694
rect 230492 94692 230498 94756
rect 169661 94618 169727 94621
rect 229093 94618 229159 94621
rect 169661 94616 229159 94618
rect 169661 94560 169666 94616
rect 169722 94560 229098 94616
rect 229154 94560 229159 94616
rect 169661 94558 229159 94560
rect 169661 94555 169727 94558
rect 229093 94555 229159 94558
rect 252502 94556 252508 94620
rect 252572 94618 252578 94620
rect 302233 94618 302299 94621
rect 252572 94616 302299 94618
rect 252572 94560 302238 94616
rect 302294 94560 302299 94616
rect 252572 94558 302299 94560
rect 252572 94556 252578 94558
rect 302233 94555 302299 94558
rect 153101 94482 153167 94485
rect 226374 94482 226380 94484
rect 153101 94480 226380 94482
rect 153101 94424 153106 94480
rect 153162 94424 226380 94480
rect 153101 94422 226380 94424
rect 153101 94419 153167 94422
rect 226374 94420 226380 94422
rect 226444 94420 226450 94484
rect 298277 94482 298343 94485
rect 583293 94482 583359 94485
rect 298277 94480 583359 94482
rect 298277 94424 298282 94480
rect 298338 94424 583298 94480
rect 583354 94424 583359 94480
rect 298277 94422 583359 94424
rect 298277 94419 298343 94422
rect 583293 94419 583359 94422
rect 125501 93394 125567 93397
rect 223614 93394 223620 93396
rect 125501 93392 223620 93394
rect 125501 93336 125506 93392
rect 125562 93336 223620 93392
rect 125501 93334 223620 93336
rect 125501 93331 125567 93334
rect 223614 93332 223620 93334
rect 223684 93332 223690 93396
rect 260414 93332 260420 93396
rect 260484 93394 260490 93396
rect 351913 93394 351979 93397
rect 260484 93392 351979 93394
rect 260484 93336 351918 93392
rect 351974 93336 351979 93392
rect 260484 93334 351979 93336
rect 260484 93332 260490 93334
rect 351913 93331 351979 93334
rect 34421 93258 34487 93261
rect 205766 93258 205772 93260
rect 34421 93256 205772 93258
rect 34421 93200 34426 93256
rect 34482 93200 205772 93256
rect 34421 93198 205772 93200
rect 34421 93195 34487 93198
rect 205766 93196 205772 93198
rect 205836 93196 205842 93260
rect 284150 93196 284156 93260
rect 284220 93258 284226 93260
rect 489913 93258 489979 93261
rect 284220 93256 489979 93258
rect 284220 93200 489918 93256
rect 489974 93200 489979 93256
rect 284220 93198 489979 93200
rect 284220 93196 284226 93198
rect 489913 93195 489979 93198
rect 26141 93122 26207 93125
rect 204294 93122 204300 93124
rect 26141 93120 204300 93122
rect 26141 93064 26146 93120
rect 26202 93064 204300 93120
rect 26141 93062 204300 93064
rect 26141 93059 26207 93062
rect 204294 93060 204300 93062
rect 204364 93060 204370 93124
rect 295006 93060 295012 93124
rect 295076 93122 295082 93124
rect 553393 93122 553459 93125
rect 295076 93120 553459 93122
rect 295076 93064 553398 93120
rect 553454 93064 553459 93120
rect 295076 93062 553459 93064
rect 295076 93060 295082 93062
rect 553393 93059 553459 93062
rect 177941 91898 178007 91901
rect 230606 91898 230612 91900
rect 177941 91896 230612 91898
rect 177941 91840 177946 91896
rect 178002 91840 230612 91896
rect 177941 91838 230612 91840
rect 177941 91835 178007 91838
rect 230606 91836 230612 91838
rect 230676 91836 230682 91900
rect 28257 91762 28323 91765
rect 202822 91762 202828 91764
rect 28257 91760 202828 91762
rect 28257 91704 28262 91760
rect 28318 91704 202828 91760
rect 28257 91702 202828 91704
rect 28257 91699 28323 91702
rect 202822 91700 202828 91702
rect 202892 91700 202898 91764
rect 264462 91700 264468 91764
rect 264532 91762 264538 91764
rect 376753 91762 376819 91765
rect 264532 91760 376819 91762
rect 264532 91704 376758 91760
rect 376814 91704 376819 91760
rect 264532 91702 376819 91704
rect 264532 91700 264538 91702
rect 376753 91699 376819 91702
rect 282126 91156 282132 91220
rect 282196 91218 282202 91220
rect 282545 91218 282611 91221
rect 282196 91216 282611 91218
rect 282196 91160 282550 91216
rect 282606 91160 282611 91216
rect 282196 91158 282611 91160
rect 282196 91156 282202 91158
rect 282545 91155 282611 91158
rect 295057 90674 295123 90677
rect 370497 90674 370563 90677
rect 295057 90672 370563 90674
rect 295057 90616 295062 90672
rect 295118 90616 370502 90672
rect 370558 90616 370563 90672
rect 295057 90614 370563 90616
rect 295057 90611 295123 90614
rect 370497 90611 370563 90614
rect 274214 90476 274220 90540
rect 274284 90538 274290 90540
rect 429837 90538 429903 90541
rect 274284 90536 429903 90538
rect 274284 90480 429842 90536
rect 429898 90480 429903 90536
rect 274284 90478 429903 90480
rect 274284 90476 274290 90478
rect 429837 90475 429903 90478
rect 194501 90402 194567 90405
rect 233182 90402 233188 90404
rect 194501 90400 233188 90402
rect 194501 90344 194506 90400
rect 194562 90344 233188 90400
rect 194501 90342 233188 90344
rect 194501 90339 194567 90342
rect 233182 90340 233188 90342
rect 233252 90340 233258 90404
rect 280705 90402 280771 90405
rect 440233 90402 440299 90405
rect 280705 90400 440299 90402
rect 280705 90344 280710 90400
rect 280766 90344 440238 90400
rect 440294 90344 440299 90400
rect 280705 90342 440299 90344
rect 280705 90339 280771 90342
rect 440233 90339 440299 90342
rect 97901 89178 97967 89181
rect 216622 89178 216628 89180
rect 97901 89176 216628 89178
rect 97901 89120 97906 89176
rect 97962 89120 216628 89176
rect 97901 89118 216628 89120
rect 97901 89115 97967 89118
rect 216622 89116 216628 89118
rect 216692 89116 216698 89180
rect 278998 89116 279004 89180
rect 279068 89178 279074 89180
rect 465073 89178 465139 89181
rect 279068 89176 465139 89178
rect 279068 89120 465078 89176
rect 465134 89120 465139 89176
rect 279068 89118 465139 89120
rect 279068 89116 279074 89118
rect 465073 89115 465139 89118
rect 79961 89042 80027 89045
rect 207749 89042 207815 89045
rect 79961 89040 207815 89042
rect 79961 88984 79966 89040
rect 80022 88984 207754 89040
rect 207810 88984 207815 89040
rect 79961 88982 207815 88984
rect 79961 88979 80027 88982
rect 207749 88979 207815 88982
rect 295190 88980 295196 89044
rect 295260 89042 295266 89044
rect 574093 89042 574159 89045
rect 295260 89040 574159 89042
rect 295260 88984 574098 89040
rect 574154 88984 574159 89040
rect 295260 88982 574159 88984
rect 295260 88980 295266 88982
rect 574093 88979 574159 88982
rect 292246 87756 292252 87820
rect 292316 87818 292322 87820
rect 538213 87818 538279 87821
rect 292316 87816 538279 87818
rect 292316 87760 538218 87816
rect 538274 87760 538279 87816
rect 292316 87758 538279 87760
rect 292316 87756 292322 87758
rect 538213 87755 538279 87758
rect 75177 87682 75243 87685
rect 212574 87682 212580 87684
rect 75177 87680 212580 87682
rect 75177 87624 75182 87680
rect 75238 87624 212580 87680
rect 75177 87622 212580 87624
rect 75177 87619 75243 87622
rect 212574 87620 212580 87622
rect 212644 87620 212650 87684
rect 290733 87682 290799 87685
rect 536833 87682 536899 87685
rect 290733 87680 536899 87682
rect 290733 87624 290738 87680
rect 290794 87624 536838 87680
rect 536894 87624 536899 87680
rect 290733 87622 536899 87624
rect 290733 87619 290799 87622
rect 536833 87619 536899 87622
rect 27521 87546 27587 87549
rect 204529 87546 204595 87549
rect 27521 87544 204595 87546
rect 27521 87488 27526 87544
rect 27582 87488 204534 87544
rect 204590 87488 204595 87544
rect 27521 87486 204595 87488
rect 27521 87483 27587 87486
rect 204529 87483 204595 87486
rect 293585 87546 293651 87549
rect 554773 87546 554839 87549
rect 293585 87544 554839 87546
rect 293585 87488 293590 87544
rect 293646 87488 554778 87544
rect 554834 87488 554839 87544
rect 293585 87486 554839 87488
rect 293585 87483 293651 87486
rect 554773 87483 554839 87486
rect 281206 86260 281212 86324
rect 281276 86322 281282 86324
rect 472617 86322 472683 86325
rect 281276 86320 472683 86322
rect 281276 86264 472622 86320
rect 472678 86264 472683 86320
rect 281276 86262 472683 86264
rect 281276 86260 281282 86262
rect 472617 86259 472683 86262
rect 188337 86186 188403 86189
rect 231894 86186 231900 86188
rect 188337 86184 231900 86186
rect 188337 86128 188342 86184
rect 188398 86128 231900 86184
rect 188337 86126 231900 86128
rect 188337 86123 188403 86126
rect 231894 86124 231900 86126
rect 231964 86124 231970 86188
rect 296437 86186 296503 86189
rect 575565 86186 575631 86189
rect 296437 86184 575631 86186
rect 296437 86128 296442 86184
rect 296498 86128 575570 86184
rect 575626 86128 575631 86184
rect 296437 86126 575631 86128
rect 296437 86123 296503 86126
rect 575565 86123 575631 86126
rect 582649 86186 582715 86189
rect 583520 86186 584960 86276
rect 582649 86184 584960 86186
rect 582649 86128 582654 86184
rect 582710 86128 584960 86184
rect 582649 86126 584960 86128
rect 582649 86123 582715 86126
rect 583520 86036 584960 86126
rect 83457 84962 83523 84965
rect 213862 84962 213868 84964
rect 83457 84960 213868 84962
rect 83457 84904 83462 84960
rect 83518 84904 213868 84960
rect 83457 84902 213868 84904
rect 83457 84899 83523 84902
rect 213862 84900 213868 84902
rect 213932 84900 213938 84964
rect 259126 84900 259132 84964
rect 259196 84962 259202 84964
rect 342253 84962 342319 84965
rect 259196 84960 342319 84962
rect 259196 84904 342258 84960
rect 342314 84904 342319 84960
rect 259196 84902 342319 84904
rect 259196 84900 259202 84902
rect 342253 84899 342319 84902
rect 57881 84826 57947 84829
rect 209814 84826 209820 84828
rect 57881 84824 209820 84826
rect -960 84690 480 84780
rect 57881 84768 57886 84824
rect 57942 84768 209820 84824
rect 57881 84766 209820 84768
rect 57881 84763 57947 84766
rect 209814 84764 209820 84766
rect 209884 84764 209890 84828
rect 267406 84764 267412 84828
rect 267476 84826 267482 84828
rect 391933 84826 391999 84829
rect 267476 84824 391999 84826
rect 267476 84768 391938 84824
rect 391994 84768 391999 84824
rect 267476 84766 391999 84768
rect 267476 84764 267482 84766
rect 391933 84763 391999 84766
rect 3141 84690 3207 84693
rect -960 84688 3207 84690
rect -960 84632 3146 84688
rect 3202 84632 3207 84688
rect -960 84630 3207 84632
rect -960 84540 480 84630
rect 3141 84627 3207 84630
rect 273110 83540 273116 83604
rect 273180 83602 273186 83604
rect 423765 83602 423831 83605
rect 273180 83600 423831 83602
rect 273180 83544 423770 83600
rect 423826 83544 423831 83600
rect 273180 83542 423831 83544
rect 273180 83540 273186 83542
rect 423765 83539 423831 83542
rect 133229 83466 133295 83469
rect 222326 83466 222332 83468
rect 133229 83464 222332 83466
rect 133229 83408 133234 83464
rect 133290 83408 222332 83464
rect 133229 83406 222332 83408
rect 133229 83403 133295 83406
rect 222326 83404 222332 83406
rect 222396 83404 222402 83468
rect 275318 83404 275324 83468
rect 275388 83466 275394 83468
rect 441613 83466 441679 83469
rect 275388 83464 441679 83466
rect 275388 83408 441618 83464
rect 441674 83408 441679 83464
rect 275388 83406 441679 83408
rect 275388 83404 275394 83406
rect 441613 83403 441679 83406
rect 35249 82106 35315 82109
rect 204437 82106 204503 82109
rect 35249 82104 204503 82106
rect 35249 82048 35254 82104
rect 35310 82048 204442 82104
rect 204498 82048 204503 82104
rect 35249 82046 204503 82048
rect 35249 82043 35315 82046
rect 204437 82043 204503 82046
rect 253606 82044 253612 82108
rect 253676 82106 253682 82108
rect 311893 82106 311959 82109
rect 253676 82104 311959 82106
rect 253676 82048 311898 82104
rect 311954 82048 311959 82104
rect 253676 82046 311959 82048
rect 253676 82044 253682 82046
rect 311893 82043 311959 82046
rect 233877 81562 233943 81565
rect 237598 81562 237604 81564
rect 233877 81560 237604 81562
rect 233877 81504 233882 81560
rect 233938 81504 237604 81560
rect 233877 81502 237604 81504
rect 233877 81499 233943 81502
rect 237598 81500 237604 81502
rect 237668 81500 237674 81564
rect 294965 80882 295031 80885
rect 522297 80882 522363 80885
rect 294965 80880 522363 80882
rect 294965 80824 294970 80880
rect 295026 80824 522302 80880
rect 522358 80824 522363 80880
rect 294965 80822 522363 80824
rect 294965 80819 295031 80822
rect 522297 80819 522363 80822
rect 49601 80746 49667 80749
rect 208342 80746 208348 80748
rect 49601 80744 208348 80746
rect 49601 80688 49606 80744
rect 49662 80688 208348 80744
rect 49601 80686 208348 80688
rect 49601 80683 49667 80686
rect 208342 80684 208348 80686
rect 208412 80684 208418 80748
rect 250846 80684 250852 80748
rect 250916 80746 250922 80748
rect 296069 80746 296135 80749
rect 250916 80744 296135 80746
rect 250916 80688 296074 80744
rect 296130 80688 296135 80744
rect 250916 80686 296135 80688
rect 250916 80684 250922 80686
rect 296069 80683 296135 80686
rect 297909 80746 297975 80749
rect 579613 80746 579679 80749
rect 297909 80744 579679 80746
rect 297909 80688 297914 80744
rect 297970 80688 579618 80744
rect 579674 80688 579679 80744
rect 297909 80686 579679 80688
rect 297909 80683 297975 80686
rect 579613 80683 579679 80686
rect 259310 79596 259316 79660
rect 259380 79658 259386 79660
rect 327717 79658 327783 79661
rect 259380 79656 327783 79658
rect 259380 79600 327722 79656
rect 327778 79600 327783 79656
rect 259380 79598 327783 79600
rect 259380 79596 259386 79598
rect 327717 79595 327783 79598
rect 122741 79522 122807 79525
rect 220854 79522 220860 79524
rect 122741 79520 220860 79522
rect 122741 79464 122746 79520
rect 122802 79464 220860 79520
rect 122741 79462 220860 79464
rect 122741 79459 122807 79462
rect 220854 79460 220860 79462
rect 220924 79460 220930 79524
rect 263174 79460 263180 79524
rect 263244 79522 263250 79524
rect 363597 79522 363663 79525
rect 263244 79520 363663 79522
rect 263244 79464 363602 79520
rect 363658 79464 363663 79520
rect 263244 79462 363663 79464
rect 263244 79460 263250 79462
rect 363597 79459 363663 79462
rect 101489 79386 101555 79389
rect 211654 79386 211660 79388
rect 101489 79384 211660 79386
rect 101489 79328 101494 79384
rect 101550 79328 211660 79384
rect 101489 79326 211660 79328
rect 101489 79323 101555 79326
rect 211654 79324 211660 79326
rect 211724 79324 211730 79388
rect 278630 79324 278636 79388
rect 278700 79386 278706 79388
rect 450537 79386 450603 79389
rect 278700 79384 450603 79386
rect 278700 79328 450542 79384
rect 450598 79328 450603 79384
rect 278700 79326 450603 79328
rect 278700 79324 278706 79326
rect 450537 79323 450603 79326
rect 267590 78100 267596 78164
rect 267660 78162 267666 78164
rect 393313 78162 393379 78165
rect 267660 78160 393379 78162
rect 267660 78104 393318 78160
rect 393374 78104 393379 78160
rect 267660 78102 393379 78104
rect 267660 78100 267666 78102
rect 393313 78099 393379 78102
rect 271638 77964 271644 78028
rect 271708 78026 271714 78028
rect 415393 78026 415459 78029
rect 271708 78024 415459 78026
rect 271708 77968 415398 78024
rect 415454 77968 415459 78024
rect 271708 77966 415459 77968
rect 271708 77964 271714 77966
rect 415393 77963 415459 77966
rect 114461 77890 114527 77893
rect 219198 77890 219204 77892
rect 114461 77888 219204 77890
rect 114461 77832 114466 77888
rect 114522 77832 219204 77888
rect 114461 77830 219204 77832
rect 114461 77827 114527 77830
rect 219198 77828 219204 77830
rect 219268 77828 219274 77892
rect 277158 77828 277164 77892
rect 277228 77890 277234 77892
rect 447777 77890 447843 77893
rect 277228 77888 447843 77890
rect 277228 77832 447782 77888
rect 447838 77832 447843 77888
rect 277228 77830 447843 77832
rect 277228 77828 277234 77830
rect 447777 77827 447843 77830
rect 255078 76740 255084 76804
rect 255148 76802 255154 76804
rect 316677 76802 316743 76805
rect 255148 76800 316743 76802
rect 255148 76744 316682 76800
rect 316738 76744 316743 76800
rect 255148 76742 316743 76744
rect 255148 76740 255154 76742
rect 316677 76739 316743 76742
rect 268878 76604 268884 76668
rect 268948 76666 268954 76668
rect 403065 76666 403131 76669
rect 268948 76664 403131 76666
rect 268948 76608 403070 76664
rect 403126 76608 403131 76664
rect 268948 76606 403131 76608
rect 268948 76604 268954 76606
rect 403065 76603 403131 76606
rect 270350 76468 270356 76532
rect 270420 76530 270426 76532
rect 409965 76530 410031 76533
rect 270420 76528 410031 76530
rect 270420 76472 409970 76528
rect 410026 76472 410031 76528
rect 270420 76470 410031 76472
rect 270420 76468 270426 76470
rect 409965 76467 410031 76470
rect 266118 75244 266124 75308
rect 266188 75306 266194 75308
rect 385033 75306 385099 75309
rect 266188 75304 385099 75306
rect 266188 75248 385038 75304
rect 385094 75248 385099 75304
rect 266188 75246 385099 75248
rect 266188 75244 266194 75246
rect 385033 75243 385099 75246
rect 286910 75108 286916 75172
rect 286980 75170 286986 75172
rect 517605 75170 517671 75173
rect 286980 75168 517671 75170
rect 286980 75112 517610 75168
rect 517666 75112 517671 75168
rect 286980 75110 517671 75112
rect 286980 75108 286986 75110
rect 517605 75107 517671 75110
rect 92381 73946 92447 73949
rect 215334 73946 215340 73948
rect 92381 73944 215340 73946
rect 92381 73888 92386 73944
rect 92442 73888 215340 73944
rect 92381 73886 215340 73888
rect 92381 73883 92447 73886
rect 215334 73884 215340 73886
rect 215404 73884 215410 73948
rect 35801 73810 35867 73813
rect 205582 73810 205588 73812
rect 35801 73808 205588 73810
rect 35801 73752 35806 73808
rect 35862 73752 205588 73808
rect 35801 73750 205588 73752
rect 35801 73747 35867 73750
rect 205582 73748 205588 73750
rect 205652 73748 205658 73812
rect 257286 73748 257292 73812
rect 257356 73810 257362 73812
rect 326337 73810 326403 73813
rect 257356 73808 326403 73810
rect 257356 73752 326342 73808
rect 326398 73752 326403 73808
rect 257356 73750 326403 73752
rect 257356 73748 257362 73750
rect 326337 73747 326403 73750
rect 583753 73266 583819 73269
rect 583710 73264 583819 73266
rect 583710 73208 583758 73264
rect 583814 73208 583819 73264
rect 583710 73203 583819 73208
rect 583710 73130 583770 73203
rect 583342 73084 583770 73130
rect 583342 73070 584960 73084
rect 583342 72994 583402 73070
rect 583520 72994 584960 73070
rect 583342 72934 584960 72994
rect 583520 72844 584960 72934
rect 260598 72388 260604 72452
rect 260668 72450 260674 72452
rect 353293 72450 353359 72453
rect 260668 72448 353359 72450
rect 260668 72392 353298 72448
rect 353354 72392 353359 72448
rect 260668 72390 353359 72392
rect 260668 72388 260674 72390
rect 353293 72387 353359 72390
rect -960 71634 480 71724
rect 3417 71634 3483 71637
rect -960 71632 3483 71634
rect -960 71576 3422 71632
rect 3478 71576 3483 71632
rect -960 71574 3483 71576
rect -960 71484 480 71574
rect 3417 71571 3483 71574
rect 264646 71164 264652 71228
rect 264716 71226 264722 71228
rect 373993 71226 374059 71229
rect 264716 71224 374059 71226
rect 264716 71168 373998 71224
rect 374054 71168 374059 71224
rect 264716 71166 374059 71168
rect 264716 71164 264722 71166
rect 373993 71163 374059 71166
rect 288198 71028 288204 71092
rect 288268 71090 288274 71092
rect 514753 71090 514819 71093
rect 288268 71088 514819 71090
rect 288268 71032 514758 71088
rect 514814 71032 514819 71088
rect 288268 71030 514819 71032
rect 288268 71028 288274 71030
rect 514753 71027 514819 71030
rect 249558 62732 249564 62796
rect 249628 62794 249634 62796
rect 275277 62794 275343 62797
rect 249628 62792 275343 62794
rect 249628 62736 275282 62792
rect 275338 62736 275343 62792
rect 249628 62734 275343 62736
rect 249628 62732 249634 62734
rect 275277 62731 275343 62734
rect 583661 60210 583727 60213
rect 583526 60208 583727 60210
rect 583526 60152 583666 60208
rect 583722 60152 583727 60208
rect 583526 60150 583727 60152
rect 583526 59802 583586 60150
rect 583661 60147 583727 60150
rect 583342 59756 583586 59802
rect 583342 59742 584960 59756
rect 583342 59666 583402 59742
rect 583520 59666 584960 59742
rect 583342 59606 584960 59666
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 3049 58578 3115 58581
rect -960 58576 3115 58578
rect -960 58520 3054 58576
rect 3110 58520 3115 58576
rect -960 58518 3115 58520
rect -960 58428 480 58518
rect 3049 58515 3115 58518
rect 299238 50220 299244 50284
rect 299308 50282 299314 50284
rect 582373 50282 582439 50285
rect 299308 50280 582439 50282
rect 299308 50224 582378 50280
rect 582434 50224 582439 50280
rect 299308 50222 582439 50224
rect 299308 50220 299314 50222
rect 582373 50219 582439 50222
rect 583569 46882 583635 46885
rect 583526 46880 583635 46882
rect 583526 46824 583574 46880
rect 583630 46824 583635 46880
rect 583526 46819 583635 46824
rect 583526 46474 583586 46819
rect 583342 46428 583586 46474
rect 583342 46414 584960 46428
rect 583342 46338 583402 46414
rect 583520 46338 584960 46414
rect 583342 46278 584960 46338
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 3417 45522 3483 45525
rect -960 45520 3483 45522
rect -960 45464 3422 45520
rect 3478 45464 3483 45520
rect -960 45462 3483 45464
rect -960 45372 480 45462
rect 3417 45459 3483 45462
rect 107561 44842 107627 44845
rect 218646 44842 218652 44844
rect 107561 44840 218652 44842
rect 107561 44784 107566 44840
rect 107622 44784 218652 44840
rect 107561 44782 218652 44784
rect 107561 44779 107627 44782
rect 218646 44780 218652 44782
rect 218716 44780 218722 44844
rect 583520 33146 584960 33236
rect 583342 33086 584960 33146
rect 583342 33010 583402 33086
rect 583520 33010 584960 33086
rect 583342 32996 584960 33010
rect 583342 32950 583770 32996
rect 583710 32874 583770 32950
rect 583845 32874 583911 32877
rect 583710 32872 583911 32874
rect 583710 32816 583850 32872
rect 583906 32816 583911 32872
rect 583710 32814 583911 32816
rect 583845 32811 583911 32814
rect -960 32466 480 32556
rect 2865 32466 2931 32469
rect -960 32464 2931 32466
rect -960 32408 2870 32464
rect 2926 32408 2931 32464
rect -960 32406 2931 32408
rect -960 32316 480 32406
rect 2865 32403 2931 32406
rect 263358 30908 263364 30972
rect 263428 30970 263434 30972
rect 367737 30970 367803 30973
rect 263428 30968 367803 30970
rect 263428 30912 367742 30968
rect 367798 30912 367803 30968
rect 263428 30910 367803 30912
rect 263428 30908 263434 30910
rect 367737 30907 367803 30910
rect 582465 19818 582531 19821
rect 583520 19818 584960 19908
rect 582465 19816 584960 19818
rect 582465 19760 582470 19816
rect 582526 19760 584960 19816
rect 582465 19758 584960 19760
rect 582465 19755 582531 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3417 19410 3483 19413
rect -960 19408 3483 19410
rect -960 19352 3422 19408
rect 3478 19352 3483 19408
rect -960 19350 3483 19352
rect -960 19260 480 19350
rect 3417 19347 3483 19350
rect 256550 11868 256556 11932
rect 256620 11930 256626 11932
rect 326337 11930 326403 11933
rect 256620 11928 326403 11930
rect 256620 11872 326342 11928
rect 326398 11872 326403 11928
rect 256620 11870 326403 11872
rect 256620 11868 256626 11870
rect 326337 11867 326403 11870
rect 274398 11732 274404 11796
rect 274468 11794 274474 11796
rect 432505 11794 432571 11797
rect 274468 11792 432571 11794
rect 274468 11736 432510 11792
rect 432566 11736 432571 11792
rect 274468 11734 432571 11736
rect 274468 11732 274474 11734
rect 432505 11731 432571 11734
rect 292430 11596 292436 11660
rect 292500 11658 292506 11660
rect 545481 11658 545547 11661
rect 292500 11656 545547 11658
rect 292500 11600 545486 11656
rect 545542 11600 545547 11656
rect 292500 11598 545547 11600
rect 292500 11596 292506 11598
rect 545481 11595 545547 11598
rect 583569 6898 583635 6901
rect 583526 6896 583635 6898
rect 583526 6840 583574 6896
rect 583630 6840 583635 6896
rect 583526 6835 583635 6840
rect 583526 6762 583586 6835
rect 583342 6716 583586 6762
rect 583342 6702 584960 6716
rect 583342 6626 583402 6702
rect 583520 6626 584960 6702
rect -960 6490 480 6580
rect 583342 6566 584960 6626
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect 583520 6476 584960 6566
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
rect 246798 6156 246804 6220
rect 246868 6218 246874 6220
rect 273621 6218 273687 6221
rect 246868 6216 273687 6218
rect 246868 6160 273626 6216
rect 273682 6160 273687 6216
rect 246868 6158 273687 6160
rect 246868 6156 246874 6158
rect 273621 6155 273687 6158
rect 281390 4796 281396 4860
rect 281460 4858 281466 4860
rect 474549 4858 474615 4861
rect 281460 4856 474615 4858
rect 281460 4800 474554 4856
rect 474610 4800 474615 4856
rect 281460 4798 474615 4800
rect 281460 4796 281466 4798
rect 474549 4795 474615 4798
rect 582189 3634 582255 3637
rect 582925 3634 582991 3637
rect 582189 3632 582991 3634
rect 582189 3576 582194 3632
rect 582250 3576 582930 3632
rect 582986 3576 582991 3632
rect 582189 3574 582991 3576
rect 582189 3571 582255 3574
rect 582925 3571 582991 3574
rect 15929 3498 15995 3501
rect 201953 3498 202019 3501
rect 15929 3496 202019 3498
rect 15929 3440 15934 3496
rect 15990 3440 201958 3496
rect 202014 3440 202019 3496
rect 15929 3438 202019 3440
rect 15929 3435 15995 3438
rect 201953 3435 202019 3438
rect 580993 3498 581059 3501
rect 582649 3498 582715 3501
rect 580993 3496 582715 3498
rect 580993 3440 580998 3496
rect 581054 3440 582654 3496
rect 582710 3440 582715 3496
rect 580993 3438 582715 3440
rect 580993 3435 581059 3438
rect 582649 3435 582715 3438
rect 202689 3362 202755 3365
rect 235257 3362 235323 3365
rect 202689 3360 235323 3362
rect 202689 3304 202694 3360
rect 202750 3304 235262 3360
rect 235318 3304 235323 3360
rect 202689 3302 235323 3304
rect 202689 3299 202755 3302
rect 235257 3299 235323 3302
rect 255957 3362 256023 3365
rect 285397 3362 285463 3365
rect 255957 3360 285463 3362
rect 255957 3304 255962 3360
rect 256018 3304 285402 3360
rect 285458 3304 285463 3360
rect 255957 3302 285463 3304
rect 255957 3299 256023 3302
rect 285397 3299 285463 3302
rect 568021 3362 568087 3365
rect 579613 3362 579679 3365
rect 568021 3360 579679 3362
rect 568021 3304 568026 3360
rect 568082 3304 579618 3360
rect 579674 3304 579679 3360
rect 568021 3302 579679 3304
rect 568021 3299 568087 3302
rect 579613 3299 579679 3302
rect 252318 1940 252324 2004
rect 252388 2002 252394 2004
rect 305545 2002 305611 2005
rect 252388 2000 305611 2002
rect 252388 1944 305550 2000
rect 305606 1944 305611 2000
rect 252388 1942 305611 1944
rect 252388 1940 252394 1942
rect 305545 1939 305611 1942
<< via3 >>
rect 298140 102172 298204 102236
rect 297956 100328 298020 100332
rect 297956 100272 297970 100328
rect 297970 100272 298020 100328
rect 297956 100268 298020 100272
rect 219388 97548 219452 97612
rect 292436 97276 292500 97340
rect 271460 97140 271524 97204
rect 252508 97004 252572 97068
rect 259316 97004 259380 97068
rect 260604 97004 260668 97068
rect 264468 97004 264532 97068
rect 267412 97064 267476 97068
rect 267412 97008 267462 97064
rect 267462 97008 267476 97064
rect 267412 97004 267476 97008
rect 273116 97004 273180 97068
rect 274220 97004 274284 97068
rect 275324 97004 275388 97068
rect 279004 97004 279068 97068
rect 202828 96868 202892 96932
rect 205956 96928 206020 96932
rect 205956 96872 205970 96928
rect 205970 96872 206020 96928
rect 205956 96868 206020 96872
rect 215340 96868 215404 96932
rect 216628 96928 216692 96932
rect 216628 96872 216678 96928
rect 216678 96872 216692 96928
rect 216628 96868 216692 96872
rect 218652 96868 218716 96932
rect 220860 96868 220924 96932
rect 222332 96928 222396 96932
rect 222332 96872 222382 96928
rect 222382 96872 222396 96928
rect 222332 96868 222396 96872
rect 223620 96928 223684 96932
rect 223620 96872 223634 96928
rect 223634 96872 223684 96928
rect 223620 96868 223684 96872
rect 237604 96928 237668 96932
rect 237604 96872 237618 96928
rect 237618 96872 237668 96928
rect 237604 96868 237668 96872
rect 246804 96868 246868 96932
rect 249564 96928 249628 96932
rect 249564 96872 249578 96928
rect 249578 96872 249628 96928
rect 249564 96868 249628 96872
rect 250852 96868 250916 96932
rect 252324 96928 252388 96932
rect 252324 96872 252374 96928
rect 252374 96872 252388 96928
rect 252324 96868 252388 96872
rect 253612 96928 253676 96932
rect 253612 96872 253662 96928
rect 253662 96872 253676 96928
rect 253612 96868 253676 96872
rect 255084 96868 255148 96932
rect 256556 96868 256620 96932
rect 257292 96868 257356 96932
rect 259132 96868 259196 96932
rect 260420 96868 260484 96932
rect 263180 96868 263244 96932
rect 263364 96928 263428 96932
rect 263364 96872 263378 96928
rect 263378 96872 263428 96928
rect 263364 96868 263428 96872
rect 264652 96868 264716 96932
rect 266124 96928 266188 96932
rect 266124 96872 266174 96928
rect 266174 96872 266188 96928
rect 266124 96868 266188 96872
rect 267596 96928 267660 96932
rect 267596 96872 267646 96928
rect 267646 96872 267660 96928
rect 267596 96868 267660 96872
rect 268884 96868 268948 96932
rect 270356 96868 270420 96932
rect 271644 96868 271708 96932
rect 274404 96868 274468 96932
rect 277164 96868 277228 96932
rect 278636 96928 278700 96932
rect 278636 96872 278650 96928
rect 278650 96872 278700 96928
rect 278636 96868 278700 96872
rect 281212 96928 281276 96932
rect 281212 96872 281226 96928
rect 281226 96872 281276 96928
rect 281212 96868 281276 96872
rect 281396 96928 281460 96932
rect 281396 96872 281446 96928
rect 281446 96872 281460 96928
rect 281396 96868 281460 96872
rect 282132 96868 282196 96932
rect 284156 96868 284220 96932
rect 286916 96928 286980 96932
rect 286916 96872 286930 96928
rect 286930 96872 286980 96928
rect 286916 96868 286980 96872
rect 288204 96868 288268 96932
rect 292252 96868 292316 96932
rect 295012 96928 295076 96932
rect 295012 96872 295026 96928
rect 295026 96872 295076 96928
rect 295012 96868 295076 96872
rect 295196 96928 295260 96932
rect 295196 96872 295246 96928
rect 295246 96872 295260 96928
rect 295196 96868 295260 96872
rect 299244 96928 299308 96932
rect 299244 96872 299294 96928
rect 299294 96872 299308 96928
rect 299244 96868 299308 96872
rect 230612 96732 230676 96796
rect 204300 96656 204364 96660
rect 204300 96600 204350 96656
rect 204350 96600 204364 96656
rect 204300 96596 204364 96600
rect 205772 96656 205836 96660
rect 205772 96600 205786 96656
rect 205786 96600 205836 96656
rect 205772 96596 205836 96600
rect 208348 96656 208412 96660
rect 208348 96600 208398 96656
rect 208398 96600 208412 96656
rect 208348 96596 208412 96600
rect 209820 96656 209884 96660
rect 209820 96600 209834 96656
rect 209834 96600 209884 96656
rect 209820 96596 209884 96600
rect 211660 96596 211724 96660
rect 212580 96656 212644 96660
rect 212580 96600 212630 96656
rect 212630 96600 212644 96656
rect 212580 96596 212644 96600
rect 213868 96596 213932 96660
rect 226380 96656 226444 96660
rect 226380 96600 226430 96656
rect 226430 96600 226444 96656
rect 226380 96596 226444 96600
rect 230428 96596 230492 96660
rect 231900 96596 231964 96660
rect 233188 96596 233252 96660
rect 271460 95780 271524 95844
rect 230428 94692 230492 94756
rect 252508 94556 252572 94620
rect 226380 94420 226444 94484
rect 223620 93332 223684 93396
rect 260420 93332 260484 93396
rect 205772 93196 205836 93260
rect 284156 93196 284220 93260
rect 204300 93060 204364 93124
rect 295012 93060 295076 93124
rect 230612 91836 230676 91900
rect 202828 91700 202892 91764
rect 264468 91700 264532 91764
rect 282132 91156 282196 91220
rect 274220 90476 274284 90540
rect 233188 90340 233252 90404
rect 216628 89116 216692 89180
rect 279004 89116 279068 89180
rect 295196 88980 295260 89044
rect 292252 87756 292316 87820
rect 212580 87620 212644 87684
rect 281212 86260 281276 86324
rect 231900 86124 231964 86188
rect 213868 84900 213932 84964
rect 259132 84900 259196 84964
rect 209820 84764 209884 84828
rect 267412 84764 267476 84828
rect 273116 83540 273180 83604
rect 222332 83404 222396 83468
rect 275324 83404 275388 83468
rect 253612 82044 253676 82108
rect 237604 81500 237668 81564
rect 208348 80684 208412 80748
rect 250852 80684 250916 80748
rect 259316 79596 259380 79660
rect 220860 79460 220924 79524
rect 263180 79460 263244 79524
rect 211660 79324 211724 79388
rect 278636 79324 278700 79388
rect 267596 78100 267660 78164
rect 271644 77964 271708 78028
rect 219204 77828 219268 77892
rect 277164 77828 277228 77892
rect 255084 76740 255148 76804
rect 268884 76604 268948 76668
rect 270356 76468 270420 76532
rect 266124 75244 266188 75308
rect 286916 75108 286980 75172
rect 215340 73884 215404 73948
rect 205588 73748 205652 73812
rect 257292 73748 257356 73812
rect 260604 72388 260668 72452
rect 264652 71164 264716 71228
rect 288204 71028 288268 71092
rect 249564 62732 249628 62796
rect 299244 50220 299308 50284
rect 218652 44780 218716 44844
rect 263364 30908 263428 30972
rect 256556 11868 256620 11932
rect 274404 11732 274468 11796
rect 292436 11596 292500 11660
rect 246804 6156 246868 6220
rect 281396 4796 281460 4860
rect 252324 1940 252388 2004
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 680614 -8106 711002
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 -8106 680614
rect -8726 680294 -8106 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 -8106 680294
rect -8726 644614 -8106 680058
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 -8106 644614
rect -8726 644294 -8106 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 -8106 644294
rect -8726 608614 -8106 644058
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 -8106 608614
rect -8726 608294 -8106 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 -8106 608294
rect -8726 572614 -8106 608058
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 -8106 572614
rect -8726 572294 -8106 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 -8106 572294
rect -8726 536614 -8106 572058
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 -8106 536614
rect -8726 536294 -8106 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 -8106 536294
rect -8726 500614 -8106 536058
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 -8106 500614
rect -8726 500294 -8106 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 -8106 500294
rect -8726 464614 -8106 500058
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 -8106 464614
rect -8726 464294 -8106 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 -8106 464294
rect -8726 428614 -8106 464058
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 -8106 428614
rect -8726 428294 -8106 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 -8106 428294
rect -8726 392614 -8106 428058
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 -8106 392614
rect -8726 392294 -8106 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 -8106 392294
rect -8726 356614 -8106 392058
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 -8106 356614
rect -8726 356294 -8106 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 -8106 356294
rect -8726 320614 -8106 356058
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 -8106 320614
rect -8726 320294 -8106 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 -8106 320294
rect -8726 284614 -8106 320058
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 -8106 284614
rect -8726 284294 -8106 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 -8106 284294
rect -8726 248614 -8106 284058
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 -8106 248614
rect -8726 248294 -8106 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 -8106 248294
rect -8726 212614 -8106 248058
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 -8106 212614
rect -8726 212294 -8106 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 -8106 212294
rect -8726 176614 -8106 212058
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 -8106 176614
rect -8726 176294 -8106 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 -8106 176294
rect -8726 140614 -8106 176058
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 -8106 140614
rect -8726 140294 -8106 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 -8106 140294
rect -8726 104614 -8106 140058
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 -8106 104614
rect -8726 104294 -8106 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 -8106 104294
rect -8726 68614 -8106 104058
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 -8106 68614
rect -8726 68294 -8106 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 -8106 68294
rect -8726 32614 -8106 68058
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 -8106 32614
rect -8726 32294 -8106 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 -8106 32294
rect -8726 -7066 -8106 32058
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 698614 -7146 710042
rect 12954 710598 13574 711590
rect 12954 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 13574 710598
rect 12954 710278 13574 710362
rect 12954 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 13574 710278
rect -7766 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 -7146 698614
rect -7766 698294 -7146 698378
rect -7766 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 -7146 698294
rect -7766 662614 -7146 698058
rect -7766 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 -7146 662614
rect -7766 662294 -7146 662378
rect -7766 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 -7146 662294
rect -7766 626614 -7146 662058
rect -7766 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 -7146 626614
rect -7766 626294 -7146 626378
rect -7766 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 -7146 626294
rect -7766 590614 -7146 626058
rect -7766 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 -7146 590614
rect -7766 590294 -7146 590378
rect -7766 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 -7146 590294
rect -7766 554614 -7146 590058
rect -7766 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 -7146 554614
rect -7766 554294 -7146 554378
rect -7766 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 -7146 554294
rect -7766 518614 -7146 554058
rect -7766 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 -7146 518614
rect -7766 518294 -7146 518378
rect -7766 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 -7146 518294
rect -7766 482614 -7146 518058
rect -7766 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 -7146 482614
rect -7766 482294 -7146 482378
rect -7766 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 -7146 482294
rect -7766 446614 -7146 482058
rect -7766 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 -7146 446614
rect -7766 446294 -7146 446378
rect -7766 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 -7146 446294
rect -7766 410614 -7146 446058
rect -7766 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 -7146 410614
rect -7766 410294 -7146 410378
rect -7766 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 -7146 410294
rect -7766 374614 -7146 410058
rect -7766 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 -7146 374614
rect -7766 374294 -7146 374378
rect -7766 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 -7146 374294
rect -7766 338614 -7146 374058
rect -7766 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 -7146 338614
rect -7766 338294 -7146 338378
rect -7766 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 -7146 338294
rect -7766 302614 -7146 338058
rect -7766 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 -7146 302614
rect -7766 302294 -7146 302378
rect -7766 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 -7146 302294
rect -7766 266614 -7146 302058
rect -7766 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 -7146 266614
rect -7766 266294 -7146 266378
rect -7766 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 -7146 266294
rect -7766 230614 -7146 266058
rect -7766 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 -7146 230614
rect -7766 230294 -7146 230378
rect -7766 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 -7146 230294
rect -7766 194614 -7146 230058
rect -7766 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 -7146 194614
rect -7766 194294 -7146 194378
rect -7766 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 -7146 194294
rect -7766 158614 -7146 194058
rect -7766 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 -7146 158614
rect -7766 158294 -7146 158378
rect -7766 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 -7146 158294
rect -7766 122614 -7146 158058
rect -7766 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 -7146 122614
rect -7766 122294 -7146 122378
rect -7766 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 -7146 122294
rect -7766 86614 -7146 122058
rect -7766 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 -7146 86614
rect -7766 86294 -7146 86378
rect -7766 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 -7146 86294
rect -7766 50614 -7146 86058
rect -7766 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 -7146 50614
rect -7766 50294 -7146 50378
rect -7766 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 -7146 50294
rect -7766 14614 -7146 50058
rect -7766 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 -7146 14614
rect -7766 14294 -7146 14378
rect -7766 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 -7146 14294
rect -7766 -6106 -7146 14058
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 676894 -6186 709082
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 -6186 676894
rect -6806 676574 -6186 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 -6186 676574
rect -6806 640894 -6186 676338
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 -6186 640894
rect -6806 640574 -6186 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 -6186 640574
rect -6806 604894 -6186 640338
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 -6186 604894
rect -6806 604574 -6186 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 -6186 604574
rect -6806 568894 -6186 604338
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 -6186 568894
rect -6806 568574 -6186 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 -6186 568574
rect -6806 532894 -6186 568338
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 -6186 532894
rect -6806 532574 -6186 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 -6186 532574
rect -6806 496894 -6186 532338
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 -6186 496894
rect -6806 496574 -6186 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 -6186 496574
rect -6806 460894 -6186 496338
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 -6186 460894
rect -6806 460574 -6186 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 -6186 460574
rect -6806 424894 -6186 460338
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 -6186 424894
rect -6806 424574 -6186 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 -6186 424574
rect -6806 388894 -6186 424338
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 -6186 388894
rect -6806 388574 -6186 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 -6186 388574
rect -6806 352894 -6186 388338
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 -6186 352894
rect -6806 352574 -6186 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 -6186 352574
rect -6806 316894 -6186 352338
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 -6186 316894
rect -6806 316574 -6186 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 -6186 316574
rect -6806 280894 -6186 316338
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 -6186 280894
rect -6806 280574 -6186 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 -6186 280574
rect -6806 244894 -6186 280338
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 -6186 244894
rect -6806 244574 -6186 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 -6186 244574
rect -6806 208894 -6186 244338
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 -6186 208894
rect -6806 208574 -6186 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 -6186 208574
rect -6806 172894 -6186 208338
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 -6186 172894
rect -6806 172574 -6186 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 -6186 172574
rect -6806 136894 -6186 172338
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 -6186 136894
rect -6806 136574 -6186 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 -6186 136574
rect -6806 100894 -6186 136338
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 -6186 100894
rect -6806 100574 -6186 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 -6186 100574
rect -6806 64894 -6186 100338
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 -6186 64894
rect -6806 64574 -6186 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 -6186 64574
rect -6806 28894 -6186 64338
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 -6186 28894
rect -6806 28574 -6186 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 -6186 28574
rect -6806 -5146 -6186 28338
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 694894 -5226 708122
rect 9234 708678 9854 709670
rect 9234 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 9854 708678
rect 9234 708358 9854 708442
rect 9234 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 9854 708358
rect -5846 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 -5226 694894
rect -5846 694574 -5226 694658
rect -5846 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 -5226 694574
rect -5846 658894 -5226 694338
rect -5846 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 -5226 658894
rect -5846 658574 -5226 658658
rect -5846 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 -5226 658574
rect -5846 622894 -5226 658338
rect -5846 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 -5226 622894
rect -5846 622574 -5226 622658
rect -5846 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 -5226 622574
rect -5846 586894 -5226 622338
rect -5846 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 -5226 586894
rect -5846 586574 -5226 586658
rect -5846 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 -5226 586574
rect -5846 550894 -5226 586338
rect -5846 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 -5226 550894
rect -5846 550574 -5226 550658
rect -5846 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 -5226 550574
rect -5846 514894 -5226 550338
rect -5846 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 -5226 514894
rect -5846 514574 -5226 514658
rect -5846 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 -5226 514574
rect -5846 478894 -5226 514338
rect -5846 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 -5226 478894
rect -5846 478574 -5226 478658
rect -5846 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 -5226 478574
rect -5846 442894 -5226 478338
rect -5846 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 -5226 442894
rect -5846 442574 -5226 442658
rect -5846 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 -5226 442574
rect -5846 406894 -5226 442338
rect -5846 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 -5226 406894
rect -5846 406574 -5226 406658
rect -5846 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 -5226 406574
rect -5846 370894 -5226 406338
rect -5846 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 -5226 370894
rect -5846 370574 -5226 370658
rect -5846 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 -5226 370574
rect -5846 334894 -5226 370338
rect -5846 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 -5226 334894
rect -5846 334574 -5226 334658
rect -5846 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 -5226 334574
rect -5846 298894 -5226 334338
rect -5846 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 -5226 298894
rect -5846 298574 -5226 298658
rect -5846 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 -5226 298574
rect -5846 262894 -5226 298338
rect -5846 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 -5226 262894
rect -5846 262574 -5226 262658
rect -5846 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 -5226 262574
rect -5846 226894 -5226 262338
rect -5846 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 -5226 226894
rect -5846 226574 -5226 226658
rect -5846 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 -5226 226574
rect -5846 190894 -5226 226338
rect -5846 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 -5226 190894
rect -5846 190574 -5226 190658
rect -5846 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 -5226 190574
rect -5846 154894 -5226 190338
rect -5846 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 -5226 154894
rect -5846 154574 -5226 154658
rect -5846 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 -5226 154574
rect -5846 118894 -5226 154338
rect -5846 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 -5226 118894
rect -5846 118574 -5226 118658
rect -5846 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 -5226 118574
rect -5846 82894 -5226 118338
rect -5846 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 -5226 82894
rect -5846 82574 -5226 82658
rect -5846 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 -5226 82574
rect -5846 46894 -5226 82338
rect -5846 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 -5226 46894
rect -5846 46574 -5226 46658
rect -5846 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 -5226 46574
rect -5846 10894 -5226 46338
rect -5846 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 -5226 10894
rect -5846 10574 -5226 10658
rect -5846 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 -5226 10574
rect -5846 -4186 -5226 10338
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 673174 -4266 707162
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 -4266 673174
rect -4886 672854 -4266 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 -4266 672854
rect -4886 637174 -4266 672618
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 -4266 637174
rect -4886 636854 -4266 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 -4266 636854
rect -4886 601174 -4266 636618
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 -4266 601174
rect -4886 600854 -4266 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 -4266 600854
rect -4886 565174 -4266 600618
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 -4266 565174
rect -4886 564854 -4266 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 -4266 564854
rect -4886 529174 -4266 564618
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 -4266 529174
rect -4886 528854 -4266 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 -4266 528854
rect -4886 493174 -4266 528618
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 -4266 493174
rect -4886 492854 -4266 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 -4266 492854
rect -4886 457174 -4266 492618
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 -4266 457174
rect -4886 456854 -4266 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 -4266 456854
rect -4886 421174 -4266 456618
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 -4266 421174
rect -4886 420854 -4266 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 -4266 420854
rect -4886 385174 -4266 420618
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 -4266 385174
rect -4886 384854 -4266 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 -4266 384854
rect -4886 349174 -4266 384618
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 -4266 349174
rect -4886 348854 -4266 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 -4266 348854
rect -4886 313174 -4266 348618
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 -4266 313174
rect -4886 312854 -4266 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 -4266 312854
rect -4886 277174 -4266 312618
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 -4266 277174
rect -4886 276854 -4266 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 -4266 276854
rect -4886 241174 -4266 276618
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 -4266 241174
rect -4886 240854 -4266 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 -4266 240854
rect -4886 205174 -4266 240618
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 -4266 205174
rect -4886 204854 -4266 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 -4266 204854
rect -4886 169174 -4266 204618
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 -4266 169174
rect -4886 168854 -4266 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 -4266 168854
rect -4886 133174 -4266 168618
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 -4266 133174
rect -4886 132854 -4266 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 -4266 132854
rect -4886 97174 -4266 132618
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 -4266 97174
rect -4886 96854 -4266 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 -4266 96854
rect -4886 61174 -4266 96618
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 -4266 61174
rect -4886 60854 -4266 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 -4266 60854
rect -4886 25174 -4266 60618
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 -4266 25174
rect -4886 24854 -4266 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 -4266 24854
rect -4886 -3226 -4266 24618
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 691174 -3306 706202
rect 5514 706758 6134 707750
rect 5514 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 6134 706758
rect 5514 706438 6134 706522
rect 5514 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 6134 706438
rect -3926 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 -3306 691174
rect -3926 690854 -3306 690938
rect -3926 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 -3306 690854
rect -3926 655174 -3306 690618
rect -3926 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 -3306 655174
rect -3926 654854 -3306 654938
rect -3926 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 -3306 654854
rect -3926 619174 -3306 654618
rect -3926 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 -3306 619174
rect -3926 618854 -3306 618938
rect -3926 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 -3306 618854
rect -3926 583174 -3306 618618
rect -3926 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 -3306 583174
rect -3926 582854 -3306 582938
rect -3926 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 -3306 582854
rect -3926 547174 -3306 582618
rect -3926 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 -3306 547174
rect -3926 546854 -3306 546938
rect -3926 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 -3306 546854
rect -3926 511174 -3306 546618
rect -3926 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 -3306 511174
rect -3926 510854 -3306 510938
rect -3926 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 -3306 510854
rect -3926 475174 -3306 510618
rect -3926 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 -3306 475174
rect -3926 474854 -3306 474938
rect -3926 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 -3306 474854
rect -3926 439174 -3306 474618
rect -3926 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 -3306 439174
rect -3926 438854 -3306 438938
rect -3926 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 -3306 438854
rect -3926 403174 -3306 438618
rect -3926 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 -3306 403174
rect -3926 402854 -3306 402938
rect -3926 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 -3306 402854
rect -3926 367174 -3306 402618
rect -3926 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 -3306 367174
rect -3926 366854 -3306 366938
rect -3926 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 -3306 366854
rect -3926 331174 -3306 366618
rect -3926 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 -3306 331174
rect -3926 330854 -3306 330938
rect -3926 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 -3306 330854
rect -3926 295174 -3306 330618
rect -3926 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 -3306 295174
rect -3926 294854 -3306 294938
rect -3926 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 -3306 294854
rect -3926 259174 -3306 294618
rect -3926 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 -3306 259174
rect -3926 258854 -3306 258938
rect -3926 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 -3306 258854
rect -3926 223174 -3306 258618
rect -3926 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 -3306 223174
rect -3926 222854 -3306 222938
rect -3926 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 -3306 222854
rect -3926 187174 -3306 222618
rect -3926 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 -3306 187174
rect -3926 186854 -3306 186938
rect -3926 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 -3306 186854
rect -3926 151174 -3306 186618
rect -3926 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 -3306 151174
rect -3926 150854 -3306 150938
rect -3926 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 -3306 150854
rect -3926 115174 -3306 150618
rect -3926 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 -3306 115174
rect -3926 114854 -3306 114938
rect -3926 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 -3306 114854
rect -3926 79174 -3306 114618
rect -3926 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 -3306 79174
rect -3926 78854 -3306 78938
rect -3926 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 -3306 78854
rect -3926 43174 -3306 78618
rect -3926 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 -3306 43174
rect -3926 42854 -3306 42938
rect -3926 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 -3306 42854
rect -3926 7174 -3306 42618
rect -3926 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 -3306 7174
rect -3926 6854 -3306 6938
rect -3926 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 -3306 6854
rect -3926 -2266 -3306 6618
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 669454 -2346 705242
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 -2346 669454
rect -2966 669134 -2346 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 -2346 669134
rect -2966 633454 -2346 668898
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 -2346 633454
rect -2966 633134 -2346 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 -2346 633134
rect -2966 597454 -2346 632898
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 -2346 597454
rect -2966 597134 -2346 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 -2346 597134
rect -2966 561454 -2346 596898
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 -2346 561454
rect -2966 561134 -2346 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 -2346 561134
rect -2966 525454 -2346 560898
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 -2346 525454
rect -2966 525134 -2346 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 -2346 525134
rect -2966 489454 -2346 524898
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 -2346 489454
rect -2966 489134 -2346 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 -2346 489134
rect -2966 453454 -2346 488898
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 -2346 453454
rect -2966 453134 -2346 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 -2346 453134
rect -2966 417454 -2346 452898
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 -2346 417454
rect -2966 417134 -2346 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 -2346 417134
rect -2966 381454 -2346 416898
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 -2346 381454
rect -2966 381134 -2346 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 -2346 381134
rect -2966 345454 -2346 380898
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 -2346 345454
rect -2966 345134 -2346 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 -2346 345134
rect -2966 309454 -2346 344898
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 -2346 309454
rect -2966 309134 -2346 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 -2346 309134
rect -2966 273454 -2346 308898
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 -2346 273454
rect -2966 273134 -2346 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 -2346 273134
rect -2966 237454 -2346 272898
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 -2346 237454
rect -2966 237134 -2346 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 -2346 237134
rect -2966 201454 -2346 236898
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 -2346 201454
rect -2966 201134 -2346 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 -2346 201134
rect -2966 165454 -2346 200898
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 -2346 165454
rect -2966 165134 -2346 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 -2346 165134
rect -2966 129454 -2346 164898
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 -2346 129454
rect -2966 129134 -2346 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 -2346 129134
rect -2966 93454 -2346 128898
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 -2346 93454
rect -2966 93134 -2346 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 -2346 93134
rect -2966 57454 -2346 92898
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 -2346 57454
rect -2966 57134 -2346 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 -2346 57134
rect -2966 21454 -2346 56898
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 -2346 21454
rect -2966 21134 -2346 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 -2346 21134
rect -2966 -1306 -2346 20898
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 705830
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 1794 -1894 2414 -902
rect 5514 691174 6134 706202
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 5514 619174 6134 654618
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 5514 259174 6134 294618
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 5514 223174 6134 258618
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 5514 187174 6134 222618
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 5514 151174 6134 186618
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 5514 115174 6134 150618
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 5514 79174 6134 114618
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 5514 43174 6134 78618
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 5514 7174 6134 42618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect 5514 -2266 6134 6618
rect 5514 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 6134 -2266
rect 5514 -2586 6134 -2502
rect 5514 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 6134 -2586
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect 5514 -3814 6134 -2822
rect 9234 694894 9854 708122
rect 9234 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 9854 694894
rect 9234 694574 9854 694658
rect 9234 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 9854 694574
rect 9234 658894 9854 694338
rect 9234 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 9854 658894
rect 9234 658574 9854 658658
rect 9234 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 9854 658574
rect 9234 622894 9854 658338
rect 9234 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 9854 622894
rect 9234 622574 9854 622658
rect 9234 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 9854 622574
rect 9234 586894 9854 622338
rect 9234 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 9854 586894
rect 9234 586574 9854 586658
rect 9234 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 9854 586574
rect 9234 550894 9854 586338
rect 9234 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 9854 550894
rect 9234 550574 9854 550658
rect 9234 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 9854 550574
rect 9234 514894 9854 550338
rect 9234 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 9854 514894
rect 9234 514574 9854 514658
rect 9234 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 9854 514574
rect 9234 478894 9854 514338
rect 9234 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 9854 478894
rect 9234 478574 9854 478658
rect 9234 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 9854 478574
rect 9234 442894 9854 478338
rect 9234 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 9854 442894
rect 9234 442574 9854 442658
rect 9234 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 9854 442574
rect 9234 406894 9854 442338
rect 9234 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 9854 406894
rect 9234 406574 9854 406658
rect 9234 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 9854 406574
rect 9234 370894 9854 406338
rect 9234 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 9854 370894
rect 9234 370574 9854 370658
rect 9234 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 9854 370574
rect 9234 334894 9854 370338
rect 9234 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 9854 334894
rect 9234 334574 9854 334658
rect 9234 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 9854 334574
rect 9234 298894 9854 334338
rect 9234 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 9854 298894
rect 9234 298574 9854 298658
rect 9234 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 9854 298574
rect 9234 262894 9854 298338
rect 9234 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 9854 262894
rect 9234 262574 9854 262658
rect 9234 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 9854 262574
rect 9234 226894 9854 262338
rect 9234 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 9854 226894
rect 9234 226574 9854 226658
rect 9234 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 9854 226574
rect 9234 190894 9854 226338
rect 9234 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 9854 190894
rect 9234 190574 9854 190658
rect 9234 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 9854 190574
rect 9234 154894 9854 190338
rect 9234 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 9854 154894
rect 9234 154574 9854 154658
rect 9234 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 9854 154574
rect 9234 118894 9854 154338
rect 9234 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 9854 118894
rect 9234 118574 9854 118658
rect 9234 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 9854 118574
rect 9234 82894 9854 118338
rect 9234 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 9854 82894
rect 9234 82574 9854 82658
rect 9234 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 9854 82574
rect 9234 46894 9854 82338
rect 9234 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 9854 46894
rect 9234 46574 9854 46658
rect 9234 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 9854 46574
rect 9234 10894 9854 46338
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect 9234 -4186 9854 10338
rect 9234 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 9854 -4186
rect 9234 -4506 9854 -4422
rect 9234 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 9854 -4506
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect 9234 -5734 9854 -4742
rect 12954 698614 13574 710042
rect 30954 711558 31574 711590
rect 30954 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 31574 711558
rect 30954 711238 31574 711322
rect 30954 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 31574 711238
rect 27234 709638 27854 709670
rect 27234 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 27854 709638
rect 27234 709318 27854 709402
rect 27234 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 27854 709318
rect 23514 707718 24134 707750
rect 23514 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 24134 707718
rect 23514 707398 24134 707482
rect 23514 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 24134 707398
rect 12954 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 13574 698614
rect 12954 698294 13574 698378
rect 12954 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 13574 698294
rect 12954 662614 13574 698058
rect 12954 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 13574 662614
rect 12954 662294 13574 662378
rect 12954 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 13574 662294
rect 12954 626614 13574 662058
rect 12954 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 13574 626614
rect 12954 626294 13574 626378
rect 12954 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 13574 626294
rect 12954 590614 13574 626058
rect 12954 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 13574 590614
rect 12954 590294 13574 590378
rect 12954 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 13574 590294
rect 12954 554614 13574 590058
rect 12954 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 13574 554614
rect 12954 554294 13574 554378
rect 12954 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 13574 554294
rect 12954 518614 13574 554058
rect 12954 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 13574 518614
rect 12954 518294 13574 518378
rect 12954 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 13574 518294
rect 12954 482614 13574 518058
rect 12954 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 13574 482614
rect 12954 482294 13574 482378
rect 12954 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 13574 482294
rect 12954 446614 13574 482058
rect 12954 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 13574 446614
rect 12954 446294 13574 446378
rect 12954 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 13574 446294
rect 12954 410614 13574 446058
rect 12954 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 13574 410614
rect 12954 410294 13574 410378
rect 12954 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 13574 410294
rect 12954 374614 13574 410058
rect 12954 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 13574 374614
rect 12954 374294 13574 374378
rect 12954 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 13574 374294
rect 12954 338614 13574 374058
rect 12954 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 13574 338614
rect 12954 338294 13574 338378
rect 12954 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 13574 338294
rect 12954 302614 13574 338058
rect 12954 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 13574 302614
rect 12954 302294 13574 302378
rect 12954 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 13574 302294
rect 12954 266614 13574 302058
rect 12954 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 13574 266614
rect 12954 266294 13574 266378
rect 12954 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 13574 266294
rect 12954 230614 13574 266058
rect 12954 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 13574 230614
rect 12954 230294 13574 230378
rect 12954 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 13574 230294
rect 12954 194614 13574 230058
rect 12954 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 13574 194614
rect 12954 194294 13574 194378
rect 12954 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 13574 194294
rect 12954 158614 13574 194058
rect 12954 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 13574 158614
rect 12954 158294 13574 158378
rect 12954 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 13574 158294
rect 12954 122614 13574 158058
rect 12954 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 13574 122614
rect 12954 122294 13574 122378
rect 12954 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 13574 122294
rect 12954 86614 13574 122058
rect 12954 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 13574 86614
rect 12954 86294 13574 86378
rect 12954 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 13574 86294
rect 12954 50614 13574 86058
rect 12954 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 13574 50614
rect 12954 50294 13574 50378
rect 12954 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 13574 50294
rect 12954 14614 13574 50058
rect 12954 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 13574 14614
rect 12954 14294 13574 14378
rect 12954 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 13574 14294
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect 12954 -6106 13574 14058
rect 19794 705798 20414 705830
rect 19794 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 20414 705798
rect 19794 705478 20414 705562
rect 19794 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 20414 705478
rect 19794 669454 20414 705242
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -1306 20414 20898
rect 19794 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 20414 -1306
rect 19794 -1626 20414 -1542
rect 19794 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 20414 -1626
rect 19794 -1894 20414 -1862
rect 23514 673174 24134 707162
rect 23514 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 24134 673174
rect 23514 672854 24134 672938
rect 23514 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 24134 672854
rect 23514 637174 24134 672618
rect 23514 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 24134 637174
rect 23514 636854 24134 636938
rect 23514 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 24134 636854
rect 23514 601174 24134 636618
rect 23514 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 24134 601174
rect 23514 600854 24134 600938
rect 23514 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 24134 600854
rect 23514 565174 24134 600618
rect 23514 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 24134 565174
rect 23514 564854 24134 564938
rect 23514 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 24134 564854
rect 23514 529174 24134 564618
rect 23514 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 24134 529174
rect 23514 528854 24134 528938
rect 23514 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 24134 528854
rect 23514 493174 24134 528618
rect 23514 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 24134 493174
rect 23514 492854 24134 492938
rect 23514 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 24134 492854
rect 23514 457174 24134 492618
rect 23514 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 24134 457174
rect 23514 456854 24134 456938
rect 23514 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 24134 456854
rect 23514 421174 24134 456618
rect 23514 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 24134 421174
rect 23514 420854 24134 420938
rect 23514 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 24134 420854
rect 23514 385174 24134 420618
rect 23514 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 24134 385174
rect 23514 384854 24134 384938
rect 23514 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 24134 384854
rect 23514 349174 24134 384618
rect 23514 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 24134 349174
rect 23514 348854 24134 348938
rect 23514 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 24134 348854
rect 23514 313174 24134 348618
rect 23514 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 24134 313174
rect 23514 312854 24134 312938
rect 23514 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 24134 312854
rect 23514 277174 24134 312618
rect 23514 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 24134 277174
rect 23514 276854 24134 276938
rect 23514 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 24134 276854
rect 23514 241174 24134 276618
rect 23514 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 24134 241174
rect 23514 240854 24134 240938
rect 23514 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 24134 240854
rect 23514 205174 24134 240618
rect 23514 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 24134 205174
rect 23514 204854 24134 204938
rect 23514 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 24134 204854
rect 23514 169174 24134 204618
rect 23514 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 24134 169174
rect 23514 168854 24134 168938
rect 23514 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 24134 168854
rect 23514 133174 24134 168618
rect 23514 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 24134 133174
rect 23514 132854 24134 132938
rect 23514 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 24134 132854
rect 23514 97174 24134 132618
rect 23514 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 24134 97174
rect 23514 96854 24134 96938
rect 23514 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 24134 96854
rect 23514 61174 24134 96618
rect 23514 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 24134 61174
rect 23514 60854 24134 60938
rect 23514 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 24134 60854
rect 23514 25174 24134 60618
rect 23514 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 24134 25174
rect 23514 24854 24134 24938
rect 23514 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 24134 24854
rect 23514 -3226 24134 24618
rect 23514 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 24134 -3226
rect 23514 -3546 24134 -3462
rect 23514 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 24134 -3546
rect 23514 -3814 24134 -3782
rect 27234 676894 27854 709082
rect 27234 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 27854 676894
rect 27234 676574 27854 676658
rect 27234 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 27854 676574
rect 27234 640894 27854 676338
rect 27234 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 27854 640894
rect 27234 640574 27854 640658
rect 27234 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 27854 640574
rect 27234 604894 27854 640338
rect 27234 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 27854 604894
rect 27234 604574 27854 604658
rect 27234 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 27854 604574
rect 27234 568894 27854 604338
rect 27234 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 27854 568894
rect 27234 568574 27854 568658
rect 27234 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 27854 568574
rect 27234 532894 27854 568338
rect 27234 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 27854 532894
rect 27234 532574 27854 532658
rect 27234 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 27854 532574
rect 27234 496894 27854 532338
rect 27234 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 27854 496894
rect 27234 496574 27854 496658
rect 27234 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 27854 496574
rect 27234 460894 27854 496338
rect 27234 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 27854 460894
rect 27234 460574 27854 460658
rect 27234 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 27854 460574
rect 27234 424894 27854 460338
rect 27234 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 27854 424894
rect 27234 424574 27854 424658
rect 27234 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 27854 424574
rect 27234 388894 27854 424338
rect 27234 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 27854 388894
rect 27234 388574 27854 388658
rect 27234 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 27854 388574
rect 27234 352894 27854 388338
rect 27234 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 27854 352894
rect 27234 352574 27854 352658
rect 27234 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 27854 352574
rect 27234 316894 27854 352338
rect 27234 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 27854 316894
rect 27234 316574 27854 316658
rect 27234 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 27854 316574
rect 27234 280894 27854 316338
rect 27234 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 27854 280894
rect 27234 280574 27854 280658
rect 27234 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 27854 280574
rect 27234 244894 27854 280338
rect 27234 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 27854 244894
rect 27234 244574 27854 244658
rect 27234 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 27854 244574
rect 27234 208894 27854 244338
rect 27234 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 27854 208894
rect 27234 208574 27854 208658
rect 27234 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 27854 208574
rect 27234 172894 27854 208338
rect 27234 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 27854 172894
rect 27234 172574 27854 172658
rect 27234 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 27854 172574
rect 27234 136894 27854 172338
rect 27234 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 27854 136894
rect 27234 136574 27854 136658
rect 27234 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 27854 136574
rect 27234 100894 27854 136338
rect 27234 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 27854 100894
rect 27234 100574 27854 100658
rect 27234 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 27854 100574
rect 27234 64894 27854 100338
rect 27234 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 27854 64894
rect 27234 64574 27854 64658
rect 27234 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 27854 64574
rect 27234 28894 27854 64338
rect 27234 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 27854 28894
rect 27234 28574 27854 28658
rect 27234 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 27854 28574
rect 27234 -5146 27854 28338
rect 27234 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 27854 -5146
rect 27234 -5466 27854 -5382
rect 27234 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 27854 -5466
rect 27234 -5734 27854 -5702
rect 30954 680614 31574 711002
rect 48954 710598 49574 711590
rect 48954 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 49574 710598
rect 48954 710278 49574 710362
rect 48954 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 49574 710278
rect 45234 708678 45854 709670
rect 45234 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 45854 708678
rect 45234 708358 45854 708442
rect 45234 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 45854 708358
rect 41514 706758 42134 707750
rect 41514 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 42134 706758
rect 41514 706438 42134 706522
rect 41514 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 42134 706438
rect 30954 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 31574 680614
rect 30954 680294 31574 680378
rect 30954 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 31574 680294
rect 30954 644614 31574 680058
rect 30954 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 31574 644614
rect 30954 644294 31574 644378
rect 30954 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 31574 644294
rect 30954 608614 31574 644058
rect 30954 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 31574 608614
rect 30954 608294 31574 608378
rect 30954 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 31574 608294
rect 30954 572614 31574 608058
rect 30954 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 31574 572614
rect 30954 572294 31574 572378
rect 30954 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 31574 572294
rect 30954 536614 31574 572058
rect 30954 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 31574 536614
rect 30954 536294 31574 536378
rect 30954 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 31574 536294
rect 30954 500614 31574 536058
rect 30954 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 31574 500614
rect 30954 500294 31574 500378
rect 30954 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 31574 500294
rect 30954 464614 31574 500058
rect 30954 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 31574 464614
rect 30954 464294 31574 464378
rect 30954 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 31574 464294
rect 30954 428614 31574 464058
rect 30954 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 31574 428614
rect 30954 428294 31574 428378
rect 30954 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 31574 428294
rect 30954 392614 31574 428058
rect 30954 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 31574 392614
rect 30954 392294 31574 392378
rect 30954 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 31574 392294
rect 30954 356614 31574 392058
rect 30954 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 31574 356614
rect 30954 356294 31574 356378
rect 30954 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 31574 356294
rect 30954 320614 31574 356058
rect 30954 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 31574 320614
rect 30954 320294 31574 320378
rect 30954 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 31574 320294
rect 30954 284614 31574 320058
rect 30954 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 31574 284614
rect 30954 284294 31574 284378
rect 30954 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 31574 284294
rect 30954 248614 31574 284058
rect 30954 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 31574 248614
rect 30954 248294 31574 248378
rect 30954 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 31574 248294
rect 30954 212614 31574 248058
rect 30954 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 31574 212614
rect 30954 212294 31574 212378
rect 30954 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 31574 212294
rect 30954 176614 31574 212058
rect 30954 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 31574 176614
rect 30954 176294 31574 176378
rect 30954 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 31574 176294
rect 30954 140614 31574 176058
rect 30954 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 31574 140614
rect 30954 140294 31574 140378
rect 30954 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 31574 140294
rect 30954 104614 31574 140058
rect 30954 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 31574 104614
rect 30954 104294 31574 104378
rect 30954 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 31574 104294
rect 30954 68614 31574 104058
rect 30954 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 31574 68614
rect 30954 68294 31574 68378
rect 30954 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 31574 68294
rect 30954 32614 31574 68058
rect 30954 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 31574 32614
rect 30954 32294 31574 32378
rect 30954 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 31574 32294
rect 12954 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 13574 -6106
rect 12954 -6426 13574 -6342
rect 12954 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 13574 -6426
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 12954 -7654 13574 -6662
rect 30954 -7066 31574 32058
rect 37794 704838 38414 705830
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -1894 38414 -902
rect 41514 691174 42134 706202
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 41514 655174 42134 690618
rect 41514 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 42134 655174
rect 41514 654854 42134 654938
rect 41514 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 42134 654854
rect 41514 619174 42134 654618
rect 41514 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 42134 619174
rect 41514 618854 42134 618938
rect 41514 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 42134 618854
rect 41514 583174 42134 618618
rect 41514 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 42134 583174
rect 41514 582854 42134 582938
rect 41514 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 42134 582854
rect 41514 547174 42134 582618
rect 41514 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 42134 547174
rect 41514 546854 42134 546938
rect 41514 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 42134 546854
rect 41514 511174 42134 546618
rect 41514 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 42134 511174
rect 41514 510854 42134 510938
rect 41514 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 42134 510854
rect 41514 475174 42134 510618
rect 41514 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 42134 475174
rect 41514 474854 42134 474938
rect 41514 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 42134 474854
rect 41514 439174 42134 474618
rect 41514 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 42134 439174
rect 41514 438854 42134 438938
rect 41514 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 42134 438854
rect 41514 403174 42134 438618
rect 41514 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 42134 403174
rect 41514 402854 42134 402938
rect 41514 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 42134 402854
rect 41514 367174 42134 402618
rect 41514 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 42134 367174
rect 41514 366854 42134 366938
rect 41514 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 42134 366854
rect 41514 331174 42134 366618
rect 41514 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 42134 331174
rect 41514 330854 42134 330938
rect 41514 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 42134 330854
rect 41514 295174 42134 330618
rect 41514 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 42134 295174
rect 41514 294854 42134 294938
rect 41514 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 42134 294854
rect 41514 259174 42134 294618
rect 41514 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 42134 259174
rect 41514 258854 42134 258938
rect 41514 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 42134 258854
rect 41514 223174 42134 258618
rect 41514 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 42134 223174
rect 41514 222854 42134 222938
rect 41514 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 42134 222854
rect 41514 187174 42134 222618
rect 41514 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 42134 187174
rect 41514 186854 42134 186938
rect 41514 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 42134 186854
rect 41514 151174 42134 186618
rect 41514 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 42134 151174
rect 41514 150854 42134 150938
rect 41514 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 42134 150854
rect 41514 115174 42134 150618
rect 41514 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 42134 115174
rect 41514 114854 42134 114938
rect 41514 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 42134 114854
rect 41514 79174 42134 114618
rect 41514 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 42134 79174
rect 41514 78854 42134 78938
rect 41514 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 42134 78854
rect 41514 43174 42134 78618
rect 41514 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 42134 43174
rect 41514 42854 42134 42938
rect 41514 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 42134 42854
rect 41514 7174 42134 42618
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -2266 42134 6618
rect 41514 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 42134 -2266
rect 41514 -2586 42134 -2502
rect 41514 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 42134 -2586
rect 41514 -3814 42134 -2822
rect 45234 694894 45854 708122
rect 45234 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 45854 694894
rect 45234 694574 45854 694658
rect 45234 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 45854 694574
rect 45234 658894 45854 694338
rect 45234 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 45854 658894
rect 45234 658574 45854 658658
rect 45234 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 45854 658574
rect 45234 622894 45854 658338
rect 45234 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 45854 622894
rect 45234 622574 45854 622658
rect 45234 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 45854 622574
rect 45234 586894 45854 622338
rect 45234 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 45854 586894
rect 45234 586574 45854 586658
rect 45234 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 45854 586574
rect 45234 550894 45854 586338
rect 45234 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 45854 550894
rect 45234 550574 45854 550658
rect 45234 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 45854 550574
rect 45234 514894 45854 550338
rect 45234 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 45854 514894
rect 45234 514574 45854 514658
rect 45234 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 45854 514574
rect 45234 478894 45854 514338
rect 45234 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 45854 478894
rect 45234 478574 45854 478658
rect 45234 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 45854 478574
rect 45234 442894 45854 478338
rect 45234 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 45854 442894
rect 45234 442574 45854 442658
rect 45234 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 45854 442574
rect 45234 406894 45854 442338
rect 45234 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 45854 406894
rect 45234 406574 45854 406658
rect 45234 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 45854 406574
rect 45234 370894 45854 406338
rect 45234 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 45854 370894
rect 45234 370574 45854 370658
rect 45234 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 45854 370574
rect 45234 334894 45854 370338
rect 45234 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 45854 334894
rect 45234 334574 45854 334658
rect 45234 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 45854 334574
rect 45234 298894 45854 334338
rect 45234 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 45854 298894
rect 45234 298574 45854 298658
rect 45234 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 45854 298574
rect 45234 262894 45854 298338
rect 45234 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 45854 262894
rect 45234 262574 45854 262658
rect 45234 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 45854 262574
rect 45234 226894 45854 262338
rect 45234 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 45854 226894
rect 45234 226574 45854 226658
rect 45234 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 45854 226574
rect 45234 190894 45854 226338
rect 45234 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 45854 190894
rect 45234 190574 45854 190658
rect 45234 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 45854 190574
rect 45234 154894 45854 190338
rect 45234 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 45854 154894
rect 45234 154574 45854 154658
rect 45234 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 45854 154574
rect 45234 118894 45854 154338
rect 45234 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 45854 118894
rect 45234 118574 45854 118658
rect 45234 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 45854 118574
rect 45234 82894 45854 118338
rect 45234 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 45854 82894
rect 45234 82574 45854 82658
rect 45234 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 45854 82574
rect 45234 46894 45854 82338
rect 45234 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 45854 46894
rect 45234 46574 45854 46658
rect 45234 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 45854 46574
rect 45234 10894 45854 46338
rect 45234 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 45854 10894
rect 45234 10574 45854 10658
rect 45234 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 45854 10574
rect 45234 -4186 45854 10338
rect 45234 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 45854 -4186
rect 45234 -4506 45854 -4422
rect 45234 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 45854 -4506
rect 45234 -5734 45854 -4742
rect 48954 698614 49574 710042
rect 66954 711558 67574 711590
rect 66954 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 67574 711558
rect 66954 711238 67574 711322
rect 66954 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 67574 711238
rect 63234 709638 63854 709670
rect 63234 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 63854 709638
rect 63234 709318 63854 709402
rect 63234 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 63854 709318
rect 59514 707718 60134 707750
rect 59514 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 60134 707718
rect 59514 707398 60134 707482
rect 59514 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 60134 707398
rect 48954 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 49574 698614
rect 48954 698294 49574 698378
rect 48954 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 49574 698294
rect 48954 662614 49574 698058
rect 48954 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 49574 662614
rect 48954 662294 49574 662378
rect 48954 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 49574 662294
rect 48954 626614 49574 662058
rect 48954 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 49574 626614
rect 48954 626294 49574 626378
rect 48954 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 49574 626294
rect 48954 590614 49574 626058
rect 48954 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 49574 590614
rect 48954 590294 49574 590378
rect 48954 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 49574 590294
rect 48954 554614 49574 590058
rect 48954 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 49574 554614
rect 48954 554294 49574 554378
rect 48954 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 49574 554294
rect 48954 518614 49574 554058
rect 48954 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 49574 518614
rect 48954 518294 49574 518378
rect 48954 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 49574 518294
rect 48954 482614 49574 518058
rect 48954 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 49574 482614
rect 48954 482294 49574 482378
rect 48954 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 49574 482294
rect 48954 446614 49574 482058
rect 48954 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 49574 446614
rect 48954 446294 49574 446378
rect 48954 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 49574 446294
rect 48954 410614 49574 446058
rect 48954 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 49574 410614
rect 48954 410294 49574 410378
rect 48954 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 49574 410294
rect 48954 374614 49574 410058
rect 48954 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 49574 374614
rect 48954 374294 49574 374378
rect 48954 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 49574 374294
rect 48954 338614 49574 374058
rect 48954 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 49574 338614
rect 48954 338294 49574 338378
rect 48954 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 49574 338294
rect 48954 302614 49574 338058
rect 48954 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 49574 302614
rect 48954 302294 49574 302378
rect 48954 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 49574 302294
rect 48954 266614 49574 302058
rect 48954 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 49574 266614
rect 48954 266294 49574 266378
rect 48954 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 49574 266294
rect 48954 230614 49574 266058
rect 48954 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 49574 230614
rect 48954 230294 49574 230378
rect 48954 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 49574 230294
rect 48954 194614 49574 230058
rect 48954 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 49574 194614
rect 48954 194294 49574 194378
rect 48954 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 49574 194294
rect 48954 158614 49574 194058
rect 48954 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 49574 158614
rect 48954 158294 49574 158378
rect 48954 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 49574 158294
rect 48954 122614 49574 158058
rect 48954 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 49574 122614
rect 48954 122294 49574 122378
rect 48954 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 49574 122294
rect 48954 86614 49574 122058
rect 48954 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 49574 86614
rect 48954 86294 49574 86378
rect 48954 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 49574 86294
rect 48954 50614 49574 86058
rect 48954 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 49574 50614
rect 48954 50294 49574 50378
rect 48954 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 49574 50294
rect 48954 14614 49574 50058
rect 48954 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 49574 14614
rect 48954 14294 49574 14378
rect 48954 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 49574 14294
rect 30954 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 31574 -7066
rect 30954 -7386 31574 -7302
rect 30954 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 31574 -7386
rect 30954 -7654 31574 -7622
rect 48954 -6106 49574 14058
rect 55794 705798 56414 705830
rect 55794 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 56414 705798
rect 55794 705478 56414 705562
rect 55794 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 56414 705478
rect 55794 669454 56414 705242
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 273454 56414 308898
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 237454 56414 272898
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55794 201454 56414 236898
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -1306 56414 20898
rect 55794 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 56414 -1306
rect 55794 -1626 56414 -1542
rect 55794 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 56414 -1626
rect 55794 -1894 56414 -1862
rect 59514 673174 60134 707162
rect 59514 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 60134 673174
rect 59514 672854 60134 672938
rect 59514 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 60134 672854
rect 59514 637174 60134 672618
rect 59514 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 60134 637174
rect 59514 636854 60134 636938
rect 59514 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 60134 636854
rect 59514 601174 60134 636618
rect 59514 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 60134 601174
rect 59514 600854 60134 600938
rect 59514 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 60134 600854
rect 59514 565174 60134 600618
rect 59514 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 60134 565174
rect 59514 564854 60134 564938
rect 59514 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 60134 564854
rect 59514 529174 60134 564618
rect 59514 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 60134 529174
rect 59514 528854 60134 528938
rect 59514 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 60134 528854
rect 59514 493174 60134 528618
rect 59514 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 60134 493174
rect 59514 492854 60134 492938
rect 59514 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 60134 492854
rect 59514 457174 60134 492618
rect 59514 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 60134 457174
rect 59514 456854 60134 456938
rect 59514 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 60134 456854
rect 59514 421174 60134 456618
rect 59514 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 60134 421174
rect 59514 420854 60134 420938
rect 59514 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 60134 420854
rect 59514 385174 60134 420618
rect 59514 384938 59546 385174
rect 59782 384938 59866 385174
rect 60102 384938 60134 385174
rect 59514 384854 60134 384938
rect 59514 384618 59546 384854
rect 59782 384618 59866 384854
rect 60102 384618 60134 384854
rect 59514 349174 60134 384618
rect 59514 348938 59546 349174
rect 59782 348938 59866 349174
rect 60102 348938 60134 349174
rect 59514 348854 60134 348938
rect 59514 348618 59546 348854
rect 59782 348618 59866 348854
rect 60102 348618 60134 348854
rect 59514 313174 60134 348618
rect 59514 312938 59546 313174
rect 59782 312938 59866 313174
rect 60102 312938 60134 313174
rect 59514 312854 60134 312938
rect 59514 312618 59546 312854
rect 59782 312618 59866 312854
rect 60102 312618 60134 312854
rect 59514 277174 60134 312618
rect 59514 276938 59546 277174
rect 59782 276938 59866 277174
rect 60102 276938 60134 277174
rect 59514 276854 60134 276938
rect 59514 276618 59546 276854
rect 59782 276618 59866 276854
rect 60102 276618 60134 276854
rect 59514 241174 60134 276618
rect 59514 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 60134 241174
rect 59514 240854 60134 240938
rect 59514 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 60134 240854
rect 59514 205174 60134 240618
rect 59514 204938 59546 205174
rect 59782 204938 59866 205174
rect 60102 204938 60134 205174
rect 59514 204854 60134 204938
rect 59514 204618 59546 204854
rect 59782 204618 59866 204854
rect 60102 204618 60134 204854
rect 59514 169174 60134 204618
rect 59514 168938 59546 169174
rect 59782 168938 59866 169174
rect 60102 168938 60134 169174
rect 59514 168854 60134 168938
rect 59514 168618 59546 168854
rect 59782 168618 59866 168854
rect 60102 168618 60134 168854
rect 59514 133174 60134 168618
rect 59514 132938 59546 133174
rect 59782 132938 59866 133174
rect 60102 132938 60134 133174
rect 59514 132854 60134 132938
rect 59514 132618 59546 132854
rect 59782 132618 59866 132854
rect 60102 132618 60134 132854
rect 59514 97174 60134 132618
rect 59514 96938 59546 97174
rect 59782 96938 59866 97174
rect 60102 96938 60134 97174
rect 59514 96854 60134 96938
rect 59514 96618 59546 96854
rect 59782 96618 59866 96854
rect 60102 96618 60134 96854
rect 59514 61174 60134 96618
rect 59514 60938 59546 61174
rect 59782 60938 59866 61174
rect 60102 60938 60134 61174
rect 59514 60854 60134 60938
rect 59514 60618 59546 60854
rect 59782 60618 59866 60854
rect 60102 60618 60134 60854
rect 59514 25174 60134 60618
rect 59514 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 60134 25174
rect 59514 24854 60134 24938
rect 59514 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 60134 24854
rect 59514 -3226 60134 24618
rect 59514 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 60134 -3226
rect 59514 -3546 60134 -3462
rect 59514 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 60134 -3546
rect 59514 -3814 60134 -3782
rect 63234 676894 63854 709082
rect 63234 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 63854 676894
rect 63234 676574 63854 676658
rect 63234 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 63854 676574
rect 63234 640894 63854 676338
rect 63234 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 63854 640894
rect 63234 640574 63854 640658
rect 63234 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 63854 640574
rect 63234 604894 63854 640338
rect 63234 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 63854 604894
rect 63234 604574 63854 604658
rect 63234 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 63854 604574
rect 63234 568894 63854 604338
rect 63234 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 63854 568894
rect 63234 568574 63854 568658
rect 63234 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 63854 568574
rect 63234 532894 63854 568338
rect 63234 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 63854 532894
rect 63234 532574 63854 532658
rect 63234 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 63854 532574
rect 63234 496894 63854 532338
rect 63234 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 63854 496894
rect 63234 496574 63854 496658
rect 63234 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 63854 496574
rect 63234 460894 63854 496338
rect 63234 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 63854 460894
rect 63234 460574 63854 460658
rect 63234 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 63854 460574
rect 63234 424894 63854 460338
rect 63234 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 63854 424894
rect 63234 424574 63854 424658
rect 63234 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 63854 424574
rect 63234 388894 63854 424338
rect 63234 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 63854 388894
rect 63234 388574 63854 388658
rect 63234 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 63854 388574
rect 63234 352894 63854 388338
rect 63234 352658 63266 352894
rect 63502 352658 63586 352894
rect 63822 352658 63854 352894
rect 63234 352574 63854 352658
rect 63234 352338 63266 352574
rect 63502 352338 63586 352574
rect 63822 352338 63854 352574
rect 63234 316894 63854 352338
rect 63234 316658 63266 316894
rect 63502 316658 63586 316894
rect 63822 316658 63854 316894
rect 63234 316574 63854 316658
rect 63234 316338 63266 316574
rect 63502 316338 63586 316574
rect 63822 316338 63854 316574
rect 63234 280894 63854 316338
rect 63234 280658 63266 280894
rect 63502 280658 63586 280894
rect 63822 280658 63854 280894
rect 63234 280574 63854 280658
rect 63234 280338 63266 280574
rect 63502 280338 63586 280574
rect 63822 280338 63854 280574
rect 63234 244894 63854 280338
rect 63234 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 63854 244894
rect 63234 244574 63854 244658
rect 63234 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 63854 244574
rect 63234 208894 63854 244338
rect 63234 208658 63266 208894
rect 63502 208658 63586 208894
rect 63822 208658 63854 208894
rect 63234 208574 63854 208658
rect 63234 208338 63266 208574
rect 63502 208338 63586 208574
rect 63822 208338 63854 208574
rect 63234 172894 63854 208338
rect 63234 172658 63266 172894
rect 63502 172658 63586 172894
rect 63822 172658 63854 172894
rect 63234 172574 63854 172658
rect 63234 172338 63266 172574
rect 63502 172338 63586 172574
rect 63822 172338 63854 172574
rect 63234 136894 63854 172338
rect 63234 136658 63266 136894
rect 63502 136658 63586 136894
rect 63822 136658 63854 136894
rect 63234 136574 63854 136658
rect 63234 136338 63266 136574
rect 63502 136338 63586 136574
rect 63822 136338 63854 136574
rect 63234 100894 63854 136338
rect 63234 100658 63266 100894
rect 63502 100658 63586 100894
rect 63822 100658 63854 100894
rect 63234 100574 63854 100658
rect 63234 100338 63266 100574
rect 63502 100338 63586 100574
rect 63822 100338 63854 100574
rect 63234 64894 63854 100338
rect 63234 64658 63266 64894
rect 63502 64658 63586 64894
rect 63822 64658 63854 64894
rect 63234 64574 63854 64658
rect 63234 64338 63266 64574
rect 63502 64338 63586 64574
rect 63822 64338 63854 64574
rect 63234 28894 63854 64338
rect 63234 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 63854 28894
rect 63234 28574 63854 28658
rect 63234 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 63854 28574
rect 63234 -5146 63854 28338
rect 63234 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 63854 -5146
rect 63234 -5466 63854 -5382
rect 63234 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 63854 -5466
rect 63234 -5734 63854 -5702
rect 66954 680614 67574 711002
rect 84954 710598 85574 711590
rect 84954 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 85574 710598
rect 84954 710278 85574 710362
rect 84954 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 85574 710278
rect 81234 708678 81854 709670
rect 81234 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 81854 708678
rect 81234 708358 81854 708442
rect 81234 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 81854 708358
rect 77514 706758 78134 707750
rect 77514 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 78134 706758
rect 77514 706438 78134 706522
rect 77514 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 78134 706438
rect 66954 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 67574 680614
rect 66954 680294 67574 680378
rect 66954 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 67574 680294
rect 66954 644614 67574 680058
rect 66954 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 67574 644614
rect 66954 644294 67574 644378
rect 66954 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 67574 644294
rect 66954 608614 67574 644058
rect 66954 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 67574 608614
rect 66954 608294 67574 608378
rect 66954 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 67574 608294
rect 66954 572614 67574 608058
rect 66954 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 67574 572614
rect 66954 572294 67574 572378
rect 66954 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 67574 572294
rect 66954 536614 67574 572058
rect 66954 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 67574 536614
rect 66954 536294 67574 536378
rect 66954 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 67574 536294
rect 66954 500614 67574 536058
rect 66954 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 67574 500614
rect 66954 500294 67574 500378
rect 66954 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 67574 500294
rect 66954 464614 67574 500058
rect 66954 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 67574 464614
rect 66954 464294 67574 464378
rect 66954 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 67574 464294
rect 66954 428614 67574 464058
rect 66954 428378 66986 428614
rect 67222 428378 67306 428614
rect 67542 428378 67574 428614
rect 66954 428294 67574 428378
rect 66954 428058 66986 428294
rect 67222 428058 67306 428294
rect 67542 428058 67574 428294
rect 66954 392614 67574 428058
rect 66954 392378 66986 392614
rect 67222 392378 67306 392614
rect 67542 392378 67574 392614
rect 66954 392294 67574 392378
rect 66954 392058 66986 392294
rect 67222 392058 67306 392294
rect 67542 392058 67574 392294
rect 66954 356614 67574 392058
rect 66954 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 67574 356614
rect 66954 356294 67574 356378
rect 66954 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 67574 356294
rect 66954 320614 67574 356058
rect 66954 320378 66986 320614
rect 67222 320378 67306 320614
rect 67542 320378 67574 320614
rect 66954 320294 67574 320378
rect 66954 320058 66986 320294
rect 67222 320058 67306 320294
rect 67542 320058 67574 320294
rect 66954 284614 67574 320058
rect 66954 284378 66986 284614
rect 67222 284378 67306 284614
rect 67542 284378 67574 284614
rect 66954 284294 67574 284378
rect 66954 284058 66986 284294
rect 67222 284058 67306 284294
rect 67542 284058 67574 284294
rect 66954 248614 67574 284058
rect 66954 248378 66986 248614
rect 67222 248378 67306 248614
rect 67542 248378 67574 248614
rect 66954 248294 67574 248378
rect 66954 248058 66986 248294
rect 67222 248058 67306 248294
rect 67542 248058 67574 248294
rect 66954 212614 67574 248058
rect 66954 212378 66986 212614
rect 67222 212378 67306 212614
rect 67542 212378 67574 212614
rect 66954 212294 67574 212378
rect 66954 212058 66986 212294
rect 67222 212058 67306 212294
rect 67542 212058 67574 212294
rect 66954 176614 67574 212058
rect 66954 176378 66986 176614
rect 67222 176378 67306 176614
rect 67542 176378 67574 176614
rect 66954 176294 67574 176378
rect 66954 176058 66986 176294
rect 67222 176058 67306 176294
rect 67542 176058 67574 176294
rect 66954 140614 67574 176058
rect 66954 140378 66986 140614
rect 67222 140378 67306 140614
rect 67542 140378 67574 140614
rect 66954 140294 67574 140378
rect 66954 140058 66986 140294
rect 67222 140058 67306 140294
rect 67542 140058 67574 140294
rect 66954 104614 67574 140058
rect 66954 104378 66986 104614
rect 67222 104378 67306 104614
rect 67542 104378 67574 104614
rect 66954 104294 67574 104378
rect 66954 104058 66986 104294
rect 67222 104058 67306 104294
rect 67542 104058 67574 104294
rect 66954 68614 67574 104058
rect 66954 68378 66986 68614
rect 67222 68378 67306 68614
rect 67542 68378 67574 68614
rect 66954 68294 67574 68378
rect 66954 68058 66986 68294
rect 67222 68058 67306 68294
rect 67542 68058 67574 68294
rect 66954 32614 67574 68058
rect 66954 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 67574 32614
rect 66954 32294 67574 32378
rect 66954 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 67574 32294
rect 48954 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 49574 -6106
rect 48954 -6426 49574 -6342
rect 48954 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 49574 -6426
rect 48954 -7654 49574 -6662
rect 66954 -7066 67574 32058
rect 73794 704838 74414 705830
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 579454 74414 614898
rect 73794 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 74414 579454
rect 73794 579134 74414 579218
rect 73794 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 74414 579134
rect 73794 543454 74414 578898
rect 73794 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 74414 543454
rect 73794 543134 74414 543218
rect 73794 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 74414 543134
rect 73794 507454 74414 542898
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 471454 74414 506898
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73794 435454 74414 470898
rect 73794 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 74414 435454
rect 73794 435134 74414 435218
rect 73794 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 74414 435134
rect 73794 399454 74414 434898
rect 73794 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 74414 399454
rect 73794 399134 74414 399218
rect 73794 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 74414 399134
rect 73794 363454 74414 398898
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 73794 327454 74414 362898
rect 73794 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 74414 327454
rect 73794 327134 74414 327218
rect 73794 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 74414 327134
rect 73794 291454 74414 326898
rect 73794 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 74414 291454
rect 73794 291134 74414 291218
rect 73794 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 74414 291134
rect 73794 255454 74414 290898
rect 73794 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 74414 255454
rect 73794 255134 74414 255218
rect 73794 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 74414 255134
rect 73794 219454 74414 254898
rect 73794 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 74414 219454
rect 73794 219134 74414 219218
rect 73794 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 74414 219134
rect 73794 183454 74414 218898
rect 73794 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 74414 183454
rect 73794 183134 74414 183218
rect 73794 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 74414 183134
rect 73794 147454 74414 182898
rect 73794 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 74414 147454
rect 73794 147134 74414 147218
rect 73794 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 74414 147134
rect 73794 111454 74414 146898
rect 73794 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 74414 111454
rect 73794 111134 74414 111218
rect 73794 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 74414 111134
rect 73794 75454 74414 110898
rect 73794 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 74414 75454
rect 73794 75134 74414 75218
rect 73794 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 74414 75134
rect 73794 39454 74414 74898
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -1894 74414 -902
rect 77514 691174 78134 706202
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 655174 78134 690618
rect 77514 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 78134 655174
rect 77514 654854 78134 654938
rect 77514 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 78134 654854
rect 77514 619174 78134 654618
rect 77514 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 78134 619174
rect 77514 618854 78134 618938
rect 77514 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 78134 618854
rect 77514 583174 78134 618618
rect 77514 582938 77546 583174
rect 77782 582938 77866 583174
rect 78102 582938 78134 583174
rect 77514 582854 78134 582938
rect 77514 582618 77546 582854
rect 77782 582618 77866 582854
rect 78102 582618 78134 582854
rect 77514 547174 78134 582618
rect 77514 546938 77546 547174
rect 77782 546938 77866 547174
rect 78102 546938 78134 547174
rect 77514 546854 78134 546938
rect 77514 546618 77546 546854
rect 77782 546618 77866 546854
rect 78102 546618 78134 546854
rect 77514 511174 78134 546618
rect 77514 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 78134 511174
rect 77514 510854 78134 510938
rect 77514 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 78134 510854
rect 77514 475174 78134 510618
rect 77514 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 78134 475174
rect 77514 474854 78134 474938
rect 77514 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 78134 474854
rect 77514 439174 78134 474618
rect 77514 438938 77546 439174
rect 77782 438938 77866 439174
rect 78102 438938 78134 439174
rect 77514 438854 78134 438938
rect 77514 438618 77546 438854
rect 77782 438618 77866 438854
rect 78102 438618 78134 438854
rect 77514 403174 78134 438618
rect 77514 402938 77546 403174
rect 77782 402938 77866 403174
rect 78102 402938 78134 403174
rect 77514 402854 78134 402938
rect 77514 402618 77546 402854
rect 77782 402618 77866 402854
rect 78102 402618 78134 402854
rect 77514 367174 78134 402618
rect 77514 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 78134 367174
rect 77514 366854 78134 366938
rect 77514 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 78134 366854
rect 77514 331174 78134 366618
rect 77514 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 78134 331174
rect 77514 330854 78134 330938
rect 77514 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 78134 330854
rect 77514 295174 78134 330618
rect 77514 294938 77546 295174
rect 77782 294938 77866 295174
rect 78102 294938 78134 295174
rect 77514 294854 78134 294938
rect 77514 294618 77546 294854
rect 77782 294618 77866 294854
rect 78102 294618 78134 294854
rect 77514 259174 78134 294618
rect 77514 258938 77546 259174
rect 77782 258938 77866 259174
rect 78102 258938 78134 259174
rect 77514 258854 78134 258938
rect 77514 258618 77546 258854
rect 77782 258618 77866 258854
rect 78102 258618 78134 258854
rect 77514 223174 78134 258618
rect 77514 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 78134 223174
rect 77514 222854 78134 222938
rect 77514 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 78134 222854
rect 77514 187174 78134 222618
rect 77514 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 78134 187174
rect 77514 186854 78134 186938
rect 77514 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 78134 186854
rect 77514 151174 78134 186618
rect 77514 150938 77546 151174
rect 77782 150938 77866 151174
rect 78102 150938 78134 151174
rect 77514 150854 78134 150938
rect 77514 150618 77546 150854
rect 77782 150618 77866 150854
rect 78102 150618 78134 150854
rect 77514 115174 78134 150618
rect 77514 114938 77546 115174
rect 77782 114938 77866 115174
rect 78102 114938 78134 115174
rect 77514 114854 78134 114938
rect 77514 114618 77546 114854
rect 77782 114618 77866 114854
rect 78102 114618 78134 114854
rect 77514 79174 78134 114618
rect 77514 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 78134 79174
rect 77514 78854 78134 78938
rect 77514 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 78134 78854
rect 77514 43174 78134 78618
rect 77514 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 78134 43174
rect 77514 42854 78134 42938
rect 77514 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 78134 42854
rect 77514 7174 78134 42618
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 77514 -2266 78134 6618
rect 77514 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 78134 -2266
rect 77514 -2586 78134 -2502
rect 77514 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 78134 -2586
rect 77514 -3814 78134 -2822
rect 81234 694894 81854 708122
rect 81234 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 81854 694894
rect 81234 694574 81854 694658
rect 81234 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 81854 694574
rect 81234 658894 81854 694338
rect 81234 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 81854 658894
rect 81234 658574 81854 658658
rect 81234 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 81854 658574
rect 81234 622894 81854 658338
rect 81234 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 81854 622894
rect 81234 622574 81854 622658
rect 81234 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 81854 622574
rect 81234 586894 81854 622338
rect 81234 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 81854 586894
rect 81234 586574 81854 586658
rect 81234 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 81854 586574
rect 81234 550894 81854 586338
rect 81234 550658 81266 550894
rect 81502 550658 81586 550894
rect 81822 550658 81854 550894
rect 81234 550574 81854 550658
rect 81234 550338 81266 550574
rect 81502 550338 81586 550574
rect 81822 550338 81854 550574
rect 81234 514894 81854 550338
rect 81234 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 81854 514894
rect 81234 514574 81854 514658
rect 81234 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 81854 514574
rect 81234 478894 81854 514338
rect 81234 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 81854 478894
rect 81234 478574 81854 478658
rect 81234 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 81854 478574
rect 81234 442894 81854 478338
rect 81234 442658 81266 442894
rect 81502 442658 81586 442894
rect 81822 442658 81854 442894
rect 81234 442574 81854 442658
rect 81234 442338 81266 442574
rect 81502 442338 81586 442574
rect 81822 442338 81854 442574
rect 81234 406894 81854 442338
rect 81234 406658 81266 406894
rect 81502 406658 81586 406894
rect 81822 406658 81854 406894
rect 81234 406574 81854 406658
rect 81234 406338 81266 406574
rect 81502 406338 81586 406574
rect 81822 406338 81854 406574
rect 81234 370894 81854 406338
rect 81234 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 81854 370894
rect 81234 370574 81854 370658
rect 81234 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 81854 370574
rect 81234 334894 81854 370338
rect 81234 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 81854 334894
rect 81234 334574 81854 334658
rect 81234 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 81854 334574
rect 81234 298894 81854 334338
rect 81234 298658 81266 298894
rect 81502 298658 81586 298894
rect 81822 298658 81854 298894
rect 81234 298574 81854 298658
rect 81234 298338 81266 298574
rect 81502 298338 81586 298574
rect 81822 298338 81854 298574
rect 81234 262894 81854 298338
rect 81234 262658 81266 262894
rect 81502 262658 81586 262894
rect 81822 262658 81854 262894
rect 81234 262574 81854 262658
rect 81234 262338 81266 262574
rect 81502 262338 81586 262574
rect 81822 262338 81854 262574
rect 81234 226894 81854 262338
rect 81234 226658 81266 226894
rect 81502 226658 81586 226894
rect 81822 226658 81854 226894
rect 81234 226574 81854 226658
rect 81234 226338 81266 226574
rect 81502 226338 81586 226574
rect 81822 226338 81854 226574
rect 81234 190894 81854 226338
rect 81234 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 81854 190894
rect 81234 190574 81854 190658
rect 81234 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 81854 190574
rect 81234 154894 81854 190338
rect 81234 154658 81266 154894
rect 81502 154658 81586 154894
rect 81822 154658 81854 154894
rect 81234 154574 81854 154658
rect 81234 154338 81266 154574
rect 81502 154338 81586 154574
rect 81822 154338 81854 154574
rect 81234 118894 81854 154338
rect 81234 118658 81266 118894
rect 81502 118658 81586 118894
rect 81822 118658 81854 118894
rect 81234 118574 81854 118658
rect 81234 118338 81266 118574
rect 81502 118338 81586 118574
rect 81822 118338 81854 118574
rect 81234 82894 81854 118338
rect 81234 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 81854 82894
rect 81234 82574 81854 82658
rect 81234 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 81854 82574
rect 81234 46894 81854 82338
rect 81234 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 81854 46894
rect 81234 46574 81854 46658
rect 81234 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 81854 46574
rect 81234 10894 81854 46338
rect 81234 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 81854 10894
rect 81234 10574 81854 10658
rect 81234 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 81854 10574
rect 81234 -4186 81854 10338
rect 81234 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 81854 -4186
rect 81234 -4506 81854 -4422
rect 81234 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 81854 -4506
rect 81234 -5734 81854 -4742
rect 84954 698614 85574 710042
rect 102954 711558 103574 711590
rect 102954 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 103574 711558
rect 102954 711238 103574 711322
rect 102954 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 103574 711238
rect 99234 709638 99854 709670
rect 99234 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 99854 709638
rect 99234 709318 99854 709402
rect 99234 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 99854 709318
rect 95514 707718 96134 707750
rect 95514 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 96134 707718
rect 95514 707398 96134 707482
rect 95514 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 96134 707398
rect 84954 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 85574 698614
rect 84954 698294 85574 698378
rect 84954 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 85574 698294
rect 84954 662614 85574 698058
rect 84954 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 85574 662614
rect 84954 662294 85574 662378
rect 84954 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 85574 662294
rect 84954 626614 85574 662058
rect 84954 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 85574 626614
rect 84954 626294 85574 626378
rect 84954 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 85574 626294
rect 84954 590614 85574 626058
rect 84954 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 85574 590614
rect 84954 590294 85574 590378
rect 84954 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 85574 590294
rect 84954 554614 85574 590058
rect 84954 554378 84986 554614
rect 85222 554378 85306 554614
rect 85542 554378 85574 554614
rect 84954 554294 85574 554378
rect 84954 554058 84986 554294
rect 85222 554058 85306 554294
rect 85542 554058 85574 554294
rect 84954 518614 85574 554058
rect 84954 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 85574 518614
rect 84954 518294 85574 518378
rect 84954 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 85574 518294
rect 84954 482614 85574 518058
rect 84954 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 85574 482614
rect 84954 482294 85574 482378
rect 84954 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 85574 482294
rect 84954 446614 85574 482058
rect 84954 446378 84986 446614
rect 85222 446378 85306 446614
rect 85542 446378 85574 446614
rect 84954 446294 85574 446378
rect 84954 446058 84986 446294
rect 85222 446058 85306 446294
rect 85542 446058 85574 446294
rect 84954 410614 85574 446058
rect 84954 410378 84986 410614
rect 85222 410378 85306 410614
rect 85542 410378 85574 410614
rect 84954 410294 85574 410378
rect 84954 410058 84986 410294
rect 85222 410058 85306 410294
rect 85542 410058 85574 410294
rect 84954 374614 85574 410058
rect 84954 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 85574 374614
rect 84954 374294 85574 374378
rect 84954 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 85574 374294
rect 84954 338614 85574 374058
rect 84954 338378 84986 338614
rect 85222 338378 85306 338614
rect 85542 338378 85574 338614
rect 84954 338294 85574 338378
rect 84954 338058 84986 338294
rect 85222 338058 85306 338294
rect 85542 338058 85574 338294
rect 84954 302614 85574 338058
rect 84954 302378 84986 302614
rect 85222 302378 85306 302614
rect 85542 302378 85574 302614
rect 84954 302294 85574 302378
rect 84954 302058 84986 302294
rect 85222 302058 85306 302294
rect 85542 302058 85574 302294
rect 84954 266614 85574 302058
rect 84954 266378 84986 266614
rect 85222 266378 85306 266614
rect 85542 266378 85574 266614
rect 84954 266294 85574 266378
rect 84954 266058 84986 266294
rect 85222 266058 85306 266294
rect 85542 266058 85574 266294
rect 84954 230614 85574 266058
rect 84954 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 85574 230614
rect 84954 230294 85574 230378
rect 84954 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 85574 230294
rect 84954 194614 85574 230058
rect 84954 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 85574 194614
rect 84954 194294 85574 194378
rect 84954 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 85574 194294
rect 84954 158614 85574 194058
rect 84954 158378 84986 158614
rect 85222 158378 85306 158614
rect 85542 158378 85574 158614
rect 84954 158294 85574 158378
rect 84954 158058 84986 158294
rect 85222 158058 85306 158294
rect 85542 158058 85574 158294
rect 84954 122614 85574 158058
rect 84954 122378 84986 122614
rect 85222 122378 85306 122614
rect 85542 122378 85574 122614
rect 84954 122294 85574 122378
rect 84954 122058 84986 122294
rect 85222 122058 85306 122294
rect 85542 122058 85574 122294
rect 84954 86614 85574 122058
rect 84954 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 85574 86614
rect 84954 86294 85574 86378
rect 84954 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 85574 86294
rect 84954 50614 85574 86058
rect 84954 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 85574 50614
rect 84954 50294 85574 50378
rect 84954 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 85574 50294
rect 84954 14614 85574 50058
rect 84954 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 85574 14614
rect 84954 14294 85574 14378
rect 84954 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 85574 14294
rect 66954 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 67574 -7066
rect 66954 -7386 67574 -7302
rect 66954 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 67574 -7386
rect 66954 -7654 67574 -7622
rect 84954 -6106 85574 14058
rect 91794 705798 92414 705830
rect 91794 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 92414 705798
rect 91794 705478 92414 705562
rect 91794 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 92414 705478
rect 91794 669454 92414 705242
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 91794 561454 92414 596898
rect 91794 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 92414 561454
rect 91794 561134 92414 561218
rect 91794 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 92414 561134
rect 91794 525454 92414 560898
rect 91794 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 92414 525454
rect 91794 525134 92414 525218
rect 91794 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 92414 525134
rect 91794 489454 92414 524898
rect 91794 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 92414 489454
rect 91794 489134 92414 489218
rect 91794 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 92414 489134
rect 91794 453454 92414 488898
rect 91794 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 92414 453454
rect 91794 453134 92414 453218
rect 91794 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 92414 453134
rect 91794 417454 92414 452898
rect 91794 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 92414 417454
rect 91794 417134 92414 417218
rect 91794 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 92414 417134
rect 91794 381454 92414 416898
rect 91794 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 92414 381454
rect 91794 381134 92414 381218
rect 91794 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 92414 381134
rect 91794 345454 92414 380898
rect 91794 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 92414 345454
rect 91794 345134 92414 345218
rect 91794 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 92414 345134
rect 91794 309454 92414 344898
rect 91794 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 92414 309454
rect 91794 309134 92414 309218
rect 91794 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 92414 309134
rect 91794 273454 92414 308898
rect 91794 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 92414 273454
rect 91794 273134 92414 273218
rect 91794 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 92414 273134
rect 91794 237454 92414 272898
rect 91794 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 92414 237454
rect 91794 237134 92414 237218
rect 91794 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 92414 237134
rect 91794 201454 92414 236898
rect 91794 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 92414 201454
rect 91794 201134 92414 201218
rect 91794 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 92414 201134
rect 91794 165454 92414 200898
rect 91794 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 92414 165454
rect 91794 165134 92414 165218
rect 91794 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 92414 165134
rect 91794 129454 92414 164898
rect 91794 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 92414 129454
rect 91794 129134 92414 129218
rect 91794 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 92414 129134
rect 91794 93454 92414 128898
rect 91794 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 92414 93454
rect 91794 93134 92414 93218
rect 91794 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 92414 93134
rect 91794 57454 92414 92898
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -1306 92414 20898
rect 91794 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 92414 -1306
rect 91794 -1626 92414 -1542
rect 91794 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 92414 -1626
rect 91794 -1894 92414 -1862
rect 95514 673174 96134 707162
rect 95514 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 96134 673174
rect 95514 672854 96134 672938
rect 95514 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 96134 672854
rect 95514 637174 96134 672618
rect 95514 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 96134 637174
rect 95514 636854 96134 636938
rect 95514 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 96134 636854
rect 95514 601174 96134 636618
rect 95514 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 96134 601174
rect 95514 600854 96134 600938
rect 95514 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 96134 600854
rect 95514 565174 96134 600618
rect 95514 564938 95546 565174
rect 95782 564938 95866 565174
rect 96102 564938 96134 565174
rect 95514 564854 96134 564938
rect 95514 564618 95546 564854
rect 95782 564618 95866 564854
rect 96102 564618 96134 564854
rect 95514 529174 96134 564618
rect 95514 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 96134 529174
rect 95514 528854 96134 528938
rect 95514 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 96134 528854
rect 95514 493174 96134 528618
rect 95514 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 96134 493174
rect 95514 492854 96134 492938
rect 95514 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 96134 492854
rect 95514 457174 96134 492618
rect 95514 456938 95546 457174
rect 95782 456938 95866 457174
rect 96102 456938 96134 457174
rect 95514 456854 96134 456938
rect 95514 456618 95546 456854
rect 95782 456618 95866 456854
rect 96102 456618 96134 456854
rect 95514 421174 96134 456618
rect 95514 420938 95546 421174
rect 95782 420938 95866 421174
rect 96102 420938 96134 421174
rect 95514 420854 96134 420938
rect 95514 420618 95546 420854
rect 95782 420618 95866 420854
rect 96102 420618 96134 420854
rect 95514 385174 96134 420618
rect 95514 384938 95546 385174
rect 95782 384938 95866 385174
rect 96102 384938 96134 385174
rect 95514 384854 96134 384938
rect 95514 384618 95546 384854
rect 95782 384618 95866 384854
rect 96102 384618 96134 384854
rect 95514 349174 96134 384618
rect 95514 348938 95546 349174
rect 95782 348938 95866 349174
rect 96102 348938 96134 349174
rect 95514 348854 96134 348938
rect 95514 348618 95546 348854
rect 95782 348618 95866 348854
rect 96102 348618 96134 348854
rect 95514 313174 96134 348618
rect 95514 312938 95546 313174
rect 95782 312938 95866 313174
rect 96102 312938 96134 313174
rect 95514 312854 96134 312938
rect 95514 312618 95546 312854
rect 95782 312618 95866 312854
rect 96102 312618 96134 312854
rect 95514 277174 96134 312618
rect 95514 276938 95546 277174
rect 95782 276938 95866 277174
rect 96102 276938 96134 277174
rect 95514 276854 96134 276938
rect 95514 276618 95546 276854
rect 95782 276618 95866 276854
rect 96102 276618 96134 276854
rect 95514 241174 96134 276618
rect 95514 240938 95546 241174
rect 95782 240938 95866 241174
rect 96102 240938 96134 241174
rect 95514 240854 96134 240938
rect 95514 240618 95546 240854
rect 95782 240618 95866 240854
rect 96102 240618 96134 240854
rect 95514 205174 96134 240618
rect 95514 204938 95546 205174
rect 95782 204938 95866 205174
rect 96102 204938 96134 205174
rect 95514 204854 96134 204938
rect 95514 204618 95546 204854
rect 95782 204618 95866 204854
rect 96102 204618 96134 204854
rect 95514 169174 96134 204618
rect 95514 168938 95546 169174
rect 95782 168938 95866 169174
rect 96102 168938 96134 169174
rect 95514 168854 96134 168938
rect 95514 168618 95546 168854
rect 95782 168618 95866 168854
rect 96102 168618 96134 168854
rect 95514 133174 96134 168618
rect 95514 132938 95546 133174
rect 95782 132938 95866 133174
rect 96102 132938 96134 133174
rect 95514 132854 96134 132938
rect 95514 132618 95546 132854
rect 95782 132618 95866 132854
rect 96102 132618 96134 132854
rect 95514 97174 96134 132618
rect 95514 96938 95546 97174
rect 95782 96938 95866 97174
rect 96102 96938 96134 97174
rect 95514 96854 96134 96938
rect 95514 96618 95546 96854
rect 95782 96618 95866 96854
rect 96102 96618 96134 96854
rect 95514 61174 96134 96618
rect 95514 60938 95546 61174
rect 95782 60938 95866 61174
rect 96102 60938 96134 61174
rect 95514 60854 96134 60938
rect 95514 60618 95546 60854
rect 95782 60618 95866 60854
rect 96102 60618 96134 60854
rect 95514 25174 96134 60618
rect 95514 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 96134 25174
rect 95514 24854 96134 24938
rect 95514 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 96134 24854
rect 95514 -3226 96134 24618
rect 95514 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 96134 -3226
rect 95514 -3546 96134 -3462
rect 95514 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 96134 -3546
rect 95514 -3814 96134 -3782
rect 99234 676894 99854 709082
rect 99234 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 99854 676894
rect 99234 676574 99854 676658
rect 99234 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 99854 676574
rect 99234 640894 99854 676338
rect 99234 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 99854 640894
rect 99234 640574 99854 640658
rect 99234 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 99854 640574
rect 99234 604894 99854 640338
rect 99234 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 99854 604894
rect 99234 604574 99854 604658
rect 99234 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 99854 604574
rect 99234 568894 99854 604338
rect 99234 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 99854 568894
rect 99234 568574 99854 568658
rect 99234 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 99854 568574
rect 99234 532894 99854 568338
rect 99234 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 99854 532894
rect 99234 532574 99854 532658
rect 99234 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 99854 532574
rect 99234 496894 99854 532338
rect 99234 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 99854 496894
rect 99234 496574 99854 496658
rect 99234 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 99854 496574
rect 99234 460894 99854 496338
rect 99234 460658 99266 460894
rect 99502 460658 99586 460894
rect 99822 460658 99854 460894
rect 99234 460574 99854 460658
rect 99234 460338 99266 460574
rect 99502 460338 99586 460574
rect 99822 460338 99854 460574
rect 99234 424894 99854 460338
rect 99234 424658 99266 424894
rect 99502 424658 99586 424894
rect 99822 424658 99854 424894
rect 99234 424574 99854 424658
rect 99234 424338 99266 424574
rect 99502 424338 99586 424574
rect 99822 424338 99854 424574
rect 99234 388894 99854 424338
rect 99234 388658 99266 388894
rect 99502 388658 99586 388894
rect 99822 388658 99854 388894
rect 99234 388574 99854 388658
rect 99234 388338 99266 388574
rect 99502 388338 99586 388574
rect 99822 388338 99854 388574
rect 99234 352894 99854 388338
rect 99234 352658 99266 352894
rect 99502 352658 99586 352894
rect 99822 352658 99854 352894
rect 99234 352574 99854 352658
rect 99234 352338 99266 352574
rect 99502 352338 99586 352574
rect 99822 352338 99854 352574
rect 99234 316894 99854 352338
rect 99234 316658 99266 316894
rect 99502 316658 99586 316894
rect 99822 316658 99854 316894
rect 99234 316574 99854 316658
rect 99234 316338 99266 316574
rect 99502 316338 99586 316574
rect 99822 316338 99854 316574
rect 99234 280894 99854 316338
rect 99234 280658 99266 280894
rect 99502 280658 99586 280894
rect 99822 280658 99854 280894
rect 99234 280574 99854 280658
rect 99234 280338 99266 280574
rect 99502 280338 99586 280574
rect 99822 280338 99854 280574
rect 99234 244894 99854 280338
rect 99234 244658 99266 244894
rect 99502 244658 99586 244894
rect 99822 244658 99854 244894
rect 99234 244574 99854 244658
rect 99234 244338 99266 244574
rect 99502 244338 99586 244574
rect 99822 244338 99854 244574
rect 99234 208894 99854 244338
rect 99234 208658 99266 208894
rect 99502 208658 99586 208894
rect 99822 208658 99854 208894
rect 99234 208574 99854 208658
rect 99234 208338 99266 208574
rect 99502 208338 99586 208574
rect 99822 208338 99854 208574
rect 99234 172894 99854 208338
rect 99234 172658 99266 172894
rect 99502 172658 99586 172894
rect 99822 172658 99854 172894
rect 99234 172574 99854 172658
rect 99234 172338 99266 172574
rect 99502 172338 99586 172574
rect 99822 172338 99854 172574
rect 99234 136894 99854 172338
rect 99234 136658 99266 136894
rect 99502 136658 99586 136894
rect 99822 136658 99854 136894
rect 99234 136574 99854 136658
rect 99234 136338 99266 136574
rect 99502 136338 99586 136574
rect 99822 136338 99854 136574
rect 99234 100894 99854 136338
rect 99234 100658 99266 100894
rect 99502 100658 99586 100894
rect 99822 100658 99854 100894
rect 99234 100574 99854 100658
rect 99234 100338 99266 100574
rect 99502 100338 99586 100574
rect 99822 100338 99854 100574
rect 99234 64894 99854 100338
rect 99234 64658 99266 64894
rect 99502 64658 99586 64894
rect 99822 64658 99854 64894
rect 99234 64574 99854 64658
rect 99234 64338 99266 64574
rect 99502 64338 99586 64574
rect 99822 64338 99854 64574
rect 99234 28894 99854 64338
rect 99234 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 99854 28894
rect 99234 28574 99854 28658
rect 99234 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 99854 28574
rect 99234 -5146 99854 28338
rect 99234 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 99854 -5146
rect 99234 -5466 99854 -5382
rect 99234 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 99854 -5466
rect 99234 -5734 99854 -5702
rect 102954 680614 103574 711002
rect 120954 710598 121574 711590
rect 120954 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 121574 710598
rect 120954 710278 121574 710362
rect 120954 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 121574 710278
rect 117234 708678 117854 709670
rect 117234 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 117854 708678
rect 117234 708358 117854 708442
rect 117234 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 117854 708358
rect 113514 706758 114134 707750
rect 113514 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 114134 706758
rect 113514 706438 114134 706522
rect 113514 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 114134 706438
rect 102954 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 103574 680614
rect 102954 680294 103574 680378
rect 102954 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 103574 680294
rect 102954 644614 103574 680058
rect 102954 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 103574 644614
rect 102954 644294 103574 644378
rect 102954 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 103574 644294
rect 102954 608614 103574 644058
rect 102954 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 103574 608614
rect 102954 608294 103574 608378
rect 102954 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 103574 608294
rect 102954 572614 103574 608058
rect 102954 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 103574 572614
rect 102954 572294 103574 572378
rect 102954 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 103574 572294
rect 102954 536614 103574 572058
rect 102954 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 103574 536614
rect 102954 536294 103574 536378
rect 102954 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 103574 536294
rect 102954 500614 103574 536058
rect 102954 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 103574 500614
rect 102954 500294 103574 500378
rect 102954 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 103574 500294
rect 102954 464614 103574 500058
rect 102954 464378 102986 464614
rect 103222 464378 103306 464614
rect 103542 464378 103574 464614
rect 102954 464294 103574 464378
rect 102954 464058 102986 464294
rect 103222 464058 103306 464294
rect 103542 464058 103574 464294
rect 102954 428614 103574 464058
rect 102954 428378 102986 428614
rect 103222 428378 103306 428614
rect 103542 428378 103574 428614
rect 102954 428294 103574 428378
rect 102954 428058 102986 428294
rect 103222 428058 103306 428294
rect 103542 428058 103574 428294
rect 102954 392614 103574 428058
rect 102954 392378 102986 392614
rect 103222 392378 103306 392614
rect 103542 392378 103574 392614
rect 102954 392294 103574 392378
rect 102954 392058 102986 392294
rect 103222 392058 103306 392294
rect 103542 392058 103574 392294
rect 102954 356614 103574 392058
rect 102954 356378 102986 356614
rect 103222 356378 103306 356614
rect 103542 356378 103574 356614
rect 102954 356294 103574 356378
rect 102954 356058 102986 356294
rect 103222 356058 103306 356294
rect 103542 356058 103574 356294
rect 102954 320614 103574 356058
rect 102954 320378 102986 320614
rect 103222 320378 103306 320614
rect 103542 320378 103574 320614
rect 102954 320294 103574 320378
rect 102954 320058 102986 320294
rect 103222 320058 103306 320294
rect 103542 320058 103574 320294
rect 102954 284614 103574 320058
rect 102954 284378 102986 284614
rect 103222 284378 103306 284614
rect 103542 284378 103574 284614
rect 102954 284294 103574 284378
rect 102954 284058 102986 284294
rect 103222 284058 103306 284294
rect 103542 284058 103574 284294
rect 102954 248614 103574 284058
rect 102954 248378 102986 248614
rect 103222 248378 103306 248614
rect 103542 248378 103574 248614
rect 102954 248294 103574 248378
rect 102954 248058 102986 248294
rect 103222 248058 103306 248294
rect 103542 248058 103574 248294
rect 102954 212614 103574 248058
rect 102954 212378 102986 212614
rect 103222 212378 103306 212614
rect 103542 212378 103574 212614
rect 102954 212294 103574 212378
rect 102954 212058 102986 212294
rect 103222 212058 103306 212294
rect 103542 212058 103574 212294
rect 102954 176614 103574 212058
rect 102954 176378 102986 176614
rect 103222 176378 103306 176614
rect 103542 176378 103574 176614
rect 102954 176294 103574 176378
rect 102954 176058 102986 176294
rect 103222 176058 103306 176294
rect 103542 176058 103574 176294
rect 102954 140614 103574 176058
rect 102954 140378 102986 140614
rect 103222 140378 103306 140614
rect 103542 140378 103574 140614
rect 102954 140294 103574 140378
rect 102954 140058 102986 140294
rect 103222 140058 103306 140294
rect 103542 140058 103574 140294
rect 102954 104614 103574 140058
rect 102954 104378 102986 104614
rect 103222 104378 103306 104614
rect 103542 104378 103574 104614
rect 102954 104294 103574 104378
rect 102954 104058 102986 104294
rect 103222 104058 103306 104294
rect 103542 104058 103574 104294
rect 102954 68614 103574 104058
rect 102954 68378 102986 68614
rect 103222 68378 103306 68614
rect 103542 68378 103574 68614
rect 102954 68294 103574 68378
rect 102954 68058 102986 68294
rect 103222 68058 103306 68294
rect 103542 68058 103574 68294
rect 102954 32614 103574 68058
rect 102954 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 103574 32614
rect 102954 32294 103574 32378
rect 102954 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 103574 32294
rect 84954 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 85574 -6106
rect 84954 -6426 85574 -6342
rect 84954 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 85574 -6426
rect 84954 -7654 85574 -6662
rect 102954 -7066 103574 32058
rect 109794 704838 110414 705830
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 109794 543454 110414 578898
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 109794 507454 110414 542898
rect 109794 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 110414 507454
rect 109794 507134 110414 507218
rect 109794 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 110414 507134
rect 109794 471454 110414 506898
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 109794 435454 110414 470898
rect 109794 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 110414 435454
rect 109794 435134 110414 435218
rect 109794 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 110414 435134
rect 109794 399454 110414 434898
rect 109794 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 110414 399454
rect 109794 399134 110414 399218
rect 109794 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 110414 399134
rect 109794 363454 110414 398898
rect 109794 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 110414 363454
rect 109794 363134 110414 363218
rect 109794 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 110414 363134
rect 109794 327454 110414 362898
rect 109794 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 110414 327454
rect 109794 327134 110414 327218
rect 109794 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 110414 327134
rect 109794 291454 110414 326898
rect 109794 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 110414 291454
rect 109794 291134 110414 291218
rect 109794 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 110414 291134
rect 109794 255454 110414 290898
rect 109794 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 110414 255454
rect 109794 255134 110414 255218
rect 109794 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 110414 255134
rect 109794 219454 110414 254898
rect 109794 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 110414 219454
rect 109794 219134 110414 219218
rect 109794 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 110414 219134
rect 109794 183454 110414 218898
rect 109794 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 110414 183454
rect 109794 183134 110414 183218
rect 109794 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 110414 183134
rect 109794 147454 110414 182898
rect 109794 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 110414 147454
rect 109794 147134 110414 147218
rect 109794 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 110414 147134
rect 109794 111454 110414 146898
rect 109794 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 110414 111454
rect 109794 111134 110414 111218
rect 109794 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 110414 111134
rect 109794 75454 110414 110898
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 109794 75134 110414 75218
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 109794 39454 110414 74898
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -1894 110414 -902
rect 113514 691174 114134 706202
rect 113514 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 114134 691174
rect 113514 690854 114134 690938
rect 113514 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 114134 690854
rect 113514 655174 114134 690618
rect 113514 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 114134 655174
rect 113514 654854 114134 654938
rect 113514 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 114134 654854
rect 113514 619174 114134 654618
rect 113514 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 114134 619174
rect 113514 618854 114134 618938
rect 113514 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 114134 618854
rect 113514 583174 114134 618618
rect 113514 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 114134 583174
rect 113514 582854 114134 582938
rect 113514 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 114134 582854
rect 113514 547174 114134 582618
rect 113514 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 114134 547174
rect 113514 546854 114134 546938
rect 113514 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 114134 546854
rect 113514 511174 114134 546618
rect 113514 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 114134 511174
rect 113514 510854 114134 510938
rect 113514 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 114134 510854
rect 113514 475174 114134 510618
rect 113514 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 114134 475174
rect 113514 474854 114134 474938
rect 113514 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 114134 474854
rect 113514 439174 114134 474618
rect 113514 438938 113546 439174
rect 113782 438938 113866 439174
rect 114102 438938 114134 439174
rect 113514 438854 114134 438938
rect 113514 438618 113546 438854
rect 113782 438618 113866 438854
rect 114102 438618 114134 438854
rect 113514 403174 114134 438618
rect 113514 402938 113546 403174
rect 113782 402938 113866 403174
rect 114102 402938 114134 403174
rect 113514 402854 114134 402938
rect 113514 402618 113546 402854
rect 113782 402618 113866 402854
rect 114102 402618 114134 402854
rect 113514 367174 114134 402618
rect 113514 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 114134 367174
rect 113514 366854 114134 366938
rect 113514 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 114134 366854
rect 113514 331174 114134 366618
rect 113514 330938 113546 331174
rect 113782 330938 113866 331174
rect 114102 330938 114134 331174
rect 113514 330854 114134 330938
rect 113514 330618 113546 330854
rect 113782 330618 113866 330854
rect 114102 330618 114134 330854
rect 113514 295174 114134 330618
rect 113514 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 114134 295174
rect 113514 294854 114134 294938
rect 113514 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 114134 294854
rect 113514 259174 114134 294618
rect 113514 258938 113546 259174
rect 113782 258938 113866 259174
rect 114102 258938 114134 259174
rect 113514 258854 114134 258938
rect 113514 258618 113546 258854
rect 113782 258618 113866 258854
rect 114102 258618 114134 258854
rect 113514 223174 114134 258618
rect 113514 222938 113546 223174
rect 113782 222938 113866 223174
rect 114102 222938 114134 223174
rect 113514 222854 114134 222938
rect 113514 222618 113546 222854
rect 113782 222618 113866 222854
rect 114102 222618 114134 222854
rect 113514 187174 114134 222618
rect 113514 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 114134 187174
rect 113514 186854 114134 186938
rect 113514 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 114134 186854
rect 113514 151174 114134 186618
rect 113514 150938 113546 151174
rect 113782 150938 113866 151174
rect 114102 150938 114134 151174
rect 113514 150854 114134 150938
rect 113514 150618 113546 150854
rect 113782 150618 113866 150854
rect 114102 150618 114134 150854
rect 113514 115174 114134 150618
rect 113514 114938 113546 115174
rect 113782 114938 113866 115174
rect 114102 114938 114134 115174
rect 113514 114854 114134 114938
rect 113514 114618 113546 114854
rect 113782 114618 113866 114854
rect 114102 114618 114134 114854
rect 113514 79174 114134 114618
rect 113514 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 114134 79174
rect 113514 78854 114134 78938
rect 113514 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 114134 78854
rect 113514 43174 114134 78618
rect 113514 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 114134 43174
rect 113514 42854 114134 42938
rect 113514 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 114134 42854
rect 113514 7174 114134 42618
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 113514 -2266 114134 6618
rect 113514 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 114134 -2266
rect 113514 -2586 114134 -2502
rect 113514 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 114134 -2586
rect 113514 -3814 114134 -2822
rect 117234 694894 117854 708122
rect 117234 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 117854 694894
rect 117234 694574 117854 694658
rect 117234 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 117854 694574
rect 117234 658894 117854 694338
rect 117234 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 117854 658894
rect 117234 658574 117854 658658
rect 117234 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 117854 658574
rect 117234 622894 117854 658338
rect 117234 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 117854 622894
rect 117234 622574 117854 622658
rect 117234 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 117854 622574
rect 117234 586894 117854 622338
rect 117234 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 117854 586894
rect 117234 586574 117854 586658
rect 117234 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 117854 586574
rect 117234 550894 117854 586338
rect 117234 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 117854 550894
rect 117234 550574 117854 550658
rect 117234 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 117854 550574
rect 117234 514894 117854 550338
rect 117234 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 117854 514894
rect 117234 514574 117854 514658
rect 117234 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 117854 514574
rect 117234 478894 117854 514338
rect 117234 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 117854 478894
rect 117234 478574 117854 478658
rect 117234 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 117854 478574
rect 117234 442894 117854 478338
rect 117234 442658 117266 442894
rect 117502 442658 117586 442894
rect 117822 442658 117854 442894
rect 117234 442574 117854 442658
rect 117234 442338 117266 442574
rect 117502 442338 117586 442574
rect 117822 442338 117854 442574
rect 117234 406894 117854 442338
rect 117234 406658 117266 406894
rect 117502 406658 117586 406894
rect 117822 406658 117854 406894
rect 117234 406574 117854 406658
rect 117234 406338 117266 406574
rect 117502 406338 117586 406574
rect 117822 406338 117854 406574
rect 117234 370894 117854 406338
rect 117234 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 117854 370894
rect 117234 370574 117854 370658
rect 117234 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 117854 370574
rect 117234 334894 117854 370338
rect 117234 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 117854 334894
rect 117234 334574 117854 334658
rect 117234 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 117854 334574
rect 117234 298894 117854 334338
rect 117234 298658 117266 298894
rect 117502 298658 117586 298894
rect 117822 298658 117854 298894
rect 117234 298574 117854 298658
rect 117234 298338 117266 298574
rect 117502 298338 117586 298574
rect 117822 298338 117854 298574
rect 117234 262894 117854 298338
rect 117234 262658 117266 262894
rect 117502 262658 117586 262894
rect 117822 262658 117854 262894
rect 117234 262574 117854 262658
rect 117234 262338 117266 262574
rect 117502 262338 117586 262574
rect 117822 262338 117854 262574
rect 117234 226894 117854 262338
rect 117234 226658 117266 226894
rect 117502 226658 117586 226894
rect 117822 226658 117854 226894
rect 117234 226574 117854 226658
rect 117234 226338 117266 226574
rect 117502 226338 117586 226574
rect 117822 226338 117854 226574
rect 117234 190894 117854 226338
rect 117234 190658 117266 190894
rect 117502 190658 117586 190894
rect 117822 190658 117854 190894
rect 117234 190574 117854 190658
rect 117234 190338 117266 190574
rect 117502 190338 117586 190574
rect 117822 190338 117854 190574
rect 117234 154894 117854 190338
rect 117234 154658 117266 154894
rect 117502 154658 117586 154894
rect 117822 154658 117854 154894
rect 117234 154574 117854 154658
rect 117234 154338 117266 154574
rect 117502 154338 117586 154574
rect 117822 154338 117854 154574
rect 117234 118894 117854 154338
rect 117234 118658 117266 118894
rect 117502 118658 117586 118894
rect 117822 118658 117854 118894
rect 117234 118574 117854 118658
rect 117234 118338 117266 118574
rect 117502 118338 117586 118574
rect 117822 118338 117854 118574
rect 117234 82894 117854 118338
rect 117234 82658 117266 82894
rect 117502 82658 117586 82894
rect 117822 82658 117854 82894
rect 117234 82574 117854 82658
rect 117234 82338 117266 82574
rect 117502 82338 117586 82574
rect 117822 82338 117854 82574
rect 117234 46894 117854 82338
rect 117234 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 117854 46894
rect 117234 46574 117854 46658
rect 117234 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 117854 46574
rect 117234 10894 117854 46338
rect 117234 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 117854 10894
rect 117234 10574 117854 10658
rect 117234 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 117854 10574
rect 117234 -4186 117854 10338
rect 117234 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 117854 -4186
rect 117234 -4506 117854 -4422
rect 117234 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 117854 -4506
rect 117234 -5734 117854 -4742
rect 120954 698614 121574 710042
rect 138954 711558 139574 711590
rect 138954 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 139574 711558
rect 138954 711238 139574 711322
rect 138954 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 139574 711238
rect 135234 709638 135854 709670
rect 135234 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 135854 709638
rect 135234 709318 135854 709402
rect 135234 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 135854 709318
rect 131514 707718 132134 707750
rect 131514 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 132134 707718
rect 131514 707398 132134 707482
rect 131514 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 132134 707398
rect 120954 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 121574 698614
rect 120954 698294 121574 698378
rect 120954 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 121574 698294
rect 120954 662614 121574 698058
rect 120954 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 121574 662614
rect 120954 662294 121574 662378
rect 120954 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 121574 662294
rect 120954 626614 121574 662058
rect 120954 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 121574 626614
rect 120954 626294 121574 626378
rect 120954 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 121574 626294
rect 120954 590614 121574 626058
rect 120954 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 121574 590614
rect 120954 590294 121574 590378
rect 120954 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 121574 590294
rect 120954 554614 121574 590058
rect 120954 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 121574 554614
rect 120954 554294 121574 554378
rect 120954 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 121574 554294
rect 120954 518614 121574 554058
rect 120954 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 121574 518614
rect 120954 518294 121574 518378
rect 120954 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 121574 518294
rect 120954 482614 121574 518058
rect 120954 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 121574 482614
rect 120954 482294 121574 482378
rect 120954 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 121574 482294
rect 120954 446614 121574 482058
rect 120954 446378 120986 446614
rect 121222 446378 121306 446614
rect 121542 446378 121574 446614
rect 120954 446294 121574 446378
rect 120954 446058 120986 446294
rect 121222 446058 121306 446294
rect 121542 446058 121574 446294
rect 120954 410614 121574 446058
rect 120954 410378 120986 410614
rect 121222 410378 121306 410614
rect 121542 410378 121574 410614
rect 120954 410294 121574 410378
rect 120954 410058 120986 410294
rect 121222 410058 121306 410294
rect 121542 410058 121574 410294
rect 120954 374614 121574 410058
rect 120954 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 121574 374614
rect 120954 374294 121574 374378
rect 120954 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 121574 374294
rect 120954 338614 121574 374058
rect 120954 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 121574 338614
rect 120954 338294 121574 338378
rect 120954 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 121574 338294
rect 120954 302614 121574 338058
rect 120954 302378 120986 302614
rect 121222 302378 121306 302614
rect 121542 302378 121574 302614
rect 120954 302294 121574 302378
rect 120954 302058 120986 302294
rect 121222 302058 121306 302294
rect 121542 302058 121574 302294
rect 120954 266614 121574 302058
rect 120954 266378 120986 266614
rect 121222 266378 121306 266614
rect 121542 266378 121574 266614
rect 120954 266294 121574 266378
rect 120954 266058 120986 266294
rect 121222 266058 121306 266294
rect 121542 266058 121574 266294
rect 120954 230614 121574 266058
rect 120954 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 121574 230614
rect 120954 230294 121574 230378
rect 120954 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 121574 230294
rect 120954 194614 121574 230058
rect 120954 194378 120986 194614
rect 121222 194378 121306 194614
rect 121542 194378 121574 194614
rect 120954 194294 121574 194378
rect 120954 194058 120986 194294
rect 121222 194058 121306 194294
rect 121542 194058 121574 194294
rect 120954 158614 121574 194058
rect 120954 158378 120986 158614
rect 121222 158378 121306 158614
rect 121542 158378 121574 158614
rect 120954 158294 121574 158378
rect 120954 158058 120986 158294
rect 121222 158058 121306 158294
rect 121542 158058 121574 158294
rect 120954 122614 121574 158058
rect 120954 122378 120986 122614
rect 121222 122378 121306 122614
rect 121542 122378 121574 122614
rect 120954 122294 121574 122378
rect 120954 122058 120986 122294
rect 121222 122058 121306 122294
rect 121542 122058 121574 122294
rect 120954 86614 121574 122058
rect 120954 86378 120986 86614
rect 121222 86378 121306 86614
rect 121542 86378 121574 86614
rect 120954 86294 121574 86378
rect 120954 86058 120986 86294
rect 121222 86058 121306 86294
rect 121542 86058 121574 86294
rect 120954 50614 121574 86058
rect 120954 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 121574 50614
rect 120954 50294 121574 50378
rect 120954 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 121574 50294
rect 120954 14614 121574 50058
rect 120954 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 121574 14614
rect 120954 14294 121574 14378
rect 120954 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 121574 14294
rect 102954 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 103574 -7066
rect 102954 -7386 103574 -7302
rect 102954 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 103574 -7386
rect 102954 -7654 103574 -7622
rect 120954 -6106 121574 14058
rect 127794 705798 128414 705830
rect 127794 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 128414 705798
rect 127794 705478 128414 705562
rect 127794 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 128414 705478
rect 127794 669454 128414 705242
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 127794 561454 128414 596898
rect 127794 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 128414 561454
rect 127794 561134 128414 561218
rect 127794 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 128414 561134
rect 127794 525454 128414 560898
rect 127794 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 128414 525454
rect 127794 525134 128414 525218
rect 127794 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 128414 525134
rect 127794 489454 128414 524898
rect 127794 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 128414 489454
rect 127794 489134 128414 489218
rect 127794 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 128414 489134
rect 127794 453454 128414 488898
rect 127794 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 128414 453454
rect 127794 453134 128414 453218
rect 127794 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 128414 453134
rect 127794 417454 128414 452898
rect 127794 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 128414 417454
rect 127794 417134 128414 417218
rect 127794 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 128414 417134
rect 127794 381454 128414 416898
rect 127794 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 128414 381454
rect 127794 381134 128414 381218
rect 127794 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 128414 381134
rect 127794 345454 128414 380898
rect 127794 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 128414 345454
rect 127794 345134 128414 345218
rect 127794 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 128414 345134
rect 127794 309454 128414 344898
rect 127794 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 128414 309454
rect 127794 309134 128414 309218
rect 127794 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 128414 309134
rect 127794 273454 128414 308898
rect 127794 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 128414 273454
rect 127794 273134 128414 273218
rect 127794 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 128414 273134
rect 127794 237454 128414 272898
rect 127794 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 128414 237454
rect 127794 237134 128414 237218
rect 127794 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 128414 237134
rect 127794 201454 128414 236898
rect 127794 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 128414 201454
rect 127794 201134 128414 201218
rect 127794 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 128414 201134
rect 127794 165454 128414 200898
rect 127794 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 128414 165454
rect 127794 165134 128414 165218
rect 127794 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 128414 165134
rect 127794 129454 128414 164898
rect 127794 129218 127826 129454
rect 128062 129218 128146 129454
rect 128382 129218 128414 129454
rect 127794 129134 128414 129218
rect 127794 128898 127826 129134
rect 128062 128898 128146 129134
rect 128382 128898 128414 129134
rect 127794 93454 128414 128898
rect 127794 93218 127826 93454
rect 128062 93218 128146 93454
rect 128382 93218 128414 93454
rect 127794 93134 128414 93218
rect 127794 92898 127826 93134
rect 128062 92898 128146 93134
rect 128382 92898 128414 93134
rect 127794 57454 128414 92898
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -1306 128414 20898
rect 127794 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 128414 -1306
rect 127794 -1626 128414 -1542
rect 127794 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 128414 -1626
rect 127794 -1894 128414 -1862
rect 131514 673174 132134 707162
rect 131514 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 132134 673174
rect 131514 672854 132134 672938
rect 131514 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 132134 672854
rect 131514 637174 132134 672618
rect 131514 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 132134 637174
rect 131514 636854 132134 636938
rect 131514 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 132134 636854
rect 131514 601174 132134 636618
rect 131514 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 132134 601174
rect 131514 600854 132134 600938
rect 131514 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 132134 600854
rect 131514 565174 132134 600618
rect 131514 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 132134 565174
rect 131514 564854 132134 564938
rect 131514 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 132134 564854
rect 131514 529174 132134 564618
rect 131514 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 132134 529174
rect 131514 528854 132134 528938
rect 131514 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 132134 528854
rect 131514 493174 132134 528618
rect 131514 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 132134 493174
rect 131514 492854 132134 492938
rect 131514 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 132134 492854
rect 131514 457174 132134 492618
rect 131514 456938 131546 457174
rect 131782 456938 131866 457174
rect 132102 456938 132134 457174
rect 131514 456854 132134 456938
rect 131514 456618 131546 456854
rect 131782 456618 131866 456854
rect 132102 456618 132134 456854
rect 131514 421174 132134 456618
rect 131514 420938 131546 421174
rect 131782 420938 131866 421174
rect 132102 420938 132134 421174
rect 131514 420854 132134 420938
rect 131514 420618 131546 420854
rect 131782 420618 131866 420854
rect 132102 420618 132134 420854
rect 131514 385174 132134 420618
rect 131514 384938 131546 385174
rect 131782 384938 131866 385174
rect 132102 384938 132134 385174
rect 131514 384854 132134 384938
rect 131514 384618 131546 384854
rect 131782 384618 131866 384854
rect 132102 384618 132134 384854
rect 131514 349174 132134 384618
rect 131514 348938 131546 349174
rect 131782 348938 131866 349174
rect 132102 348938 132134 349174
rect 131514 348854 132134 348938
rect 131514 348618 131546 348854
rect 131782 348618 131866 348854
rect 132102 348618 132134 348854
rect 131514 313174 132134 348618
rect 131514 312938 131546 313174
rect 131782 312938 131866 313174
rect 132102 312938 132134 313174
rect 131514 312854 132134 312938
rect 131514 312618 131546 312854
rect 131782 312618 131866 312854
rect 132102 312618 132134 312854
rect 131514 277174 132134 312618
rect 131514 276938 131546 277174
rect 131782 276938 131866 277174
rect 132102 276938 132134 277174
rect 131514 276854 132134 276938
rect 131514 276618 131546 276854
rect 131782 276618 131866 276854
rect 132102 276618 132134 276854
rect 131514 241174 132134 276618
rect 131514 240938 131546 241174
rect 131782 240938 131866 241174
rect 132102 240938 132134 241174
rect 131514 240854 132134 240938
rect 131514 240618 131546 240854
rect 131782 240618 131866 240854
rect 132102 240618 132134 240854
rect 131514 205174 132134 240618
rect 131514 204938 131546 205174
rect 131782 204938 131866 205174
rect 132102 204938 132134 205174
rect 131514 204854 132134 204938
rect 131514 204618 131546 204854
rect 131782 204618 131866 204854
rect 132102 204618 132134 204854
rect 131514 169174 132134 204618
rect 131514 168938 131546 169174
rect 131782 168938 131866 169174
rect 132102 168938 132134 169174
rect 131514 168854 132134 168938
rect 131514 168618 131546 168854
rect 131782 168618 131866 168854
rect 132102 168618 132134 168854
rect 131514 133174 132134 168618
rect 131514 132938 131546 133174
rect 131782 132938 131866 133174
rect 132102 132938 132134 133174
rect 131514 132854 132134 132938
rect 131514 132618 131546 132854
rect 131782 132618 131866 132854
rect 132102 132618 132134 132854
rect 131514 97174 132134 132618
rect 131514 96938 131546 97174
rect 131782 96938 131866 97174
rect 132102 96938 132134 97174
rect 131514 96854 132134 96938
rect 131514 96618 131546 96854
rect 131782 96618 131866 96854
rect 132102 96618 132134 96854
rect 131514 61174 132134 96618
rect 131514 60938 131546 61174
rect 131782 60938 131866 61174
rect 132102 60938 132134 61174
rect 131514 60854 132134 60938
rect 131514 60618 131546 60854
rect 131782 60618 131866 60854
rect 132102 60618 132134 60854
rect 131514 25174 132134 60618
rect 131514 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 132134 25174
rect 131514 24854 132134 24938
rect 131514 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 132134 24854
rect 131514 -3226 132134 24618
rect 131514 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 132134 -3226
rect 131514 -3546 132134 -3462
rect 131514 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 132134 -3546
rect 131514 -3814 132134 -3782
rect 135234 676894 135854 709082
rect 135234 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 135854 676894
rect 135234 676574 135854 676658
rect 135234 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 135854 676574
rect 135234 640894 135854 676338
rect 135234 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 135854 640894
rect 135234 640574 135854 640658
rect 135234 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 135854 640574
rect 135234 604894 135854 640338
rect 135234 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 135854 604894
rect 135234 604574 135854 604658
rect 135234 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 135854 604574
rect 135234 568894 135854 604338
rect 135234 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 135854 568894
rect 135234 568574 135854 568658
rect 135234 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 135854 568574
rect 135234 532894 135854 568338
rect 135234 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 135854 532894
rect 135234 532574 135854 532658
rect 135234 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 135854 532574
rect 135234 496894 135854 532338
rect 135234 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 135854 496894
rect 135234 496574 135854 496658
rect 135234 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 135854 496574
rect 135234 460894 135854 496338
rect 135234 460658 135266 460894
rect 135502 460658 135586 460894
rect 135822 460658 135854 460894
rect 135234 460574 135854 460658
rect 135234 460338 135266 460574
rect 135502 460338 135586 460574
rect 135822 460338 135854 460574
rect 135234 424894 135854 460338
rect 135234 424658 135266 424894
rect 135502 424658 135586 424894
rect 135822 424658 135854 424894
rect 135234 424574 135854 424658
rect 135234 424338 135266 424574
rect 135502 424338 135586 424574
rect 135822 424338 135854 424574
rect 135234 388894 135854 424338
rect 135234 388658 135266 388894
rect 135502 388658 135586 388894
rect 135822 388658 135854 388894
rect 135234 388574 135854 388658
rect 135234 388338 135266 388574
rect 135502 388338 135586 388574
rect 135822 388338 135854 388574
rect 135234 352894 135854 388338
rect 135234 352658 135266 352894
rect 135502 352658 135586 352894
rect 135822 352658 135854 352894
rect 135234 352574 135854 352658
rect 135234 352338 135266 352574
rect 135502 352338 135586 352574
rect 135822 352338 135854 352574
rect 135234 316894 135854 352338
rect 135234 316658 135266 316894
rect 135502 316658 135586 316894
rect 135822 316658 135854 316894
rect 135234 316574 135854 316658
rect 135234 316338 135266 316574
rect 135502 316338 135586 316574
rect 135822 316338 135854 316574
rect 135234 280894 135854 316338
rect 135234 280658 135266 280894
rect 135502 280658 135586 280894
rect 135822 280658 135854 280894
rect 135234 280574 135854 280658
rect 135234 280338 135266 280574
rect 135502 280338 135586 280574
rect 135822 280338 135854 280574
rect 135234 244894 135854 280338
rect 135234 244658 135266 244894
rect 135502 244658 135586 244894
rect 135822 244658 135854 244894
rect 135234 244574 135854 244658
rect 135234 244338 135266 244574
rect 135502 244338 135586 244574
rect 135822 244338 135854 244574
rect 135234 208894 135854 244338
rect 135234 208658 135266 208894
rect 135502 208658 135586 208894
rect 135822 208658 135854 208894
rect 135234 208574 135854 208658
rect 135234 208338 135266 208574
rect 135502 208338 135586 208574
rect 135822 208338 135854 208574
rect 135234 172894 135854 208338
rect 135234 172658 135266 172894
rect 135502 172658 135586 172894
rect 135822 172658 135854 172894
rect 135234 172574 135854 172658
rect 135234 172338 135266 172574
rect 135502 172338 135586 172574
rect 135822 172338 135854 172574
rect 135234 136894 135854 172338
rect 135234 136658 135266 136894
rect 135502 136658 135586 136894
rect 135822 136658 135854 136894
rect 135234 136574 135854 136658
rect 135234 136338 135266 136574
rect 135502 136338 135586 136574
rect 135822 136338 135854 136574
rect 135234 100894 135854 136338
rect 135234 100658 135266 100894
rect 135502 100658 135586 100894
rect 135822 100658 135854 100894
rect 135234 100574 135854 100658
rect 135234 100338 135266 100574
rect 135502 100338 135586 100574
rect 135822 100338 135854 100574
rect 135234 64894 135854 100338
rect 135234 64658 135266 64894
rect 135502 64658 135586 64894
rect 135822 64658 135854 64894
rect 135234 64574 135854 64658
rect 135234 64338 135266 64574
rect 135502 64338 135586 64574
rect 135822 64338 135854 64574
rect 135234 28894 135854 64338
rect 135234 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 135854 28894
rect 135234 28574 135854 28658
rect 135234 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 135854 28574
rect 135234 -5146 135854 28338
rect 135234 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 135854 -5146
rect 135234 -5466 135854 -5382
rect 135234 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 135854 -5466
rect 135234 -5734 135854 -5702
rect 138954 680614 139574 711002
rect 156954 710598 157574 711590
rect 156954 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 157574 710598
rect 156954 710278 157574 710362
rect 156954 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 157574 710278
rect 153234 708678 153854 709670
rect 153234 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 153854 708678
rect 153234 708358 153854 708442
rect 153234 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 153854 708358
rect 149514 706758 150134 707750
rect 149514 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 150134 706758
rect 149514 706438 150134 706522
rect 149514 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 150134 706438
rect 138954 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 139574 680614
rect 138954 680294 139574 680378
rect 138954 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 139574 680294
rect 138954 644614 139574 680058
rect 138954 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 139574 644614
rect 138954 644294 139574 644378
rect 138954 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 139574 644294
rect 138954 608614 139574 644058
rect 138954 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 139574 608614
rect 138954 608294 139574 608378
rect 138954 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 139574 608294
rect 138954 572614 139574 608058
rect 138954 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 139574 572614
rect 138954 572294 139574 572378
rect 138954 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 139574 572294
rect 138954 536614 139574 572058
rect 138954 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 139574 536614
rect 138954 536294 139574 536378
rect 138954 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 139574 536294
rect 138954 500614 139574 536058
rect 138954 500378 138986 500614
rect 139222 500378 139306 500614
rect 139542 500378 139574 500614
rect 138954 500294 139574 500378
rect 138954 500058 138986 500294
rect 139222 500058 139306 500294
rect 139542 500058 139574 500294
rect 138954 464614 139574 500058
rect 138954 464378 138986 464614
rect 139222 464378 139306 464614
rect 139542 464378 139574 464614
rect 138954 464294 139574 464378
rect 138954 464058 138986 464294
rect 139222 464058 139306 464294
rect 139542 464058 139574 464294
rect 138954 428614 139574 464058
rect 138954 428378 138986 428614
rect 139222 428378 139306 428614
rect 139542 428378 139574 428614
rect 138954 428294 139574 428378
rect 138954 428058 138986 428294
rect 139222 428058 139306 428294
rect 139542 428058 139574 428294
rect 138954 392614 139574 428058
rect 138954 392378 138986 392614
rect 139222 392378 139306 392614
rect 139542 392378 139574 392614
rect 138954 392294 139574 392378
rect 138954 392058 138986 392294
rect 139222 392058 139306 392294
rect 139542 392058 139574 392294
rect 138954 356614 139574 392058
rect 138954 356378 138986 356614
rect 139222 356378 139306 356614
rect 139542 356378 139574 356614
rect 138954 356294 139574 356378
rect 138954 356058 138986 356294
rect 139222 356058 139306 356294
rect 139542 356058 139574 356294
rect 138954 320614 139574 356058
rect 138954 320378 138986 320614
rect 139222 320378 139306 320614
rect 139542 320378 139574 320614
rect 138954 320294 139574 320378
rect 138954 320058 138986 320294
rect 139222 320058 139306 320294
rect 139542 320058 139574 320294
rect 138954 284614 139574 320058
rect 138954 284378 138986 284614
rect 139222 284378 139306 284614
rect 139542 284378 139574 284614
rect 138954 284294 139574 284378
rect 138954 284058 138986 284294
rect 139222 284058 139306 284294
rect 139542 284058 139574 284294
rect 138954 248614 139574 284058
rect 138954 248378 138986 248614
rect 139222 248378 139306 248614
rect 139542 248378 139574 248614
rect 138954 248294 139574 248378
rect 138954 248058 138986 248294
rect 139222 248058 139306 248294
rect 139542 248058 139574 248294
rect 138954 212614 139574 248058
rect 138954 212378 138986 212614
rect 139222 212378 139306 212614
rect 139542 212378 139574 212614
rect 138954 212294 139574 212378
rect 138954 212058 138986 212294
rect 139222 212058 139306 212294
rect 139542 212058 139574 212294
rect 138954 176614 139574 212058
rect 138954 176378 138986 176614
rect 139222 176378 139306 176614
rect 139542 176378 139574 176614
rect 138954 176294 139574 176378
rect 138954 176058 138986 176294
rect 139222 176058 139306 176294
rect 139542 176058 139574 176294
rect 138954 140614 139574 176058
rect 138954 140378 138986 140614
rect 139222 140378 139306 140614
rect 139542 140378 139574 140614
rect 138954 140294 139574 140378
rect 138954 140058 138986 140294
rect 139222 140058 139306 140294
rect 139542 140058 139574 140294
rect 138954 104614 139574 140058
rect 138954 104378 138986 104614
rect 139222 104378 139306 104614
rect 139542 104378 139574 104614
rect 138954 104294 139574 104378
rect 138954 104058 138986 104294
rect 139222 104058 139306 104294
rect 139542 104058 139574 104294
rect 138954 68614 139574 104058
rect 138954 68378 138986 68614
rect 139222 68378 139306 68614
rect 139542 68378 139574 68614
rect 138954 68294 139574 68378
rect 138954 68058 138986 68294
rect 139222 68058 139306 68294
rect 139542 68058 139574 68294
rect 138954 32614 139574 68058
rect 138954 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 139574 32614
rect 138954 32294 139574 32378
rect 138954 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 139574 32294
rect 120954 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 121574 -6106
rect 120954 -6426 121574 -6342
rect 120954 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 121574 -6426
rect 120954 -7654 121574 -6662
rect 138954 -7066 139574 32058
rect 145794 704838 146414 705830
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 543454 146414 578898
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 507454 146414 542898
rect 145794 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 146414 507454
rect 145794 507134 146414 507218
rect 145794 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 146414 507134
rect 145794 471454 146414 506898
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 435454 146414 470898
rect 145794 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 146414 435454
rect 145794 435134 146414 435218
rect 145794 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 146414 435134
rect 145794 399454 146414 434898
rect 145794 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 146414 399454
rect 145794 399134 146414 399218
rect 145794 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 146414 399134
rect 145794 363454 146414 398898
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 145794 327454 146414 362898
rect 145794 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 146414 327454
rect 145794 327134 146414 327218
rect 145794 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 146414 327134
rect 145794 291454 146414 326898
rect 145794 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 146414 291454
rect 145794 291134 146414 291218
rect 145794 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 146414 291134
rect 145794 255454 146414 290898
rect 145794 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 146414 255454
rect 145794 255134 146414 255218
rect 145794 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 146414 255134
rect 145794 219454 146414 254898
rect 145794 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 146414 219454
rect 145794 219134 146414 219218
rect 145794 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 146414 219134
rect 145794 183454 146414 218898
rect 145794 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 146414 183454
rect 145794 183134 146414 183218
rect 145794 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 146414 183134
rect 145794 147454 146414 182898
rect 145794 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 146414 147454
rect 145794 147134 146414 147218
rect 145794 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 146414 147134
rect 145794 111454 146414 146898
rect 145794 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 146414 111454
rect 145794 111134 146414 111218
rect 145794 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 146414 111134
rect 145794 75454 146414 110898
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145794 75134 146414 75218
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 145794 39454 146414 74898
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -1894 146414 -902
rect 149514 691174 150134 706202
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 655174 150134 690618
rect 149514 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 150134 655174
rect 149514 654854 150134 654938
rect 149514 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 150134 654854
rect 149514 619174 150134 654618
rect 149514 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 150134 619174
rect 149514 618854 150134 618938
rect 149514 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 150134 618854
rect 149514 583174 150134 618618
rect 149514 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 150134 583174
rect 149514 582854 150134 582938
rect 149514 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 150134 582854
rect 149514 547174 150134 582618
rect 149514 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 150134 547174
rect 149514 546854 150134 546938
rect 149514 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 150134 546854
rect 149514 511174 150134 546618
rect 149514 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 150134 511174
rect 149514 510854 150134 510938
rect 149514 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 150134 510854
rect 149514 475174 150134 510618
rect 149514 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 150134 475174
rect 149514 474854 150134 474938
rect 149514 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 150134 474854
rect 149514 439174 150134 474618
rect 149514 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 150134 439174
rect 149514 438854 150134 438938
rect 149514 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 150134 438854
rect 149514 403174 150134 438618
rect 149514 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 150134 403174
rect 149514 402854 150134 402938
rect 149514 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 150134 402854
rect 149514 367174 150134 402618
rect 149514 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 150134 367174
rect 149514 366854 150134 366938
rect 149514 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 150134 366854
rect 149514 331174 150134 366618
rect 149514 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 150134 331174
rect 149514 330854 150134 330938
rect 149514 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 150134 330854
rect 149514 295174 150134 330618
rect 149514 294938 149546 295174
rect 149782 294938 149866 295174
rect 150102 294938 150134 295174
rect 149514 294854 150134 294938
rect 149514 294618 149546 294854
rect 149782 294618 149866 294854
rect 150102 294618 150134 294854
rect 149514 259174 150134 294618
rect 149514 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 150134 259174
rect 149514 258854 150134 258938
rect 149514 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 150134 258854
rect 149514 223174 150134 258618
rect 149514 222938 149546 223174
rect 149782 222938 149866 223174
rect 150102 222938 150134 223174
rect 149514 222854 150134 222938
rect 149514 222618 149546 222854
rect 149782 222618 149866 222854
rect 150102 222618 150134 222854
rect 149514 187174 150134 222618
rect 149514 186938 149546 187174
rect 149782 186938 149866 187174
rect 150102 186938 150134 187174
rect 149514 186854 150134 186938
rect 149514 186618 149546 186854
rect 149782 186618 149866 186854
rect 150102 186618 150134 186854
rect 149514 151174 150134 186618
rect 149514 150938 149546 151174
rect 149782 150938 149866 151174
rect 150102 150938 150134 151174
rect 149514 150854 150134 150938
rect 149514 150618 149546 150854
rect 149782 150618 149866 150854
rect 150102 150618 150134 150854
rect 149514 115174 150134 150618
rect 149514 114938 149546 115174
rect 149782 114938 149866 115174
rect 150102 114938 150134 115174
rect 149514 114854 150134 114938
rect 149514 114618 149546 114854
rect 149782 114618 149866 114854
rect 150102 114618 150134 114854
rect 149514 79174 150134 114618
rect 149514 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 150134 79174
rect 149514 78854 150134 78938
rect 149514 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 150134 78854
rect 149514 43174 150134 78618
rect 149514 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 150134 43174
rect 149514 42854 150134 42938
rect 149514 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 150134 42854
rect 149514 7174 150134 42618
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 149514 -2266 150134 6618
rect 149514 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 150134 -2266
rect 149514 -2586 150134 -2502
rect 149514 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 150134 -2586
rect 149514 -3814 150134 -2822
rect 153234 694894 153854 708122
rect 153234 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 153854 694894
rect 153234 694574 153854 694658
rect 153234 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 153854 694574
rect 153234 658894 153854 694338
rect 153234 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 153854 658894
rect 153234 658574 153854 658658
rect 153234 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 153854 658574
rect 153234 622894 153854 658338
rect 153234 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 153854 622894
rect 153234 622574 153854 622658
rect 153234 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 153854 622574
rect 153234 586894 153854 622338
rect 153234 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 153854 586894
rect 153234 586574 153854 586658
rect 153234 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 153854 586574
rect 153234 550894 153854 586338
rect 153234 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 153854 550894
rect 153234 550574 153854 550658
rect 153234 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 153854 550574
rect 153234 514894 153854 550338
rect 153234 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 153854 514894
rect 153234 514574 153854 514658
rect 153234 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 153854 514574
rect 153234 478894 153854 514338
rect 153234 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 153854 478894
rect 153234 478574 153854 478658
rect 153234 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 153854 478574
rect 153234 442894 153854 478338
rect 153234 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 153854 442894
rect 153234 442574 153854 442658
rect 153234 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 153854 442574
rect 153234 406894 153854 442338
rect 153234 406658 153266 406894
rect 153502 406658 153586 406894
rect 153822 406658 153854 406894
rect 153234 406574 153854 406658
rect 153234 406338 153266 406574
rect 153502 406338 153586 406574
rect 153822 406338 153854 406574
rect 153234 370894 153854 406338
rect 153234 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 153854 370894
rect 153234 370574 153854 370658
rect 153234 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 153854 370574
rect 153234 334894 153854 370338
rect 153234 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 153854 334894
rect 153234 334574 153854 334658
rect 153234 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 153854 334574
rect 153234 298894 153854 334338
rect 153234 298658 153266 298894
rect 153502 298658 153586 298894
rect 153822 298658 153854 298894
rect 153234 298574 153854 298658
rect 153234 298338 153266 298574
rect 153502 298338 153586 298574
rect 153822 298338 153854 298574
rect 153234 262894 153854 298338
rect 153234 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 153854 262894
rect 153234 262574 153854 262658
rect 153234 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 153854 262574
rect 153234 226894 153854 262338
rect 153234 226658 153266 226894
rect 153502 226658 153586 226894
rect 153822 226658 153854 226894
rect 153234 226574 153854 226658
rect 153234 226338 153266 226574
rect 153502 226338 153586 226574
rect 153822 226338 153854 226574
rect 153234 190894 153854 226338
rect 153234 190658 153266 190894
rect 153502 190658 153586 190894
rect 153822 190658 153854 190894
rect 153234 190574 153854 190658
rect 153234 190338 153266 190574
rect 153502 190338 153586 190574
rect 153822 190338 153854 190574
rect 153234 154894 153854 190338
rect 153234 154658 153266 154894
rect 153502 154658 153586 154894
rect 153822 154658 153854 154894
rect 153234 154574 153854 154658
rect 153234 154338 153266 154574
rect 153502 154338 153586 154574
rect 153822 154338 153854 154574
rect 153234 118894 153854 154338
rect 153234 118658 153266 118894
rect 153502 118658 153586 118894
rect 153822 118658 153854 118894
rect 153234 118574 153854 118658
rect 153234 118338 153266 118574
rect 153502 118338 153586 118574
rect 153822 118338 153854 118574
rect 153234 82894 153854 118338
rect 153234 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 153854 82894
rect 153234 82574 153854 82658
rect 153234 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 153854 82574
rect 153234 46894 153854 82338
rect 153234 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 153854 46894
rect 153234 46574 153854 46658
rect 153234 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 153854 46574
rect 153234 10894 153854 46338
rect 153234 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 153854 10894
rect 153234 10574 153854 10658
rect 153234 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 153854 10574
rect 153234 -4186 153854 10338
rect 153234 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 153854 -4186
rect 153234 -4506 153854 -4422
rect 153234 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 153854 -4506
rect 153234 -5734 153854 -4742
rect 156954 698614 157574 710042
rect 174954 711558 175574 711590
rect 174954 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 175574 711558
rect 174954 711238 175574 711322
rect 174954 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 175574 711238
rect 171234 709638 171854 709670
rect 171234 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 171854 709638
rect 171234 709318 171854 709402
rect 171234 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 171854 709318
rect 167514 707718 168134 707750
rect 167514 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 168134 707718
rect 167514 707398 168134 707482
rect 167514 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 168134 707398
rect 156954 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 157574 698614
rect 156954 698294 157574 698378
rect 156954 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 157574 698294
rect 156954 662614 157574 698058
rect 156954 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 157574 662614
rect 156954 662294 157574 662378
rect 156954 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 157574 662294
rect 156954 626614 157574 662058
rect 156954 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 157574 626614
rect 156954 626294 157574 626378
rect 156954 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 157574 626294
rect 156954 590614 157574 626058
rect 156954 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 157574 590614
rect 156954 590294 157574 590378
rect 156954 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 157574 590294
rect 156954 554614 157574 590058
rect 156954 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 157574 554614
rect 156954 554294 157574 554378
rect 156954 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 157574 554294
rect 156954 518614 157574 554058
rect 156954 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 157574 518614
rect 156954 518294 157574 518378
rect 156954 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 157574 518294
rect 156954 482614 157574 518058
rect 156954 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 157574 482614
rect 156954 482294 157574 482378
rect 156954 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 157574 482294
rect 156954 446614 157574 482058
rect 156954 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 157574 446614
rect 156954 446294 157574 446378
rect 156954 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 157574 446294
rect 156954 410614 157574 446058
rect 156954 410378 156986 410614
rect 157222 410378 157306 410614
rect 157542 410378 157574 410614
rect 156954 410294 157574 410378
rect 156954 410058 156986 410294
rect 157222 410058 157306 410294
rect 157542 410058 157574 410294
rect 156954 374614 157574 410058
rect 156954 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 157574 374614
rect 156954 374294 157574 374378
rect 156954 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 157574 374294
rect 156954 338614 157574 374058
rect 156954 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 157574 338614
rect 156954 338294 157574 338378
rect 156954 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 157574 338294
rect 156954 302614 157574 338058
rect 156954 302378 156986 302614
rect 157222 302378 157306 302614
rect 157542 302378 157574 302614
rect 156954 302294 157574 302378
rect 156954 302058 156986 302294
rect 157222 302058 157306 302294
rect 157542 302058 157574 302294
rect 156954 266614 157574 302058
rect 156954 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 157574 266614
rect 156954 266294 157574 266378
rect 156954 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 157574 266294
rect 156954 230614 157574 266058
rect 156954 230378 156986 230614
rect 157222 230378 157306 230614
rect 157542 230378 157574 230614
rect 156954 230294 157574 230378
rect 156954 230058 156986 230294
rect 157222 230058 157306 230294
rect 157542 230058 157574 230294
rect 156954 194614 157574 230058
rect 156954 194378 156986 194614
rect 157222 194378 157306 194614
rect 157542 194378 157574 194614
rect 156954 194294 157574 194378
rect 156954 194058 156986 194294
rect 157222 194058 157306 194294
rect 157542 194058 157574 194294
rect 156954 158614 157574 194058
rect 163794 705798 164414 705830
rect 163794 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 164414 705798
rect 163794 705478 164414 705562
rect 163794 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 164414 705478
rect 163794 669454 164414 705242
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 163794 561454 164414 596898
rect 163794 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 164414 561454
rect 163794 561134 164414 561218
rect 163794 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 164414 561134
rect 163794 525454 164414 560898
rect 163794 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 164414 525454
rect 163794 525134 164414 525218
rect 163794 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 164414 525134
rect 163794 489454 164414 524898
rect 163794 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 164414 489454
rect 163794 489134 164414 489218
rect 163794 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 164414 489134
rect 163794 453454 164414 488898
rect 163794 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 164414 453454
rect 163794 453134 164414 453218
rect 163794 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 164414 453134
rect 163794 417454 164414 452898
rect 163794 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 164414 417454
rect 163794 417134 164414 417218
rect 163794 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 164414 417134
rect 163794 381454 164414 416898
rect 163794 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 164414 381454
rect 163794 381134 164414 381218
rect 163794 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 164414 381134
rect 163794 345454 164414 380898
rect 163794 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 164414 345454
rect 163794 345134 164414 345218
rect 163794 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 164414 345134
rect 163794 309454 164414 344898
rect 163794 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 164414 309454
rect 163794 309134 164414 309218
rect 163794 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 164414 309134
rect 163794 273454 164414 308898
rect 163794 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 164414 273454
rect 163794 273134 164414 273218
rect 163794 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 164414 273134
rect 163794 237454 164414 272898
rect 163794 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 164414 237454
rect 163794 237134 164414 237218
rect 163794 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 164414 237134
rect 163794 201454 164414 236898
rect 163794 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 164414 201454
rect 163794 201134 164414 201218
rect 163794 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 164414 201134
rect 163794 192000 164414 200898
rect 167514 673174 168134 707162
rect 167514 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 168134 673174
rect 167514 672854 168134 672938
rect 167514 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 168134 672854
rect 167514 637174 168134 672618
rect 167514 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 168134 637174
rect 167514 636854 168134 636938
rect 167514 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 168134 636854
rect 167514 601174 168134 636618
rect 167514 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 168134 601174
rect 167514 600854 168134 600938
rect 167514 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 168134 600854
rect 167514 565174 168134 600618
rect 167514 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 168134 565174
rect 167514 564854 168134 564938
rect 167514 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 168134 564854
rect 167514 529174 168134 564618
rect 167514 528938 167546 529174
rect 167782 528938 167866 529174
rect 168102 528938 168134 529174
rect 167514 528854 168134 528938
rect 167514 528618 167546 528854
rect 167782 528618 167866 528854
rect 168102 528618 168134 528854
rect 167514 493174 168134 528618
rect 167514 492938 167546 493174
rect 167782 492938 167866 493174
rect 168102 492938 168134 493174
rect 167514 492854 168134 492938
rect 167514 492618 167546 492854
rect 167782 492618 167866 492854
rect 168102 492618 168134 492854
rect 167514 457174 168134 492618
rect 167514 456938 167546 457174
rect 167782 456938 167866 457174
rect 168102 456938 168134 457174
rect 167514 456854 168134 456938
rect 167514 456618 167546 456854
rect 167782 456618 167866 456854
rect 168102 456618 168134 456854
rect 167514 421174 168134 456618
rect 167514 420938 167546 421174
rect 167782 420938 167866 421174
rect 168102 420938 168134 421174
rect 167514 420854 168134 420938
rect 167514 420618 167546 420854
rect 167782 420618 167866 420854
rect 168102 420618 168134 420854
rect 167514 385174 168134 420618
rect 167514 384938 167546 385174
rect 167782 384938 167866 385174
rect 168102 384938 168134 385174
rect 167514 384854 168134 384938
rect 167514 384618 167546 384854
rect 167782 384618 167866 384854
rect 168102 384618 168134 384854
rect 167514 349174 168134 384618
rect 167514 348938 167546 349174
rect 167782 348938 167866 349174
rect 168102 348938 168134 349174
rect 167514 348854 168134 348938
rect 167514 348618 167546 348854
rect 167782 348618 167866 348854
rect 168102 348618 168134 348854
rect 167514 313174 168134 348618
rect 167514 312938 167546 313174
rect 167782 312938 167866 313174
rect 168102 312938 168134 313174
rect 167514 312854 168134 312938
rect 167514 312618 167546 312854
rect 167782 312618 167866 312854
rect 168102 312618 168134 312854
rect 167514 277174 168134 312618
rect 167514 276938 167546 277174
rect 167782 276938 167866 277174
rect 168102 276938 168134 277174
rect 167514 276854 168134 276938
rect 167514 276618 167546 276854
rect 167782 276618 167866 276854
rect 168102 276618 168134 276854
rect 167514 241174 168134 276618
rect 167514 240938 167546 241174
rect 167782 240938 167866 241174
rect 168102 240938 168134 241174
rect 167514 240854 168134 240938
rect 167514 240618 167546 240854
rect 167782 240618 167866 240854
rect 168102 240618 168134 240854
rect 167514 205174 168134 240618
rect 167514 204938 167546 205174
rect 167782 204938 167866 205174
rect 168102 204938 168134 205174
rect 167514 204854 168134 204938
rect 167514 204618 167546 204854
rect 167782 204618 167866 204854
rect 168102 204618 168134 204854
rect 167514 192000 168134 204618
rect 171234 676894 171854 709082
rect 171234 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 171854 676894
rect 171234 676574 171854 676658
rect 171234 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 171854 676574
rect 171234 640894 171854 676338
rect 171234 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 171854 640894
rect 171234 640574 171854 640658
rect 171234 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 171854 640574
rect 171234 604894 171854 640338
rect 171234 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 171854 604894
rect 171234 604574 171854 604658
rect 171234 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 171854 604574
rect 171234 568894 171854 604338
rect 171234 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 171854 568894
rect 171234 568574 171854 568658
rect 171234 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 171854 568574
rect 171234 532894 171854 568338
rect 171234 532658 171266 532894
rect 171502 532658 171586 532894
rect 171822 532658 171854 532894
rect 171234 532574 171854 532658
rect 171234 532338 171266 532574
rect 171502 532338 171586 532574
rect 171822 532338 171854 532574
rect 171234 496894 171854 532338
rect 171234 496658 171266 496894
rect 171502 496658 171586 496894
rect 171822 496658 171854 496894
rect 171234 496574 171854 496658
rect 171234 496338 171266 496574
rect 171502 496338 171586 496574
rect 171822 496338 171854 496574
rect 171234 460894 171854 496338
rect 171234 460658 171266 460894
rect 171502 460658 171586 460894
rect 171822 460658 171854 460894
rect 171234 460574 171854 460658
rect 171234 460338 171266 460574
rect 171502 460338 171586 460574
rect 171822 460338 171854 460574
rect 171234 424894 171854 460338
rect 171234 424658 171266 424894
rect 171502 424658 171586 424894
rect 171822 424658 171854 424894
rect 171234 424574 171854 424658
rect 171234 424338 171266 424574
rect 171502 424338 171586 424574
rect 171822 424338 171854 424574
rect 171234 388894 171854 424338
rect 171234 388658 171266 388894
rect 171502 388658 171586 388894
rect 171822 388658 171854 388894
rect 171234 388574 171854 388658
rect 171234 388338 171266 388574
rect 171502 388338 171586 388574
rect 171822 388338 171854 388574
rect 171234 352894 171854 388338
rect 171234 352658 171266 352894
rect 171502 352658 171586 352894
rect 171822 352658 171854 352894
rect 171234 352574 171854 352658
rect 171234 352338 171266 352574
rect 171502 352338 171586 352574
rect 171822 352338 171854 352574
rect 171234 316894 171854 352338
rect 171234 316658 171266 316894
rect 171502 316658 171586 316894
rect 171822 316658 171854 316894
rect 171234 316574 171854 316658
rect 171234 316338 171266 316574
rect 171502 316338 171586 316574
rect 171822 316338 171854 316574
rect 171234 280894 171854 316338
rect 171234 280658 171266 280894
rect 171502 280658 171586 280894
rect 171822 280658 171854 280894
rect 171234 280574 171854 280658
rect 171234 280338 171266 280574
rect 171502 280338 171586 280574
rect 171822 280338 171854 280574
rect 171234 244894 171854 280338
rect 171234 244658 171266 244894
rect 171502 244658 171586 244894
rect 171822 244658 171854 244894
rect 171234 244574 171854 244658
rect 171234 244338 171266 244574
rect 171502 244338 171586 244574
rect 171822 244338 171854 244574
rect 171234 208894 171854 244338
rect 171234 208658 171266 208894
rect 171502 208658 171586 208894
rect 171822 208658 171854 208894
rect 171234 208574 171854 208658
rect 171234 208338 171266 208574
rect 171502 208338 171586 208574
rect 171822 208338 171854 208574
rect 171234 192000 171854 208338
rect 174954 680614 175574 711002
rect 192954 710598 193574 711590
rect 192954 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 193574 710598
rect 192954 710278 193574 710362
rect 192954 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 193574 710278
rect 189234 708678 189854 709670
rect 189234 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 189854 708678
rect 189234 708358 189854 708442
rect 189234 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 189854 708358
rect 185514 706758 186134 707750
rect 185514 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 186134 706758
rect 185514 706438 186134 706522
rect 185514 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 186134 706438
rect 174954 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 175574 680614
rect 174954 680294 175574 680378
rect 174954 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 175574 680294
rect 174954 644614 175574 680058
rect 174954 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 175574 644614
rect 174954 644294 175574 644378
rect 174954 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 175574 644294
rect 174954 608614 175574 644058
rect 174954 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 175574 608614
rect 174954 608294 175574 608378
rect 174954 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 175574 608294
rect 174954 572614 175574 608058
rect 174954 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 175574 572614
rect 174954 572294 175574 572378
rect 174954 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 175574 572294
rect 174954 536614 175574 572058
rect 174954 536378 174986 536614
rect 175222 536378 175306 536614
rect 175542 536378 175574 536614
rect 174954 536294 175574 536378
rect 174954 536058 174986 536294
rect 175222 536058 175306 536294
rect 175542 536058 175574 536294
rect 174954 500614 175574 536058
rect 174954 500378 174986 500614
rect 175222 500378 175306 500614
rect 175542 500378 175574 500614
rect 174954 500294 175574 500378
rect 174954 500058 174986 500294
rect 175222 500058 175306 500294
rect 175542 500058 175574 500294
rect 174954 464614 175574 500058
rect 174954 464378 174986 464614
rect 175222 464378 175306 464614
rect 175542 464378 175574 464614
rect 174954 464294 175574 464378
rect 174954 464058 174986 464294
rect 175222 464058 175306 464294
rect 175542 464058 175574 464294
rect 174954 428614 175574 464058
rect 174954 428378 174986 428614
rect 175222 428378 175306 428614
rect 175542 428378 175574 428614
rect 174954 428294 175574 428378
rect 174954 428058 174986 428294
rect 175222 428058 175306 428294
rect 175542 428058 175574 428294
rect 174954 392614 175574 428058
rect 174954 392378 174986 392614
rect 175222 392378 175306 392614
rect 175542 392378 175574 392614
rect 174954 392294 175574 392378
rect 174954 392058 174986 392294
rect 175222 392058 175306 392294
rect 175542 392058 175574 392294
rect 174954 356614 175574 392058
rect 174954 356378 174986 356614
rect 175222 356378 175306 356614
rect 175542 356378 175574 356614
rect 174954 356294 175574 356378
rect 174954 356058 174986 356294
rect 175222 356058 175306 356294
rect 175542 356058 175574 356294
rect 174954 320614 175574 356058
rect 174954 320378 174986 320614
rect 175222 320378 175306 320614
rect 175542 320378 175574 320614
rect 174954 320294 175574 320378
rect 174954 320058 174986 320294
rect 175222 320058 175306 320294
rect 175542 320058 175574 320294
rect 174954 284614 175574 320058
rect 174954 284378 174986 284614
rect 175222 284378 175306 284614
rect 175542 284378 175574 284614
rect 174954 284294 175574 284378
rect 174954 284058 174986 284294
rect 175222 284058 175306 284294
rect 175542 284058 175574 284294
rect 174954 248614 175574 284058
rect 174954 248378 174986 248614
rect 175222 248378 175306 248614
rect 175542 248378 175574 248614
rect 174954 248294 175574 248378
rect 174954 248058 174986 248294
rect 175222 248058 175306 248294
rect 175542 248058 175574 248294
rect 174954 212614 175574 248058
rect 174954 212378 174986 212614
rect 175222 212378 175306 212614
rect 175542 212378 175574 212614
rect 174954 212294 175574 212378
rect 174954 212058 174986 212294
rect 175222 212058 175306 212294
rect 175542 212058 175574 212294
rect 162243 183454 162563 183486
rect 162243 183218 162285 183454
rect 162521 183218 162563 183454
rect 162243 183134 162563 183218
rect 162243 182898 162285 183134
rect 162521 182898 162563 183134
rect 162243 182866 162563 182898
rect 164840 183454 165160 183486
rect 164840 183218 164882 183454
rect 165118 183218 165160 183454
rect 164840 183134 165160 183218
rect 164840 182898 164882 183134
rect 165118 182898 165160 183134
rect 164840 182866 165160 182898
rect 167437 183454 167757 183486
rect 167437 183218 167479 183454
rect 167715 183218 167757 183454
rect 167437 183134 167757 183218
rect 167437 182898 167479 183134
rect 167715 182898 167757 183134
rect 167437 182866 167757 182898
rect 174954 176614 175574 212058
rect 174954 176378 174986 176614
rect 175222 176378 175306 176614
rect 175542 176378 175574 176614
rect 174954 176294 175574 176378
rect 174954 176058 174986 176294
rect 175222 176058 175306 176294
rect 175542 176058 175574 176294
rect 163541 165454 163861 165486
rect 163541 165218 163583 165454
rect 163819 165218 163861 165454
rect 163541 165134 163861 165218
rect 163541 164898 163583 165134
rect 163819 164898 163861 165134
rect 163541 164866 163861 164898
rect 166138 165454 166458 165486
rect 166138 165218 166180 165454
rect 166416 165218 166458 165454
rect 166138 165134 166458 165218
rect 166138 164898 166180 165134
rect 166416 164898 166458 165134
rect 166138 164866 166458 164898
rect 156954 158378 156986 158614
rect 157222 158378 157306 158614
rect 157542 158378 157574 158614
rect 156954 158294 157574 158378
rect 156954 158058 156986 158294
rect 157222 158058 157306 158294
rect 157542 158058 157574 158294
rect 156954 122614 157574 158058
rect 163794 156000 164414 158000
rect 167514 156000 168134 158000
rect 171234 156000 171854 158000
rect 162243 147454 162563 147486
rect 162243 147218 162285 147454
rect 162521 147218 162563 147454
rect 162243 147134 162563 147218
rect 162243 146898 162285 147134
rect 162521 146898 162563 147134
rect 162243 146866 162563 146898
rect 164840 147454 165160 147486
rect 164840 147218 164882 147454
rect 165118 147218 165160 147454
rect 164840 147134 165160 147218
rect 164840 146898 164882 147134
rect 165118 146898 165160 147134
rect 164840 146866 165160 146898
rect 167437 147454 167757 147486
rect 167437 147218 167479 147454
rect 167715 147218 167757 147454
rect 167437 147134 167757 147218
rect 167437 146898 167479 147134
rect 167715 146898 167757 147134
rect 167437 146866 167757 146898
rect 174954 140614 175574 176058
rect 174954 140378 174986 140614
rect 175222 140378 175306 140614
rect 175542 140378 175574 140614
rect 174954 140294 175574 140378
rect 174954 140058 174986 140294
rect 175222 140058 175306 140294
rect 175542 140058 175574 140294
rect 163541 129454 163861 129486
rect 163541 129218 163583 129454
rect 163819 129218 163861 129454
rect 163541 129134 163861 129218
rect 163541 128898 163583 129134
rect 163819 128898 163861 129134
rect 163541 128866 163861 128898
rect 166138 129454 166458 129486
rect 166138 129218 166180 129454
rect 166416 129218 166458 129454
rect 166138 129134 166458 129218
rect 166138 128898 166180 129134
rect 166416 128898 166458 129134
rect 166138 128866 166458 128898
rect 156954 122378 156986 122614
rect 157222 122378 157306 122614
rect 157542 122378 157574 122614
rect 156954 122294 157574 122378
rect 156954 122058 156986 122294
rect 157222 122058 157306 122294
rect 157542 122058 157574 122294
rect 156954 86614 157574 122058
rect 156954 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 157574 86614
rect 156954 86294 157574 86378
rect 156954 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 157574 86294
rect 156954 50614 157574 86058
rect 156954 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 157574 50614
rect 156954 50294 157574 50378
rect 156954 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 157574 50294
rect 156954 14614 157574 50058
rect 156954 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 157574 14614
rect 156954 14294 157574 14378
rect 156954 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 157574 14294
rect 138954 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 139574 -7066
rect 138954 -7386 139574 -7302
rect 138954 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 139574 -7386
rect 138954 -7654 139574 -7622
rect 156954 -6106 157574 14058
rect 163794 93454 164414 122000
rect 163794 93218 163826 93454
rect 164062 93218 164146 93454
rect 164382 93218 164414 93454
rect 163794 93134 164414 93218
rect 163794 92898 163826 93134
rect 164062 92898 164146 93134
rect 164382 92898 164414 93134
rect 163794 57454 164414 92898
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -1306 164414 20898
rect 163794 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 164414 -1306
rect 163794 -1626 164414 -1542
rect 163794 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 164414 -1626
rect 163794 -1894 164414 -1862
rect 167514 97174 168134 122000
rect 167514 96938 167546 97174
rect 167782 96938 167866 97174
rect 168102 96938 168134 97174
rect 167514 96854 168134 96938
rect 167514 96618 167546 96854
rect 167782 96618 167866 96854
rect 168102 96618 168134 96854
rect 167514 61174 168134 96618
rect 167514 60938 167546 61174
rect 167782 60938 167866 61174
rect 168102 60938 168134 61174
rect 167514 60854 168134 60938
rect 167514 60618 167546 60854
rect 167782 60618 167866 60854
rect 168102 60618 168134 60854
rect 167514 25174 168134 60618
rect 167514 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 168134 25174
rect 167514 24854 168134 24938
rect 167514 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 168134 24854
rect 167514 -3226 168134 24618
rect 167514 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 168134 -3226
rect 167514 -3546 168134 -3462
rect 167514 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 168134 -3546
rect 167514 -3814 168134 -3782
rect 171234 100894 171854 122000
rect 171234 100658 171266 100894
rect 171502 100658 171586 100894
rect 171822 100658 171854 100894
rect 171234 100574 171854 100658
rect 171234 100338 171266 100574
rect 171502 100338 171586 100574
rect 171822 100338 171854 100574
rect 171234 64894 171854 100338
rect 171234 64658 171266 64894
rect 171502 64658 171586 64894
rect 171822 64658 171854 64894
rect 171234 64574 171854 64658
rect 171234 64338 171266 64574
rect 171502 64338 171586 64574
rect 171822 64338 171854 64574
rect 171234 28894 171854 64338
rect 171234 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 171854 28894
rect 171234 28574 171854 28658
rect 171234 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 171854 28574
rect 171234 -5146 171854 28338
rect 171234 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 171854 -5146
rect 171234 -5466 171854 -5382
rect 171234 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 171854 -5466
rect 171234 -5734 171854 -5702
rect 174954 104614 175574 140058
rect 174954 104378 174986 104614
rect 175222 104378 175306 104614
rect 175542 104378 175574 104614
rect 174954 104294 175574 104378
rect 174954 104058 174986 104294
rect 175222 104058 175306 104294
rect 175542 104058 175574 104294
rect 174954 68614 175574 104058
rect 174954 68378 174986 68614
rect 175222 68378 175306 68614
rect 175542 68378 175574 68614
rect 174954 68294 175574 68378
rect 174954 68058 174986 68294
rect 175222 68058 175306 68294
rect 175542 68058 175574 68294
rect 174954 32614 175574 68058
rect 174954 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 175574 32614
rect 174954 32294 175574 32378
rect 174954 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 175574 32294
rect 156954 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 157574 -6106
rect 156954 -6426 157574 -6342
rect 156954 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 157574 -6426
rect 156954 -7654 157574 -6662
rect 174954 -7066 175574 32058
rect 181794 704838 182414 705830
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 543454 182414 578898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 507454 182414 542898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 181794 471454 182414 506898
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 181794 435454 182414 470898
rect 181794 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 182414 435454
rect 181794 435134 182414 435218
rect 181794 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 182414 435134
rect 181794 399454 182414 434898
rect 181794 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 182414 399454
rect 181794 399134 182414 399218
rect 181794 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 182414 399134
rect 181794 363454 182414 398898
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 181794 327454 182414 362898
rect 181794 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 182414 327454
rect 181794 327134 182414 327218
rect 181794 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 182414 327134
rect 181794 291454 182414 326898
rect 181794 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 182414 291454
rect 181794 291134 182414 291218
rect 181794 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 182414 291134
rect 181794 255454 182414 290898
rect 181794 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 182414 255454
rect 181794 255134 182414 255218
rect 181794 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 182414 255134
rect 181794 219454 182414 254898
rect 181794 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 182414 219454
rect 181794 219134 182414 219218
rect 181794 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 182414 219134
rect 181794 183454 182414 218898
rect 181794 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 182414 183454
rect 181794 183134 182414 183218
rect 181794 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 182414 183134
rect 181794 147454 182414 182898
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 111454 182414 146898
rect 181794 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 182414 111454
rect 181794 111134 182414 111218
rect 181794 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 182414 111134
rect 181794 75454 182414 110898
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 181794 39454 182414 74898
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -1894 182414 -902
rect 185514 691174 186134 706202
rect 185514 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 186134 691174
rect 185514 690854 186134 690938
rect 185514 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 186134 690854
rect 185514 655174 186134 690618
rect 185514 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 186134 655174
rect 185514 654854 186134 654938
rect 185514 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 186134 654854
rect 185514 619174 186134 654618
rect 185514 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 186134 619174
rect 185514 618854 186134 618938
rect 185514 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 186134 618854
rect 185514 583174 186134 618618
rect 185514 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 186134 583174
rect 185514 582854 186134 582938
rect 185514 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 186134 582854
rect 185514 547174 186134 582618
rect 185514 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 186134 547174
rect 185514 546854 186134 546938
rect 185514 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 186134 546854
rect 185514 511174 186134 546618
rect 185514 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 186134 511174
rect 185514 510854 186134 510938
rect 185514 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 186134 510854
rect 185514 475174 186134 510618
rect 185514 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 186134 475174
rect 185514 474854 186134 474938
rect 185514 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 186134 474854
rect 185514 439174 186134 474618
rect 185514 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 186134 439174
rect 185514 438854 186134 438938
rect 185514 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 186134 438854
rect 185514 403174 186134 438618
rect 185514 402938 185546 403174
rect 185782 402938 185866 403174
rect 186102 402938 186134 403174
rect 185514 402854 186134 402938
rect 185514 402618 185546 402854
rect 185782 402618 185866 402854
rect 186102 402618 186134 402854
rect 185514 367174 186134 402618
rect 185514 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 186134 367174
rect 185514 366854 186134 366938
rect 185514 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 186134 366854
rect 185514 331174 186134 366618
rect 185514 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 186134 331174
rect 185514 330854 186134 330938
rect 185514 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 186134 330854
rect 185514 295174 186134 330618
rect 185514 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 186134 295174
rect 185514 294854 186134 294938
rect 185514 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 186134 294854
rect 185514 259174 186134 294618
rect 185514 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 186134 259174
rect 185514 258854 186134 258938
rect 185514 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 186134 258854
rect 185514 223174 186134 258618
rect 185514 222938 185546 223174
rect 185782 222938 185866 223174
rect 186102 222938 186134 223174
rect 185514 222854 186134 222938
rect 185514 222618 185546 222854
rect 185782 222618 185866 222854
rect 186102 222618 186134 222854
rect 185514 187174 186134 222618
rect 185514 186938 185546 187174
rect 185782 186938 185866 187174
rect 186102 186938 186134 187174
rect 185514 186854 186134 186938
rect 185514 186618 185546 186854
rect 185782 186618 185866 186854
rect 186102 186618 186134 186854
rect 185514 151174 186134 186618
rect 185514 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 186134 151174
rect 185514 150854 186134 150938
rect 185514 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 186134 150854
rect 185514 115174 186134 150618
rect 185514 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 186134 115174
rect 185514 114854 186134 114938
rect 185514 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 186134 114854
rect 185514 79174 186134 114618
rect 185514 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 186134 79174
rect 185514 78854 186134 78938
rect 185514 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 186134 78854
rect 185514 43174 186134 78618
rect 185514 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 186134 43174
rect 185514 42854 186134 42938
rect 185514 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 186134 42854
rect 185514 7174 186134 42618
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 185514 -2266 186134 6618
rect 185514 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 186134 -2266
rect 185514 -2586 186134 -2502
rect 185514 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 186134 -2586
rect 185514 -3814 186134 -2822
rect 189234 694894 189854 708122
rect 189234 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 189854 694894
rect 189234 694574 189854 694658
rect 189234 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 189854 694574
rect 189234 658894 189854 694338
rect 189234 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 189854 658894
rect 189234 658574 189854 658658
rect 189234 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 189854 658574
rect 189234 622894 189854 658338
rect 189234 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 189854 622894
rect 189234 622574 189854 622658
rect 189234 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 189854 622574
rect 189234 586894 189854 622338
rect 189234 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 189854 586894
rect 189234 586574 189854 586658
rect 189234 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 189854 586574
rect 189234 550894 189854 586338
rect 189234 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 189854 550894
rect 189234 550574 189854 550658
rect 189234 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 189854 550574
rect 189234 514894 189854 550338
rect 189234 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 189854 514894
rect 189234 514574 189854 514658
rect 189234 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 189854 514574
rect 189234 478894 189854 514338
rect 189234 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 189854 478894
rect 189234 478574 189854 478658
rect 189234 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 189854 478574
rect 189234 442894 189854 478338
rect 189234 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 189854 442894
rect 189234 442574 189854 442658
rect 189234 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 189854 442574
rect 189234 406894 189854 442338
rect 189234 406658 189266 406894
rect 189502 406658 189586 406894
rect 189822 406658 189854 406894
rect 189234 406574 189854 406658
rect 189234 406338 189266 406574
rect 189502 406338 189586 406574
rect 189822 406338 189854 406574
rect 189234 370894 189854 406338
rect 189234 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 189854 370894
rect 189234 370574 189854 370658
rect 189234 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 189854 370574
rect 189234 334894 189854 370338
rect 189234 334658 189266 334894
rect 189502 334658 189586 334894
rect 189822 334658 189854 334894
rect 189234 334574 189854 334658
rect 189234 334338 189266 334574
rect 189502 334338 189586 334574
rect 189822 334338 189854 334574
rect 189234 298894 189854 334338
rect 189234 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 189854 298894
rect 189234 298574 189854 298658
rect 189234 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 189854 298574
rect 189234 262894 189854 298338
rect 189234 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 189854 262894
rect 189234 262574 189854 262658
rect 189234 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 189854 262574
rect 189234 226894 189854 262338
rect 189234 226658 189266 226894
rect 189502 226658 189586 226894
rect 189822 226658 189854 226894
rect 189234 226574 189854 226658
rect 189234 226338 189266 226574
rect 189502 226338 189586 226574
rect 189822 226338 189854 226574
rect 189234 190894 189854 226338
rect 189234 190658 189266 190894
rect 189502 190658 189586 190894
rect 189822 190658 189854 190894
rect 189234 190574 189854 190658
rect 189234 190338 189266 190574
rect 189502 190338 189586 190574
rect 189822 190338 189854 190574
rect 189234 154894 189854 190338
rect 189234 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 189854 154894
rect 189234 154574 189854 154658
rect 189234 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 189854 154574
rect 189234 118894 189854 154338
rect 189234 118658 189266 118894
rect 189502 118658 189586 118894
rect 189822 118658 189854 118894
rect 189234 118574 189854 118658
rect 189234 118338 189266 118574
rect 189502 118338 189586 118574
rect 189822 118338 189854 118574
rect 189234 82894 189854 118338
rect 189234 82658 189266 82894
rect 189502 82658 189586 82894
rect 189822 82658 189854 82894
rect 189234 82574 189854 82658
rect 189234 82338 189266 82574
rect 189502 82338 189586 82574
rect 189822 82338 189854 82574
rect 189234 46894 189854 82338
rect 189234 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 189854 46894
rect 189234 46574 189854 46658
rect 189234 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 189854 46574
rect 189234 10894 189854 46338
rect 189234 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 189854 10894
rect 189234 10574 189854 10658
rect 189234 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 189854 10574
rect 189234 -4186 189854 10338
rect 189234 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 189854 -4186
rect 189234 -4506 189854 -4422
rect 189234 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 189854 -4506
rect 189234 -5734 189854 -4742
rect 192954 698614 193574 710042
rect 210954 711558 211574 711590
rect 210954 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 211574 711558
rect 210954 711238 211574 711322
rect 210954 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 211574 711238
rect 207234 709638 207854 709670
rect 207234 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 207854 709638
rect 207234 709318 207854 709402
rect 207234 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 207854 709318
rect 203514 707718 204134 707750
rect 203514 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 204134 707718
rect 203514 707398 204134 707482
rect 203514 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 204134 707398
rect 192954 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 193574 698614
rect 192954 698294 193574 698378
rect 192954 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 193574 698294
rect 192954 662614 193574 698058
rect 192954 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 193574 662614
rect 192954 662294 193574 662378
rect 192954 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 193574 662294
rect 192954 626614 193574 662058
rect 192954 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 193574 626614
rect 192954 626294 193574 626378
rect 192954 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 193574 626294
rect 192954 590614 193574 626058
rect 192954 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 193574 590614
rect 192954 590294 193574 590378
rect 192954 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 193574 590294
rect 192954 554614 193574 590058
rect 192954 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 193574 554614
rect 192954 554294 193574 554378
rect 192954 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 193574 554294
rect 192954 518614 193574 554058
rect 192954 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 193574 518614
rect 192954 518294 193574 518378
rect 192954 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 193574 518294
rect 192954 482614 193574 518058
rect 192954 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 193574 482614
rect 192954 482294 193574 482378
rect 192954 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 193574 482294
rect 192954 446614 193574 482058
rect 192954 446378 192986 446614
rect 193222 446378 193306 446614
rect 193542 446378 193574 446614
rect 192954 446294 193574 446378
rect 192954 446058 192986 446294
rect 193222 446058 193306 446294
rect 193542 446058 193574 446294
rect 192954 410614 193574 446058
rect 192954 410378 192986 410614
rect 193222 410378 193306 410614
rect 193542 410378 193574 410614
rect 192954 410294 193574 410378
rect 192954 410058 192986 410294
rect 193222 410058 193306 410294
rect 193542 410058 193574 410294
rect 192954 374614 193574 410058
rect 192954 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 193574 374614
rect 192954 374294 193574 374378
rect 192954 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 193574 374294
rect 192954 338614 193574 374058
rect 192954 338378 192986 338614
rect 193222 338378 193306 338614
rect 193542 338378 193574 338614
rect 192954 338294 193574 338378
rect 192954 338058 192986 338294
rect 193222 338058 193306 338294
rect 193542 338058 193574 338294
rect 192954 302614 193574 338058
rect 192954 302378 192986 302614
rect 193222 302378 193306 302614
rect 193542 302378 193574 302614
rect 192954 302294 193574 302378
rect 192954 302058 192986 302294
rect 193222 302058 193306 302294
rect 193542 302058 193574 302294
rect 192954 266614 193574 302058
rect 192954 266378 192986 266614
rect 193222 266378 193306 266614
rect 193542 266378 193574 266614
rect 192954 266294 193574 266378
rect 192954 266058 192986 266294
rect 193222 266058 193306 266294
rect 193542 266058 193574 266294
rect 192954 230614 193574 266058
rect 192954 230378 192986 230614
rect 193222 230378 193306 230614
rect 193542 230378 193574 230614
rect 192954 230294 193574 230378
rect 192954 230058 192986 230294
rect 193222 230058 193306 230294
rect 193542 230058 193574 230294
rect 192954 194614 193574 230058
rect 199794 705798 200414 705830
rect 199794 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 200414 705798
rect 199794 705478 200414 705562
rect 199794 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 200414 705478
rect 199794 669454 200414 705242
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 561454 200414 596898
rect 199794 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 200414 561454
rect 199794 561134 200414 561218
rect 199794 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 200414 561134
rect 199794 525454 200414 560898
rect 199794 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 200414 525454
rect 199794 525134 200414 525218
rect 199794 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 200414 525134
rect 199794 489454 200414 524898
rect 199794 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 200414 489454
rect 199794 489134 200414 489218
rect 199794 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 200414 489134
rect 199794 453454 200414 488898
rect 199794 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 200414 453454
rect 199794 453134 200414 453218
rect 199794 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 200414 453134
rect 199794 417454 200414 452898
rect 199794 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 200414 417454
rect 199794 417134 200414 417218
rect 199794 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 200414 417134
rect 199794 381454 200414 416898
rect 199794 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 200414 381454
rect 199794 381134 200414 381218
rect 199794 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 200414 381134
rect 199794 345454 200414 380898
rect 199794 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 200414 345454
rect 199794 345134 200414 345218
rect 199794 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 200414 345134
rect 199794 309454 200414 344898
rect 199794 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 200414 309454
rect 199794 309134 200414 309218
rect 199794 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 200414 309134
rect 199794 273454 200414 308898
rect 199794 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 200414 273454
rect 199794 273134 200414 273218
rect 199794 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 200414 273134
rect 199794 237454 200414 272898
rect 199794 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 200414 237454
rect 199794 237134 200414 237218
rect 199794 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 200414 237134
rect 199794 202000 200414 236898
rect 203514 673174 204134 707162
rect 203514 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 204134 673174
rect 203514 672854 204134 672938
rect 203514 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 204134 672854
rect 203514 637174 204134 672618
rect 203514 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 204134 637174
rect 203514 636854 204134 636938
rect 203514 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 204134 636854
rect 203514 601174 204134 636618
rect 203514 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 204134 601174
rect 203514 600854 204134 600938
rect 203514 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 204134 600854
rect 203514 565174 204134 600618
rect 203514 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 204134 565174
rect 203514 564854 204134 564938
rect 203514 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 204134 564854
rect 203514 529174 204134 564618
rect 203514 528938 203546 529174
rect 203782 528938 203866 529174
rect 204102 528938 204134 529174
rect 203514 528854 204134 528938
rect 203514 528618 203546 528854
rect 203782 528618 203866 528854
rect 204102 528618 204134 528854
rect 203514 493174 204134 528618
rect 203514 492938 203546 493174
rect 203782 492938 203866 493174
rect 204102 492938 204134 493174
rect 203514 492854 204134 492938
rect 203514 492618 203546 492854
rect 203782 492618 203866 492854
rect 204102 492618 204134 492854
rect 203514 457174 204134 492618
rect 203514 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 204134 457174
rect 203514 456854 204134 456938
rect 203514 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 204134 456854
rect 203514 421174 204134 456618
rect 203514 420938 203546 421174
rect 203782 420938 203866 421174
rect 204102 420938 204134 421174
rect 203514 420854 204134 420938
rect 203514 420618 203546 420854
rect 203782 420618 203866 420854
rect 204102 420618 204134 420854
rect 203514 385174 204134 420618
rect 203514 384938 203546 385174
rect 203782 384938 203866 385174
rect 204102 384938 204134 385174
rect 203514 384854 204134 384938
rect 203514 384618 203546 384854
rect 203782 384618 203866 384854
rect 204102 384618 204134 384854
rect 203514 349174 204134 384618
rect 203514 348938 203546 349174
rect 203782 348938 203866 349174
rect 204102 348938 204134 349174
rect 203514 348854 204134 348938
rect 203514 348618 203546 348854
rect 203782 348618 203866 348854
rect 204102 348618 204134 348854
rect 203514 313174 204134 348618
rect 203514 312938 203546 313174
rect 203782 312938 203866 313174
rect 204102 312938 204134 313174
rect 203514 312854 204134 312938
rect 203514 312618 203546 312854
rect 203782 312618 203866 312854
rect 204102 312618 204134 312854
rect 203514 277174 204134 312618
rect 203514 276938 203546 277174
rect 203782 276938 203866 277174
rect 204102 276938 204134 277174
rect 203514 276854 204134 276938
rect 203514 276618 203546 276854
rect 203782 276618 203866 276854
rect 204102 276618 204134 276854
rect 203514 241174 204134 276618
rect 203514 240938 203546 241174
rect 203782 240938 203866 241174
rect 204102 240938 204134 241174
rect 203514 240854 204134 240938
rect 203514 240618 203546 240854
rect 203782 240618 203866 240854
rect 204102 240618 204134 240854
rect 203514 205174 204134 240618
rect 203514 204938 203546 205174
rect 203782 204938 203866 205174
rect 204102 204938 204134 205174
rect 203514 204854 204134 204938
rect 203514 204618 203546 204854
rect 203782 204618 203866 204854
rect 204102 204618 204134 204854
rect 203514 202000 204134 204618
rect 207234 676894 207854 709082
rect 207234 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 207854 676894
rect 207234 676574 207854 676658
rect 207234 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 207854 676574
rect 207234 640894 207854 676338
rect 207234 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 207854 640894
rect 207234 640574 207854 640658
rect 207234 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 207854 640574
rect 207234 604894 207854 640338
rect 207234 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 207854 604894
rect 207234 604574 207854 604658
rect 207234 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 207854 604574
rect 207234 568894 207854 604338
rect 207234 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 207854 568894
rect 207234 568574 207854 568658
rect 207234 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 207854 568574
rect 207234 532894 207854 568338
rect 207234 532658 207266 532894
rect 207502 532658 207586 532894
rect 207822 532658 207854 532894
rect 207234 532574 207854 532658
rect 207234 532338 207266 532574
rect 207502 532338 207586 532574
rect 207822 532338 207854 532574
rect 207234 496894 207854 532338
rect 207234 496658 207266 496894
rect 207502 496658 207586 496894
rect 207822 496658 207854 496894
rect 207234 496574 207854 496658
rect 207234 496338 207266 496574
rect 207502 496338 207586 496574
rect 207822 496338 207854 496574
rect 207234 460894 207854 496338
rect 207234 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 207854 460894
rect 207234 460574 207854 460658
rect 207234 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 207854 460574
rect 207234 424894 207854 460338
rect 207234 424658 207266 424894
rect 207502 424658 207586 424894
rect 207822 424658 207854 424894
rect 207234 424574 207854 424658
rect 207234 424338 207266 424574
rect 207502 424338 207586 424574
rect 207822 424338 207854 424574
rect 207234 388894 207854 424338
rect 207234 388658 207266 388894
rect 207502 388658 207586 388894
rect 207822 388658 207854 388894
rect 207234 388574 207854 388658
rect 207234 388338 207266 388574
rect 207502 388338 207586 388574
rect 207822 388338 207854 388574
rect 207234 352894 207854 388338
rect 207234 352658 207266 352894
rect 207502 352658 207586 352894
rect 207822 352658 207854 352894
rect 207234 352574 207854 352658
rect 207234 352338 207266 352574
rect 207502 352338 207586 352574
rect 207822 352338 207854 352574
rect 207234 316894 207854 352338
rect 207234 316658 207266 316894
rect 207502 316658 207586 316894
rect 207822 316658 207854 316894
rect 207234 316574 207854 316658
rect 207234 316338 207266 316574
rect 207502 316338 207586 316574
rect 207822 316338 207854 316574
rect 207234 280894 207854 316338
rect 207234 280658 207266 280894
rect 207502 280658 207586 280894
rect 207822 280658 207854 280894
rect 207234 280574 207854 280658
rect 207234 280338 207266 280574
rect 207502 280338 207586 280574
rect 207822 280338 207854 280574
rect 207234 244894 207854 280338
rect 207234 244658 207266 244894
rect 207502 244658 207586 244894
rect 207822 244658 207854 244894
rect 207234 244574 207854 244658
rect 207234 244338 207266 244574
rect 207502 244338 207586 244574
rect 207822 244338 207854 244574
rect 207234 208894 207854 244338
rect 207234 208658 207266 208894
rect 207502 208658 207586 208894
rect 207822 208658 207854 208894
rect 207234 208574 207854 208658
rect 207234 208338 207266 208574
rect 207502 208338 207586 208574
rect 207822 208338 207854 208574
rect 207234 202000 207854 208338
rect 210954 680614 211574 711002
rect 228954 710598 229574 711590
rect 228954 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 229574 710598
rect 228954 710278 229574 710362
rect 228954 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 229574 710278
rect 225234 708678 225854 709670
rect 225234 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 225854 708678
rect 225234 708358 225854 708442
rect 225234 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 225854 708358
rect 221514 706758 222134 707750
rect 221514 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 222134 706758
rect 221514 706438 222134 706522
rect 221514 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 222134 706438
rect 210954 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 211574 680614
rect 210954 680294 211574 680378
rect 210954 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 211574 680294
rect 210954 644614 211574 680058
rect 210954 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 211574 644614
rect 210954 644294 211574 644378
rect 210954 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 211574 644294
rect 210954 608614 211574 644058
rect 210954 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 211574 608614
rect 210954 608294 211574 608378
rect 210954 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 211574 608294
rect 210954 572614 211574 608058
rect 210954 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 211574 572614
rect 210954 572294 211574 572378
rect 210954 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 211574 572294
rect 210954 536614 211574 572058
rect 210954 536378 210986 536614
rect 211222 536378 211306 536614
rect 211542 536378 211574 536614
rect 210954 536294 211574 536378
rect 210954 536058 210986 536294
rect 211222 536058 211306 536294
rect 211542 536058 211574 536294
rect 210954 500614 211574 536058
rect 210954 500378 210986 500614
rect 211222 500378 211306 500614
rect 211542 500378 211574 500614
rect 210954 500294 211574 500378
rect 210954 500058 210986 500294
rect 211222 500058 211306 500294
rect 211542 500058 211574 500294
rect 210954 464614 211574 500058
rect 210954 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 211574 464614
rect 210954 464294 211574 464378
rect 210954 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 211574 464294
rect 210954 428614 211574 464058
rect 210954 428378 210986 428614
rect 211222 428378 211306 428614
rect 211542 428378 211574 428614
rect 210954 428294 211574 428378
rect 210954 428058 210986 428294
rect 211222 428058 211306 428294
rect 211542 428058 211574 428294
rect 210954 392614 211574 428058
rect 210954 392378 210986 392614
rect 211222 392378 211306 392614
rect 211542 392378 211574 392614
rect 210954 392294 211574 392378
rect 210954 392058 210986 392294
rect 211222 392058 211306 392294
rect 211542 392058 211574 392294
rect 210954 356614 211574 392058
rect 210954 356378 210986 356614
rect 211222 356378 211306 356614
rect 211542 356378 211574 356614
rect 210954 356294 211574 356378
rect 210954 356058 210986 356294
rect 211222 356058 211306 356294
rect 211542 356058 211574 356294
rect 210954 320614 211574 356058
rect 210954 320378 210986 320614
rect 211222 320378 211306 320614
rect 211542 320378 211574 320614
rect 210954 320294 211574 320378
rect 210954 320058 210986 320294
rect 211222 320058 211306 320294
rect 211542 320058 211574 320294
rect 210954 284614 211574 320058
rect 210954 284378 210986 284614
rect 211222 284378 211306 284614
rect 211542 284378 211574 284614
rect 210954 284294 211574 284378
rect 210954 284058 210986 284294
rect 211222 284058 211306 284294
rect 211542 284058 211574 284294
rect 210954 248614 211574 284058
rect 210954 248378 210986 248614
rect 211222 248378 211306 248614
rect 211542 248378 211574 248614
rect 210954 248294 211574 248378
rect 210954 248058 210986 248294
rect 211222 248058 211306 248294
rect 211542 248058 211574 248294
rect 210954 212614 211574 248058
rect 210954 212378 210986 212614
rect 211222 212378 211306 212614
rect 211542 212378 211574 212614
rect 210954 212294 211574 212378
rect 210954 212058 210986 212294
rect 211222 212058 211306 212294
rect 211542 212058 211574 212294
rect 210954 202000 211574 212058
rect 217794 704838 218414 705830
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 543454 218414 578898
rect 217794 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 218414 543454
rect 217794 543134 218414 543218
rect 217794 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 218414 543134
rect 217794 507454 218414 542898
rect 217794 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 218414 507454
rect 217794 507134 218414 507218
rect 217794 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 218414 507134
rect 217794 471454 218414 506898
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 217794 435454 218414 470898
rect 217794 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 218414 435454
rect 217794 435134 218414 435218
rect 217794 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 218414 435134
rect 217794 399454 218414 434898
rect 217794 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 218414 399454
rect 217794 399134 218414 399218
rect 217794 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 218414 399134
rect 217794 363454 218414 398898
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 217794 327454 218414 362898
rect 217794 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 218414 327454
rect 217794 327134 218414 327218
rect 217794 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 218414 327134
rect 217794 291454 218414 326898
rect 217794 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 218414 291454
rect 217794 291134 218414 291218
rect 217794 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 218414 291134
rect 217794 255454 218414 290898
rect 217794 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 218414 255454
rect 217794 255134 218414 255218
rect 217794 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 218414 255134
rect 217794 219454 218414 254898
rect 217794 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 218414 219454
rect 217794 219134 218414 219218
rect 217794 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 218414 219134
rect 217794 202000 218414 218898
rect 221514 691174 222134 706202
rect 221514 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 222134 691174
rect 221514 690854 222134 690938
rect 221514 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 222134 690854
rect 221514 655174 222134 690618
rect 221514 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 222134 655174
rect 221514 654854 222134 654938
rect 221514 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 222134 654854
rect 221514 619174 222134 654618
rect 221514 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 222134 619174
rect 221514 618854 222134 618938
rect 221514 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 222134 618854
rect 221514 583174 222134 618618
rect 221514 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 222134 583174
rect 221514 582854 222134 582938
rect 221514 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 222134 582854
rect 221514 547174 222134 582618
rect 221514 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 222134 547174
rect 221514 546854 222134 546938
rect 221514 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 222134 546854
rect 221514 511174 222134 546618
rect 221514 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 222134 511174
rect 221514 510854 222134 510938
rect 221514 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 222134 510854
rect 221514 475174 222134 510618
rect 221514 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 222134 475174
rect 221514 474854 222134 474938
rect 221514 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 222134 474854
rect 221514 439174 222134 474618
rect 221514 438938 221546 439174
rect 221782 438938 221866 439174
rect 222102 438938 222134 439174
rect 221514 438854 222134 438938
rect 221514 438618 221546 438854
rect 221782 438618 221866 438854
rect 222102 438618 222134 438854
rect 221514 403174 222134 438618
rect 221514 402938 221546 403174
rect 221782 402938 221866 403174
rect 222102 402938 222134 403174
rect 221514 402854 222134 402938
rect 221514 402618 221546 402854
rect 221782 402618 221866 402854
rect 222102 402618 222134 402854
rect 221514 367174 222134 402618
rect 221514 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 222134 367174
rect 221514 366854 222134 366938
rect 221514 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 222134 366854
rect 221514 331174 222134 366618
rect 221514 330938 221546 331174
rect 221782 330938 221866 331174
rect 222102 330938 222134 331174
rect 221514 330854 222134 330938
rect 221514 330618 221546 330854
rect 221782 330618 221866 330854
rect 222102 330618 222134 330854
rect 221514 295174 222134 330618
rect 221514 294938 221546 295174
rect 221782 294938 221866 295174
rect 222102 294938 222134 295174
rect 221514 294854 222134 294938
rect 221514 294618 221546 294854
rect 221782 294618 221866 294854
rect 222102 294618 222134 294854
rect 221514 259174 222134 294618
rect 221514 258938 221546 259174
rect 221782 258938 221866 259174
rect 222102 258938 222134 259174
rect 221514 258854 222134 258938
rect 221514 258618 221546 258854
rect 221782 258618 221866 258854
rect 222102 258618 222134 258854
rect 221514 223174 222134 258618
rect 221514 222938 221546 223174
rect 221782 222938 221866 223174
rect 222102 222938 222134 223174
rect 221514 222854 222134 222938
rect 221514 222618 221546 222854
rect 221782 222618 221866 222854
rect 222102 222618 222134 222854
rect 221514 202000 222134 222618
rect 225234 694894 225854 708122
rect 225234 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 225854 694894
rect 225234 694574 225854 694658
rect 225234 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 225854 694574
rect 225234 658894 225854 694338
rect 225234 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 225854 658894
rect 225234 658574 225854 658658
rect 225234 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 225854 658574
rect 225234 622894 225854 658338
rect 225234 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 225854 622894
rect 225234 622574 225854 622658
rect 225234 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 225854 622574
rect 225234 586894 225854 622338
rect 225234 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 225854 586894
rect 225234 586574 225854 586658
rect 225234 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 225854 586574
rect 225234 550894 225854 586338
rect 225234 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 225854 550894
rect 225234 550574 225854 550658
rect 225234 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 225854 550574
rect 225234 514894 225854 550338
rect 225234 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 225854 514894
rect 225234 514574 225854 514658
rect 225234 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 225854 514574
rect 225234 478894 225854 514338
rect 225234 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 225854 478894
rect 225234 478574 225854 478658
rect 225234 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 225854 478574
rect 225234 442894 225854 478338
rect 225234 442658 225266 442894
rect 225502 442658 225586 442894
rect 225822 442658 225854 442894
rect 225234 442574 225854 442658
rect 225234 442338 225266 442574
rect 225502 442338 225586 442574
rect 225822 442338 225854 442574
rect 225234 406894 225854 442338
rect 225234 406658 225266 406894
rect 225502 406658 225586 406894
rect 225822 406658 225854 406894
rect 225234 406574 225854 406658
rect 225234 406338 225266 406574
rect 225502 406338 225586 406574
rect 225822 406338 225854 406574
rect 225234 370894 225854 406338
rect 225234 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 225854 370894
rect 225234 370574 225854 370658
rect 225234 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 225854 370574
rect 225234 334894 225854 370338
rect 225234 334658 225266 334894
rect 225502 334658 225586 334894
rect 225822 334658 225854 334894
rect 225234 334574 225854 334658
rect 225234 334338 225266 334574
rect 225502 334338 225586 334574
rect 225822 334338 225854 334574
rect 225234 298894 225854 334338
rect 225234 298658 225266 298894
rect 225502 298658 225586 298894
rect 225822 298658 225854 298894
rect 225234 298574 225854 298658
rect 225234 298338 225266 298574
rect 225502 298338 225586 298574
rect 225822 298338 225854 298574
rect 225234 262894 225854 298338
rect 225234 262658 225266 262894
rect 225502 262658 225586 262894
rect 225822 262658 225854 262894
rect 225234 262574 225854 262658
rect 225234 262338 225266 262574
rect 225502 262338 225586 262574
rect 225822 262338 225854 262574
rect 225234 226894 225854 262338
rect 225234 226658 225266 226894
rect 225502 226658 225586 226894
rect 225822 226658 225854 226894
rect 225234 226574 225854 226658
rect 225234 226338 225266 226574
rect 225502 226338 225586 226574
rect 225822 226338 225854 226574
rect 225234 202000 225854 226338
rect 228954 698614 229574 710042
rect 246954 711558 247574 711590
rect 246954 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 247574 711558
rect 246954 711238 247574 711322
rect 246954 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 247574 711238
rect 243234 709638 243854 709670
rect 243234 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 243854 709638
rect 243234 709318 243854 709402
rect 243234 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 243854 709318
rect 239514 707718 240134 707750
rect 239514 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 240134 707718
rect 239514 707398 240134 707482
rect 239514 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 240134 707398
rect 228954 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 229574 698614
rect 228954 698294 229574 698378
rect 228954 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 229574 698294
rect 228954 662614 229574 698058
rect 228954 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 229574 662614
rect 228954 662294 229574 662378
rect 228954 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 229574 662294
rect 228954 626614 229574 662058
rect 228954 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 229574 626614
rect 228954 626294 229574 626378
rect 228954 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 229574 626294
rect 228954 590614 229574 626058
rect 228954 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 229574 590614
rect 228954 590294 229574 590378
rect 228954 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 229574 590294
rect 228954 554614 229574 590058
rect 228954 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 229574 554614
rect 228954 554294 229574 554378
rect 228954 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 229574 554294
rect 228954 518614 229574 554058
rect 228954 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 229574 518614
rect 228954 518294 229574 518378
rect 228954 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 229574 518294
rect 228954 482614 229574 518058
rect 228954 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 229574 482614
rect 228954 482294 229574 482378
rect 228954 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 229574 482294
rect 228954 446614 229574 482058
rect 228954 446378 228986 446614
rect 229222 446378 229306 446614
rect 229542 446378 229574 446614
rect 228954 446294 229574 446378
rect 228954 446058 228986 446294
rect 229222 446058 229306 446294
rect 229542 446058 229574 446294
rect 228954 410614 229574 446058
rect 228954 410378 228986 410614
rect 229222 410378 229306 410614
rect 229542 410378 229574 410614
rect 228954 410294 229574 410378
rect 228954 410058 228986 410294
rect 229222 410058 229306 410294
rect 229542 410058 229574 410294
rect 228954 374614 229574 410058
rect 228954 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 229574 374614
rect 228954 374294 229574 374378
rect 228954 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 229574 374294
rect 228954 338614 229574 374058
rect 228954 338378 228986 338614
rect 229222 338378 229306 338614
rect 229542 338378 229574 338614
rect 228954 338294 229574 338378
rect 228954 338058 228986 338294
rect 229222 338058 229306 338294
rect 229542 338058 229574 338294
rect 228954 302614 229574 338058
rect 228954 302378 228986 302614
rect 229222 302378 229306 302614
rect 229542 302378 229574 302614
rect 228954 302294 229574 302378
rect 228954 302058 228986 302294
rect 229222 302058 229306 302294
rect 229542 302058 229574 302294
rect 228954 266614 229574 302058
rect 228954 266378 228986 266614
rect 229222 266378 229306 266614
rect 229542 266378 229574 266614
rect 228954 266294 229574 266378
rect 228954 266058 228986 266294
rect 229222 266058 229306 266294
rect 229542 266058 229574 266294
rect 228954 230614 229574 266058
rect 228954 230378 228986 230614
rect 229222 230378 229306 230614
rect 229542 230378 229574 230614
rect 228954 230294 229574 230378
rect 228954 230058 228986 230294
rect 229222 230058 229306 230294
rect 229542 230058 229574 230294
rect 228954 202000 229574 230058
rect 235794 705798 236414 705830
rect 235794 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 236414 705798
rect 235794 705478 236414 705562
rect 235794 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 236414 705478
rect 235794 669454 236414 705242
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 597454 236414 632898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 561454 236414 596898
rect 235794 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 236414 561454
rect 235794 561134 236414 561218
rect 235794 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 236414 561134
rect 235794 525454 236414 560898
rect 235794 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 236414 525454
rect 235794 525134 236414 525218
rect 235794 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 236414 525134
rect 235794 489454 236414 524898
rect 235794 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 236414 489454
rect 235794 489134 236414 489218
rect 235794 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 236414 489134
rect 235794 453454 236414 488898
rect 235794 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 236414 453454
rect 235794 453134 236414 453218
rect 235794 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 236414 453134
rect 235794 417454 236414 452898
rect 235794 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 236414 417454
rect 235794 417134 236414 417218
rect 235794 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 236414 417134
rect 235794 381454 236414 416898
rect 235794 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 236414 381454
rect 235794 381134 236414 381218
rect 235794 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 236414 381134
rect 235794 345454 236414 380898
rect 235794 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 236414 345454
rect 235794 345134 236414 345218
rect 235794 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 236414 345134
rect 235794 309454 236414 344898
rect 235794 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 236414 309454
rect 235794 309134 236414 309218
rect 235794 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 236414 309134
rect 235794 273454 236414 308898
rect 235794 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 236414 273454
rect 235794 273134 236414 273218
rect 235794 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 236414 273134
rect 235794 237454 236414 272898
rect 235794 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 236414 237454
rect 235794 237134 236414 237218
rect 235794 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 236414 237134
rect 235794 202000 236414 236898
rect 239514 673174 240134 707162
rect 239514 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 240134 673174
rect 239514 672854 240134 672938
rect 239514 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 240134 672854
rect 239514 637174 240134 672618
rect 239514 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 240134 637174
rect 239514 636854 240134 636938
rect 239514 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 240134 636854
rect 239514 601174 240134 636618
rect 239514 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 240134 601174
rect 239514 600854 240134 600938
rect 239514 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 240134 600854
rect 239514 565174 240134 600618
rect 239514 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 240134 565174
rect 239514 564854 240134 564938
rect 239514 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 240134 564854
rect 239514 529174 240134 564618
rect 239514 528938 239546 529174
rect 239782 528938 239866 529174
rect 240102 528938 240134 529174
rect 239514 528854 240134 528938
rect 239514 528618 239546 528854
rect 239782 528618 239866 528854
rect 240102 528618 240134 528854
rect 239514 493174 240134 528618
rect 239514 492938 239546 493174
rect 239782 492938 239866 493174
rect 240102 492938 240134 493174
rect 239514 492854 240134 492938
rect 239514 492618 239546 492854
rect 239782 492618 239866 492854
rect 240102 492618 240134 492854
rect 239514 457174 240134 492618
rect 239514 456938 239546 457174
rect 239782 456938 239866 457174
rect 240102 456938 240134 457174
rect 239514 456854 240134 456938
rect 239514 456618 239546 456854
rect 239782 456618 239866 456854
rect 240102 456618 240134 456854
rect 239514 421174 240134 456618
rect 239514 420938 239546 421174
rect 239782 420938 239866 421174
rect 240102 420938 240134 421174
rect 239514 420854 240134 420938
rect 239514 420618 239546 420854
rect 239782 420618 239866 420854
rect 240102 420618 240134 420854
rect 239514 385174 240134 420618
rect 239514 384938 239546 385174
rect 239782 384938 239866 385174
rect 240102 384938 240134 385174
rect 239514 384854 240134 384938
rect 239514 384618 239546 384854
rect 239782 384618 239866 384854
rect 240102 384618 240134 384854
rect 239514 349174 240134 384618
rect 239514 348938 239546 349174
rect 239782 348938 239866 349174
rect 240102 348938 240134 349174
rect 239514 348854 240134 348938
rect 239514 348618 239546 348854
rect 239782 348618 239866 348854
rect 240102 348618 240134 348854
rect 239514 313174 240134 348618
rect 239514 312938 239546 313174
rect 239782 312938 239866 313174
rect 240102 312938 240134 313174
rect 239514 312854 240134 312938
rect 239514 312618 239546 312854
rect 239782 312618 239866 312854
rect 240102 312618 240134 312854
rect 239514 277174 240134 312618
rect 239514 276938 239546 277174
rect 239782 276938 239866 277174
rect 240102 276938 240134 277174
rect 239514 276854 240134 276938
rect 239514 276618 239546 276854
rect 239782 276618 239866 276854
rect 240102 276618 240134 276854
rect 239514 241174 240134 276618
rect 239514 240938 239546 241174
rect 239782 240938 239866 241174
rect 240102 240938 240134 241174
rect 239514 240854 240134 240938
rect 239514 240618 239546 240854
rect 239782 240618 239866 240854
rect 240102 240618 240134 240854
rect 239514 205174 240134 240618
rect 239514 204938 239546 205174
rect 239782 204938 239866 205174
rect 240102 204938 240134 205174
rect 239514 204854 240134 204938
rect 239514 204618 239546 204854
rect 239782 204618 239866 204854
rect 240102 204618 240134 204854
rect 239514 202000 240134 204618
rect 243234 676894 243854 709082
rect 243234 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 243854 676894
rect 243234 676574 243854 676658
rect 243234 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 243854 676574
rect 243234 640894 243854 676338
rect 243234 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 243854 640894
rect 243234 640574 243854 640658
rect 243234 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 243854 640574
rect 243234 604894 243854 640338
rect 243234 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 243854 604894
rect 243234 604574 243854 604658
rect 243234 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 243854 604574
rect 243234 568894 243854 604338
rect 243234 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 243854 568894
rect 243234 568574 243854 568658
rect 243234 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 243854 568574
rect 243234 532894 243854 568338
rect 243234 532658 243266 532894
rect 243502 532658 243586 532894
rect 243822 532658 243854 532894
rect 243234 532574 243854 532658
rect 243234 532338 243266 532574
rect 243502 532338 243586 532574
rect 243822 532338 243854 532574
rect 243234 496894 243854 532338
rect 243234 496658 243266 496894
rect 243502 496658 243586 496894
rect 243822 496658 243854 496894
rect 243234 496574 243854 496658
rect 243234 496338 243266 496574
rect 243502 496338 243586 496574
rect 243822 496338 243854 496574
rect 243234 460894 243854 496338
rect 243234 460658 243266 460894
rect 243502 460658 243586 460894
rect 243822 460658 243854 460894
rect 243234 460574 243854 460658
rect 243234 460338 243266 460574
rect 243502 460338 243586 460574
rect 243822 460338 243854 460574
rect 243234 424894 243854 460338
rect 243234 424658 243266 424894
rect 243502 424658 243586 424894
rect 243822 424658 243854 424894
rect 243234 424574 243854 424658
rect 243234 424338 243266 424574
rect 243502 424338 243586 424574
rect 243822 424338 243854 424574
rect 243234 388894 243854 424338
rect 243234 388658 243266 388894
rect 243502 388658 243586 388894
rect 243822 388658 243854 388894
rect 243234 388574 243854 388658
rect 243234 388338 243266 388574
rect 243502 388338 243586 388574
rect 243822 388338 243854 388574
rect 243234 352894 243854 388338
rect 243234 352658 243266 352894
rect 243502 352658 243586 352894
rect 243822 352658 243854 352894
rect 243234 352574 243854 352658
rect 243234 352338 243266 352574
rect 243502 352338 243586 352574
rect 243822 352338 243854 352574
rect 243234 316894 243854 352338
rect 243234 316658 243266 316894
rect 243502 316658 243586 316894
rect 243822 316658 243854 316894
rect 243234 316574 243854 316658
rect 243234 316338 243266 316574
rect 243502 316338 243586 316574
rect 243822 316338 243854 316574
rect 243234 280894 243854 316338
rect 243234 280658 243266 280894
rect 243502 280658 243586 280894
rect 243822 280658 243854 280894
rect 243234 280574 243854 280658
rect 243234 280338 243266 280574
rect 243502 280338 243586 280574
rect 243822 280338 243854 280574
rect 243234 244894 243854 280338
rect 243234 244658 243266 244894
rect 243502 244658 243586 244894
rect 243822 244658 243854 244894
rect 243234 244574 243854 244658
rect 243234 244338 243266 244574
rect 243502 244338 243586 244574
rect 243822 244338 243854 244574
rect 243234 208894 243854 244338
rect 243234 208658 243266 208894
rect 243502 208658 243586 208894
rect 243822 208658 243854 208894
rect 243234 208574 243854 208658
rect 243234 208338 243266 208574
rect 243502 208338 243586 208574
rect 243822 208338 243854 208574
rect 243234 202000 243854 208338
rect 246954 680614 247574 711002
rect 264954 710598 265574 711590
rect 264954 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 265574 710598
rect 264954 710278 265574 710362
rect 264954 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 265574 710278
rect 261234 708678 261854 709670
rect 261234 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 261854 708678
rect 261234 708358 261854 708442
rect 261234 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 261854 708358
rect 257514 706758 258134 707750
rect 257514 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 258134 706758
rect 257514 706438 258134 706522
rect 257514 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 258134 706438
rect 246954 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 247574 680614
rect 246954 680294 247574 680378
rect 246954 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 247574 680294
rect 246954 644614 247574 680058
rect 246954 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 247574 644614
rect 246954 644294 247574 644378
rect 246954 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 247574 644294
rect 246954 608614 247574 644058
rect 246954 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 247574 608614
rect 246954 608294 247574 608378
rect 246954 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 247574 608294
rect 246954 572614 247574 608058
rect 246954 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 247574 572614
rect 246954 572294 247574 572378
rect 246954 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 247574 572294
rect 246954 536614 247574 572058
rect 246954 536378 246986 536614
rect 247222 536378 247306 536614
rect 247542 536378 247574 536614
rect 246954 536294 247574 536378
rect 246954 536058 246986 536294
rect 247222 536058 247306 536294
rect 247542 536058 247574 536294
rect 246954 500614 247574 536058
rect 246954 500378 246986 500614
rect 247222 500378 247306 500614
rect 247542 500378 247574 500614
rect 246954 500294 247574 500378
rect 246954 500058 246986 500294
rect 247222 500058 247306 500294
rect 247542 500058 247574 500294
rect 246954 464614 247574 500058
rect 246954 464378 246986 464614
rect 247222 464378 247306 464614
rect 247542 464378 247574 464614
rect 246954 464294 247574 464378
rect 246954 464058 246986 464294
rect 247222 464058 247306 464294
rect 247542 464058 247574 464294
rect 246954 428614 247574 464058
rect 246954 428378 246986 428614
rect 247222 428378 247306 428614
rect 247542 428378 247574 428614
rect 246954 428294 247574 428378
rect 246954 428058 246986 428294
rect 247222 428058 247306 428294
rect 247542 428058 247574 428294
rect 246954 392614 247574 428058
rect 246954 392378 246986 392614
rect 247222 392378 247306 392614
rect 247542 392378 247574 392614
rect 246954 392294 247574 392378
rect 246954 392058 246986 392294
rect 247222 392058 247306 392294
rect 247542 392058 247574 392294
rect 246954 356614 247574 392058
rect 246954 356378 246986 356614
rect 247222 356378 247306 356614
rect 247542 356378 247574 356614
rect 246954 356294 247574 356378
rect 246954 356058 246986 356294
rect 247222 356058 247306 356294
rect 247542 356058 247574 356294
rect 246954 320614 247574 356058
rect 246954 320378 246986 320614
rect 247222 320378 247306 320614
rect 247542 320378 247574 320614
rect 246954 320294 247574 320378
rect 246954 320058 246986 320294
rect 247222 320058 247306 320294
rect 247542 320058 247574 320294
rect 246954 284614 247574 320058
rect 246954 284378 246986 284614
rect 247222 284378 247306 284614
rect 247542 284378 247574 284614
rect 246954 284294 247574 284378
rect 246954 284058 246986 284294
rect 247222 284058 247306 284294
rect 247542 284058 247574 284294
rect 246954 248614 247574 284058
rect 246954 248378 246986 248614
rect 247222 248378 247306 248614
rect 247542 248378 247574 248614
rect 246954 248294 247574 248378
rect 246954 248058 246986 248294
rect 247222 248058 247306 248294
rect 247542 248058 247574 248294
rect 246954 212614 247574 248058
rect 246954 212378 246986 212614
rect 247222 212378 247306 212614
rect 247542 212378 247574 212614
rect 246954 212294 247574 212378
rect 246954 212058 246986 212294
rect 247222 212058 247306 212294
rect 247542 212058 247574 212294
rect 246954 202000 247574 212058
rect 253794 704838 254414 705830
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 543454 254414 578898
rect 253794 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 254414 543454
rect 253794 543134 254414 543218
rect 253794 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 254414 543134
rect 253794 507454 254414 542898
rect 253794 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 254414 507454
rect 253794 507134 254414 507218
rect 253794 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 254414 507134
rect 253794 471454 254414 506898
rect 253794 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 254414 471454
rect 253794 471134 254414 471218
rect 253794 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 254414 471134
rect 253794 435454 254414 470898
rect 253794 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 254414 435454
rect 253794 435134 254414 435218
rect 253794 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 254414 435134
rect 253794 399454 254414 434898
rect 253794 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 254414 399454
rect 253794 399134 254414 399218
rect 253794 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 254414 399134
rect 253794 363454 254414 398898
rect 253794 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 254414 363454
rect 253794 363134 254414 363218
rect 253794 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 254414 363134
rect 253794 327454 254414 362898
rect 253794 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 254414 327454
rect 253794 327134 254414 327218
rect 253794 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 254414 327134
rect 253794 291454 254414 326898
rect 253794 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 254414 291454
rect 253794 291134 254414 291218
rect 253794 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 254414 291134
rect 253794 255454 254414 290898
rect 253794 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 254414 255454
rect 253794 255134 254414 255218
rect 253794 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 254414 255134
rect 253794 219454 254414 254898
rect 253794 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 254414 219454
rect 253794 219134 254414 219218
rect 253794 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 254414 219134
rect 253794 202000 254414 218898
rect 257514 691174 258134 706202
rect 257514 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 258134 691174
rect 257514 690854 258134 690938
rect 257514 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 258134 690854
rect 257514 655174 258134 690618
rect 257514 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 258134 655174
rect 257514 654854 258134 654938
rect 257514 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 258134 654854
rect 257514 619174 258134 654618
rect 257514 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 258134 619174
rect 257514 618854 258134 618938
rect 257514 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 258134 618854
rect 257514 583174 258134 618618
rect 257514 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 258134 583174
rect 257514 582854 258134 582938
rect 257514 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 258134 582854
rect 257514 547174 258134 582618
rect 257514 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 258134 547174
rect 257514 546854 258134 546938
rect 257514 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 258134 546854
rect 257514 511174 258134 546618
rect 257514 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 258134 511174
rect 257514 510854 258134 510938
rect 257514 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 258134 510854
rect 257514 475174 258134 510618
rect 257514 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 258134 475174
rect 257514 474854 258134 474938
rect 257514 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 258134 474854
rect 257514 439174 258134 474618
rect 257514 438938 257546 439174
rect 257782 438938 257866 439174
rect 258102 438938 258134 439174
rect 257514 438854 258134 438938
rect 257514 438618 257546 438854
rect 257782 438618 257866 438854
rect 258102 438618 258134 438854
rect 257514 403174 258134 438618
rect 257514 402938 257546 403174
rect 257782 402938 257866 403174
rect 258102 402938 258134 403174
rect 257514 402854 258134 402938
rect 257514 402618 257546 402854
rect 257782 402618 257866 402854
rect 258102 402618 258134 402854
rect 257514 367174 258134 402618
rect 257514 366938 257546 367174
rect 257782 366938 257866 367174
rect 258102 366938 258134 367174
rect 257514 366854 258134 366938
rect 257514 366618 257546 366854
rect 257782 366618 257866 366854
rect 258102 366618 258134 366854
rect 257514 331174 258134 366618
rect 257514 330938 257546 331174
rect 257782 330938 257866 331174
rect 258102 330938 258134 331174
rect 257514 330854 258134 330938
rect 257514 330618 257546 330854
rect 257782 330618 257866 330854
rect 258102 330618 258134 330854
rect 257514 295174 258134 330618
rect 257514 294938 257546 295174
rect 257782 294938 257866 295174
rect 258102 294938 258134 295174
rect 257514 294854 258134 294938
rect 257514 294618 257546 294854
rect 257782 294618 257866 294854
rect 258102 294618 258134 294854
rect 257514 259174 258134 294618
rect 257514 258938 257546 259174
rect 257782 258938 257866 259174
rect 258102 258938 258134 259174
rect 257514 258854 258134 258938
rect 257514 258618 257546 258854
rect 257782 258618 257866 258854
rect 258102 258618 258134 258854
rect 257514 223174 258134 258618
rect 257514 222938 257546 223174
rect 257782 222938 257866 223174
rect 258102 222938 258134 223174
rect 257514 222854 258134 222938
rect 257514 222618 257546 222854
rect 257782 222618 257866 222854
rect 258102 222618 258134 222854
rect 257514 202000 258134 222618
rect 261234 694894 261854 708122
rect 261234 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 261854 694894
rect 261234 694574 261854 694658
rect 261234 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 261854 694574
rect 261234 658894 261854 694338
rect 261234 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 261854 658894
rect 261234 658574 261854 658658
rect 261234 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 261854 658574
rect 261234 622894 261854 658338
rect 261234 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 261854 622894
rect 261234 622574 261854 622658
rect 261234 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 261854 622574
rect 261234 586894 261854 622338
rect 261234 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 261854 586894
rect 261234 586574 261854 586658
rect 261234 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 261854 586574
rect 261234 550894 261854 586338
rect 261234 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 261854 550894
rect 261234 550574 261854 550658
rect 261234 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 261854 550574
rect 261234 514894 261854 550338
rect 261234 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 261854 514894
rect 261234 514574 261854 514658
rect 261234 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 261854 514574
rect 261234 478894 261854 514338
rect 261234 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 261854 478894
rect 261234 478574 261854 478658
rect 261234 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 261854 478574
rect 261234 442894 261854 478338
rect 261234 442658 261266 442894
rect 261502 442658 261586 442894
rect 261822 442658 261854 442894
rect 261234 442574 261854 442658
rect 261234 442338 261266 442574
rect 261502 442338 261586 442574
rect 261822 442338 261854 442574
rect 261234 406894 261854 442338
rect 261234 406658 261266 406894
rect 261502 406658 261586 406894
rect 261822 406658 261854 406894
rect 261234 406574 261854 406658
rect 261234 406338 261266 406574
rect 261502 406338 261586 406574
rect 261822 406338 261854 406574
rect 261234 370894 261854 406338
rect 261234 370658 261266 370894
rect 261502 370658 261586 370894
rect 261822 370658 261854 370894
rect 261234 370574 261854 370658
rect 261234 370338 261266 370574
rect 261502 370338 261586 370574
rect 261822 370338 261854 370574
rect 261234 334894 261854 370338
rect 261234 334658 261266 334894
rect 261502 334658 261586 334894
rect 261822 334658 261854 334894
rect 261234 334574 261854 334658
rect 261234 334338 261266 334574
rect 261502 334338 261586 334574
rect 261822 334338 261854 334574
rect 261234 298894 261854 334338
rect 261234 298658 261266 298894
rect 261502 298658 261586 298894
rect 261822 298658 261854 298894
rect 261234 298574 261854 298658
rect 261234 298338 261266 298574
rect 261502 298338 261586 298574
rect 261822 298338 261854 298574
rect 261234 262894 261854 298338
rect 261234 262658 261266 262894
rect 261502 262658 261586 262894
rect 261822 262658 261854 262894
rect 261234 262574 261854 262658
rect 261234 262338 261266 262574
rect 261502 262338 261586 262574
rect 261822 262338 261854 262574
rect 261234 226894 261854 262338
rect 261234 226658 261266 226894
rect 261502 226658 261586 226894
rect 261822 226658 261854 226894
rect 261234 226574 261854 226658
rect 261234 226338 261266 226574
rect 261502 226338 261586 226574
rect 261822 226338 261854 226574
rect 261234 202000 261854 226338
rect 264954 698614 265574 710042
rect 282954 711558 283574 711590
rect 282954 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 283574 711558
rect 282954 711238 283574 711322
rect 282954 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 283574 711238
rect 279234 709638 279854 709670
rect 279234 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 279854 709638
rect 279234 709318 279854 709402
rect 279234 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 279854 709318
rect 275514 707718 276134 707750
rect 275514 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 276134 707718
rect 275514 707398 276134 707482
rect 275514 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 276134 707398
rect 264954 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 265574 698614
rect 264954 698294 265574 698378
rect 264954 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 265574 698294
rect 264954 662614 265574 698058
rect 264954 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 265574 662614
rect 264954 662294 265574 662378
rect 264954 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 265574 662294
rect 264954 626614 265574 662058
rect 264954 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 265574 626614
rect 264954 626294 265574 626378
rect 264954 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 265574 626294
rect 264954 590614 265574 626058
rect 264954 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 265574 590614
rect 264954 590294 265574 590378
rect 264954 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 265574 590294
rect 264954 554614 265574 590058
rect 264954 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 265574 554614
rect 264954 554294 265574 554378
rect 264954 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 265574 554294
rect 264954 518614 265574 554058
rect 264954 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 265574 518614
rect 264954 518294 265574 518378
rect 264954 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 265574 518294
rect 264954 482614 265574 518058
rect 264954 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 265574 482614
rect 264954 482294 265574 482378
rect 264954 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 265574 482294
rect 264954 446614 265574 482058
rect 264954 446378 264986 446614
rect 265222 446378 265306 446614
rect 265542 446378 265574 446614
rect 264954 446294 265574 446378
rect 264954 446058 264986 446294
rect 265222 446058 265306 446294
rect 265542 446058 265574 446294
rect 264954 410614 265574 446058
rect 264954 410378 264986 410614
rect 265222 410378 265306 410614
rect 265542 410378 265574 410614
rect 264954 410294 265574 410378
rect 264954 410058 264986 410294
rect 265222 410058 265306 410294
rect 265542 410058 265574 410294
rect 264954 374614 265574 410058
rect 264954 374378 264986 374614
rect 265222 374378 265306 374614
rect 265542 374378 265574 374614
rect 264954 374294 265574 374378
rect 264954 374058 264986 374294
rect 265222 374058 265306 374294
rect 265542 374058 265574 374294
rect 264954 338614 265574 374058
rect 264954 338378 264986 338614
rect 265222 338378 265306 338614
rect 265542 338378 265574 338614
rect 264954 338294 265574 338378
rect 264954 338058 264986 338294
rect 265222 338058 265306 338294
rect 265542 338058 265574 338294
rect 264954 302614 265574 338058
rect 264954 302378 264986 302614
rect 265222 302378 265306 302614
rect 265542 302378 265574 302614
rect 264954 302294 265574 302378
rect 264954 302058 264986 302294
rect 265222 302058 265306 302294
rect 265542 302058 265574 302294
rect 264954 266614 265574 302058
rect 264954 266378 264986 266614
rect 265222 266378 265306 266614
rect 265542 266378 265574 266614
rect 264954 266294 265574 266378
rect 264954 266058 264986 266294
rect 265222 266058 265306 266294
rect 265542 266058 265574 266294
rect 264954 230614 265574 266058
rect 264954 230378 264986 230614
rect 265222 230378 265306 230614
rect 265542 230378 265574 230614
rect 264954 230294 265574 230378
rect 264954 230058 264986 230294
rect 265222 230058 265306 230294
rect 265542 230058 265574 230294
rect 264954 202000 265574 230058
rect 271794 705798 272414 705830
rect 271794 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 272414 705798
rect 271794 705478 272414 705562
rect 271794 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 272414 705478
rect 271794 669454 272414 705242
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 561454 272414 596898
rect 271794 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 272414 561454
rect 271794 561134 272414 561218
rect 271794 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 272414 561134
rect 271794 525454 272414 560898
rect 271794 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 272414 525454
rect 271794 525134 272414 525218
rect 271794 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 272414 525134
rect 271794 489454 272414 524898
rect 271794 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 272414 489454
rect 271794 489134 272414 489218
rect 271794 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 272414 489134
rect 271794 453454 272414 488898
rect 271794 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 272414 453454
rect 271794 453134 272414 453218
rect 271794 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 272414 453134
rect 271794 417454 272414 452898
rect 271794 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 272414 417454
rect 271794 417134 272414 417218
rect 271794 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 272414 417134
rect 271794 381454 272414 416898
rect 271794 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 272414 381454
rect 271794 381134 272414 381218
rect 271794 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 272414 381134
rect 271794 345454 272414 380898
rect 271794 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 272414 345454
rect 271794 345134 272414 345218
rect 271794 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 272414 345134
rect 271794 309454 272414 344898
rect 271794 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 272414 309454
rect 271794 309134 272414 309218
rect 271794 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 272414 309134
rect 271794 273454 272414 308898
rect 271794 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 272414 273454
rect 271794 273134 272414 273218
rect 271794 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 272414 273134
rect 271794 237454 272414 272898
rect 271794 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 272414 237454
rect 271794 237134 272414 237218
rect 271794 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 272414 237134
rect 271794 202000 272414 236898
rect 275514 673174 276134 707162
rect 275514 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 276134 673174
rect 275514 672854 276134 672938
rect 275514 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 276134 672854
rect 275514 637174 276134 672618
rect 275514 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 276134 637174
rect 275514 636854 276134 636938
rect 275514 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 276134 636854
rect 275514 601174 276134 636618
rect 275514 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 276134 601174
rect 275514 600854 276134 600938
rect 275514 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 276134 600854
rect 275514 565174 276134 600618
rect 275514 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 276134 565174
rect 275514 564854 276134 564938
rect 275514 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 276134 564854
rect 275514 529174 276134 564618
rect 275514 528938 275546 529174
rect 275782 528938 275866 529174
rect 276102 528938 276134 529174
rect 275514 528854 276134 528938
rect 275514 528618 275546 528854
rect 275782 528618 275866 528854
rect 276102 528618 276134 528854
rect 275514 493174 276134 528618
rect 275514 492938 275546 493174
rect 275782 492938 275866 493174
rect 276102 492938 276134 493174
rect 275514 492854 276134 492938
rect 275514 492618 275546 492854
rect 275782 492618 275866 492854
rect 276102 492618 276134 492854
rect 275514 457174 276134 492618
rect 275514 456938 275546 457174
rect 275782 456938 275866 457174
rect 276102 456938 276134 457174
rect 275514 456854 276134 456938
rect 275514 456618 275546 456854
rect 275782 456618 275866 456854
rect 276102 456618 276134 456854
rect 275514 421174 276134 456618
rect 275514 420938 275546 421174
rect 275782 420938 275866 421174
rect 276102 420938 276134 421174
rect 275514 420854 276134 420938
rect 275514 420618 275546 420854
rect 275782 420618 275866 420854
rect 276102 420618 276134 420854
rect 275514 385174 276134 420618
rect 275514 384938 275546 385174
rect 275782 384938 275866 385174
rect 276102 384938 276134 385174
rect 275514 384854 276134 384938
rect 275514 384618 275546 384854
rect 275782 384618 275866 384854
rect 276102 384618 276134 384854
rect 275514 349174 276134 384618
rect 275514 348938 275546 349174
rect 275782 348938 275866 349174
rect 276102 348938 276134 349174
rect 275514 348854 276134 348938
rect 275514 348618 275546 348854
rect 275782 348618 275866 348854
rect 276102 348618 276134 348854
rect 275514 313174 276134 348618
rect 275514 312938 275546 313174
rect 275782 312938 275866 313174
rect 276102 312938 276134 313174
rect 275514 312854 276134 312938
rect 275514 312618 275546 312854
rect 275782 312618 275866 312854
rect 276102 312618 276134 312854
rect 275514 277174 276134 312618
rect 275514 276938 275546 277174
rect 275782 276938 275866 277174
rect 276102 276938 276134 277174
rect 275514 276854 276134 276938
rect 275514 276618 275546 276854
rect 275782 276618 275866 276854
rect 276102 276618 276134 276854
rect 275514 241174 276134 276618
rect 275514 240938 275546 241174
rect 275782 240938 275866 241174
rect 276102 240938 276134 241174
rect 275514 240854 276134 240938
rect 275514 240618 275546 240854
rect 275782 240618 275866 240854
rect 276102 240618 276134 240854
rect 275514 205174 276134 240618
rect 275514 204938 275546 205174
rect 275782 204938 275866 205174
rect 276102 204938 276134 205174
rect 275514 204854 276134 204938
rect 275514 204618 275546 204854
rect 275782 204618 275866 204854
rect 276102 204618 276134 204854
rect 275514 202000 276134 204618
rect 279234 676894 279854 709082
rect 279234 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 279854 676894
rect 279234 676574 279854 676658
rect 279234 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 279854 676574
rect 279234 640894 279854 676338
rect 279234 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 279854 640894
rect 279234 640574 279854 640658
rect 279234 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 279854 640574
rect 279234 604894 279854 640338
rect 279234 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 279854 604894
rect 279234 604574 279854 604658
rect 279234 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 279854 604574
rect 279234 568894 279854 604338
rect 279234 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 279854 568894
rect 279234 568574 279854 568658
rect 279234 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 279854 568574
rect 279234 532894 279854 568338
rect 279234 532658 279266 532894
rect 279502 532658 279586 532894
rect 279822 532658 279854 532894
rect 279234 532574 279854 532658
rect 279234 532338 279266 532574
rect 279502 532338 279586 532574
rect 279822 532338 279854 532574
rect 279234 496894 279854 532338
rect 279234 496658 279266 496894
rect 279502 496658 279586 496894
rect 279822 496658 279854 496894
rect 279234 496574 279854 496658
rect 279234 496338 279266 496574
rect 279502 496338 279586 496574
rect 279822 496338 279854 496574
rect 279234 460894 279854 496338
rect 279234 460658 279266 460894
rect 279502 460658 279586 460894
rect 279822 460658 279854 460894
rect 279234 460574 279854 460658
rect 279234 460338 279266 460574
rect 279502 460338 279586 460574
rect 279822 460338 279854 460574
rect 279234 424894 279854 460338
rect 279234 424658 279266 424894
rect 279502 424658 279586 424894
rect 279822 424658 279854 424894
rect 279234 424574 279854 424658
rect 279234 424338 279266 424574
rect 279502 424338 279586 424574
rect 279822 424338 279854 424574
rect 279234 388894 279854 424338
rect 279234 388658 279266 388894
rect 279502 388658 279586 388894
rect 279822 388658 279854 388894
rect 279234 388574 279854 388658
rect 279234 388338 279266 388574
rect 279502 388338 279586 388574
rect 279822 388338 279854 388574
rect 279234 352894 279854 388338
rect 279234 352658 279266 352894
rect 279502 352658 279586 352894
rect 279822 352658 279854 352894
rect 279234 352574 279854 352658
rect 279234 352338 279266 352574
rect 279502 352338 279586 352574
rect 279822 352338 279854 352574
rect 279234 316894 279854 352338
rect 279234 316658 279266 316894
rect 279502 316658 279586 316894
rect 279822 316658 279854 316894
rect 279234 316574 279854 316658
rect 279234 316338 279266 316574
rect 279502 316338 279586 316574
rect 279822 316338 279854 316574
rect 279234 280894 279854 316338
rect 279234 280658 279266 280894
rect 279502 280658 279586 280894
rect 279822 280658 279854 280894
rect 279234 280574 279854 280658
rect 279234 280338 279266 280574
rect 279502 280338 279586 280574
rect 279822 280338 279854 280574
rect 279234 244894 279854 280338
rect 279234 244658 279266 244894
rect 279502 244658 279586 244894
rect 279822 244658 279854 244894
rect 279234 244574 279854 244658
rect 279234 244338 279266 244574
rect 279502 244338 279586 244574
rect 279822 244338 279854 244574
rect 279234 208894 279854 244338
rect 279234 208658 279266 208894
rect 279502 208658 279586 208894
rect 279822 208658 279854 208894
rect 279234 208574 279854 208658
rect 279234 208338 279266 208574
rect 279502 208338 279586 208574
rect 279822 208338 279854 208574
rect 279234 202000 279854 208338
rect 282954 680614 283574 711002
rect 300954 710598 301574 711590
rect 300954 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 301574 710598
rect 300954 710278 301574 710362
rect 300954 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 301574 710278
rect 297234 708678 297854 709670
rect 297234 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 297854 708678
rect 297234 708358 297854 708442
rect 297234 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 297854 708358
rect 293514 706758 294134 707750
rect 293514 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 294134 706758
rect 293514 706438 294134 706522
rect 293514 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 294134 706438
rect 282954 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 283574 680614
rect 282954 680294 283574 680378
rect 282954 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 283574 680294
rect 282954 644614 283574 680058
rect 282954 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 283574 644614
rect 282954 644294 283574 644378
rect 282954 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 283574 644294
rect 282954 608614 283574 644058
rect 282954 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 283574 608614
rect 282954 608294 283574 608378
rect 282954 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 283574 608294
rect 282954 572614 283574 608058
rect 282954 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 283574 572614
rect 282954 572294 283574 572378
rect 282954 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 283574 572294
rect 282954 536614 283574 572058
rect 282954 536378 282986 536614
rect 283222 536378 283306 536614
rect 283542 536378 283574 536614
rect 282954 536294 283574 536378
rect 282954 536058 282986 536294
rect 283222 536058 283306 536294
rect 283542 536058 283574 536294
rect 282954 500614 283574 536058
rect 282954 500378 282986 500614
rect 283222 500378 283306 500614
rect 283542 500378 283574 500614
rect 282954 500294 283574 500378
rect 282954 500058 282986 500294
rect 283222 500058 283306 500294
rect 283542 500058 283574 500294
rect 282954 464614 283574 500058
rect 282954 464378 282986 464614
rect 283222 464378 283306 464614
rect 283542 464378 283574 464614
rect 282954 464294 283574 464378
rect 282954 464058 282986 464294
rect 283222 464058 283306 464294
rect 283542 464058 283574 464294
rect 282954 428614 283574 464058
rect 282954 428378 282986 428614
rect 283222 428378 283306 428614
rect 283542 428378 283574 428614
rect 282954 428294 283574 428378
rect 282954 428058 282986 428294
rect 283222 428058 283306 428294
rect 283542 428058 283574 428294
rect 282954 392614 283574 428058
rect 282954 392378 282986 392614
rect 283222 392378 283306 392614
rect 283542 392378 283574 392614
rect 282954 392294 283574 392378
rect 282954 392058 282986 392294
rect 283222 392058 283306 392294
rect 283542 392058 283574 392294
rect 282954 356614 283574 392058
rect 282954 356378 282986 356614
rect 283222 356378 283306 356614
rect 283542 356378 283574 356614
rect 282954 356294 283574 356378
rect 282954 356058 282986 356294
rect 283222 356058 283306 356294
rect 283542 356058 283574 356294
rect 282954 320614 283574 356058
rect 282954 320378 282986 320614
rect 283222 320378 283306 320614
rect 283542 320378 283574 320614
rect 282954 320294 283574 320378
rect 282954 320058 282986 320294
rect 283222 320058 283306 320294
rect 283542 320058 283574 320294
rect 282954 284614 283574 320058
rect 282954 284378 282986 284614
rect 283222 284378 283306 284614
rect 283542 284378 283574 284614
rect 282954 284294 283574 284378
rect 282954 284058 282986 284294
rect 283222 284058 283306 284294
rect 283542 284058 283574 284294
rect 282954 248614 283574 284058
rect 282954 248378 282986 248614
rect 283222 248378 283306 248614
rect 283542 248378 283574 248614
rect 282954 248294 283574 248378
rect 282954 248058 282986 248294
rect 283222 248058 283306 248294
rect 283542 248058 283574 248294
rect 282954 212614 283574 248058
rect 282954 212378 282986 212614
rect 283222 212378 283306 212614
rect 283542 212378 283574 212614
rect 282954 212294 283574 212378
rect 282954 212058 282986 212294
rect 283222 212058 283306 212294
rect 283542 212058 283574 212294
rect 282954 202000 283574 212058
rect 289794 704838 290414 705830
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 543454 290414 578898
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289794 507454 290414 542898
rect 289794 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 290414 507454
rect 289794 507134 290414 507218
rect 289794 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 290414 507134
rect 289794 471454 290414 506898
rect 289794 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 290414 471454
rect 289794 471134 290414 471218
rect 289794 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 290414 471134
rect 289794 435454 290414 470898
rect 289794 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 290414 435454
rect 289794 435134 290414 435218
rect 289794 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 290414 435134
rect 289794 399454 290414 434898
rect 289794 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 290414 399454
rect 289794 399134 290414 399218
rect 289794 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 290414 399134
rect 289794 363454 290414 398898
rect 289794 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 290414 363454
rect 289794 363134 290414 363218
rect 289794 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 290414 363134
rect 289794 327454 290414 362898
rect 289794 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 290414 327454
rect 289794 327134 290414 327218
rect 289794 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 290414 327134
rect 289794 291454 290414 326898
rect 289794 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 290414 291454
rect 289794 291134 290414 291218
rect 289794 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 290414 291134
rect 289794 255454 290414 290898
rect 289794 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 290414 255454
rect 289794 255134 290414 255218
rect 289794 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 290414 255134
rect 289794 219454 290414 254898
rect 289794 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 290414 219454
rect 289794 219134 290414 219218
rect 289794 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 290414 219134
rect 289794 202000 290414 218898
rect 293514 691174 294134 706202
rect 293514 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 294134 691174
rect 293514 690854 294134 690938
rect 293514 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 294134 690854
rect 293514 655174 294134 690618
rect 293514 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 294134 655174
rect 293514 654854 294134 654938
rect 293514 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 294134 654854
rect 293514 619174 294134 654618
rect 293514 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 294134 619174
rect 293514 618854 294134 618938
rect 293514 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 294134 618854
rect 293514 583174 294134 618618
rect 293514 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 294134 583174
rect 293514 582854 294134 582938
rect 293514 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 294134 582854
rect 293514 547174 294134 582618
rect 293514 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 294134 547174
rect 293514 546854 294134 546938
rect 293514 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 294134 546854
rect 293514 511174 294134 546618
rect 293514 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 294134 511174
rect 293514 510854 294134 510938
rect 293514 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 294134 510854
rect 293514 475174 294134 510618
rect 293514 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 294134 475174
rect 293514 474854 294134 474938
rect 293514 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 294134 474854
rect 293514 439174 294134 474618
rect 293514 438938 293546 439174
rect 293782 438938 293866 439174
rect 294102 438938 294134 439174
rect 293514 438854 294134 438938
rect 293514 438618 293546 438854
rect 293782 438618 293866 438854
rect 294102 438618 294134 438854
rect 293514 403174 294134 438618
rect 293514 402938 293546 403174
rect 293782 402938 293866 403174
rect 294102 402938 294134 403174
rect 293514 402854 294134 402938
rect 293514 402618 293546 402854
rect 293782 402618 293866 402854
rect 294102 402618 294134 402854
rect 293514 367174 294134 402618
rect 293514 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 294134 367174
rect 293514 366854 294134 366938
rect 293514 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 294134 366854
rect 293514 331174 294134 366618
rect 293514 330938 293546 331174
rect 293782 330938 293866 331174
rect 294102 330938 294134 331174
rect 293514 330854 294134 330938
rect 293514 330618 293546 330854
rect 293782 330618 293866 330854
rect 294102 330618 294134 330854
rect 293514 295174 294134 330618
rect 293514 294938 293546 295174
rect 293782 294938 293866 295174
rect 294102 294938 294134 295174
rect 293514 294854 294134 294938
rect 293514 294618 293546 294854
rect 293782 294618 293866 294854
rect 294102 294618 294134 294854
rect 293514 259174 294134 294618
rect 293514 258938 293546 259174
rect 293782 258938 293866 259174
rect 294102 258938 294134 259174
rect 293514 258854 294134 258938
rect 293514 258618 293546 258854
rect 293782 258618 293866 258854
rect 294102 258618 294134 258854
rect 293514 223174 294134 258618
rect 293514 222938 293546 223174
rect 293782 222938 293866 223174
rect 294102 222938 294134 223174
rect 293514 222854 294134 222938
rect 293514 222618 293546 222854
rect 293782 222618 293866 222854
rect 294102 222618 294134 222854
rect 293514 202000 294134 222618
rect 297234 694894 297854 708122
rect 297234 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 297854 694894
rect 297234 694574 297854 694658
rect 297234 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 297854 694574
rect 297234 658894 297854 694338
rect 297234 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 297854 658894
rect 297234 658574 297854 658658
rect 297234 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 297854 658574
rect 297234 622894 297854 658338
rect 297234 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 297854 622894
rect 297234 622574 297854 622658
rect 297234 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 297854 622574
rect 297234 586894 297854 622338
rect 297234 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 297854 586894
rect 297234 586574 297854 586658
rect 297234 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 297854 586574
rect 297234 550894 297854 586338
rect 297234 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 297854 550894
rect 297234 550574 297854 550658
rect 297234 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 297854 550574
rect 297234 514894 297854 550338
rect 297234 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 297854 514894
rect 297234 514574 297854 514658
rect 297234 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 297854 514574
rect 297234 478894 297854 514338
rect 297234 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 297854 478894
rect 297234 478574 297854 478658
rect 297234 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 297854 478574
rect 297234 442894 297854 478338
rect 297234 442658 297266 442894
rect 297502 442658 297586 442894
rect 297822 442658 297854 442894
rect 297234 442574 297854 442658
rect 297234 442338 297266 442574
rect 297502 442338 297586 442574
rect 297822 442338 297854 442574
rect 297234 406894 297854 442338
rect 297234 406658 297266 406894
rect 297502 406658 297586 406894
rect 297822 406658 297854 406894
rect 297234 406574 297854 406658
rect 297234 406338 297266 406574
rect 297502 406338 297586 406574
rect 297822 406338 297854 406574
rect 297234 370894 297854 406338
rect 297234 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 297854 370894
rect 297234 370574 297854 370658
rect 297234 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 297854 370574
rect 297234 334894 297854 370338
rect 297234 334658 297266 334894
rect 297502 334658 297586 334894
rect 297822 334658 297854 334894
rect 297234 334574 297854 334658
rect 297234 334338 297266 334574
rect 297502 334338 297586 334574
rect 297822 334338 297854 334574
rect 297234 298894 297854 334338
rect 297234 298658 297266 298894
rect 297502 298658 297586 298894
rect 297822 298658 297854 298894
rect 297234 298574 297854 298658
rect 297234 298338 297266 298574
rect 297502 298338 297586 298574
rect 297822 298338 297854 298574
rect 297234 262894 297854 298338
rect 297234 262658 297266 262894
rect 297502 262658 297586 262894
rect 297822 262658 297854 262894
rect 297234 262574 297854 262658
rect 297234 262338 297266 262574
rect 297502 262338 297586 262574
rect 297822 262338 297854 262574
rect 297234 226894 297854 262338
rect 297234 226658 297266 226894
rect 297502 226658 297586 226894
rect 297822 226658 297854 226894
rect 297234 226574 297854 226658
rect 297234 226338 297266 226574
rect 297502 226338 297586 226574
rect 297822 226338 297854 226574
rect 297234 202000 297854 226338
rect 300954 698614 301574 710042
rect 318954 711558 319574 711590
rect 318954 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 319574 711558
rect 318954 711238 319574 711322
rect 318954 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 319574 711238
rect 315234 709638 315854 709670
rect 315234 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 315854 709638
rect 315234 709318 315854 709402
rect 315234 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 315854 709318
rect 311514 707718 312134 707750
rect 311514 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 312134 707718
rect 311514 707398 312134 707482
rect 311514 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 312134 707398
rect 300954 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 301574 698614
rect 300954 698294 301574 698378
rect 300954 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 301574 698294
rect 300954 662614 301574 698058
rect 300954 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 301574 662614
rect 300954 662294 301574 662378
rect 300954 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 301574 662294
rect 300954 626614 301574 662058
rect 300954 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 301574 626614
rect 300954 626294 301574 626378
rect 300954 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 301574 626294
rect 300954 590614 301574 626058
rect 300954 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 301574 590614
rect 300954 590294 301574 590378
rect 300954 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 301574 590294
rect 300954 554614 301574 590058
rect 300954 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 301574 554614
rect 300954 554294 301574 554378
rect 300954 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 301574 554294
rect 300954 518614 301574 554058
rect 300954 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 301574 518614
rect 300954 518294 301574 518378
rect 300954 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 301574 518294
rect 300954 482614 301574 518058
rect 300954 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 301574 482614
rect 300954 482294 301574 482378
rect 300954 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 301574 482294
rect 300954 446614 301574 482058
rect 300954 446378 300986 446614
rect 301222 446378 301306 446614
rect 301542 446378 301574 446614
rect 300954 446294 301574 446378
rect 300954 446058 300986 446294
rect 301222 446058 301306 446294
rect 301542 446058 301574 446294
rect 300954 410614 301574 446058
rect 300954 410378 300986 410614
rect 301222 410378 301306 410614
rect 301542 410378 301574 410614
rect 300954 410294 301574 410378
rect 300954 410058 300986 410294
rect 301222 410058 301306 410294
rect 301542 410058 301574 410294
rect 300954 374614 301574 410058
rect 300954 374378 300986 374614
rect 301222 374378 301306 374614
rect 301542 374378 301574 374614
rect 300954 374294 301574 374378
rect 300954 374058 300986 374294
rect 301222 374058 301306 374294
rect 301542 374058 301574 374294
rect 300954 338614 301574 374058
rect 300954 338378 300986 338614
rect 301222 338378 301306 338614
rect 301542 338378 301574 338614
rect 300954 338294 301574 338378
rect 300954 338058 300986 338294
rect 301222 338058 301306 338294
rect 301542 338058 301574 338294
rect 300954 302614 301574 338058
rect 300954 302378 300986 302614
rect 301222 302378 301306 302614
rect 301542 302378 301574 302614
rect 300954 302294 301574 302378
rect 300954 302058 300986 302294
rect 301222 302058 301306 302294
rect 301542 302058 301574 302294
rect 300954 266614 301574 302058
rect 300954 266378 300986 266614
rect 301222 266378 301306 266614
rect 301542 266378 301574 266614
rect 300954 266294 301574 266378
rect 300954 266058 300986 266294
rect 301222 266058 301306 266294
rect 301542 266058 301574 266294
rect 300954 230614 301574 266058
rect 300954 230378 300986 230614
rect 301222 230378 301306 230614
rect 301542 230378 301574 230614
rect 300954 230294 301574 230378
rect 300954 230058 300986 230294
rect 301222 230058 301306 230294
rect 301542 230058 301574 230294
rect 300954 202000 301574 230058
rect 307794 705798 308414 705830
rect 307794 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 308414 705798
rect 307794 705478 308414 705562
rect 307794 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 308414 705478
rect 307794 669454 308414 705242
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 561454 308414 596898
rect 307794 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 308414 561454
rect 307794 561134 308414 561218
rect 307794 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 308414 561134
rect 307794 525454 308414 560898
rect 307794 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 308414 525454
rect 307794 525134 308414 525218
rect 307794 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 308414 525134
rect 307794 489454 308414 524898
rect 307794 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 308414 489454
rect 307794 489134 308414 489218
rect 307794 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 308414 489134
rect 307794 453454 308414 488898
rect 307794 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 308414 453454
rect 307794 453134 308414 453218
rect 307794 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 308414 453134
rect 307794 417454 308414 452898
rect 307794 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 308414 417454
rect 307794 417134 308414 417218
rect 307794 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 308414 417134
rect 307794 381454 308414 416898
rect 307794 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 308414 381454
rect 307794 381134 308414 381218
rect 307794 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 308414 381134
rect 307794 345454 308414 380898
rect 307794 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 308414 345454
rect 307794 345134 308414 345218
rect 307794 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 308414 345134
rect 307794 309454 308414 344898
rect 307794 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 308414 309454
rect 307794 309134 308414 309218
rect 307794 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 308414 309134
rect 307794 273454 308414 308898
rect 307794 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 308414 273454
rect 307794 273134 308414 273218
rect 307794 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 308414 273134
rect 307794 237454 308414 272898
rect 307794 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 308414 237454
rect 307794 237134 308414 237218
rect 307794 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 308414 237134
rect 192954 194378 192986 194614
rect 193222 194378 193306 194614
rect 193542 194378 193574 194614
rect 192954 194294 193574 194378
rect 192954 194058 192986 194294
rect 193222 194058 193306 194294
rect 193542 194058 193574 194294
rect 192954 158614 193574 194058
rect 307794 201454 308414 236898
rect 307794 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 308414 201454
rect 307794 201134 308414 201218
rect 307794 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 308414 201134
rect 204208 183454 204528 183486
rect 204208 183218 204250 183454
rect 204486 183218 204528 183454
rect 204208 183134 204528 183218
rect 204208 182898 204250 183134
rect 204486 182898 204528 183134
rect 204208 182866 204528 182898
rect 234928 183454 235248 183486
rect 234928 183218 234970 183454
rect 235206 183218 235248 183454
rect 234928 183134 235248 183218
rect 234928 182898 234970 183134
rect 235206 182898 235248 183134
rect 234928 182866 235248 182898
rect 265648 183454 265968 183486
rect 265648 183218 265690 183454
rect 265926 183218 265968 183454
rect 265648 183134 265968 183218
rect 265648 182898 265690 183134
rect 265926 182898 265968 183134
rect 265648 182866 265968 182898
rect 296368 183454 296688 183486
rect 296368 183218 296410 183454
rect 296646 183218 296688 183454
rect 296368 183134 296688 183218
rect 296368 182898 296410 183134
rect 296646 182898 296688 183134
rect 296368 182866 296688 182898
rect 219568 165454 219888 165486
rect 219568 165218 219610 165454
rect 219846 165218 219888 165454
rect 219568 165134 219888 165218
rect 219568 164898 219610 165134
rect 219846 164898 219888 165134
rect 219568 164866 219888 164898
rect 250288 165454 250608 165486
rect 250288 165218 250330 165454
rect 250566 165218 250608 165454
rect 250288 165134 250608 165218
rect 250288 164898 250330 165134
rect 250566 164898 250608 165134
rect 250288 164866 250608 164898
rect 281008 165454 281328 165486
rect 281008 165218 281050 165454
rect 281286 165218 281328 165454
rect 281008 165134 281328 165218
rect 281008 164898 281050 165134
rect 281286 164898 281328 165134
rect 281008 164866 281328 164898
rect 307794 165454 308414 200898
rect 307794 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 308414 165454
rect 307794 165134 308414 165218
rect 307794 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 308414 165134
rect 192954 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 193574 158614
rect 192954 158294 193574 158378
rect 192954 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 193574 158294
rect 192954 122614 193574 158058
rect 204208 147454 204528 147486
rect 204208 147218 204250 147454
rect 204486 147218 204528 147454
rect 204208 147134 204528 147218
rect 204208 146898 204250 147134
rect 204486 146898 204528 147134
rect 204208 146866 204528 146898
rect 234928 147454 235248 147486
rect 234928 147218 234970 147454
rect 235206 147218 235248 147454
rect 234928 147134 235248 147218
rect 234928 146898 234970 147134
rect 235206 146898 235248 147134
rect 234928 146866 235248 146898
rect 265648 147454 265968 147486
rect 265648 147218 265690 147454
rect 265926 147218 265968 147454
rect 265648 147134 265968 147218
rect 265648 146898 265690 147134
rect 265926 146898 265968 147134
rect 265648 146866 265968 146898
rect 296368 147454 296688 147486
rect 296368 147218 296410 147454
rect 296646 147218 296688 147454
rect 296368 147134 296688 147218
rect 296368 146898 296410 147134
rect 296646 146898 296688 147134
rect 296368 146866 296688 146898
rect 219568 129454 219888 129486
rect 219568 129218 219610 129454
rect 219846 129218 219888 129454
rect 219568 129134 219888 129218
rect 219568 128898 219610 129134
rect 219846 128898 219888 129134
rect 219568 128866 219888 128898
rect 250288 129454 250608 129486
rect 250288 129218 250330 129454
rect 250566 129218 250608 129454
rect 250288 129134 250608 129218
rect 250288 128898 250330 129134
rect 250566 128898 250608 129134
rect 250288 128866 250608 128898
rect 281008 129454 281328 129486
rect 281008 129218 281050 129454
rect 281286 129218 281328 129454
rect 281008 129134 281328 129218
rect 281008 128898 281050 129134
rect 281286 128898 281328 129134
rect 281008 128866 281328 128898
rect 307794 129454 308414 164898
rect 307794 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 308414 129454
rect 307794 129134 308414 129218
rect 307794 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 308414 129134
rect 192954 122378 192986 122614
rect 193222 122378 193306 122614
rect 193542 122378 193574 122614
rect 192954 122294 193574 122378
rect 192954 122058 192986 122294
rect 193222 122058 193306 122294
rect 193542 122058 193574 122294
rect 192954 86614 193574 122058
rect 204208 111454 204528 111486
rect 204208 111218 204250 111454
rect 204486 111218 204528 111454
rect 204208 111134 204528 111218
rect 204208 110898 204250 111134
rect 204486 110898 204528 111134
rect 204208 110866 204528 110898
rect 234928 111454 235248 111486
rect 234928 111218 234970 111454
rect 235206 111218 235248 111454
rect 234928 111134 235248 111218
rect 234928 110898 234970 111134
rect 235206 110898 235248 111134
rect 234928 110866 235248 110898
rect 265648 111454 265968 111486
rect 265648 111218 265690 111454
rect 265926 111218 265968 111454
rect 265648 111134 265968 111218
rect 265648 110898 265690 111134
rect 265926 110898 265968 111134
rect 265648 110866 265968 110898
rect 296368 111454 296688 111486
rect 296368 111218 296410 111454
rect 296646 111218 296688 111454
rect 296368 111134 296688 111218
rect 296368 110898 296410 111134
rect 296646 110898 296688 111134
rect 296368 110866 296688 110898
rect 297958 102310 298202 102370
rect 297958 100333 298018 102310
rect 298142 102237 298202 102310
rect 298139 102236 298205 102237
rect 298139 102172 298140 102236
rect 298204 102172 298205 102236
rect 298139 102171 298205 102172
rect 297955 100332 298021 100333
rect 297955 100268 297956 100332
rect 298020 100268 298021 100332
rect 297955 100267 298021 100268
rect 192954 86378 192986 86614
rect 193222 86378 193306 86614
rect 193542 86378 193574 86614
rect 192954 86294 193574 86378
rect 192954 86058 192986 86294
rect 193222 86058 193306 86294
rect 193542 86058 193574 86294
rect 192954 50614 193574 86058
rect 192954 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 193574 50614
rect 192954 50294 193574 50378
rect 192954 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 193574 50294
rect 192954 14614 193574 50058
rect 192954 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 193574 14614
rect 192954 14294 193574 14378
rect 192954 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 193574 14294
rect 174954 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 175574 -7066
rect 174954 -7386 175574 -7302
rect 174954 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 175574 -7386
rect 174954 -7654 175574 -7622
rect 192954 -6106 193574 14058
rect 199794 93454 200414 98000
rect 203514 97174 204134 98000
rect 203514 96938 203546 97174
rect 203782 96938 203866 97174
rect 204102 96938 204134 97174
rect 202827 96932 202893 96933
rect 202827 96868 202828 96932
rect 202892 96868 202893 96932
rect 202827 96867 202893 96868
rect 199794 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 200414 93454
rect 199794 93134 200414 93218
rect 199794 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 200414 93134
rect 199794 57454 200414 92898
rect 202830 91765 202890 96867
rect 203514 96854 204134 96938
rect 205955 96932 206021 96933
rect 205955 96868 205956 96932
rect 206020 96868 206021 96932
rect 205955 96867 206021 96868
rect 203514 96618 203546 96854
rect 203782 96618 203866 96854
rect 204102 96618 204134 96854
rect 202827 91764 202893 91765
rect 202827 91700 202828 91764
rect 202892 91700 202893 91764
rect 202827 91699 202893 91700
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 21454 200414 56898
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -1306 200414 20898
rect 199794 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 200414 -1306
rect 199794 -1626 200414 -1542
rect 199794 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 200414 -1626
rect 199794 -1894 200414 -1862
rect 203514 61174 204134 96618
rect 204299 96660 204365 96661
rect 204299 96596 204300 96660
rect 204364 96596 204365 96660
rect 204299 96595 204365 96596
rect 205771 96660 205837 96661
rect 205771 96596 205772 96660
rect 205836 96596 205837 96660
rect 205771 96595 205837 96596
rect 204302 93125 204362 96595
rect 205774 93261 205834 96595
rect 205771 93260 205837 93261
rect 205771 93196 205772 93260
rect 205836 93196 205837 93260
rect 205771 93195 205837 93196
rect 204299 93124 204365 93125
rect 204299 93060 204300 93124
rect 204364 93060 204365 93124
rect 204299 93059 204365 93060
rect 205958 89730 206018 96867
rect 205590 89670 206018 89730
rect 205590 73813 205650 89670
rect 205587 73812 205653 73813
rect 205587 73748 205588 73812
rect 205652 73748 205653 73812
rect 205587 73747 205653 73748
rect 203514 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 204134 61174
rect 203514 60854 204134 60938
rect 203514 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 204134 60854
rect 203514 25174 204134 60618
rect 203514 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 204134 25174
rect 203514 24854 204134 24938
rect 203514 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 204134 24854
rect 203514 -3226 204134 24618
rect 203514 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 204134 -3226
rect 203514 -3546 204134 -3462
rect 203514 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 204134 -3546
rect 203514 -3814 204134 -3782
rect 207234 64894 207854 98000
rect 208347 96660 208413 96661
rect 208347 96596 208348 96660
rect 208412 96596 208413 96660
rect 208347 96595 208413 96596
rect 209819 96660 209885 96661
rect 209819 96596 209820 96660
rect 209884 96596 209885 96660
rect 209819 96595 209885 96596
rect 208350 80749 208410 96595
rect 209822 84829 209882 96595
rect 209819 84828 209885 84829
rect 209819 84764 209820 84828
rect 209884 84764 209885 84828
rect 209819 84763 209885 84764
rect 208347 80748 208413 80749
rect 208347 80684 208348 80748
rect 208412 80684 208413 80748
rect 208347 80683 208413 80684
rect 207234 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 207854 64894
rect 207234 64574 207854 64658
rect 207234 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 207854 64574
rect 207234 28894 207854 64338
rect 207234 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 207854 28894
rect 207234 28574 207854 28658
rect 207234 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 207854 28574
rect 207234 -5146 207854 28338
rect 207234 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 207854 -5146
rect 207234 -5466 207854 -5382
rect 207234 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 207854 -5466
rect 207234 -5734 207854 -5702
rect 210954 68614 211574 98000
rect 215339 96932 215405 96933
rect 215339 96868 215340 96932
rect 215404 96868 215405 96932
rect 215339 96867 215405 96868
rect 216627 96932 216693 96933
rect 216627 96868 216628 96932
rect 216692 96868 216693 96932
rect 216627 96867 216693 96868
rect 211659 96660 211725 96661
rect 211659 96596 211660 96660
rect 211724 96596 211725 96660
rect 211659 96595 211725 96596
rect 212579 96660 212645 96661
rect 212579 96596 212580 96660
rect 212644 96596 212645 96660
rect 212579 96595 212645 96596
rect 213867 96660 213933 96661
rect 213867 96596 213868 96660
rect 213932 96596 213933 96660
rect 213867 96595 213933 96596
rect 211662 79389 211722 96595
rect 212582 87685 212642 96595
rect 212579 87684 212645 87685
rect 212579 87620 212580 87684
rect 212644 87620 212645 87684
rect 212579 87619 212645 87620
rect 213870 84965 213930 96595
rect 213867 84964 213933 84965
rect 213867 84900 213868 84964
rect 213932 84900 213933 84964
rect 213867 84899 213933 84900
rect 211659 79388 211725 79389
rect 211659 79324 211660 79388
rect 211724 79324 211725 79388
rect 211659 79323 211725 79324
rect 215342 73949 215402 96867
rect 216630 89181 216690 96867
rect 216627 89180 216693 89181
rect 216627 89116 216628 89180
rect 216692 89116 216693 89180
rect 216627 89115 216693 89116
rect 217794 75454 218414 98000
rect 219387 97612 219453 97613
rect 219387 97610 219388 97612
rect 219206 97550 219388 97610
rect 218651 96932 218717 96933
rect 218651 96868 218652 96932
rect 218716 96868 218717 96932
rect 218651 96867 218717 96868
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 215339 73948 215405 73949
rect 215339 73884 215340 73948
rect 215404 73884 215405 73948
rect 215339 73883 215405 73884
rect 210954 68378 210986 68614
rect 211222 68378 211306 68614
rect 211542 68378 211574 68614
rect 210954 68294 211574 68378
rect 210954 68058 210986 68294
rect 211222 68058 211306 68294
rect 211542 68058 211574 68294
rect 210954 32614 211574 68058
rect 210954 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 211574 32614
rect 210954 32294 211574 32378
rect 210954 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 211574 32294
rect 192954 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 193574 -6106
rect 192954 -6426 193574 -6342
rect 192954 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 193574 -6426
rect 192954 -7654 193574 -6662
rect 210954 -7066 211574 32058
rect 217794 39454 218414 74898
rect 218654 44845 218714 96867
rect 219206 77893 219266 97550
rect 219387 97548 219388 97550
rect 219452 97548 219453 97612
rect 219387 97547 219453 97548
rect 220859 96932 220925 96933
rect 220859 96868 220860 96932
rect 220924 96868 220925 96932
rect 220859 96867 220925 96868
rect 220862 79525 220922 96867
rect 220859 79524 220925 79525
rect 220859 79460 220860 79524
rect 220924 79460 220925 79524
rect 220859 79459 220925 79460
rect 221514 79174 222134 98000
rect 222331 96932 222397 96933
rect 222331 96868 222332 96932
rect 222396 96868 222397 96932
rect 222331 96867 222397 96868
rect 223619 96932 223685 96933
rect 223619 96868 223620 96932
rect 223684 96868 223685 96932
rect 223619 96867 223685 96868
rect 222334 83469 222394 96867
rect 223622 93397 223682 96867
rect 223619 93396 223685 93397
rect 223619 93332 223620 93396
rect 223684 93332 223685 93396
rect 223619 93331 223685 93332
rect 222331 83468 222397 83469
rect 222331 83404 222332 83468
rect 222396 83404 222397 83468
rect 222331 83403 222397 83404
rect 221514 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 222134 79174
rect 221514 78854 222134 78938
rect 221514 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 222134 78854
rect 219203 77892 219269 77893
rect 219203 77828 219204 77892
rect 219268 77828 219269 77892
rect 219203 77827 219269 77828
rect 218651 44844 218717 44845
rect 218651 44780 218652 44844
rect 218716 44780 218717 44844
rect 218651 44779 218717 44780
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -1894 218414 -902
rect 221514 43174 222134 78618
rect 221514 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 222134 43174
rect 221514 42854 222134 42938
rect 221514 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 222134 42854
rect 221514 7174 222134 42618
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -2266 222134 6618
rect 221514 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 222134 -2266
rect 221514 -2586 222134 -2502
rect 221514 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 222134 -2586
rect 221514 -3814 222134 -2822
rect 225234 82894 225854 98000
rect 226379 96660 226445 96661
rect 226379 96596 226380 96660
rect 226444 96596 226445 96660
rect 226379 96595 226445 96596
rect 226382 94485 226442 96595
rect 226379 94484 226445 94485
rect 226379 94420 226380 94484
rect 226444 94420 226445 94484
rect 226379 94419 226445 94420
rect 225234 82658 225266 82894
rect 225502 82658 225586 82894
rect 225822 82658 225854 82894
rect 225234 82574 225854 82658
rect 225234 82338 225266 82574
rect 225502 82338 225586 82574
rect 225822 82338 225854 82574
rect 225234 46894 225854 82338
rect 225234 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 225854 46894
rect 225234 46574 225854 46658
rect 225234 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 225854 46574
rect 225234 10894 225854 46338
rect 225234 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 225854 10894
rect 225234 10574 225854 10658
rect 225234 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 225854 10574
rect 225234 -4186 225854 10338
rect 225234 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 225854 -4186
rect 225234 -4506 225854 -4422
rect 225234 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 225854 -4506
rect 225234 -5734 225854 -4742
rect 228954 86614 229574 98000
rect 230611 96796 230677 96797
rect 230611 96732 230612 96796
rect 230676 96732 230677 96796
rect 230611 96731 230677 96732
rect 230427 96660 230493 96661
rect 230427 96596 230428 96660
rect 230492 96596 230493 96660
rect 230427 96595 230493 96596
rect 230430 94757 230490 96595
rect 230427 94756 230493 94757
rect 230427 94692 230428 94756
rect 230492 94692 230493 94756
rect 230427 94691 230493 94692
rect 230614 91901 230674 96731
rect 231899 96660 231965 96661
rect 231899 96596 231900 96660
rect 231964 96596 231965 96660
rect 231899 96595 231965 96596
rect 233187 96660 233253 96661
rect 233187 96596 233188 96660
rect 233252 96596 233253 96660
rect 233187 96595 233253 96596
rect 230611 91900 230677 91901
rect 230611 91836 230612 91900
rect 230676 91836 230677 91900
rect 230611 91835 230677 91836
rect 228954 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 229574 86614
rect 228954 86294 229574 86378
rect 228954 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 229574 86294
rect 231902 86189 231962 96595
rect 233190 90405 233250 96595
rect 235794 93454 236414 98000
rect 239514 97174 240134 98000
rect 239514 96938 239546 97174
rect 239782 96938 239866 97174
rect 240102 96938 240134 97174
rect 237603 96932 237669 96933
rect 237603 96868 237604 96932
rect 237668 96868 237669 96932
rect 237603 96867 237669 96868
rect 235794 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 236414 93454
rect 235794 93134 236414 93218
rect 235794 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 236414 93134
rect 233187 90404 233253 90405
rect 233187 90340 233188 90404
rect 233252 90340 233253 90404
rect 233187 90339 233253 90340
rect 231899 86188 231965 86189
rect 231899 86124 231900 86188
rect 231964 86124 231965 86188
rect 231899 86123 231965 86124
rect 228954 50614 229574 86058
rect 228954 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 229574 50614
rect 228954 50294 229574 50378
rect 228954 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 229574 50294
rect 228954 14614 229574 50058
rect 228954 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 229574 14614
rect 228954 14294 229574 14378
rect 228954 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 229574 14294
rect 210954 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 211574 -7066
rect 210954 -7386 211574 -7302
rect 210954 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 211574 -7386
rect 210954 -7654 211574 -7622
rect 228954 -6106 229574 14058
rect 235794 57454 236414 92898
rect 237606 81565 237666 96867
rect 239514 96854 240134 96938
rect 239514 96618 239546 96854
rect 239782 96618 239866 96854
rect 240102 96618 240134 96854
rect 237603 81564 237669 81565
rect 237603 81500 237604 81564
rect 237668 81500 237669 81564
rect 237603 81499 237669 81500
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -1306 236414 20898
rect 235794 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 236414 -1306
rect 235794 -1626 236414 -1542
rect 235794 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 236414 -1626
rect 235794 -1894 236414 -1862
rect 239514 61174 240134 96618
rect 239514 60938 239546 61174
rect 239782 60938 239866 61174
rect 240102 60938 240134 61174
rect 239514 60854 240134 60938
rect 239514 60618 239546 60854
rect 239782 60618 239866 60854
rect 240102 60618 240134 60854
rect 239514 25174 240134 60618
rect 239514 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 240134 25174
rect 239514 24854 240134 24938
rect 239514 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 240134 24854
rect 239514 -3226 240134 24618
rect 239514 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 240134 -3226
rect 239514 -3546 240134 -3462
rect 239514 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 240134 -3546
rect 239514 -3814 240134 -3782
rect 243234 64894 243854 98000
rect 246803 96932 246869 96933
rect 246803 96868 246804 96932
rect 246868 96868 246869 96932
rect 246803 96867 246869 96868
rect 243234 64658 243266 64894
rect 243502 64658 243586 64894
rect 243822 64658 243854 64894
rect 243234 64574 243854 64658
rect 243234 64338 243266 64574
rect 243502 64338 243586 64574
rect 243822 64338 243854 64574
rect 243234 28894 243854 64338
rect 243234 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 243854 28894
rect 243234 28574 243854 28658
rect 243234 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 243854 28574
rect 243234 -5146 243854 28338
rect 246806 6221 246866 96867
rect 246954 68614 247574 98000
rect 252507 97068 252573 97069
rect 252507 97004 252508 97068
rect 252572 97004 252573 97068
rect 252507 97003 252573 97004
rect 249563 96932 249629 96933
rect 249563 96868 249564 96932
rect 249628 96868 249629 96932
rect 249563 96867 249629 96868
rect 250851 96932 250917 96933
rect 250851 96868 250852 96932
rect 250916 96868 250917 96932
rect 250851 96867 250917 96868
rect 252323 96932 252389 96933
rect 252323 96868 252324 96932
rect 252388 96868 252389 96932
rect 252323 96867 252389 96868
rect 246954 68378 246986 68614
rect 247222 68378 247306 68614
rect 247542 68378 247574 68614
rect 246954 68294 247574 68378
rect 246954 68058 246986 68294
rect 247222 68058 247306 68294
rect 247542 68058 247574 68294
rect 246954 32614 247574 68058
rect 249566 62797 249626 96867
rect 250854 80749 250914 96867
rect 250851 80748 250917 80749
rect 250851 80684 250852 80748
rect 250916 80684 250917 80748
rect 250851 80683 250917 80684
rect 249563 62796 249629 62797
rect 249563 62732 249564 62796
rect 249628 62732 249629 62796
rect 249563 62731 249629 62732
rect 246954 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 247574 32614
rect 246954 32294 247574 32378
rect 246954 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 247574 32294
rect 246803 6220 246869 6221
rect 246803 6156 246804 6220
rect 246868 6156 246869 6220
rect 246803 6155 246869 6156
rect 243234 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 243854 -5146
rect 243234 -5466 243854 -5382
rect 243234 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 243854 -5466
rect 243234 -5734 243854 -5702
rect 228954 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 229574 -6106
rect 228954 -6426 229574 -6342
rect 228954 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 229574 -6426
rect 228954 -7654 229574 -6662
rect 246954 -7066 247574 32058
rect 252326 2005 252386 96867
rect 252510 94621 252570 97003
rect 253611 96932 253677 96933
rect 253611 96868 253612 96932
rect 253676 96868 253677 96932
rect 253611 96867 253677 96868
rect 252507 94620 252573 94621
rect 252507 94556 252508 94620
rect 252572 94556 252573 94620
rect 252507 94555 252573 94556
rect 253614 82109 253674 96867
rect 253611 82108 253677 82109
rect 253611 82044 253612 82108
rect 253676 82044 253677 82108
rect 253611 82043 253677 82044
rect 253794 75454 254414 98000
rect 255083 96932 255149 96933
rect 255083 96868 255084 96932
rect 255148 96868 255149 96932
rect 255083 96867 255149 96868
rect 256555 96932 256621 96933
rect 256555 96868 256556 96932
rect 256620 96868 256621 96932
rect 256555 96867 256621 96868
rect 257291 96932 257357 96933
rect 257291 96868 257292 96932
rect 257356 96868 257357 96932
rect 257291 96867 257357 96868
rect 255086 76805 255146 96867
rect 255083 76804 255149 76805
rect 255083 76740 255084 76804
rect 255148 76740 255149 76804
rect 255083 76739 255149 76740
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253794 39454 254414 74898
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 256558 11933 256618 96867
rect 257294 73813 257354 96867
rect 257514 79174 258134 98000
rect 259315 97068 259381 97069
rect 259315 97004 259316 97068
rect 259380 97004 259381 97068
rect 259315 97003 259381 97004
rect 260603 97068 260669 97069
rect 260603 97004 260604 97068
rect 260668 97004 260669 97068
rect 260603 97003 260669 97004
rect 259131 96932 259197 96933
rect 259131 96868 259132 96932
rect 259196 96868 259197 96932
rect 259131 96867 259197 96868
rect 259134 84965 259194 96867
rect 259131 84964 259197 84965
rect 259131 84900 259132 84964
rect 259196 84900 259197 84964
rect 259131 84899 259197 84900
rect 259318 79661 259378 97003
rect 260419 96932 260485 96933
rect 260419 96868 260420 96932
rect 260484 96868 260485 96932
rect 260419 96867 260485 96868
rect 260422 93397 260482 96867
rect 260419 93396 260485 93397
rect 260419 93332 260420 93396
rect 260484 93332 260485 93396
rect 260419 93331 260485 93332
rect 259315 79660 259381 79661
rect 259315 79596 259316 79660
rect 259380 79596 259381 79660
rect 259315 79595 259381 79596
rect 257514 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 258134 79174
rect 257514 78854 258134 78938
rect 257514 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 258134 78854
rect 257291 73812 257357 73813
rect 257291 73748 257292 73812
rect 257356 73748 257357 73812
rect 257291 73747 257357 73748
rect 257514 43174 258134 78618
rect 260606 72453 260666 97003
rect 261234 82894 261854 98000
rect 264467 97068 264533 97069
rect 264467 97004 264468 97068
rect 264532 97004 264533 97068
rect 264467 97003 264533 97004
rect 263179 96932 263245 96933
rect 263179 96868 263180 96932
rect 263244 96868 263245 96932
rect 263179 96867 263245 96868
rect 263363 96932 263429 96933
rect 263363 96868 263364 96932
rect 263428 96868 263429 96932
rect 263363 96867 263429 96868
rect 261234 82658 261266 82894
rect 261502 82658 261586 82894
rect 261822 82658 261854 82894
rect 261234 82574 261854 82658
rect 261234 82338 261266 82574
rect 261502 82338 261586 82574
rect 261822 82338 261854 82574
rect 260603 72452 260669 72453
rect 260603 72388 260604 72452
rect 260668 72388 260669 72452
rect 260603 72387 260669 72388
rect 257514 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 258134 43174
rect 257514 42854 258134 42938
rect 257514 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 258134 42854
rect 256555 11932 256621 11933
rect 256555 11868 256556 11932
rect 256620 11868 256621 11932
rect 256555 11867 256621 11868
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 252323 2004 252389 2005
rect 252323 1940 252324 2004
rect 252388 1940 252389 2004
rect 252323 1939 252389 1940
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -1894 254414 -902
rect 257514 7174 258134 42618
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 257514 -2266 258134 6618
rect 257514 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 258134 -2266
rect 257514 -2586 258134 -2502
rect 257514 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 258134 -2586
rect 257514 -3814 258134 -2822
rect 261234 46894 261854 82338
rect 263182 79525 263242 96867
rect 263179 79524 263245 79525
rect 263179 79460 263180 79524
rect 263244 79460 263245 79524
rect 263179 79459 263245 79460
rect 261234 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 261854 46894
rect 261234 46574 261854 46658
rect 261234 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 261854 46574
rect 261234 10894 261854 46338
rect 263366 30973 263426 96867
rect 264470 91765 264530 97003
rect 264651 96932 264717 96933
rect 264651 96868 264652 96932
rect 264716 96868 264717 96932
rect 264651 96867 264717 96868
rect 264467 91764 264533 91765
rect 264467 91700 264468 91764
rect 264532 91700 264533 91764
rect 264467 91699 264533 91700
rect 264654 71229 264714 96867
rect 264954 86614 265574 98000
rect 271459 97204 271525 97205
rect 271459 97140 271460 97204
rect 271524 97140 271525 97204
rect 271459 97139 271525 97140
rect 267411 97068 267477 97069
rect 267411 97004 267412 97068
rect 267476 97004 267477 97068
rect 267411 97003 267477 97004
rect 266123 96932 266189 96933
rect 266123 96868 266124 96932
rect 266188 96868 266189 96932
rect 266123 96867 266189 96868
rect 264954 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 265574 86614
rect 264954 86294 265574 86378
rect 264954 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 265574 86294
rect 264651 71228 264717 71229
rect 264651 71164 264652 71228
rect 264716 71164 264717 71228
rect 264651 71163 264717 71164
rect 264954 50614 265574 86058
rect 266126 75309 266186 96867
rect 267414 84829 267474 97003
rect 267595 96932 267661 96933
rect 267595 96868 267596 96932
rect 267660 96868 267661 96932
rect 267595 96867 267661 96868
rect 268883 96932 268949 96933
rect 268883 96868 268884 96932
rect 268948 96868 268949 96932
rect 268883 96867 268949 96868
rect 270355 96932 270421 96933
rect 270355 96868 270356 96932
rect 270420 96868 270421 96932
rect 270355 96867 270421 96868
rect 267411 84828 267477 84829
rect 267411 84764 267412 84828
rect 267476 84764 267477 84828
rect 267411 84763 267477 84764
rect 267598 78165 267658 96867
rect 267595 78164 267661 78165
rect 267595 78100 267596 78164
rect 267660 78100 267661 78164
rect 267595 78099 267661 78100
rect 268886 76669 268946 96867
rect 268883 76668 268949 76669
rect 268883 76604 268884 76668
rect 268948 76604 268949 76668
rect 268883 76603 268949 76604
rect 270358 76533 270418 96867
rect 271462 95845 271522 97139
rect 271643 96932 271709 96933
rect 271643 96868 271644 96932
rect 271708 96868 271709 96932
rect 271643 96867 271709 96868
rect 271459 95844 271525 95845
rect 271459 95780 271460 95844
rect 271524 95780 271525 95844
rect 271459 95779 271525 95780
rect 271646 78029 271706 96867
rect 271794 93454 272414 98000
rect 275514 97174 276134 98000
rect 273115 97068 273181 97069
rect 273115 97004 273116 97068
rect 273180 97004 273181 97068
rect 273115 97003 273181 97004
rect 274219 97068 274285 97069
rect 274219 97004 274220 97068
rect 274284 97004 274285 97068
rect 274219 97003 274285 97004
rect 275323 97068 275389 97069
rect 275323 97004 275324 97068
rect 275388 97004 275389 97068
rect 275323 97003 275389 97004
rect 271794 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 272414 93454
rect 271794 93134 272414 93218
rect 271794 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 272414 93134
rect 271643 78028 271709 78029
rect 271643 77964 271644 78028
rect 271708 77964 271709 78028
rect 271643 77963 271709 77964
rect 270355 76532 270421 76533
rect 270355 76468 270356 76532
rect 270420 76468 270421 76532
rect 270355 76467 270421 76468
rect 266123 75308 266189 75309
rect 266123 75244 266124 75308
rect 266188 75244 266189 75308
rect 266123 75243 266189 75244
rect 264954 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 265574 50614
rect 264954 50294 265574 50378
rect 264954 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 265574 50294
rect 263363 30972 263429 30973
rect 263363 30908 263364 30972
rect 263428 30908 263429 30972
rect 263363 30907 263429 30908
rect 261234 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 261854 10894
rect 261234 10574 261854 10658
rect 261234 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 261854 10574
rect 261234 -4186 261854 10338
rect 261234 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 261854 -4186
rect 261234 -4506 261854 -4422
rect 261234 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 261854 -4506
rect 261234 -5734 261854 -4742
rect 264954 14614 265574 50058
rect 264954 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 265574 14614
rect 264954 14294 265574 14378
rect 264954 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 265574 14294
rect 246954 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 247574 -7066
rect 246954 -7386 247574 -7302
rect 246954 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 247574 -7386
rect 246954 -7654 247574 -7622
rect 264954 -6106 265574 14058
rect 271794 57454 272414 92898
rect 273118 83605 273178 97003
rect 274222 90541 274282 97003
rect 274403 96932 274469 96933
rect 274403 96868 274404 96932
rect 274468 96868 274469 96932
rect 274403 96867 274469 96868
rect 274219 90540 274285 90541
rect 274219 90476 274220 90540
rect 274284 90476 274285 90540
rect 274219 90475 274285 90476
rect 273115 83604 273181 83605
rect 273115 83540 273116 83604
rect 273180 83540 273181 83604
rect 273115 83539 273181 83540
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -1306 272414 20898
rect 274406 11797 274466 96867
rect 275326 83469 275386 97003
rect 275514 96938 275546 97174
rect 275782 96938 275866 97174
rect 276102 96938 276134 97174
rect 279003 97068 279069 97069
rect 279003 97004 279004 97068
rect 279068 97004 279069 97068
rect 279003 97003 279069 97004
rect 275514 96854 276134 96938
rect 277163 96932 277229 96933
rect 277163 96868 277164 96932
rect 277228 96868 277229 96932
rect 277163 96867 277229 96868
rect 278635 96932 278701 96933
rect 278635 96868 278636 96932
rect 278700 96868 278701 96932
rect 278635 96867 278701 96868
rect 275514 96618 275546 96854
rect 275782 96618 275866 96854
rect 276102 96618 276134 96854
rect 275323 83468 275389 83469
rect 275323 83404 275324 83468
rect 275388 83404 275389 83468
rect 275323 83403 275389 83404
rect 275514 61174 276134 96618
rect 277166 77893 277226 96867
rect 278638 79389 278698 96867
rect 279006 89181 279066 97003
rect 279003 89180 279069 89181
rect 279003 89116 279004 89180
rect 279068 89116 279069 89180
rect 279003 89115 279069 89116
rect 278635 79388 278701 79389
rect 278635 79324 278636 79388
rect 278700 79324 278701 79388
rect 278635 79323 278701 79324
rect 277163 77892 277229 77893
rect 277163 77828 277164 77892
rect 277228 77828 277229 77892
rect 277163 77827 277229 77828
rect 275514 60938 275546 61174
rect 275782 60938 275866 61174
rect 276102 60938 276134 61174
rect 275514 60854 276134 60938
rect 275514 60618 275546 60854
rect 275782 60618 275866 60854
rect 276102 60618 276134 60854
rect 275514 25174 276134 60618
rect 275514 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 276134 25174
rect 275514 24854 276134 24938
rect 275514 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 276134 24854
rect 274403 11796 274469 11797
rect 274403 11732 274404 11796
rect 274468 11732 274469 11796
rect 274403 11731 274469 11732
rect 271794 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 272414 -1306
rect 271794 -1626 272414 -1542
rect 271794 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 272414 -1626
rect 271794 -1894 272414 -1862
rect 275514 -3226 276134 24618
rect 275514 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 276134 -3226
rect 275514 -3546 276134 -3462
rect 275514 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 276134 -3546
rect 275514 -3814 276134 -3782
rect 279234 64894 279854 98000
rect 281211 96932 281277 96933
rect 281211 96868 281212 96932
rect 281276 96868 281277 96932
rect 281211 96867 281277 96868
rect 281395 96932 281461 96933
rect 281395 96868 281396 96932
rect 281460 96868 281461 96932
rect 281395 96867 281461 96868
rect 282131 96932 282197 96933
rect 282131 96868 282132 96932
rect 282196 96868 282197 96932
rect 282131 96867 282197 96868
rect 281214 86325 281274 96867
rect 281211 86324 281277 86325
rect 281211 86260 281212 86324
rect 281276 86260 281277 86324
rect 281211 86259 281277 86260
rect 279234 64658 279266 64894
rect 279502 64658 279586 64894
rect 279822 64658 279854 64894
rect 279234 64574 279854 64658
rect 279234 64338 279266 64574
rect 279502 64338 279586 64574
rect 279822 64338 279854 64574
rect 279234 28894 279854 64338
rect 279234 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 279854 28894
rect 279234 28574 279854 28658
rect 279234 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 279854 28574
rect 279234 -5146 279854 28338
rect 281398 4861 281458 96867
rect 282134 91221 282194 96867
rect 282131 91220 282197 91221
rect 282131 91156 282132 91220
rect 282196 91156 282197 91220
rect 282131 91155 282197 91156
rect 282954 68614 283574 98000
rect 284155 96932 284221 96933
rect 284155 96868 284156 96932
rect 284220 96868 284221 96932
rect 284155 96867 284221 96868
rect 286915 96932 286981 96933
rect 286915 96868 286916 96932
rect 286980 96868 286981 96932
rect 286915 96867 286981 96868
rect 288203 96932 288269 96933
rect 288203 96868 288204 96932
rect 288268 96868 288269 96932
rect 288203 96867 288269 96868
rect 284158 93261 284218 96867
rect 284155 93260 284221 93261
rect 284155 93196 284156 93260
rect 284220 93196 284221 93260
rect 284155 93195 284221 93196
rect 286918 75173 286978 96867
rect 286915 75172 286981 75173
rect 286915 75108 286916 75172
rect 286980 75108 286981 75172
rect 286915 75107 286981 75108
rect 288206 71093 288266 96867
rect 289794 75454 290414 98000
rect 292435 97340 292501 97341
rect 292435 97276 292436 97340
rect 292500 97276 292501 97340
rect 292435 97275 292501 97276
rect 292251 96932 292317 96933
rect 292251 96868 292252 96932
rect 292316 96868 292317 96932
rect 292251 96867 292317 96868
rect 292254 87821 292314 96867
rect 292251 87820 292317 87821
rect 292251 87756 292252 87820
rect 292316 87756 292317 87820
rect 292251 87755 292317 87756
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 288203 71092 288269 71093
rect 288203 71028 288204 71092
rect 288268 71028 288269 71092
rect 288203 71027 288269 71028
rect 282954 68378 282986 68614
rect 283222 68378 283306 68614
rect 283542 68378 283574 68614
rect 282954 68294 283574 68378
rect 282954 68058 282986 68294
rect 283222 68058 283306 68294
rect 283542 68058 283574 68294
rect 282954 32614 283574 68058
rect 282954 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 283574 32614
rect 282954 32294 283574 32378
rect 282954 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 283574 32294
rect 281395 4860 281461 4861
rect 281395 4796 281396 4860
rect 281460 4796 281461 4860
rect 281395 4795 281461 4796
rect 279234 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 279854 -5146
rect 279234 -5466 279854 -5382
rect 279234 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 279854 -5466
rect 279234 -5734 279854 -5702
rect 264954 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 265574 -6106
rect 264954 -6426 265574 -6342
rect 264954 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 265574 -6426
rect 264954 -7654 265574 -6662
rect 282954 -7066 283574 32058
rect 289794 39454 290414 74898
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 292438 11661 292498 97275
rect 293514 79174 294134 98000
rect 295011 96932 295077 96933
rect 295011 96868 295012 96932
rect 295076 96868 295077 96932
rect 295011 96867 295077 96868
rect 295195 96932 295261 96933
rect 295195 96868 295196 96932
rect 295260 96868 295261 96932
rect 295195 96867 295261 96868
rect 295014 93125 295074 96867
rect 295011 93124 295077 93125
rect 295011 93060 295012 93124
rect 295076 93060 295077 93124
rect 295011 93059 295077 93060
rect 295198 89045 295258 96867
rect 295195 89044 295261 89045
rect 295195 88980 295196 89044
rect 295260 88980 295261 89044
rect 295195 88979 295261 88980
rect 293514 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 294134 79174
rect 293514 78854 294134 78938
rect 293514 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 294134 78854
rect 293514 43174 294134 78618
rect 293514 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 294134 43174
rect 293514 42854 294134 42938
rect 293514 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 294134 42854
rect 292435 11660 292501 11661
rect 292435 11596 292436 11660
rect 292500 11596 292501 11660
rect 292435 11595 292501 11596
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -1894 290414 -902
rect 293514 7174 294134 42618
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 293514 -2266 294134 6618
rect 293514 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 294134 -2266
rect 293514 -2586 294134 -2502
rect 293514 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 294134 -2586
rect 293514 -3814 294134 -2822
rect 297234 82894 297854 98000
rect 299243 96932 299309 96933
rect 299243 96868 299244 96932
rect 299308 96868 299309 96932
rect 299243 96867 299309 96868
rect 297234 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 297854 82894
rect 297234 82574 297854 82658
rect 297234 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 297854 82574
rect 297234 46894 297854 82338
rect 299246 50285 299306 96867
rect 300954 86614 301574 98000
rect 300954 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 301574 86614
rect 300954 86294 301574 86378
rect 300954 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 301574 86294
rect 300954 50614 301574 86058
rect 300954 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 301574 50614
rect 300954 50294 301574 50378
rect 299243 50284 299309 50285
rect 299243 50220 299244 50284
rect 299308 50220 299309 50284
rect 299243 50219 299309 50220
rect 297234 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 297854 46894
rect 297234 46574 297854 46658
rect 297234 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 297854 46574
rect 297234 10894 297854 46338
rect 297234 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 297854 10894
rect 297234 10574 297854 10658
rect 297234 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 297854 10574
rect 297234 -4186 297854 10338
rect 297234 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 297854 -4186
rect 297234 -4506 297854 -4422
rect 297234 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 297854 -4506
rect 297234 -5734 297854 -4742
rect 300954 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 301574 50294
rect 300954 14614 301574 50058
rect 300954 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 301574 14614
rect 300954 14294 301574 14378
rect 300954 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 301574 14294
rect 282954 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 283574 -7066
rect 282954 -7386 283574 -7302
rect 282954 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 283574 -7386
rect 282954 -7654 283574 -7622
rect 300954 -6106 301574 14058
rect 307794 93454 308414 128898
rect 307794 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 308414 93454
rect 307794 93134 308414 93218
rect 307794 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 308414 93134
rect 307794 57454 308414 92898
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -1306 308414 20898
rect 307794 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 308414 -1306
rect 307794 -1626 308414 -1542
rect 307794 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 308414 -1626
rect 307794 -1894 308414 -1862
rect 311514 673174 312134 707162
rect 311514 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 312134 673174
rect 311514 672854 312134 672938
rect 311514 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 312134 672854
rect 311514 637174 312134 672618
rect 311514 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 312134 637174
rect 311514 636854 312134 636938
rect 311514 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 312134 636854
rect 311514 601174 312134 636618
rect 311514 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 312134 601174
rect 311514 600854 312134 600938
rect 311514 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 312134 600854
rect 311514 565174 312134 600618
rect 311514 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 312134 565174
rect 311514 564854 312134 564938
rect 311514 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 312134 564854
rect 311514 529174 312134 564618
rect 311514 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 312134 529174
rect 311514 528854 312134 528938
rect 311514 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 312134 528854
rect 311514 493174 312134 528618
rect 311514 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 312134 493174
rect 311514 492854 312134 492938
rect 311514 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 312134 492854
rect 311514 457174 312134 492618
rect 311514 456938 311546 457174
rect 311782 456938 311866 457174
rect 312102 456938 312134 457174
rect 311514 456854 312134 456938
rect 311514 456618 311546 456854
rect 311782 456618 311866 456854
rect 312102 456618 312134 456854
rect 311514 421174 312134 456618
rect 311514 420938 311546 421174
rect 311782 420938 311866 421174
rect 312102 420938 312134 421174
rect 311514 420854 312134 420938
rect 311514 420618 311546 420854
rect 311782 420618 311866 420854
rect 312102 420618 312134 420854
rect 311514 385174 312134 420618
rect 311514 384938 311546 385174
rect 311782 384938 311866 385174
rect 312102 384938 312134 385174
rect 311514 384854 312134 384938
rect 311514 384618 311546 384854
rect 311782 384618 311866 384854
rect 312102 384618 312134 384854
rect 311514 349174 312134 384618
rect 311514 348938 311546 349174
rect 311782 348938 311866 349174
rect 312102 348938 312134 349174
rect 311514 348854 312134 348938
rect 311514 348618 311546 348854
rect 311782 348618 311866 348854
rect 312102 348618 312134 348854
rect 311514 313174 312134 348618
rect 311514 312938 311546 313174
rect 311782 312938 311866 313174
rect 312102 312938 312134 313174
rect 311514 312854 312134 312938
rect 311514 312618 311546 312854
rect 311782 312618 311866 312854
rect 312102 312618 312134 312854
rect 311514 277174 312134 312618
rect 311514 276938 311546 277174
rect 311782 276938 311866 277174
rect 312102 276938 312134 277174
rect 311514 276854 312134 276938
rect 311514 276618 311546 276854
rect 311782 276618 311866 276854
rect 312102 276618 312134 276854
rect 311514 241174 312134 276618
rect 311514 240938 311546 241174
rect 311782 240938 311866 241174
rect 312102 240938 312134 241174
rect 311514 240854 312134 240938
rect 311514 240618 311546 240854
rect 311782 240618 311866 240854
rect 312102 240618 312134 240854
rect 311514 205174 312134 240618
rect 311514 204938 311546 205174
rect 311782 204938 311866 205174
rect 312102 204938 312134 205174
rect 311514 204854 312134 204938
rect 311514 204618 311546 204854
rect 311782 204618 311866 204854
rect 312102 204618 312134 204854
rect 311514 169174 312134 204618
rect 311514 168938 311546 169174
rect 311782 168938 311866 169174
rect 312102 168938 312134 169174
rect 311514 168854 312134 168938
rect 311514 168618 311546 168854
rect 311782 168618 311866 168854
rect 312102 168618 312134 168854
rect 311514 133174 312134 168618
rect 311514 132938 311546 133174
rect 311782 132938 311866 133174
rect 312102 132938 312134 133174
rect 311514 132854 312134 132938
rect 311514 132618 311546 132854
rect 311782 132618 311866 132854
rect 312102 132618 312134 132854
rect 311514 97174 312134 132618
rect 311514 96938 311546 97174
rect 311782 96938 311866 97174
rect 312102 96938 312134 97174
rect 311514 96854 312134 96938
rect 311514 96618 311546 96854
rect 311782 96618 311866 96854
rect 312102 96618 312134 96854
rect 311514 61174 312134 96618
rect 311514 60938 311546 61174
rect 311782 60938 311866 61174
rect 312102 60938 312134 61174
rect 311514 60854 312134 60938
rect 311514 60618 311546 60854
rect 311782 60618 311866 60854
rect 312102 60618 312134 60854
rect 311514 25174 312134 60618
rect 311514 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 312134 25174
rect 311514 24854 312134 24938
rect 311514 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 312134 24854
rect 311514 -3226 312134 24618
rect 311514 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 312134 -3226
rect 311514 -3546 312134 -3462
rect 311514 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 312134 -3546
rect 311514 -3814 312134 -3782
rect 315234 676894 315854 709082
rect 315234 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 315854 676894
rect 315234 676574 315854 676658
rect 315234 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 315854 676574
rect 315234 640894 315854 676338
rect 315234 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 315854 640894
rect 315234 640574 315854 640658
rect 315234 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 315854 640574
rect 315234 604894 315854 640338
rect 315234 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 315854 604894
rect 315234 604574 315854 604658
rect 315234 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 315854 604574
rect 315234 568894 315854 604338
rect 315234 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 315854 568894
rect 315234 568574 315854 568658
rect 315234 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 315854 568574
rect 315234 532894 315854 568338
rect 315234 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 315854 532894
rect 315234 532574 315854 532658
rect 315234 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 315854 532574
rect 315234 496894 315854 532338
rect 315234 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 315854 496894
rect 315234 496574 315854 496658
rect 315234 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 315854 496574
rect 315234 460894 315854 496338
rect 315234 460658 315266 460894
rect 315502 460658 315586 460894
rect 315822 460658 315854 460894
rect 315234 460574 315854 460658
rect 315234 460338 315266 460574
rect 315502 460338 315586 460574
rect 315822 460338 315854 460574
rect 315234 424894 315854 460338
rect 315234 424658 315266 424894
rect 315502 424658 315586 424894
rect 315822 424658 315854 424894
rect 315234 424574 315854 424658
rect 315234 424338 315266 424574
rect 315502 424338 315586 424574
rect 315822 424338 315854 424574
rect 315234 388894 315854 424338
rect 315234 388658 315266 388894
rect 315502 388658 315586 388894
rect 315822 388658 315854 388894
rect 315234 388574 315854 388658
rect 315234 388338 315266 388574
rect 315502 388338 315586 388574
rect 315822 388338 315854 388574
rect 315234 352894 315854 388338
rect 315234 352658 315266 352894
rect 315502 352658 315586 352894
rect 315822 352658 315854 352894
rect 315234 352574 315854 352658
rect 315234 352338 315266 352574
rect 315502 352338 315586 352574
rect 315822 352338 315854 352574
rect 315234 316894 315854 352338
rect 315234 316658 315266 316894
rect 315502 316658 315586 316894
rect 315822 316658 315854 316894
rect 315234 316574 315854 316658
rect 315234 316338 315266 316574
rect 315502 316338 315586 316574
rect 315822 316338 315854 316574
rect 315234 280894 315854 316338
rect 315234 280658 315266 280894
rect 315502 280658 315586 280894
rect 315822 280658 315854 280894
rect 315234 280574 315854 280658
rect 315234 280338 315266 280574
rect 315502 280338 315586 280574
rect 315822 280338 315854 280574
rect 315234 244894 315854 280338
rect 315234 244658 315266 244894
rect 315502 244658 315586 244894
rect 315822 244658 315854 244894
rect 315234 244574 315854 244658
rect 315234 244338 315266 244574
rect 315502 244338 315586 244574
rect 315822 244338 315854 244574
rect 315234 208894 315854 244338
rect 315234 208658 315266 208894
rect 315502 208658 315586 208894
rect 315822 208658 315854 208894
rect 315234 208574 315854 208658
rect 315234 208338 315266 208574
rect 315502 208338 315586 208574
rect 315822 208338 315854 208574
rect 315234 172894 315854 208338
rect 315234 172658 315266 172894
rect 315502 172658 315586 172894
rect 315822 172658 315854 172894
rect 315234 172574 315854 172658
rect 315234 172338 315266 172574
rect 315502 172338 315586 172574
rect 315822 172338 315854 172574
rect 315234 136894 315854 172338
rect 315234 136658 315266 136894
rect 315502 136658 315586 136894
rect 315822 136658 315854 136894
rect 315234 136574 315854 136658
rect 315234 136338 315266 136574
rect 315502 136338 315586 136574
rect 315822 136338 315854 136574
rect 315234 100894 315854 136338
rect 315234 100658 315266 100894
rect 315502 100658 315586 100894
rect 315822 100658 315854 100894
rect 315234 100574 315854 100658
rect 315234 100338 315266 100574
rect 315502 100338 315586 100574
rect 315822 100338 315854 100574
rect 315234 64894 315854 100338
rect 315234 64658 315266 64894
rect 315502 64658 315586 64894
rect 315822 64658 315854 64894
rect 315234 64574 315854 64658
rect 315234 64338 315266 64574
rect 315502 64338 315586 64574
rect 315822 64338 315854 64574
rect 315234 28894 315854 64338
rect 315234 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 315854 28894
rect 315234 28574 315854 28658
rect 315234 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 315854 28574
rect 315234 -5146 315854 28338
rect 315234 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 315854 -5146
rect 315234 -5466 315854 -5382
rect 315234 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 315854 -5466
rect 315234 -5734 315854 -5702
rect 318954 680614 319574 711002
rect 336954 710598 337574 711590
rect 336954 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 337574 710598
rect 336954 710278 337574 710362
rect 336954 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 337574 710278
rect 333234 708678 333854 709670
rect 333234 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 333854 708678
rect 333234 708358 333854 708442
rect 333234 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 333854 708358
rect 329514 706758 330134 707750
rect 329514 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 330134 706758
rect 329514 706438 330134 706522
rect 329514 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 330134 706438
rect 318954 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 319574 680614
rect 318954 680294 319574 680378
rect 318954 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 319574 680294
rect 318954 644614 319574 680058
rect 318954 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 319574 644614
rect 318954 644294 319574 644378
rect 318954 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 319574 644294
rect 318954 608614 319574 644058
rect 318954 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 319574 608614
rect 318954 608294 319574 608378
rect 318954 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 319574 608294
rect 318954 572614 319574 608058
rect 318954 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 319574 572614
rect 318954 572294 319574 572378
rect 318954 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 319574 572294
rect 318954 536614 319574 572058
rect 318954 536378 318986 536614
rect 319222 536378 319306 536614
rect 319542 536378 319574 536614
rect 318954 536294 319574 536378
rect 318954 536058 318986 536294
rect 319222 536058 319306 536294
rect 319542 536058 319574 536294
rect 318954 500614 319574 536058
rect 318954 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 319574 500614
rect 318954 500294 319574 500378
rect 318954 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 319574 500294
rect 318954 464614 319574 500058
rect 318954 464378 318986 464614
rect 319222 464378 319306 464614
rect 319542 464378 319574 464614
rect 318954 464294 319574 464378
rect 318954 464058 318986 464294
rect 319222 464058 319306 464294
rect 319542 464058 319574 464294
rect 318954 428614 319574 464058
rect 318954 428378 318986 428614
rect 319222 428378 319306 428614
rect 319542 428378 319574 428614
rect 318954 428294 319574 428378
rect 318954 428058 318986 428294
rect 319222 428058 319306 428294
rect 319542 428058 319574 428294
rect 318954 392614 319574 428058
rect 318954 392378 318986 392614
rect 319222 392378 319306 392614
rect 319542 392378 319574 392614
rect 318954 392294 319574 392378
rect 318954 392058 318986 392294
rect 319222 392058 319306 392294
rect 319542 392058 319574 392294
rect 318954 356614 319574 392058
rect 318954 356378 318986 356614
rect 319222 356378 319306 356614
rect 319542 356378 319574 356614
rect 318954 356294 319574 356378
rect 318954 356058 318986 356294
rect 319222 356058 319306 356294
rect 319542 356058 319574 356294
rect 318954 320614 319574 356058
rect 318954 320378 318986 320614
rect 319222 320378 319306 320614
rect 319542 320378 319574 320614
rect 318954 320294 319574 320378
rect 318954 320058 318986 320294
rect 319222 320058 319306 320294
rect 319542 320058 319574 320294
rect 318954 284614 319574 320058
rect 318954 284378 318986 284614
rect 319222 284378 319306 284614
rect 319542 284378 319574 284614
rect 318954 284294 319574 284378
rect 318954 284058 318986 284294
rect 319222 284058 319306 284294
rect 319542 284058 319574 284294
rect 318954 248614 319574 284058
rect 318954 248378 318986 248614
rect 319222 248378 319306 248614
rect 319542 248378 319574 248614
rect 318954 248294 319574 248378
rect 318954 248058 318986 248294
rect 319222 248058 319306 248294
rect 319542 248058 319574 248294
rect 318954 212614 319574 248058
rect 318954 212378 318986 212614
rect 319222 212378 319306 212614
rect 319542 212378 319574 212614
rect 318954 212294 319574 212378
rect 318954 212058 318986 212294
rect 319222 212058 319306 212294
rect 319542 212058 319574 212294
rect 318954 176614 319574 212058
rect 318954 176378 318986 176614
rect 319222 176378 319306 176614
rect 319542 176378 319574 176614
rect 318954 176294 319574 176378
rect 318954 176058 318986 176294
rect 319222 176058 319306 176294
rect 319542 176058 319574 176294
rect 318954 140614 319574 176058
rect 318954 140378 318986 140614
rect 319222 140378 319306 140614
rect 319542 140378 319574 140614
rect 318954 140294 319574 140378
rect 318954 140058 318986 140294
rect 319222 140058 319306 140294
rect 319542 140058 319574 140294
rect 318954 104614 319574 140058
rect 318954 104378 318986 104614
rect 319222 104378 319306 104614
rect 319542 104378 319574 104614
rect 318954 104294 319574 104378
rect 318954 104058 318986 104294
rect 319222 104058 319306 104294
rect 319542 104058 319574 104294
rect 318954 68614 319574 104058
rect 318954 68378 318986 68614
rect 319222 68378 319306 68614
rect 319542 68378 319574 68614
rect 318954 68294 319574 68378
rect 318954 68058 318986 68294
rect 319222 68058 319306 68294
rect 319542 68058 319574 68294
rect 318954 32614 319574 68058
rect 318954 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 319574 32614
rect 318954 32294 319574 32378
rect 318954 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 319574 32294
rect 300954 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 301574 -6106
rect 300954 -6426 301574 -6342
rect 300954 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 301574 -6426
rect 300954 -7654 301574 -6662
rect 318954 -7066 319574 32058
rect 325794 704838 326414 705830
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 543454 326414 578898
rect 325794 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 326414 543454
rect 325794 543134 326414 543218
rect 325794 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 326414 543134
rect 325794 507454 326414 542898
rect 325794 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 326414 507454
rect 325794 507134 326414 507218
rect 325794 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 326414 507134
rect 325794 471454 326414 506898
rect 325794 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 326414 471454
rect 325794 471134 326414 471218
rect 325794 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 326414 471134
rect 325794 435454 326414 470898
rect 325794 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 326414 435454
rect 325794 435134 326414 435218
rect 325794 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 326414 435134
rect 325794 399454 326414 434898
rect 325794 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 326414 399454
rect 325794 399134 326414 399218
rect 325794 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 326414 399134
rect 325794 363454 326414 398898
rect 325794 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 326414 363454
rect 325794 363134 326414 363218
rect 325794 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 326414 363134
rect 325794 327454 326414 362898
rect 325794 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 326414 327454
rect 325794 327134 326414 327218
rect 325794 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 326414 327134
rect 325794 291454 326414 326898
rect 325794 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 326414 291454
rect 325794 291134 326414 291218
rect 325794 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 326414 291134
rect 325794 255454 326414 290898
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 325794 219454 326414 254898
rect 325794 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 326414 219454
rect 325794 219134 326414 219218
rect 325794 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 326414 219134
rect 325794 183454 326414 218898
rect 325794 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 326414 183454
rect 325794 183134 326414 183218
rect 325794 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 326414 183134
rect 325794 147454 326414 182898
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 325794 111454 326414 146898
rect 325794 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 326414 111454
rect 325794 111134 326414 111218
rect 325794 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 326414 111134
rect 325794 75454 326414 110898
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -1894 326414 -902
rect 329514 691174 330134 706202
rect 329514 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 330134 691174
rect 329514 690854 330134 690938
rect 329514 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 330134 690854
rect 329514 655174 330134 690618
rect 329514 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 330134 655174
rect 329514 654854 330134 654938
rect 329514 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 330134 654854
rect 329514 619174 330134 654618
rect 329514 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 330134 619174
rect 329514 618854 330134 618938
rect 329514 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 330134 618854
rect 329514 583174 330134 618618
rect 329514 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 330134 583174
rect 329514 582854 330134 582938
rect 329514 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 330134 582854
rect 329514 547174 330134 582618
rect 329514 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 330134 547174
rect 329514 546854 330134 546938
rect 329514 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 330134 546854
rect 329514 511174 330134 546618
rect 329514 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 330134 511174
rect 329514 510854 330134 510938
rect 329514 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 330134 510854
rect 329514 475174 330134 510618
rect 329514 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 330134 475174
rect 329514 474854 330134 474938
rect 329514 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 330134 474854
rect 329514 439174 330134 474618
rect 329514 438938 329546 439174
rect 329782 438938 329866 439174
rect 330102 438938 330134 439174
rect 329514 438854 330134 438938
rect 329514 438618 329546 438854
rect 329782 438618 329866 438854
rect 330102 438618 330134 438854
rect 329514 403174 330134 438618
rect 329514 402938 329546 403174
rect 329782 402938 329866 403174
rect 330102 402938 330134 403174
rect 329514 402854 330134 402938
rect 329514 402618 329546 402854
rect 329782 402618 329866 402854
rect 330102 402618 330134 402854
rect 329514 367174 330134 402618
rect 329514 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 330134 367174
rect 329514 366854 330134 366938
rect 329514 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 330134 366854
rect 329514 331174 330134 366618
rect 329514 330938 329546 331174
rect 329782 330938 329866 331174
rect 330102 330938 330134 331174
rect 329514 330854 330134 330938
rect 329514 330618 329546 330854
rect 329782 330618 329866 330854
rect 330102 330618 330134 330854
rect 329514 295174 330134 330618
rect 329514 294938 329546 295174
rect 329782 294938 329866 295174
rect 330102 294938 330134 295174
rect 329514 294854 330134 294938
rect 329514 294618 329546 294854
rect 329782 294618 329866 294854
rect 330102 294618 330134 294854
rect 329514 259174 330134 294618
rect 329514 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 330134 259174
rect 329514 258854 330134 258938
rect 329514 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 330134 258854
rect 329514 223174 330134 258618
rect 329514 222938 329546 223174
rect 329782 222938 329866 223174
rect 330102 222938 330134 223174
rect 329514 222854 330134 222938
rect 329514 222618 329546 222854
rect 329782 222618 329866 222854
rect 330102 222618 330134 222854
rect 329514 187174 330134 222618
rect 329514 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 330134 187174
rect 329514 186854 330134 186938
rect 329514 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 330134 186854
rect 329514 151174 330134 186618
rect 329514 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 330134 151174
rect 329514 150854 330134 150938
rect 329514 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 330134 150854
rect 329514 115174 330134 150618
rect 329514 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 330134 115174
rect 329514 114854 330134 114938
rect 329514 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 330134 114854
rect 329514 79174 330134 114618
rect 329514 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 330134 79174
rect 329514 78854 330134 78938
rect 329514 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 330134 78854
rect 329514 43174 330134 78618
rect 329514 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 330134 43174
rect 329514 42854 330134 42938
rect 329514 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 330134 42854
rect 329514 7174 330134 42618
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 329514 -2266 330134 6618
rect 329514 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 330134 -2266
rect 329514 -2586 330134 -2502
rect 329514 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 330134 -2586
rect 329514 -3814 330134 -2822
rect 333234 694894 333854 708122
rect 333234 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 333854 694894
rect 333234 694574 333854 694658
rect 333234 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 333854 694574
rect 333234 658894 333854 694338
rect 333234 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 333854 658894
rect 333234 658574 333854 658658
rect 333234 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 333854 658574
rect 333234 622894 333854 658338
rect 333234 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 333854 622894
rect 333234 622574 333854 622658
rect 333234 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 333854 622574
rect 333234 586894 333854 622338
rect 333234 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 333854 586894
rect 333234 586574 333854 586658
rect 333234 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 333854 586574
rect 333234 550894 333854 586338
rect 333234 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 333854 550894
rect 333234 550574 333854 550658
rect 333234 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 333854 550574
rect 333234 514894 333854 550338
rect 333234 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 333854 514894
rect 333234 514574 333854 514658
rect 333234 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 333854 514574
rect 333234 478894 333854 514338
rect 333234 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 333854 478894
rect 333234 478574 333854 478658
rect 333234 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 333854 478574
rect 333234 442894 333854 478338
rect 333234 442658 333266 442894
rect 333502 442658 333586 442894
rect 333822 442658 333854 442894
rect 333234 442574 333854 442658
rect 333234 442338 333266 442574
rect 333502 442338 333586 442574
rect 333822 442338 333854 442574
rect 333234 406894 333854 442338
rect 333234 406658 333266 406894
rect 333502 406658 333586 406894
rect 333822 406658 333854 406894
rect 333234 406574 333854 406658
rect 333234 406338 333266 406574
rect 333502 406338 333586 406574
rect 333822 406338 333854 406574
rect 333234 370894 333854 406338
rect 333234 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 333854 370894
rect 333234 370574 333854 370658
rect 333234 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 333854 370574
rect 333234 334894 333854 370338
rect 333234 334658 333266 334894
rect 333502 334658 333586 334894
rect 333822 334658 333854 334894
rect 333234 334574 333854 334658
rect 333234 334338 333266 334574
rect 333502 334338 333586 334574
rect 333822 334338 333854 334574
rect 333234 298894 333854 334338
rect 333234 298658 333266 298894
rect 333502 298658 333586 298894
rect 333822 298658 333854 298894
rect 333234 298574 333854 298658
rect 333234 298338 333266 298574
rect 333502 298338 333586 298574
rect 333822 298338 333854 298574
rect 333234 262894 333854 298338
rect 333234 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 333854 262894
rect 333234 262574 333854 262658
rect 333234 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 333854 262574
rect 333234 226894 333854 262338
rect 333234 226658 333266 226894
rect 333502 226658 333586 226894
rect 333822 226658 333854 226894
rect 333234 226574 333854 226658
rect 333234 226338 333266 226574
rect 333502 226338 333586 226574
rect 333822 226338 333854 226574
rect 333234 190894 333854 226338
rect 333234 190658 333266 190894
rect 333502 190658 333586 190894
rect 333822 190658 333854 190894
rect 333234 190574 333854 190658
rect 333234 190338 333266 190574
rect 333502 190338 333586 190574
rect 333822 190338 333854 190574
rect 333234 154894 333854 190338
rect 333234 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 333854 154894
rect 333234 154574 333854 154658
rect 333234 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 333854 154574
rect 333234 118894 333854 154338
rect 333234 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 333854 118894
rect 333234 118574 333854 118658
rect 333234 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 333854 118574
rect 333234 82894 333854 118338
rect 333234 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 333854 82894
rect 333234 82574 333854 82658
rect 333234 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 333854 82574
rect 333234 46894 333854 82338
rect 333234 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 333854 46894
rect 333234 46574 333854 46658
rect 333234 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 333854 46574
rect 333234 10894 333854 46338
rect 333234 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 333854 10894
rect 333234 10574 333854 10658
rect 333234 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 333854 10574
rect 333234 -4186 333854 10338
rect 333234 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 333854 -4186
rect 333234 -4506 333854 -4422
rect 333234 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 333854 -4506
rect 333234 -5734 333854 -4742
rect 336954 698614 337574 710042
rect 354954 711558 355574 711590
rect 354954 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 355574 711558
rect 354954 711238 355574 711322
rect 354954 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 355574 711238
rect 351234 709638 351854 709670
rect 351234 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 351854 709638
rect 351234 709318 351854 709402
rect 351234 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 351854 709318
rect 347514 707718 348134 707750
rect 347514 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 348134 707718
rect 347514 707398 348134 707482
rect 347514 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 348134 707398
rect 336954 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 337574 698614
rect 336954 698294 337574 698378
rect 336954 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 337574 698294
rect 336954 662614 337574 698058
rect 336954 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 337574 662614
rect 336954 662294 337574 662378
rect 336954 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 337574 662294
rect 336954 626614 337574 662058
rect 336954 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 337574 626614
rect 336954 626294 337574 626378
rect 336954 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 337574 626294
rect 336954 590614 337574 626058
rect 336954 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 337574 590614
rect 336954 590294 337574 590378
rect 336954 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 337574 590294
rect 336954 554614 337574 590058
rect 336954 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 337574 554614
rect 336954 554294 337574 554378
rect 336954 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 337574 554294
rect 336954 518614 337574 554058
rect 336954 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 337574 518614
rect 336954 518294 337574 518378
rect 336954 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 337574 518294
rect 336954 482614 337574 518058
rect 336954 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 337574 482614
rect 336954 482294 337574 482378
rect 336954 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 337574 482294
rect 336954 446614 337574 482058
rect 336954 446378 336986 446614
rect 337222 446378 337306 446614
rect 337542 446378 337574 446614
rect 336954 446294 337574 446378
rect 336954 446058 336986 446294
rect 337222 446058 337306 446294
rect 337542 446058 337574 446294
rect 336954 410614 337574 446058
rect 336954 410378 336986 410614
rect 337222 410378 337306 410614
rect 337542 410378 337574 410614
rect 336954 410294 337574 410378
rect 336954 410058 336986 410294
rect 337222 410058 337306 410294
rect 337542 410058 337574 410294
rect 336954 374614 337574 410058
rect 336954 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 337574 374614
rect 336954 374294 337574 374378
rect 336954 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 337574 374294
rect 336954 338614 337574 374058
rect 336954 338378 336986 338614
rect 337222 338378 337306 338614
rect 337542 338378 337574 338614
rect 336954 338294 337574 338378
rect 336954 338058 336986 338294
rect 337222 338058 337306 338294
rect 337542 338058 337574 338294
rect 336954 302614 337574 338058
rect 336954 302378 336986 302614
rect 337222 302378 337306 302614
rect 337542 302378 337574 302614
rect 336954 302294 337574 302378
rect 336954 302058 336986 302294
rect 337222 302058 337306 302294
rect 337542 302058 337574 302294
rect 336954 266614 337574 302058
rect 336954 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 337574 266614
rect 336954 266294 337574 266378
rect 336954 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 337574 266294
rect 336954 230614 337574 266058
rect 336954 230378 336986 230614
rect 337222 230378 337306 230614
rect 337542 230378 337574 230614
rect 336954 230294 337574 230378
rect 336954 230058 336986 230294
rect 337222 230058 337306 230294
rect 337542 230058 337574 230294
rect 336954 194614 337574 230058
rect 336954 194378 336986 194614
rect 337222 194378 337306 194614
rect 337542 194378 337574 194614
rect 336954 194294 337574 194378
rect 336954 194058 336986 194294
rect 337222 194058 337306 194294
rect 337542 194058 337574 194294
rect 336954 158614 337574 194058
rect 336954 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 337574 158614
rect 336954 158294 337574 158378
rect 336954 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 337574 158294
rect 336954 122614 337574 158058
rect 336954 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 337574 122614
rect 336954 122294 337574 122378
rect 336954 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 337574 122294
rect 336954 86614 337574 122058
rect 336954 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 337574 86614
rect 336954 86294 337574 86378
rect 336954 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 337574 86294
rect 336954 50614 337574 86058
rect 336954 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 337574 50614
rect 336954 50294 337574 50378
rect 336954 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 337574 50294
rect 336954 14614 337574 50058
rect 336954 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 337574 14614
rect 336954 14294 337574 14378
rect 336954 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 337574 14294
rect 318954 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 319574 -7066
rect 318954 -7386 319574 -7302
rect 318954 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 319574 -7386
rect 318954 -7654 319574 -7622
rect 336954 -6106 337574 14058
rect 343794 705798 344414 705830
rect 343794 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 344414 705798
rect 343794 705478 344414 705562
rect 343794 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 344414 705478
rect 343794 669454 344414 705242
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 561454 344414 596898
rect 343794 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 344414 561454
rect 343794 561134 344414 561218
rect 343794 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 344414 561134
rect 343794 525454 344414 560898
rect 343794 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 344414 525454
rect 343794 525134 344414 525218
rect 343794 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 344414 525134
rect 343794 489454 344414 524898
rect 343794 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 344414 489454
rect 343794 489134 344414 489218
rect 343794 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 344414 489134
rect 343794 453454 344414 488898
rect 343794 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 344414 453454
rect 343794 453134 344414 453218
rect 343794 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 344414 453134
rect 343794 417454 344414 452898
rect 343794 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 344414 417454
rect 343794 417134 344414 417218
rect 343794 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 344414 417134
rect 343794 381454 344414 416898
rect 343794 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 344414 381454
rect 343794 381134 344414 381218
rect 343794 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 344414 381134
rect 343794 345454 344414 380898
rect 343794 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 344414 345454
rect 343794 345134 344414 345218
rect 343794 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 344414 345134
rect 343794 309454 344414 344898
rect 343794 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 344414 309454
rect 343794 309134 344414 309218
rect 343794 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 344414 309134
rect 343794 273454 344414 308898
rect 343794 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 344414 273454
rect 343794 273134 344414 273218
rect 343794 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 344414 273134
rect 343794 237454 344414 272898
rect 343794 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 344414 237454
rect 343794 237134 344414 237218
rect 343794 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 344414 237134
rect 343794 201454 344414 236898
rect 343794 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 344414 201454
rect 343794 201134 344414 201218
rect 343794 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 344414 201134
rect 343794 165454 344414 200898
rect 343794 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 344414 165454
rect 343794 165134 344414 165218
rect 343794 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 344414 165134
rect 343794 129454 344414 164898
rect 343794 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 344414 129454
rect 343794 129134 344414 129218
rect 343794 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 344414 129134
rect 343794 93454 344414 128898
rect 343794 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 344414 93454
rect 343794 93134 344414 93218
rect 343794 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 344414 93134
rect 343794 57454 344414 92898
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -1306 344414 20898
rect 343794 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 344414 -1306
rect 343794 -1626 344414 -1542
rect 343794 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 344414 -1626
rect 343794 -1894 344414 -1862
rect 347514 673174 348134 707162
rect 347514 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 348134 673174
rect 347514 672854 348134 672938
rect 347514 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 348134 672854
rect 347514 637174 348134 672618
rect 347514 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 348134 637174
rect 347514 636854 348134 636938
rect 347514 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 348134 636854
rect 347514 601174 348134 636618
rect 347514 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 348134 601174
rect 347514 600854 348134 600938
rect 347514 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 348134 600854
rect 347514 565174 348134 600618
rect 347514 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 348134 565174
rect 347514 564854 348134 564938
rect 347514 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 348134 564854
rect 347514 529174 348134 564618
rect 347514 528938 347546 529174
rect 347782 528938 347866 529174
rect 348102 528938 348134 529174
rect 347514 528854 348134 528938
rect 347514 528618 347546 528854
rect 347782 528618 347866 528854
rect 348102 528618 348134 528854
rect 347514 493174 348134 528618
rect 347514 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 348134 493174
rect 347514 492854 348134 492938
rect 347514 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 348134 492854
rect 347514 457174 348134 492618
rect 347514 456938 347546 457174
rect 347782 456938 347866 457174
rect 348102 456938 348134 457174
rect 347514 456854 348134 456938
rect 347514 456618 347546 456854
rect 347782 456618 347866 456854
rect 348102 456618 348134 456854
rect 347514 421174 348134 456618
rect 347514 420938 347546 421174
rect 347782 420938 347866 421174
rect 348102 420938 348134 421174
rect 347514 420854 348134 420938
rect 347514 420618 347546 420854
rect 347782 420618 347866 420854
rect 348102 420618 348134 420854
rect 347514 385174 348134 420618
rect 347514 384938 347546 385174
rect 347782 384938 347866 385174
rect 348102 384938 348134 385174
rect 347514 384854 348134 384938
rect 347514 384618 347546 384854
rect 347782 384618 347866 384854
rect 348102 384618 348134 384854
rect 347514 349174 348134 384618
rect 347514 348938 347546 349174
rect 347782 348938 347866 349174
rect 348102 348938 348134 349174
rect 347514 348854 348134 348938
rect 347514 348618 347546 348854
rect 347782 348618 347866 348854
rect 348102 348618 348134 348854
rect 347514 313174 348134 348618
rect 347514 312938 347546 313174
rect 347782 312938 347866 313174
rect 348102 312938 348134 313174
rect 347514 312854 348134 312938
rect 347514 312618 347546 312854
rect 347782 312618 347866 312854
rect 348102 312618 348134 312854
rect 347514 277174 348134 312618
rect 347514 276938 347546 277174
rect 347782 276938 347866 277174
rect 348102 276938 348134 277174
rect 347514 276854 348134 276938
rect 347514 276618 347546 276854
rect 347782 276618 347866 276854
rect 348102 276618 348134 276854
rect 347514 241174 348134 276618
rect 347514 240938 347546 241174
rect 347782 240938 347866 241174
rect 348102 240938 348134 241174
rect 347514 240854 348134 240938
rect 347514 240618 347546 240854
rect 347782 240618 347866 240854
rect 348102 240618 348134 240854
rect 347514 205174 348134 240618
rect 347514 204938 347546 205174
rect 347782 204938 347866 205174
rect 348102 204938 348134 205174
rect 347514 204854 348134 204938
rect 347514 204618 347546 204854
rect 347782 204618 347866 204854
rect 348102 204618 348134 204854
rect 347514 169174 348134 204618
rect 347514 168938 347546 169174
rect 347782 168938 347866 169174
rect 348102 168938 348134 169174
rect 347514 168854 348134 168938
rect 347514 168618 347546 168854
rect 347782 168618 347866 168854
rect 348102 168618 348134 168854
rect 347514 133174 348134 168618
rect 347514 132938 347546 133174
rect 347782 132938 347866 133174
rect 348102 132938 348134 133174
rect 347514 132854 348134 132938
rect 347514 132618 347546 132854
rect 347782 132618 347866 132854
rect 348102 132618 348134 132854
rect 347514 97174 348134 132618
rect 347514 96938 347546 97174
rect 347782 96938 347866 97174
rect 348102 96938 348134 97174
rect 347514 96854 348134 96938
rect 347514 96618 347546 96854
rect 347782 96618 347866 96854
rect 348102 96618 348134 96854
rect 347514 61174 348134 96618
rect 347514 60938 347546 61174
rect 347782 60938 347866 61174
rect 348102 60938 348134 61174
rect 347514 60854 348134 60938
rect 347514 60618 347546 60854
rect 347782 60618 347866 60854
rect 348102 60618 348134 60854
rect 347514 25174 348134 60618
rect 347514 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 348134 25174
rect 347514 24854 348134 24938
rect 347514 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 348134 24854
rect 347514 -3226 348134 24618
rect 347514 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 348134 -3226
rect 347514 -3546 348134 -3462
rect 347514 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 348134 -3546
rect 347514 -3814 348134 -3782
rect 351234 676894 351854 709082
rect 351234 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 351854 676894
rect 351234 676574 351854 676658
rect 351234 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 351854 676574
rect 351234 640894 351854 676338
rect 351234 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 351854 640894
rect 351234 640574 351854 640658
rect 351234 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 351854 640574
rect 351234 604894 351854 640338
rect 351234 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 351854 604894
rect 351234 604574 351854 604658
rect 351234 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 351854 604574
rect 351234 568894 351854 604338
rect 351234 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 351854 568894
rect 351234 568574 351854 568658
rect 351234 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 351854 568574
rect 351234 532894 351854 568338
rect 351234 532658 351266 532894
rect 351502 532658 351586 532894
rect 351822 532658 351854 532894
rect 351234 532574 351854 532658
rect 351234 532338 351266 532574
rect 351502 532338 351586 532574
rect 351822 532338 351854 532574
rect 351234 496894 351854 532338
rect 351234 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 351854 496894
rect 351234 496574 351854 496658
rect 351234 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 351854 496574
rect 351234 460894 351854 496338
rect 351234 460658 351266 460894
rect 351502 460658 351586 460894
rect 351822 460658 351854 460894
rect 351234 460574 351854 460658
rect 351234 460338 351266 460574
rect 351502 460338 351586 460574
rect 351822 460338 351854 460574
rect 351234 424894 351854 460338
rect 351234 424658 351266 424894
rect 351502 424658 351586 424894
rect 351822 424658 351854 424894
rect 351234 424574 351854 424658
rect 351234 424338 351266 424574
rect 351502 424338 351586 424574
rect 351822 424338 351854 424574
rect 351234 388894 351854 424338
rect 351234 388658 351266 388894
rect 351502 388658 351586 388894
rect 351822 388658 351854 388894
rect 351234 388574 351854 388658
rect 351234 388338 351266 388574
rect 351502 388338 351586 388574
rect 351822 388338 351854 388574
rect 351234 352894 351854 388338
rect 351234 352658 351266 352894
rect 351502 352658 351586 352894
rect 351822 352658 351854 352894
rect 351234 352574 351854 352658
rect 351234 352338 351266 352574
rect 351502 352338 351586 352574
rect 351822 352338 351854 352574
rect 351234 316894 351854 352338
rect 351234 316658 351266 316894
rect 351502 316658 351586 316894
rect 351822 316658 351854 316894
rect 351234 316574 351854 316658
rect 351234 316338 351266 316574
rect 351502 316338 351586 316574
rect 351822 316338 351854 316574
rect 351234 280894 351854 316338
rect 351234 280658 351266 280894
rect 351502 280658 351586 280894
rect 351822 280658 351854 280894
rect 351234 280574 351854 280658
rect 351234 280338 351266 280574
rect 351502 280338 351586 280574
rect 351822 280338 351854 280574
rect 351234 244894 351854 280338
rect 351234 244658 351266 244894
rect 351502 244658 351586 244894
rect 351822 244658 351854 244894
rect 351234 244574 351854 244658
rect 351234 244338 351266 244574
rect 351502 244338 351586 244574
rect 351822 244338 351854 244574
rect 351234 208894 351854 244338
rect 351234 208658 351266 208894
rect 351502 208658 351586 208894
rect 351822 208658 351854 208894
rect 351234 208574 351854 208658
rect 351234 208338 351266 208574
rect 351502 208338 351586 208574
rect 351822 208338 351854 208574
rect 351234 172894 351854 208338
rect 351234 172658 351266 172894
rect 351502 172658 351586 172894
rect 351822 172658 351854 172894
rect 351234 172574 351854 172658
rect 351234 172338 351266 172574
rect 351502 172338 351586 172574
rect 351822 172338 351854 172574
rect 351234 136894 351854 172338
rect 351234 136658 351266 136894
rect 351502 136658 351586 136894
rect 351822 136658 351854 136894
rect 351234 136574 351854 136658
rect 351234 136338 351266 136574
rect 351502 136338 351586 136574
rect 351822 136338 351854 136574
rect 351234 100894 351854 136338
rect 351234 100658 351266 100894
rect 351502 100658 351586 100894
rect 351822 100658 351854 100894
rect 351234 100574 351854 100658
rect 351234 100338 351266 100574
rect 351502 100338 351586 100574
rect 351822 100338 351854 100574
rect 351234 64894 351854 100338
rect 351234 64658 351266 64894
rect 351502 64658 351586 64894
rect 351822 64658 351854 64894
rect 351234 64574 351854 64658
rect 351234 64338 351266 64574
rect 351502 64338 351586 64574
rect 351822 64338 351854 64574
rect 351234 28894 351854 64338
rect 351234 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 351854 28894
rect 351234 28574 351854 28658
rect 351234 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 351854 28574
rect 351234 -5146 351854 28338
rect 351234 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 351854 -5146
rect 351234 -5466 351854 -5382
rect 351234 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 351854 -5466
rect 351234 -5734 351854 -5702
rect 354954 680614 355574 711002
rect 372954 710598 373574 711590
rect 372954 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 373574 710598
rect 372954 710278 373574 710362
rect 372954 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 373574 710278
rect 369234 708678 369854 709670
rect 369234 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 369854 708678
rect 369234 708358 369854 708442
rect 369234 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 369854 708358
rect 365514 706758 366134 707750
rect 365514 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 366134 706758
rect 365514 706438 366134 706522
rect 365514 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 366134 706438
rect 354954 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 355574 680614
rect 354954 680294 355574 680378
rect 354954 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 355574 680294
rect 354954 644614 355574 680058
rect 354954 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 355574 644614
rect 354954 644294 355574 644378
rect 354954 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 355574 644294
rect 354954 608614 355574 644058
rect 354954 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 355574 608614
rect 354954 608294 355574 608378
rect 354954 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 355574 608294
rect 354954 572614 355574 608058
rect 354954 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 355574 572614
rect 354954 572294 355574 572378
rect 354954 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 355574 572294
rect 354954 536614 355574 572058
rect 354954 536378 354986 536614
rect 355222 536378 355306 536614
rect 355542 536378 355574 536614
rect 354954 536294 355574 536378
rect 354954 536058 354986 536294
rect 355222 536058 355306 536294
rect 355542 536058 355574 536294
rect 354954 500614 355574 536058
rect 354954 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 355574 500614
rect 354954 500294 355574 500378
rect 354954 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 355574 500294
rect 354954 464614 355574 500058
rect 354954 464378 354986 464614
rect 355222 464378 355306 464614
rect 355542 464378 355574 464614
rect 354954 464294 355574 464378
rect 354954 464058 354986 464294
rect 355222 464058 355306 464294
rect 355542 464058 355574 464294
rect 354954 428614 355574 464058
rect 354954 428378 354986 428614
rect 355222 428378 355306 428614
rect 355542 428378 355574 428614
rect 354954 428294 355574 428378
rect 354954 428058 354986 428294
rect 355222 428058 355306 428294
rect 355542 428058 355574 428294
rect 354954 392614 355574 428058
rect 354954 392378 354986 392614
rect 355222 392378 355306 392614
rect 355542 392378 355574 392614
rect 354954 392294 355574 392378
rect 354954 392058 354986 392294
rect 355222 392058 355306 392294
rect 355542 392058 355574 392294
rect 354954 356614 355574 392058
rect 354954 356378 354986 356614
rect 355222 356378 355306 356614
rect 355542 356378 355574 356614
rect 354954 356294 355574 356378
rect 354954 356058 354986 356294
rect 355222 356058 355306 356294
rect 355542 356058 355574 356294
rect 354954 320614 355574 356058
rect 354954 320378 354986 320614
rect 355222 320378 355306 320614
rect 355542 320378 355574 320614
rect 354954 320294 355574 320378
rect 354954 320058 354986 320294
rect 355222 320058 355306 320294
rect 355542 320058 355574 320294
rect 354954 284614 355574 320058
rect 354954 284378 354986 284614
rect 355222 284378 355306 284614
rect 355542 284378 355574 284614
rect 354954 284294 355574 284378
rect 354954 284058 354986 284294
rect 355222 284058 355306 284294
rect 355542 284058 355574 284294
rect 354954 248614 355574 284058
rect 354954 248378 354986 248614
rect 355222 248378 355306 248614
rect 355542 248378 355574 248614
rect 354954 248294 355574 248378
rect 354954 248058 354986 248294
rect 355222 248058 355306 248294
rect 355542 248058 355574 248294
rect 354954 212614 355574 248058
rect 354954 212378 354986 212614
rect 355222 212378 355306 212614
rect 355542 212378 355574 212614
rect 354954 212294 355574 212378
rect 354954 212058 354986 212294
rect 355222 212058 355306 212294
rect 355542 212058 355574 212294
rect 354954 176614 355574 212058
rect 354954 176378 354986 176614
rect 355222 176378 355306 176614
rect 355542 176378 355574 176614
rect 354954 176294 355574 176378
rect 354954 176058 354986 176294
rect 355222 176058 355306 176294
rect 355542 176058 355574 176294
rect 354954 140614 355574 176058
rect 354954 140378 354986 140614
rect 355222 140378 355306 140614
rect 355542 140378 355574 140614
rect 354954 140294 355574 140378
rect 354954 140058 354986 140294
rect 355222 140058 355306 140294
rect 355542 140058 355574 140294
rect 354954 104614 355574 140058
rect 354954 104378 354986 104614
rect 355222 104378 355306 104614
rect 355542 104378 355574 104614
rect 354954 104294 355574 104378
rect 354954 104058 354986 104294
rect 355222 104058 355306 104294
rect 355542 104058 355574 104294
rect 354954 68614 355574 104058
rect 354954 68378 354986 68614
rect 355222 68378 355306 68614
rect 355542 68378 355574 68614
rect 354954 68294 355574 68378
rect 354954 68058 354986 68294
rect 355222 68058 355306 68294
rect 355542 68058 355574 68294
rect 354954 32614 355574 68058
rect 354954 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 355574 32614
rect 354954 32294 355574 32378
rect 354954 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 355574 32294
rect 336954 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 337574 -6106
rect 336954 -6426 337574 -6342
rect 336954 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 337574 -6426
rect 336954 -7654 337574 -6662
rect 354954 -7066 355574 32058
rect 361794 704838 362414 705830
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 435454 362414 470898
rect 361794 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 362414 435454
rect 361794 435134 362414 435218
rect 361794 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 362414 435134
rect 361794 399454 362414 434898
rect 361794 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 362414 399454
rect 361794 399134 362414 399218
rect 361794 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 362414 399134
rect 361794 363454 362414 398898
rect 361794 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 362414 363454
rect 361794 363134 362414 363218
rect 361794 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 362414 363134
rect 361794 327454 362414 362898
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 361794 291454 362414 326898
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 219454 362414 254898
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 361794 147454 362414 182898
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -1894 362414 -902
rect 365514 691174 366134 706202
rect 365514 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 366134 691174
rect 365514 690854 366134 690938
rect 365514 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 366134 690854
rect 365514 655174 366134 690618
rect 365514 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 366134 655174
rect 365514 654854 366134 654938
rect 365514 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 366134 654854
rect 365514 619174 366134 654618
rect 365514 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 366134 619174
rect 365514 618854 366134 618938
rect 365514 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 366134 618854
rect 365514 583174 366134 618618
rect 365514 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 366134 583174
rect 365514 582854 366134 582938
rect 365514 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 366134 582854
rect 365514 547174 366134 582618
rect 365514 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 366134 547174
rect 365514 546854 366134 546938
rect 365514 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 366134 546854
rect 365514 511174 366134 546618
rect 365514 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 366134 511174
rect 365514 510854 366134 510938
rect 365514 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 366134 510854
rect 365514 475174 366134 510618
rect 365514 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 366134 475174
rect 365514 474854 366134 474938
rect 365514 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 366134 474854
rect 365514 439174 366134 474618
rect 365514 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 366134 439174
rect 365514 438854 366134 438938
rect 365514 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 366134 438854
rect 365514 403174 366134 438618
rect 365514 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 366134 403174
rect 365514 402854 366134 402938
rect 365514 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 366134 402854
rect 365514 367174 366134 402618
rect 365514 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 366134 367174
rect 365514 366854 366134 366938
rect 365514 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 366134 366854
rect 365514 331174 366134 366618
rect 365514 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 366134 331174
rect 365514 330854 366134 330938
rect 365514 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 366134 330854
rect 365514 295174 366134 330618
rect 365514 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 366134 295174
rect 365514 294854 366134 294938
rect 365514 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 366134 294854
rect 365514 259174 366134 294618
rect 365514 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 366134 259174
rect 365514 258854 366134 258938
rect 365514 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 366134 258854
rect 365514 223174 366134 258618
rect 365514 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 366134 223174
rect 365514 222854 366134 222938
rect 365514 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 366134 222854
rect 365514 187174 366134 222618
rect 365514 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 366134 187174
rect 365514 186854 366134 186938
rect 365514 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 366134 186854
rect 365514 151174 366134 186618
rect 365514 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 366134 151174
rect 365514 150854 366134 150938
rect 365514 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 366134 150854
rect 365514 115174 366134 150618
rect 365514 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 366134 115174
rect 365514 114854 366134 114938
rect 365514 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 366134 114854
rect 365514 79174 366134 114618
rect 365514 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 366134 79174
rect 365514 78854 366134 78938
rect 365514 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 366134 78854
rect 365514 43174 366134 78618
rect 365514 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 366134 43174
rect 365514 42854 366134 42938
rect 365514 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 366134 42854
rect 365514 7174 366134 42618
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 365514 -2266 366134 6618
rect 365514 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 366134 -2266
rect 365514 -2586 366134 -2502
rect 365514 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 366134 -2586
rect 365514 -3814 366134 -2822
rect 369234 694894 369854 708122
rect 369234 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 369854 694894
rect 369234 694574 369854 694658
rect 369234 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 369854 694574
rect 369234 658894 369854 694338
rect 369234 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 369854 658894
rect 369234 658574 369854 658658
rect 369234 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 369854 658574
rect 369234 622894 369854 658338
rect 369234 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 369854 622894
rect 369234 622574 369854 622658
rect 369234 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 369854 622574
rect 369234 586894 369854 622338
rect 369234 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 369854 586894
rect 369234 586574 369854 586658
rect 369234 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 369854 586574
rect 369234 550894 369854 586338
rect 369234 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 369854 550894
rect 369234 550574 369854 550658
rect 369234 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 369854 550574
rect 369234 514894 369854 550338
rect 369234 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 369854 514894
rect 369234 514574 369854 514658
rect 369234 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 369854 514574
rect 369234 478894 369854 514338
rect 369234 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 369854 478894
rect 369234 478574 369854 478658
rect 369234 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 369854 478574
rect 369234 442894 369854 478338
rect 369234 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 369854 442894
rect 369234 442574 369854 442658
rect 369234 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 369854 442574
rect 369234 406894 369854 442338
rect 369234 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 369854 406894
rect 369234 406574 369854 406658
rect 369234 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 369854 406574
rect 369234 370894 369854 406338
rect 369234 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 369854 370894
rect 369234 370574 369854 370658
rect 369234 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 369854 370574
rect 369234 334894 369854 370338
rect 369234 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 369854 334894
rect 369234 334574 369854 334658
rect 369234 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 369854 334574
rect 369234 298894 369854 334338
rect 369234 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 369854 298894
rect 369234 298574 369854 298658
rect 369234 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 369854 298574
rect 369234 262894 369854 298338
rect 369234 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 369854 262894
rect 369234 262574 369854 262658
rect 369234 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 369854 262574
rect 369234 226894 369854 262338
rect 369234 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 369854 226894
rect 369234 226574 369854 226658
rect 369234 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 369854 226574
rect 369234 190894 369854 226338
rect 369234 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 369854 190894
rect 369234 190574 369854 190658
rect 369234 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 369854 190574
rect 369234 154894 369854 190338
rect 369234 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 369854 154894
rect 369234 154574 369854 154658
rect 369234 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 369854 154574
rect 369234 118894 369854 154338
rect 369234 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 369854 118894
rect 369234 118574 369854 118658
rect 369234 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 369854 118574
rect 369234 82894 369854 118338
rect 369234 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 369854 82894
rect 369234 82574 369854 82658
rect 369234 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 369854 82574
rect 369234 46894 369854 82338
rect 369234 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 369854 46894
rect 369234 46574 369854 46658
rect 369234 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 369854 46574
rect 369234 10894 369854 46338
rect 369234 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 369854 10894
rect 369234 10574 369854 10658
rect 369234 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 369854 10574
rect 369234 -4186 369854 10338
rect 369234 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 369854 -4186
rect 369234 -4506 369854 -4422
rect 369234 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 369854 -4506
rect 369234 -5734 369854 -4742
rect 372954 698614 373574 710042
rect 390954 711558 391574 711590
rect 390954 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 391574 711558
rect 390954 711238 391574 711322
rect 390954 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 391574 711238
rect 387234 709638 387854 709670
rect 387234 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 387854 709638
rect 387234 709318 387854 709402
rect 387234 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 387854 709318
rect 383514 707718 384134 707750
rect 383514 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 384134 707718
rect 383514 707398 384134 707482
rect 383514 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 384134 707398
rect 372954 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 373574 698614
rect 372954 698294 373574 698378
rect 372954 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 373574 698294
rect 372954 662614 373574 698058
rect 372954 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 373574 662614
rect 372954 662294 373574 662378
rect 372954 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 373574 662294
rect 372954 626614 373574 662058
rect 372954 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 373574 626614
rect 372954 626294 373574 626378
rect 372954 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 373574 626294
rect 372954 590614 373574 626058
rect 372954 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 373574 590614
rect 372954 590294 373574 590378
rect 372954 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 373574 590294
rect 372954 554614 373574 590058
rect 372954 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 373574 554614
rect 372954 554294 373574 554378
rect 372954 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 373574 554294
rect 372954 518614 373574 554058
rect 372954 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 373574 518614
rect 372954 518294 373574 518378
rect 372954 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 373574 518294
rect 372954 482614 373574 518058
rect 372954 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 373574 482614
rect 372954 482294 373574 482378
rect 372954 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 373574 482294
rect 372954 446614 373574 482058
rect 372954 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 373574 446614
rect 372954 446294 373574 446378
rect 372954 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 373574 446294
rect 372954 410614 373574 446058
rect 372954 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 373574 410614
rect 372954 410294 373574 410378
rect 372954 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 373574 410294
rect 372954 374614 373574 410058
rect 372954 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 373574 374614
rect 372954 374294 373574 374378
rect 372954 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 373574 374294
rect 372954 338614 373574 374058
rect 372954 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 373574 338614
rect 372954 338294 373574 338378
rect 372954 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 373574 338294
rect 372954 302614 373574 338058
rect 372954 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 373574 302614
rect 372954 302294 373574 302378
rect 372954 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 373574 302294
rect 372954 266614 373574 302058
rect 372954 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 373574 266614
rect 372954 266294 373574 266378
rect 372954 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 373574 266294
rect 372954 230614 373574 266058
rect 372954 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 373574 230614
rect 372954 230294 373574 230378
rect 372954 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 373574 230294
rect 372954 194614 373574 230058
rect 372954 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 373574 194614
rect 372954 194294 373574 194378
rect 372954 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 373574 194294
rect 372954 158614 373574 194058
rect 372954 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 373574 158614
rect 372954 158294 373574 158378
rect 372954 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 373574 158294
rect 372954 122614 373574 158058
rect 372954 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 373574 122614
rect 372954 122294 373574 122378
rect 372954 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 373574 122294
rect 372954 86614 373574 122058
rect 372954 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 373574 86614
rect 372954 86294 373574 86378
rect 372954 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 373574 86294
rect 372954 50614 373574 86058
rect 372954 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 373574 50614
rect 372954 50294 373574 50378
rect 372954 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 373574 50294
rect 372954 14614 373574 50058
rect 372954 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 373574 14614
rect 372954 14294 373574 14378
rect 372954 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 373574 14294
rect 354954 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 355574 -7066
rect 354954 -7386 355574 -7302
rect 354954 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 355574 -7386
rect 354954 -7654 355574 -7622
rect 372954 -6106 373574 14058
rect 379794 705798 380414 705830
rect 379794 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 380414 705798
rect 379794 705478 380414 705562
rect 379794 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 380414 705478
rect 379794 669454 380414 705242
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 561454 380414 596898
rect 379794 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 380414 561454
rect 379794 561134 380414 561218
rect 379794 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 380414 561134
rect 379794 525454 380414 560898
rect 379794 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 380414 525454
rect 379794 525134 380414 525218
rect 379794 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 380414 525134
rect 379794 489454 380414 524898
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 379794 489134 380414 489218
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 379794 453454 380414 488898
rect 379794 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 380414 453454
rect 379794 453134 380414 453218
rect 379794 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 380414 453134
rect 379794 417454 380414 452898
rect 379794 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 380414 417454
rect 379794 417134 380414 417218
rect 379794 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 380414 417134
rect 379794 381454 380414 416898
rect 379794 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 380414 381454
rect 379794 381134 380414 381218
rect 379794 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 380414 381134
rect 379794 345454 380414 380898
rect 379794 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 380414 345454
rect 379794 345134 380414 345218
rect 379794 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 380414 345134
rect 379794 309454 380414 344898
rect 379794 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 380414 309454
rect 379794 309134 380414 309218
rect 379794 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 380414 309134
rect 379794 273454 380414 308898
rect 379794 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 380414 273454
rect 379794 273134 380414 273218
rect 379794 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 380414 273134
rect 379794 237454 380414 272898
rect 379794 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 380414 237454
rect 379794 237134 380414 237218
rect 379794 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 380414 237134
rect 379794 201454 380414 236898
rect 379794 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 380414 201454
rect 379794 201134 380414 201218
rect 379794 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 380414 201134
rect 379794 165454 380414 200898
rect 379794 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 380414 165454
rect 379794 165134 380414 165218
rect 379794 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 380414 165134
rect 379794 129454 380414 164898
rect 379794 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 380414 129454
rect 379794 129134 380414 129218
rect 379794 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 380414 129134
rect 379794 93454 380414 128898
rect 379794 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 380414 93454
rect 379794 93134 380414 93218
rect 379794 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 380414 93134
rect 379794 57454 380414 92898
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -1306 380414 20898
rect 379794 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 380414 -1306
rect 379794 -1626 380414 -1542
rect 379794 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 380414 -1626
rect 379794 -1894 380414 -1862
rect 383514 673174 384134 707162
rect 383514 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 384134 673174
rect 383514 672854 384134 672938
rect 383514 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 384134 672854
rect 383514 637174 384134 672618
rect 383514 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 384134 637174
rect 383514 636854 384134 636938
rect 383514 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 384134 636854
rect 383514 601174 384134 636618
rect 383514 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 384134 601174
rect 383514 600854 384134 600938
rect 383514 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 384134 600854
rect 383514 565174 384134 600618
rect 383514 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 384134 565174
rect 383514 564854 384134 564938
rect 383514 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 384134 564854
rect 383514 529174 384134 564618
rect 383514 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 384134 529174
rect 383514 528854 384134 528938
rect 383514 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 384134 528854
rect 383514 493174 384134 528618
rect 383514 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 384134 493174
rect 383514 492854 384134 492938
rect 383514 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 384134 492854
rect 383514 457174 384134 492618
rect 383514 456938 383546 457174
rect 383782 456938 383866 457174
rect 384102 456938 384134 457174
rect 383514 456854 384134 456938
rect 383514 456618 383546 456854
rect 383782 456618 383866 456854
rect 384102 456618 384134 456854
rect 383514 421174 384134 456618
rect 383514 420938 383546 421174
rect 383782 420938 383866 421174
rect 384102 420938 384134 421174
rect 383514 420854 384134 420938
rect 383514 420618 383546 420854
rect 383782 420618 383866 420854
rect 384102 420618 384134 420854
rect 383514 385174 384134 420618
rect 383514 384938 383546 385174
rect 383782 384938 383866 385174
rect 384102 384938 384134 385174
rect 383514 384854 384134 384938
rect 383514 384618 383546 384854
rect 383782 384618 383866 384854
rect 384102 384618 384134 384854
rect 383514 349174 384134 384618
rect 383514 348938 383546 349174
rect 383782 348938 383866 349174
rect 384102 348938 384134 349174
rect 383514 348854 384134 348938
rect 383514 348618 383546 348854
rect 383782 348618 383866 348854
rect 384102 348618 384134 348854
rect 383514 313174 384134 348618
rect 383514 312938 383546 313174
rect 383782 312938 383866 313174
rect 384102 312938 384134 313174
rect 383514 312854 384134 312938
rect 383514 312618 383546 312854
rect 383782 312618 383866 312854
rect 384102 312618 384134 312854
rect 383514 277174 384134 312618
rect 383514 276938 383546 277174
rect 383782 276938 383866 277174
rect 384102 276938 384134 277174
rect 383514 276854 384134 276938
rect 383514 276618 383546 276854
rect 383782 276618 383866 276854
rect 384102 276618 384134 276854
rect 383514 241174 384134 276618
rect 383514 240938 383546 241174
rect 383782 240938 383866 241174
rect 384102 240938 384134 241174
rect 383514 240854 384134 240938
rect 383514 240618 383546 240854
rect 383782 240618 383866 240854
rect 384102 240618 384134 240854
rect 383514 205174 384134 240618
rect 383514 204938 383546 205174
rect 383782 204938 383866 205174
rect 384102 204938 384134 205174
rect 383514 204854 384134 204938
rect 383514 204618 383546 204854
rect 383782 204618 383866 204854
rect 384102 204618 384134 204854
rect 383514 169174 384134 204618
rect 383514 168938 383546 169174
rect 383782 168938 383866 169174
rect 384102 168938 384134 169174
rect 383514 168854 384134 168938
rect 383514 168618 383546 168854
rect 383782 168618 383866 168854
rect 384102 168618 384134 168854
rect 383514 133174 384134 168618
rect 383514 132938 383546 133174
rect 383782 132938 383866 133174
rect 384102 132938 384134 133174
rect 383514 132854 384134 132938
rect 383514 132618 383546 132854
rect 383782 132618 383866 132854
rect 384102 132618 384134 132854
rect 383514 97174 384134 132618
rect 383514 96938 383546 97174
rect 383782 96938 383866 97174
rect 384102 96938 384134 97174
rect 383514 96854 384134 96938
rect 383514 96618 383546 96854
rect 383782 96618 383866 96854
rect 384102 96618 384134 96854
rect 383514 61174 384134 96618
rect 383514 60938 383546 61174
rect 383782 60938 383866 61174
rect 384102 60938 384134 61174
rect 383514 60854 384134 60938
rect 383514 60618 383546 60854
rect 383782 60618 383866 60854
rect 384102 60618 384134 60854
rect 383514 25174 384134 60618
rect 383514 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 384134 25174
rect 383514 24854 384134 24938
rect 383514 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 384134 24854
rect 383514 -3226 384134 24618
rect 383514 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 384134 -3226
rect 383514 -3546 384134 -3462
rect 383514 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 384134 -3546
rect 383514 -3814 384134 -3782
rect 387234 676894 387854 709082
rect 387234 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 387854 676894
rect 387234 676574 387854 676658
rect 387234 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 387854 676574
rect 387234 640894 387854 676338
rect 387234 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 387854 640894
rect 387234 640574 387854 640658
rect 387234 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 387854 640574
rect 387234 604894 387854 640338
rect 387234 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 387854 604894
rect 387234 604574 387854 604658
rect 387234 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 387854 604574
rect 387234 568894 387854 604338
rect 387234 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 387854 568894
rect 387234 568574 387854 568658
rect 387234 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 387854 568574
rect 387234 532894 387854 568338
rect 387234 532658 387266 532894
rect 387502 532658 387586 532894
rect 387822 532658 387854 532894
rect 387234 532574 387854 532658
rect 387234 532338 387266 532574
rect 387502 532338 387586 532574
rect 387822 532338 387854 532574
rect 387234 496894 387854 532338
rect 387234 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 387854 496894
rect 387234 496574 387854 496658
rect 387234 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 387854 496574
rect 387234 460894 387854 496338
rect 387234 460658 387266 460894
rect 387502 460658 387586 460894
rect 387822 460658 387854 460894
rect 387234 460574 387854 460658
rect 387234 460338 387266 460574
rect 387502 460338 387586 460574
rect 387822 460338 387854 460574
rect 387234 424894 387854 460338
rect 387234 424658 387266 424894
rect 387502 424658 387586 424894
rect 387822 424658 387854 424894
rect 387234 424574 387854 424658
rect 387234 424338 387266 424574
rect 387502 424338 387586 424574
rect 387822 424338 387854 424574
rect 387234 388894 387854 424338
rect 387234 388658 387266 388894
rect 387502 388658 387586 388894
rect 387822 388658 387854 388894
rect 387234 388574 387854 388658
rect 387234 388338 387266 388574
rect 387502 388338 387586 388574
rect 387822 388338 387854 388574
rect 387234 352894 387854 388338
rect 387234 352658 387266 352894
rect 387502 352658 387586 352894
rect 387822 352658 387854 352894
rect 387234 352574 387854 352658
rect 387234 352338 387266 352574
rect 387502 352338 387586 352574
rect 387822 352338 387854 352574
rect 387234 316894 387854 352338
rect 387234 316658 387266 316894
rect 387502 316658 387586 316894
rect 387822 316658 387854 316894
rect 387234 316574 387854 316658
rect 387234 316338 387266 316574
rect 387502 316338 387586 316574
rect 387822 316338 387854 316574
rect 387234 280894 387854 316338
rect 387234 280658 387266 280894
rect 387502 280658 387586 280894
rect 387822 280658 387854 280894
rect 387234 280574 387854 280658
rect 387234 280338 387266 280574
rect 387502 280338 387586 280574
rect 387822 280338 387854 280574
rect 387234 244894 387854 280338
rect 387234 244658 387266 244894
rect 387502 244658 387586 244894
rect 387822 244658 387854 244894
rect 387234 244574 387854 244658
rect 387234 244338 387266 244574
rect 387502 244338 387586 244574
rect 387822 244338 387854 244574
rect 387234 208894 387854 244338
rect 387234 208658 387266 208894
rect 387502 208658 387586 208894
rect 387822 208658 387854 208894
rect 387234 208574 387854 208658
rect 387234 208338 387266 208574
rect 387502 208338 387586 208574
rect 387822 208338 387854 208574
rect 387234 172894 387854 208338
rect 387234 172658 387266 172894
rect 387502 172658 387586 172894
rect 387822 172658 387854 172894
rect 387234 172574 387854 172658
rect 387234 172338 387266 172574
rect 387502 172338 387586 172574
rect 387822 172338 387854 172574
rect 387234 136894 387854 172338
rect 387234 136658 387266 136894
rect 387502 136658 387586 136894
rect 387822 136658 387854 136894
rect 387234 136574 387854 136658
rect 387234 136338 387266 136574
rect 387502 136338 387586 136574
rect 387822 136338 387854 136574
rect 387234 100894 387854 136338
rect 387234 100658 387266 100894
rect 387502 100658 387586 100894
rect 387822 100658 387854 100894
rect 387234 100574 387854 100658
rect 387234 100338 387266 100574
rect 387502 100338 387586 100574
rect 387822 100338 387854 100574
rect 387234 64894 387854 100338
rect 387234 64658 387266 64894
rect 387502 64658 387586 64894
rect 387822 64658 387854 64894
rect 387234 64574 387854 64658
rect 387234 64338 387266 64574
rect 387502 64338 387586 64574
rect 387822 64338 387854 64574
rect 387234 28894 387854 64338
rect 387234 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 387854 28894
rect 387234 28574 387854 28658
rect 387234 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 387854 28574
rect 387234 -5146 387854 28338
rect 387234 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 387854 -5146
rect 387234 -5466 387854 -5382
rect 387234 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 387854 -5466
rect 387234 -5734 387854 -5702
rect 390954 680614 391574 711002
rect 408954 710598 409574 711590
rect 408954 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 409574 710598
rect 408954 710278 409574 710362
rect 408954 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 409574 710278
rect 405234 708678 405854 709670
rect 405234 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 405854 708678
rect 405234 708358 405854 708442
rect 405234 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 405854 708358
rect 401514 706758 402134 707750
rect 401514 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 402134 706758
rect 401514 706438 402134 706522
rect 401514 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 402134 706438
rect 390954 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 391574 680614
rect 390954 680294 391574 680378
rect 390954 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 391574 680294
rect 390954 644614 391574 680058
rect 390954 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 391574 644614
rect 390954 644294 391574 644378
rect 390954 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 391574 644294
rect 390954 608614 391574 644058
rect 390954 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 391574 608614
rect 390954 608294 391574 608378
rect 390954 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 391574 608294
rect 390954 572614 391574 608058
rect 390954 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 391574 572614
rect 390954 572294 391574 572378
rect 390954 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 391574 572294
rect 390954 536614 391574 572058
rect 390954 536378 390986 536614
rect 391222 536378 391306 536614
rect 391542 536378 391574 536614
rect 390954 536294 391574 536378
rect 390954 536058 390986 536294
rect 391222 536058 391306 536294
rect 391542 536058 391574 536294
rect 390954 500614 391574 536058
rect 390954 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 391574 500614
rect 390954 500294 391574 500378
rect 390954 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 391574 500294
rect 390954 464614 391574 500058
rect 390954 464378 390986 464614
rect 391222 464378 391306 464614
rect 391542 464378 391574 464614
rect 390954 464294 391574 464378
rect 390954 464058 390986 464294
rect 391222 464058 391306 464294
rect 391542 464058 391574 464294
rect 390954 428614 391574 464058
rect 390954 428378 390986 428614
rect 391222 428378 391306 428614
rect 391542 428378 391574 428614
rect 390954 428294 391574 428378
rect 390954 428058 390986 428294
rect 391222 428058 391306 428294
rect 391542 428058 391574 428294
rect 390954 392614 391574 428058
rect 390954 392378 390986 392614
rect 391222 392378 391306 392614
rect 391542 392378 391574 392614
rect 390954 392294 391574 392378
rect 390954 392058 390986 392294
rect 391222 392058 391306 392294
rect 391542 392058 391574 392294
rect 390954 356614 391574 392058
rect 390954 356378 390986 356614
rect 391222 356378 391306 356614
rect 391542 356378 391574 356614
rect 390954 356294 391574 356378
rect 390954 356058 390986 356294
rect 391222 356058 391306 356294
rect 391542 356058 391574 356294
rect 390954 320614 391574 356058
rect 390954 320378 390986 320614
rect 391222 320378 391306 320614
rect 391542 320378 391574 320614
rect 390954 320294 391574 320378
rect 390954 320058 390986 320294
rect 391222 320058 391306 320294
rect 391542 320058 391574 320294
rect 390954 284614 391574 320058
rect 390954 284378 390986 284614
rect 391222 284378 391306 284614
rect 391542 284378 391574 284614
rect 390954 284294 391574 284378
rect 390954 284058 390986 284294
rect 391222 284058 391306 284294
rect 391542 284058 391574 284294
rect 390954 248614 391574 284058
rect 390954 248378 390986 248614
rect 391222 248378 391306 248614
rect 391542 248378 391574 248614
rect 390954 248294 391574 248378
rect 390954 248058 390986 248294
rect 391222 248058 391306 248294
rect 391542 248058 391574 248294
rect 390954 212614 391574 248058
rect 390954 212378 390986 212614
rect 391222 212378 391306 212614
rect 391542 212378 391574 212614
rect 390954 212294 391574 212378
rect 390954 212058 390986 212294
rect 391222 212058 391306 212294
rect 391542 212058 391574 212294
rect 390954 176614 391574 212058
rect 390954 176378 390986 176614
rect 391222 176378 391306 176614
rect 391542 176378 391574 176614
rect 390954 176294 391574 176378
rect 390954 176058 390986 176294
rect 391222 176058 391306 176294
rect 391542 176058 391574 176294
rect 390954 140614 391574 176058
rect 390954 140378 390986 140614
rect 391222 140378 391306 140614
rect 391542 140378 391574 140614
rect 390954 140294 391574 140378
rect 390954 140058 390986 140294
rect 391222 140058 391306 140294
rect 391542 140058 391574 140294
rect 390954 104614 391574 140058
rect 390954 104378 390986 104614
rect 391222 104378 391306 104614
rect 391542 104378 391574 104614
rect 390954 104294 391574 104378
rect 390954 104058 390986 104294
rect 391222 104058 391306 104294
rect 391542 104058 391574 104294
rect 390954 68614 391574 104058
rect 390954 68378 390986 68614
rect 391222 68378 391306 68614
rect 391542 68378 391574 68614
rect 390954 68294 391574 68378
rect 390954 68058 390986 68294
rect 391222 68058 391306 68294
rect 391542 68058 391574 68294
rect 390954 32614 391574 68058
rect 390954 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 391574 32614
rect 390954 32294 391574 32378
rect 390954 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 391574 32294
rect 372954 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 373574 -6106
rect 372954 -6426 373574 -6342
rect 372954 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 373574 -6426
rect 372954 -7654 373574 -6662
rect 390954 -7066 391574 32058
rect 397794 704838 398414 705830
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 397794 363454 398414 398898
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 219454 398414 254898
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397794 147454 398414 182898
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -1894 398414 -902
rect 401514 691174 402134 706202
rect 401514 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 402134 691174
rect 401514 690854 402134 690938
rect 401514 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 402134 690854
rect 401514 655174 402134 690618
rect 401514 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 402134 655174
rect 401514 654854 402134 654938
rect 401514 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 402134 654854
rect 401514 619174 402134 654618
rect 401514 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 402134 619174
rect 401514 618854 402134 618938
rect 401514 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 402134 618854
rect 401514 583174 402134 618618
rect 401514 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 402134 583174
rect 401514 582854 402134 582938
rect 401514 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 402134 582854
rect 401514 547174 402134 582618
rect 401514 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 402134 547174
rect 401514 546854 402134 546938
rect 401514 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 402134 546854
rect 401514 511174 402134 546618
rect 401514 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 402134 511174
rect 401514 510854 402134 510938
rect 401514 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 402134 510854
rect 401514 475174 402134 510618
rect 401514 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 402134 475174
rect 401514 474854 402134 474938
rect 401514 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 402134 474854
rect 401514 439174 402134 474618
rect 401514 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 402134 439174
rect 401514 438854 402134 438938
rect 401514 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 402134 438854
rect 401514 403174 402134 438618
rect 401514 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 402134 403174
rect 401514 402854 402134 402938
rect 401514 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 402134 402854
rect 401514 367174 402134 402618
rect 401514 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 402134 367174
rect 401514 366854 402134 366938
rect 401514 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 402134 366854
rect 401514 331174 402134 366618
rect 401514 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 402134 331174
rect 401514 330854 402134 330938
rect 401514 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 402134 330854
rect 401514 295174 402134 330618
rect 401514 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 402134 295174
rect 401514 294854 402134 294938
rect 401514 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 402134 294854
rect 401514 259174 402134 294618
rect 401514 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 402134 259174
rect 401514 258854 402134 258938
rect 401514 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 402134 258854
rect 401514 223174 402134 258618
rect 401514 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 402134 223174
rect 401514 222854 402134 222938
rect 401514 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 402134 222854
rect 401514 187174 402134 222618
rect 401514 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 402134 187174
rect 401514 186854 402134 186938
rect 401514 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 402134 186854
rect 401514 151174 402134 186618
rect 401514 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 402134 151174
rect 401514 150854 402134 150938
rect 401514 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 402134 150854
rect 401514 115174 402134 150618
rect 401514 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 402134 115174
rect 401514 114854 402134 114938
rect 401514 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 402134 114854
rect 401514 79174 402134 114618
rect 401514 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 402134 79174
rect 401514 78854 402134 78938
rect 401514 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 402134 78854
rect 401514 43174 402134 78618
rect 401514 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 402134 43174
rect 401514 42854 402134 42938
rect 401514 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 402134 42854
rect 401514 7174 402134 42618
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 401514 -2266 402134 6618
rect 401514 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 402134 -2266
rect 401514 -2586 402134 -2502
rect 401514 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 402134 -2586
rect 401514 -3814 402134 -2822
rect 405234 694894 405854 708122
rect 405234 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 405854 694894
rect 405234 694574 405854 694658
rect 405234 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 405854 694574
rect 405234 658894 405854 694338
rect 405234 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 405854 658894
rect 405234 658574 405854 658658
rect 405234 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 405854 658574
rect 405234 622894 405854 658338
rect 405234 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 405854 622894
rect 405234 622574 405854 622658
rect 405234 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 405854 622574
rect 405234 586894 405854 622338
rect 405234 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 405854 586894
rect 405234 586574 405854 586658
rect 405234 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 405854 586574
rect 405234 550894 405854 586338
rect 405234 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 405854 550894
rect 405234 550574 405854 550658
rect 405234 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 405854 550574
rect 405234 514894 405854 550338
rect 405234 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 405854 514894
rect 405234 514574 405854 514658
rect 405234 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 405854 514574
rect 405234 478894 405854 514338
rect 405234 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 405854 478894
rect 405234 478574 405854 478658
rect 405234 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 405854 478574
rect 405234 442894 405854 478338
rect 405234 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 405854 442894
rect 405234 442574 405854 442658
rect 405234 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 405854 442574
rect 405234 406894 405854 442338
rect 405234 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 405854 406894
rect 405234 406574 405854 406658
rect 405234 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 405854 406574
rect 405234 370894 405854 406338
rect 405234 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 405854 370894
rect 405234 370574 405854 370658
rect 405234 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 405854 370574
rect 405234 334894 405854 370338
rect 405234 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 405854 334894
rect 405234 334574 405854 334658
rect 405234 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 405854 334574
rect 405234 298894 405854 334338
rect 405234 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 405854 298894
rect 405234 298574 405854 298658
rect 405234 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 405854 298574
rect 405234 262894 405854 298338
rect 405234 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 405854 262894
rect 405234 262574 405854 262658
rect 405234 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 405854 262574
rect 405234 226894 405854 262338
rect 405234 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 405854 226894
rect 405234 226574 405854 226658
rect 405234 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 405854 226574
rect 405234 190894 405854 226338
rect 405234 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 405854 190894
rect 405234 190574 405854 190658
rect 405234 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 405854 190574
rect 405234 154894 405854 190338
rect 405234 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 405854 154894
rect 405234 154574 405854 154658
rect 405234 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 405854 154574
rect 405234 118894 405854 154338
rect 405234 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 405854 118894
rect 405234 118574 405854 118658
rect 405234 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 405854 118574
rect 405234 82894 405854 118338
rect 405234 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 405854 82894
rect 405234 82574 405854 82658
rect 405234 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 405854 82574
rect 405234 46894 405854 82338
rect 405234 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 405854 46894
rect 405234 46574 405854 46658
rect 405234 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 405854 46574
rect 405234 10894 405854 46338
rect 405234 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 405854 10894
rect 405234 10574 405854 10658
rect 405234 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 405854 10574
rect 405234 -4186 405854 10338
rect 405234 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 405854 -4186
rect 405234 -4506 405854 -4422
rect 405234 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 405854 -4506
rect 405234 -5734 405854 -4742
rect 408954 698614 409574 710042
rect 426954 711558 427574 711590
rect 426954 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 427574 711558
rect 426954 711238 427574 711322
rect 426954 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 427574 711238
rect 423234 709638 423854 709670
rect 423234 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 423854 709638
rect 423234 709318 423854 709402
rect 423234 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 423854 709318
rect 419514 707718 420134 707750
rect 419514 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 420134 707718
rect 419514 707398 420134 707482
rect 419514 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 420134 707398
rect 408954 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 409574 698614
rect 408954 698294 409574 698378
rect 408954 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 409574 698294
rect 408954 662614 409574 698058
rect 408954 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 409574 662614
rect 408954 662294 409574 662378
rect 408954 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 409574 662294
rect 408954 626614 409574 662058
rect 408954 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 409574 626614
rect 408954 626294 409574 626378
rect 408954 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 409574 626294
rect 408954 590614 409574 626058
rect 408954 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 409574 590614
rect 408954 590294 409574 590378
rect 408954 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 409574 590294
rect 408954 554614 409574 590058
rect 408954 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 409574 554614
rect 408954 554294 409574 554378
rect 408954 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 409574 554294
rect 408954 518614 409574 554058
rect 408954 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 409574 518614
rect 408954 518294 409574 518378
rect 408954 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 409574 518294
rect 408954 482614 409574 518058
rect 408954 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 409574 482614
rect 408954 482294 409574 482378
rect 408954 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 409574 482294
rect 408954 446614 409574 482058
rect 408954 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 409574 446614
rect 408954 446294 409574 446378
rect 408954 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 409574 446294
rect 408954 410614 409574 446058
rect 408954 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 409574 410614
rect 408954 410294 409574 410378
rect 408954 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 409574 410294
rect 408954 374614 409574 410058
rect 408954 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 409574 374614
rect 408954 374294 409574 374378
rect 408954 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 409574 374294
rect 408954 338614 409574 374058
rect 408954 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 409574 338614
rect 408954 338294 409574 338378
rect 408954 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 409574 338294
rect 408954 302614 409574 338058
rect 408954 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 409574 302614
rect 408954 302294 409574 302378
rect 408954 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 409574 302294
rect 408954 266614 409574 302058
rect 408954 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 409574 266614
rect 408954 266294 409574 266378
rect 408954 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 409574 266294
rect 408954 230614 409574 266058
rect 408954 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 409574 230614
rect 408954 230294 409574 230378
rect 408954 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 409574 230294
rect 408954 194614 409574 230058
rect 408954 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 409574 194614
rect 408954 194294 409574 194378
rect 408954 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 409574 194294
rect 408954 158614 409574 194058
rect 408954 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 409574 158614
rect 408954 158294 409574 158378
rect 408954 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 409574 158294
rect 408954 122614 409574 158058
rect 408954 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 409574 122614
rect 408954 122294 409574 122378
rect 408954 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 409574 122294
rect 408954 86614 409574 122058
rect 408954 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 409574 86614
rect 408954 86294 409574 86378
rect 408954 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 409574 86294
rect 408954 50614 409574 86058
rect 408954 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 409574 50614
rect 408954 50294 409574 50378
rect 408954 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 409574 50294
rect 408954 14614 409574 50058
rect 408954 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 409574 14614
rect 408954 14294 409574 14378
rect 408954 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 409574 14294
rect 390954 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 391574 -7066
rect 390954 -7386 391574 -7302
rect 390954 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 391574 -7386
rect 390954 -7654 391574 -7622
rect 408954 -6106 409574 14058
rect 415794 705798 416414 705830
rect 415794 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 416414 705798
rect 415794 705478 416414 705562
rect 415794 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 416414 705478
rect 415794 669454 416414 705242
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 561454 416414 596898
rect 415794 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 416414 561454
rect 415794 561134 416414 561218
rect 415794 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 416414 561134
rect 415794 525454 416414 560898
rect 415794 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 416414 525454
rect 415794 525134 416414 525218
rect 415794 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 416414 525134
rect 415794 489454 416414 524898
rect 415794 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 416414 489454
rect 415794 489134 416414 489218
rect 415794 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 416414 489134
rect 415794 453454 416414 488898
rect 415794 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 416414 453454
rect 415794 453134 416414 453218
rect 415794 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 416414 453134
rect 415794 417454 416414 452898
rect 415794 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 416414 417454
rect 415794 417134 416414 417218
rect 415794 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 416414 417134
rect 415794 381454 416414 416898
rect 415794 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 416414 381454
rect 415794 381134 416414 381218
rect 415794 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 416414 381134
rect 415794 345454 416414 380898
rect 415794 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 416414 345454
rect 415794 345134 416414 345218
rect 415794 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 416414 345134
rect 415794 309454 416414 344898
rect 415794 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 416414 309454
rect 415794 309134 416414 309218
rect 415794 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 416414 309134
rect 415794 273454 416414 308898
rect 415794 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 416414 273454
rect 415794 273134 416414 273218
rect 415794 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 416414 273134
rect 415794 237454 416414 272898
rect 415794 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 416414 237454
rect 415794 237134 416414 237218
rect 415794 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 416414 237134
rect 415794 201454 416414 236898
rect 415794 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 416414 201454
rect 415794 201134 416414 201218
rect 415794 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 416414 201134
rect 415794 165454 416414 200898
rect 415794 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 416414 165454
rect 415794 165134 416414 165218
rect 415794 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 416414 165134
rect 415794 129454 416414 164898
rect 415794 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 416414 129454
rect 415794 129134 416414 129218
rect 415794 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 416414 129134
rect 415794 93454 416414 128898
rect 415794 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 416414 93454
rect 415794 93134 416414 93218
rect 415794 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 416414 93134
rect 415794 57454 416414 92898
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -1306 416414 20898
rect 415794 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 416414 -1306
rect 415794 -1626 416414 -1542
rect 415794 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 416414 -1626
rect 415794 -1894 416414 -1862
rect 419514 673174 420134 707162
rect 419514 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 420134 673174
rect 419514 672854 420134 672938
rect 419514 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 420134 672854
rect 419514 637174 420134 672618
rect 419514 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 420134 637174
rect 419514 636854 420134 636938
rect 419514 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 420134 636854
rect 419514 601174 420134 636618
rect 419514 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 420134 601174
rect 419514 600854 420134 600938
rect 419514 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 420134 600854
rect 419514 565174 420134 600618
rect 419514 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 420134 565174
rect 419514 564854 420134 564938
rect 419514 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 420134 564854
rect 419514 529174 420134 564618
rect 419514 528938 419546 529174
rect 419782 528938 419866 529174
rect 420102 528938 420134 529174
rect 419514 528854 420134 528938
rect 419514 528618 419546 528854
rect 419782 528618 419866 528854
rect 420102 528618 420134 528854
rect 419514 493174 420134 528618
rect 419514 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 420134 493174
rect 419514 492854 420134 492938
rect 419514 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 420134 492854
rect 419514 457174 420134 492618
rect 419514 456938 419546 457174
rect 419782 456938 419866 457174
rect 420102 456938 420134 457174
rect 419514 456854 420134 456938
rect 419514 456618 419546 456854
rect 419782 456618 419866 456854
rect 420102 456618 420134 456854
rect 419514 421174 420134 456618
rect 419514 420938 419546 421174
rect 419782 420938 419866 421174
rect 420102 420938 420134 421174
rect 419514 420854 420134 420938
rect 419514 420618 419546 420854
rect 419782 420618 419866 420854
rect 420102 420618 420134 420854
rect 419514 385174 420134 420618
rect 419514 384938 419546 385174
rect 419782 384938 419866 385174
rect 420102 384938 420134 385174
rect 419514 384854 420134 384938
rect 419514 384618 419546 384854
rect 419782 384618 419866 384854
rect 420102 384618 420134 384854
rect 419514 349174 420134 384618
rect 419514 348938 419546 349174
rect 419782 348938 419866 349174
rect 420102 348938 420134 349174
rect 419514 348854 420134 348938
rect 419514 348618 419546 348854
rect 419782 348618 419866 348854
rect 420102 348618 420134 348854
rect 419514 313174 420134 348618
rect 419514 312938 419546 313174
rect 419782 312938 419866 313174
rect 420102 312938 420134 313174
rect 419514 312854 420134 312938
rect 419514 312618 419546 312854
rect 419782 312618 419866 312854
rect 420102 312618 420134 312854
rect 419514 277174 420134 312618
rect 419514 276938 419546 277174
rect 419782 276938 419866 277174
rect 420102 276938 420134 277174
rect 419514 276854 420134 276938
rect 419514 276618 419546 276854
rect 419782 276618 419866 276854
rect 420102 276618 420134 276854
rect 419514 241174 420134 276618
rect 419514 240938 419546 241174
rect 419782 240938 419866 241174
rect 420102 240938 420134 241174
rect 419514 240854 420134 240938
rect 419514 240618 419546 240854
rect 419782 240618 419866 240854
rect 420102 240618 420134 240854
rect 419514 205174 420134 240618
rect 419514 204938 419546 205174
rect 419782 204938 419866 205174
rect 420102 204938 420134 205174
rect 419514 204854 420134 204938
rect 419514 204618 419546 204854
rect 419782 204618 419866 204854
rect 420102 204618 420134 204854
rect 419514 169174 420134 204618
rect 419514 168938 419546 169174
rect 419782 168938 419866 169174
rect 420102 168938 420134 169174
rect 419514 168854 420134 168938
rect 419514 168618 419546 168854
rect 419782 168618 419866 168854
rect 420102 168618 420134 168854
rect 419514 133174 420134 168618
rect 419514 132938 419546 133174
rect 419782 132938 419866 133174
rect 420102 132938 420134 133174
rect 419514 132854 420134 132938
rect 419514 132618 419546 132854
rect 419782 132618 419866 132854
rect 420102 132618 420134 132854
rect 419514 97174 420134 132618
rect 419514 96938 419546 97174
rect 419782 96938 419866 97174
rect 420102 96938 420134 97174
rect 419514 96854 420134 96938
rect 419514 96618 419546 96854
rect 419782 96618 419866 96854
rect 420102 96618 420134 96854
rect 419514 61174 420134 96618
rect 419514 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 420134 61174
rect 419514 60854 420134 60938
rect 419514 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 420134 60854
rect 419514 25174 420134 60618
rect 419514 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 420134 25174
rect 419514 24854 420134 24938
rect 419514 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 420134 24854
rect 419514 -3226 420134 24618
rect 419514 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 420134 -3226
rect 419514 -3546 420134 -3462
rect 419514 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 420134 -3546
rect 419514 -3814 420134 -3782
rect 423234 676894 423854 709082
rect 423234 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 423854 676894
rect 423234 676574 423854 676658
rect 423234 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 423854 676574
rect 423234 640894 423854 676338
rect 423234 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 423854 640894
rect 423234 640574 423854 640658
rect 423234 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 423854 640574
rect 423234 604894 423854 640338
rect 423234 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 423854 604894
rect 423234 604574 423854 604658
rect 423234 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 423854 604574
rect 423234 568894 423854 604338
rect 423234 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 423854 568894
rect 423234 568574 423854 568658
rect 423234 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 423854 568574
rect 423234 532894 423854 568338
rect 423234 532658 423266 532894
rect 423502 532658 423586 532894
rect 423822 532658 423854 532894
rect 423234 532574 423854 532658
rect 423234 532338 423266 532574
rect 423502 532338 423586 532574
rect 423822 532338 423854 532574
rect 423234 496894 423854 532338
rect 423234 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 423854 496894
rect 423234 496574 423854 496658
rect 423234 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 423854 496574
rect 423234 460894 423854 496338
rect 423234 460658 423266 460894
rect 423502 460658 423586 460894
rect 423822 460658 423854 460894
rect 423234 460574 423854 460658
rect 423234 460338 423266 460574
rect 423502 460338 423586 460574
rect 423822 460338 423854 460574
rect 423234 424894 423854 460338
rect 423234 424658 423266 424894
rect 423502 424658 423586 424894
rect 423822 424658 423854 424894
rect 423234 424574 423854 424658
rect 423234 424338 423266 424574
rect 423502 424338 423586 424574
rect 423822 424338 423854 424574
rect 423234 388894 423854 424338
rect 423234 388658 423266 388894
rect 423502 388658 423586 388894
rect 423822 388658 423854 388894
rect 423234 388574 423854 388658
rect 423234 388338 423266 388574
rect 423502 388338 423586 388574
rect 423822 388338 423854 388574
rect 423234 352894 423854 388338
rect 423234 352658 423266 352894
rect 423502 352658 423586 352894
rect 423822 352658 423854 352894
rect 423234 352574 423854 352658
rect 423234 352338 423266 352574
rect 423502 352338 423586 352574
rect 423822 352338 423854 352574
rect 423234 316894 423854 352338
rect 423234 316658 423266 316894
rect 423502 316658 423586 316894
rect 423822 316658 423854 316894
rect 423234 316574 423854 316658
rect 423234 316338 423266 316574
rect 423502 316338 423586 316574
rect 423822 316338 423854 316574
rect 423234 280894 423854 316338
rect 423234 280658 423266 280894
rect 423502 280658 423586 280894
rect 423822 280658 423854 280894
rect 423234 280574 423854 280658
rect 423234 280338 423266 280574
rect 423502 280338 423586 280574
rect 423822 280338 423854 280574
rect 423234 244894 423854 280338
rect 423234 244658 423266 244894
rect 423502 244658 423586 244894
rect 423822 244658 423854 244894
rect 423234 244574 423854 244658
rect 423234 244338 423266 244574
rect 423502 244338 423586 244574
rect 423822 244338 423854 244574
rect 423234 208894 423854 244338
rect 423234 208658 423266 208894
rect 423502 208658 423586 208894
rect 423822 208658 423854 208894
rect 423234 208574 423854 208658
rect 423234 208338 423266 208574
rect 423502 208338 423586 208574
rect 423822 208338 423854 208574
rect 423234 172894 423854 208338
rect 423234 172658 423266 172894
rect 423502 172658 423586 172894
rect 423822 172658 423854 172894
rect 423234 172574 423854 172658
rect 423234 172338 423266 172574
rect 423502 172338 423586 172574
rect 423822 172338 423854 172574
rect 423234 136894 423854 172338
rect 423234 136658 423266 136894
rect 423502 136658 423586 136894
rect 423822 136658 423854 136894
rect 423234 136574 423854 136658
rect 423234 136338 423266 136574
rect 423502 136338 423586 136574
rect 423822 136338 423854 136574
rect 423234 100894 423854 136338
rect 423234 100658 423266 100894
rect 423502 100658 423586 100894
rect 423822 100658 423854 100894
rect 423234 100574 423854 100658
rect 423234 100338 423266 100574
rect 423502 100338 423586 100574
rect 423822 100338 423854 100574
rect 423234 64894 423854 100338
rect 423234 64658 423266 64894
rect 423502 64658 423586 64894
rect 423822 64658 423854 64894
rect 423234 64574 423854 64658
rect 423234 64338 423266 64574
rect 423502 64338 423586 64574
rect 423822 64338 423854 64574
rect 423234 28894 423854 64338
rect 423234 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 423854 28894
rect 423234 28574 423854 28658
rect 423234 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 423854 28574
rect 423234 -5146 423854 28338
rect 423234 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 423854 -5146
rect 423234 -5466 423854 -5382
rect 423234 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 423854 -5466
rect 423234 -5734 423854 -5702
rect 426954 680614 427574 711002
rect 444954 710598 445574 711590
rect 444954 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 445574 710598
rect 444954 710278 445574 710362
rect 444954 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 445574 710278
rect 441234 708678 441854 709670
rect 441234 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 441854 708678
rect 441234 708358 441854 708442
rect 441234 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 441854 708358
rect 437514 706758 438134 707750
rect 437514 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 438134 706758
rect 437514 706438 438134 706522
rect 437514 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 438134 706438
rect 426954 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 427574 680614
rect 426954 680294 427574 680378
rect 426954 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 427574 680294
rect 426954 644614 427574 680058
rect 426954 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 427574 644614
rect 426954 644294 427574 644378
rect 426954 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 427574 644294
rect 426954 608614 427574 644058
rect 426954 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 427574 608614
rect 426954 608294 427574 608378
rect 426954 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 427574 608294
rect 426954 572614 427574 608058
rect 426954 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 427574 572614
rect 426954 572294 427574 572378
rect 426954 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 427574 572294
rect 426954 536614 427574 572058
rect 426954 536378 426986 536614
rect 427222 536378 427306 536614
rect 427542 536378 427574 536614
rect 426954 536294 427574 536378
rect 426954 536058 426986 536294
rect 427222 536058 427306 536294
rect 427542 536058 427574 536294
rect 426954 500614 427574 536058
rect 426954 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 427574 500614
rect 426954 500294 427574 500378
rect 426954 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 427574 500294
rect 426954 464614 427574 500058
rect 426954 464378 426986 464614
rect 427222 464378 427306 464614
rect 427542 464378 427574 464614
rect 426954 464294 427574 464378
rect 426954 464058 426986 464294
rect 427222 464058 427306 464294
rect 427542 464058 427574 464294
rect 426954 428614 427574 464058
rect 426954 428378 426986 428614
rect 427222 428378 427306 428614
rect 427542 428378 427574 428614
rect 426954 428294 427574 428378
rect 426954 428058 426986 428294
rect 427222 428058 427306 428294
rect 427542 428058 427574 428294
rect 426954 392614 427574 428058
rect 426954 392378 426986 392614
rect 427222 392378 427306 392614
rect 427542 392378 427574 392614
rect 426954 392294 427574 392378
rect 426954 392058 426986 392294
rect 427222 392058 427306 392294
rect 427542 392058 427574 392294
rect 426954 356614 427574 392058
rect 426954 356378 426986 356614
rect 427222 356378 427306 356614
rect 427542 356378 427574 356614
rect 426954 356294 427574 356378
rect 426954 356058 426986 356294
rect 427222 356058 427306 356294
rect 427542 356058 427574 356294
rect 426954 320614 427574 356058
rect 426954 320378 426986 320614
rect 427222 320378 427306 320614
rect 427542 320378 427574 320614
rect 426954 320294 427574 320378
rect 426954 320058 426986 320294
rect 427222 320058 427306 320294
rect 427542 320058 427574 320294
rect 426954 284614 427574 320058
rect 426954 284378 426986 284614
rect 427222 284378 427306 284614
rect 427542 284378 427574 284614
rect 426954 284294 427574 284378
rect 426954 284058 426986 284294
rect 427222 284058 427306 284294
rect 427542 284058 427574 284294
rect 426954 248614 427574 284058
rect 426954 248378 426986 248614
rect 427222 248378 427306 248614
rect 427542 248378 427574 248614
rect 426954 248294 427574 248378
rect 426954 248058 426986 248294
rect 427222 248058 427306 248294
rect 427542 248058 427574 248294
rect 426954 212614 427574 248058
rect 426954 212378 426986 212614
rect 427222 212378 427306 212614
rect 427542 212378 427574 212614
rect 426954 212294 427574 212378
rect 426954 212058 426986 212294
rect 427222 212058 427306 212294
rect 427542 212058 427574 212294
rect 426954 176614 427574 212058
rect 426954 176378 426986 176614
rect 427222 176378 427306 176614
rect 427542 176378 427574 176614
rect 426954 176294 427574 176378
rect 426954 176058 426986 176294
rect 427222 176058 427306 176294
rect 427542 176058 427574 176294
rect 426954 140614 427574 176058
rect 426954 140378 426986 140614
rect 427222 140378 427306 140614
rect 427542 140378 427574 140614
rect 426954 140294 427574 140378
rect 426954 140058 426986 140294
rect 427222 140058 427306 140294
rect 427542 140058 427574 140294
rect 426954 104614 427574 140058
rect 426954 104378 426986 104614
rect 427222 104378 427306 104614
rect 427542 104378 427574 104614
rect 426954 104294 427574 104378
rect 426954 104058 426986 104294
rect 427222 104058 427306 104294
rect 427542 104058 427574 104294
rect 426954 68614 427574 104058
rect 426954 68378 426986 68614
rect 427222 68378 427306 68614
rect 427542 68378 427574 68614
rect 426954 68294 427574 68378
rect 426954 68058 426986 68294
rect 427222 68058 427306 68294
rect 427542 68058 427574 68294
rect 426954 32614 427574 68058
rect 426954 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 427574 32614
rect 426954 32294 427574 32378
rect 426954 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 427574 32294
rect 408954 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 409574 -6106
rect 408954 -6426 409574 -6342
rect 408954 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 409574 -6426
rect 408954 -7654 409574 -6662
rect 426954 -7066 427574 32058
rect 433794 704838 434414 705830
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 435454 434414 470898
rect 433794 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 434414 435454
rect 433794 435134 434414 435218
rect 433794 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 434414 435134
rect 433794 399454 434414 434898
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 363454 434414 398898
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 433794 147454 434414 182898
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 111454 434414 146898
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -1894 434414 -902
rect 437514 691174 438134 706202
rect 437514 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 438134 691174
rect 437514 690854 438134 690938
rect 437514 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 438134 690854
rect 437514 655174 438134 690618
rect 437514 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 438134 655174
rect 437514 654854 438134 654938
rect 437514 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 438134 654854
rect 437514 619174 438134 654618
rect 437514 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 438134 619174
rect 437514 618854 438134 618938
rect 437514 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 438134 618854
rect 437514 583174 438134 618618
rect 437514 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 438134 583174
rect 437514 582854 438134 582938
rect 437514 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 438134 582854
rect 437514 547174 438134 582618
rect 437514 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 438134 547174
rect 437514 546854 438134 546938
rect 437514 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 438134 546854
rect 437514 511174 438134 546618
rect 437514 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 438134 511174
rect 437514 510854 438134 510938
rect 437514 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 438134 510854
rect 437514 475174 438134 510618
rect 437514 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 438134 475174
rect 437514 474854 438134 474938
rect 437514 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 438134 474854
rect 437514 439174 438134 474618
rect 437514 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 438134 439174
rect 437514 438854 438134 438938
rect 437514 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 438134 438854
rect 437514 403174 438134 438618
rect 437514 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 438134 403174
rect 437514 402854 438134 402938
rect 437514 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 438134 402854
rect 437514 367174 438134 402618
rect 437514 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 438134 367174
rect 437514 366854 438134 366938
rect 437514 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 438134 366854
rect 437514 331174 438134 366618
rect 437514 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 438134 331174
rect 437514 330854 438134 330938
rect 437514 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 438134 330854
rect 437514 295174 438134 330618
rect 437514 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 438134 295174
rect 437514 294854 438134 294938
rect 437514 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 438134 294854
rect 437514 259174 438134 294618
rect 437514 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 438134 259174
rect 437514 258854 438134 258938
rect 437514 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 438134 258854
rect 437514 223174 438134 258618
rect 437514 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 438134 223174
rect 437514 222854 438134 222938
rect 437514 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 438134 222854
rect 437514 187174 438134 222618
rect 437514 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 438134 187174
rect 437514 186854 438134 186938
rect 437514 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 438134 186854
rect 437514 151174 438134 186618
rect 437514 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 438134 151174
rect 437514 150854 438134 150938
rect 437514 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 438134 150854
rect 437514 115174 438134 150618
rect 437514 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 438134 115174
rect 437514 114854 438134 114938
rect 437514 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 438134 114854
rect 437514 79174 438134 114618
rect 437514 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 438134 79174
rect 437514 78854 438134 78938
rect 437514 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 438134 78854
rect 437514 43174 438134 78618
rect 437514 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 438134 43174
rect 437514 42854 438134 42938
rect 437514 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 438134 42854
rect 437514 7174 438134 42618
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -2266 438134 6618
rect 437514 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 438134 -2266
rect 437514 -2586 438134 -2502
rect 437514 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 438134 -2586
rect 437514 -3814 438134 -2822
rect 441234 694894 441854 708122
rect 441234 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 441854 694894
rect 441234 694574 441854 694658
rect 441234 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 441854 694574
rect 441234 658894 441854 694338
rect 441234 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 441854 658894
rect 441234 658574 441854 658658
rect 441234 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 441854 658574
rect 441234 622894 441854 658338
rect 441234 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 441854 622894
rect 441234 622574 441854 622658
rect 441234 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 441854 622574
rect 441234 586894 441854 622338
rect 441234 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 441854 586894
rect 441234 586574 441854 586658
rect 441234 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 441854 586574
rect 441234 550894 441854 586338
rect 441234 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 441854 550894
rect 441234 550574 441854 550658
rect 441234 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 441854 550574
rect 441234 514894 441854 550338
rect 441234 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 441854 514894
rect 441234 514574 441854 514658
rect 441234 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 441854 514574
rect 441234 478894 441854 514338
rect 441234 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 441854 478894
rect 441234 478574 441854 478658
rect 441234 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 441854 478574
rect 441234 442894 441854 478338
rect 441234 442658 441266 442894
rect 441502 442658 441586 442894
rect 441822 442658 441854 442894
rect 441234 442574 441854 442658
rect 441234 442338 441266 442574
rect 441502 442338 441586 442574
rect 441822 442338 441854 442574
rect 441234 406894 441854 442338
rect 441234 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 441854 406894
rect 441234 406574 441854 406658
rect 441234 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 441854 406574
rect 441234 370894 441854 406338
rect 441234 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 441854 370894
rect 441234 370574 441854 370658
rect 441234 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 441854 370574
rect 441234 334894 441854 370338
rect 441234 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 441854 334894
rect 441234 334574 441854 334658
rect 441234 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 441854 334574
rect 441234 298894 441854 334338
rect 441234 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 441854 298894
rect 441234 298574 441854 298658
rect 441234 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 441854 298574
rect 441234 262894 441854 298338
rect 441234 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 441854 262894
rect 441234 262574 441854 262658
rect 441234 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 441854 262574
rect 441234 226894 441854 262338
rect 441234 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 441854 226894
rect 441234 226574 441854 226658
rect 441234 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 441854 226574
rect 441234 190894 441854 226338
rect 441234 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 441854 190894
rect 441234 190574 441854 190658
rect 441234 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 441854 190574
rect 441234 154894 441854 190338
rect 441234 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 441854 154894
rect 441234 154574 441854 154658
rect 441234 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 441854 154574
rect 441234 118894 441854 154338
rect 441234 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 441854 118894
rect 441234 118574 441854 118658
rect 441234 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 441854 118574
rect 441234 82894 441854 118338
rect 441234 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 441854 82894
rect 441234 82574 441854 82658
rect 441234 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 441854 82574
rect 441234 46894 441854 82338
rect 441234 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 441854 46894
rect 441234 46574 441854 46658
rect 441234 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 441854 46574
rect 441234 10894 441854 46338
rect 441234 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 441854 10894
rect 441234 10574 441854 10658
rect 441234 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 441854 10574
rect 441234 -4186 441854 10338
rect 441234 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 441854 -4186
rect 441234 -4506 441854 -4422
rect 441234 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 441854 -4506
rect 441234 -5734 441854 -4742
rect 444954 698614 445574 710042
rect 462954 711558 463574 711590
rect 462954 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 463574 711558
rect 462954 711238 463574 711322
rect 462954 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 463574 711238
rect 459234 709638 459854 709670
rect 459234 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 459854 709638
rect 459234 709318 459854 709402
rect 459234 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 459854 709318
rect 455514 707718 456134 707750
rect 455514 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 456134 707718
rect 455514 707398 456134 707482
rect 455514 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 456134 707398
rect 444954 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 445574 698614
rect 444954 698294 445574 698378
rect 444954 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 445574 698294
rect 444954 662614 445574 698058
rect 444954 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 445574 662614
rect 444954 662294 445574 662378
rect 444954 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 445574 662294
rect 444954 626614 445574 662058
rect 444954 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 445574 626614
rect 444954 626294 445574 626378
rect 444954 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 445574 626294
rect 444954 590614 445574 626058
rect 444954 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 445574 590614
rect 444954 590294 445574 590378
rect 444954 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 445574 590294
rect 444954 554614 445574 590058
rect 444954 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 445574 554614
rect 444954 554294 445574 554378
rect 444954 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 445574 554294
rect 444954 518614 445574 554058
rect 444954 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 445574 518614
rect 444954 518294 445574 518378
rect 444954 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 445574 518294
rect 444954 482614 445574 518058
rect 444954 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 445574 482614
rect 444954 482294 445574 482378
rect 444954 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 445574 482294
rect 444954 446614 445574 482058
rect 444954 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 445574 446614
rect 444954 446294 445574 446378
rect 444954 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 445574 446294
rect 444954 410614 445574 446058
rect 444954 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 445574 410614
rect 444954 410294 445574 410378
rect 444954 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 445574 410294
rect 444954 374614 445574 410058
rect 444954 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 445574 374614
rect 444954 374294 445574 374378
rect 444954 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 445574 374294
rect 444954 338614 445574 374058
rect 444954 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 445574 338614
rect 444954 338294 445574 338378
rect 444954 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 445574 338294
rect 444954 302614 445574 338058
rect 444954 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 445574 302614
rect 444954 302294 445574 302378
rect 444954 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 445574 302294
rect 444954 266614 445574 302058
rect 444954 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 445574 266614
rect 444954 266294 445574 266378
rect 444954 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 445574 266294
rect 444954 230614 445574 266058
rect 444954 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 445574 230614
rect 444954 230294 445574 230378
rect 444954 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 445574 230294
rect 444954 194614 445574 230058
rect 444954 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 445574 194614
rect 444954 194294 445574 194378
rect 444954 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 445574 194294
rect 444954 158614 445574 194058
rect 444954 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 445574 158614
rect 444954 158294 445574 158378
rect 444954 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 445574 158294
rect 444954 122614 445574 158058
rect 444954 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 445574 122614
rect 444954 122294 445574 122378
rect 444954 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 445574 122294
rect 444954 86614 445574 122058
rect 444954 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 445574 86614
rect 444954 86294 445574 86378
rect 444954 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 445574 86294
rect 444954 50614 445574 86058
rect 444954 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 445574 50614
rect 444954 50294 445574 50378
rect 444954 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 445574 50294
rect 444954 14614 445574 50058
rect 444954 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 445574 14614
rect 444954 14294 445574 14378
rect 444954 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 445574 14294
rect 426954 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 427574 -7066
rect 426954 -7386 427574 -7302
rect 426954 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 427574 -7386
rect 426954 -7654 427574 -7622
rect 444954 -6106 445574 14058
rect 451794 705798 452414 705830
rect 451794 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 452414 705798
rect 451794 705478 452414 705562
rect 451794 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 452414 705478
rect 451794 669454 452414 705242
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 453454 452414 488898
rect 451794 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 452414 453454
rect 451794 453134 452414 453218
rect 451794 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 452414 453134
rect 451794 417454 452414 452898
rect 451794 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 452414 417454
rect 451794 417134 452414 417218
rect 451794 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 452414 417134
rect 451794 381454 452414 416898
rect 451794 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 452414 381454
rect 451794 381134 452414 381218
rect 451794 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 452414 381134
rect 451794 345454 452414 380898
rect 451794 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 452414 345454
rect 451794 345134 452414 345218
rect 451794 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 452414 345134
rect 451794 309454 452414 344898
rect 451794 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 452414 309454
rect 451794 309134 452414 309218
rect 451794 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 452414 309134
rect 451794 273454 452414 308898
rect 451794 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 452414 273454
rect 451794 273134 452414 273218
rect 451794 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 452414 273134
rect 451794 237454 452414 272898
rect 451794 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 452414 237454
rect 451794 237134 452414 237218
rect 451794 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 452414 237134
rect 451794 201454 452414 236898
rect 451794 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 452414 201454
rect 451794 201134 452414 201218
rect 451794 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 452414 201134
rect 451794 165454 452414 200898
rect 451794 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 452414 165454
rect 451794 165134 452414 165218
rect 451794 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 452414 165134
rect 451794 129454 452414 164898
rect 451794 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 452414 129454
rect 451794 129134 452414 129218
rect 451794 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 452414 129134
rect 451794 93454 452414 128898
rect 451794 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 452414 93454
rect 451794 93134 452414 93218
rect 451794 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 452414 93134
rect 451794 57454 452414 92898
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -1306 452414 20898
rect 451794 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 452414 -1306
rect 451794 -1626 452414 -1542
rect 451794 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 452414 -1626
rect 451794 -1894 452414 -1862
rect 455514 673174 456134 707162
rect 455514 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 456134 673174
rect 455514 672854 456134 672938
rect 455514 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 456134 672854
rect 455514 637174 456134 672618
rect 455514 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 456134 637174
rect 455514 636854 456134 636938
rect 455514 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 456134 636854
rect 455514 601174 456134 636618
rect 455514 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 456134 601174
rect 455514 600854 456134 600938
rect 455514 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 456134 600854
rect 455514 565174 456134 600618
rect 455514 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 456134 565174
rect 455514 564854 456134 564938
rect 455514 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 456134 564854
rect 455514 529174 456134 564618
rect 455514 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 456134 529174
rect 455514 528854 456134 528938
rect 455514 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 456134 528854
rect 455514 493174 456134 528618
rect 455514 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 456134 493174
rect 455514 492854 456134 492938
rect 455514 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 456134 492854
rect 455514 457174 456134 492618
rect 455514 456938 455546 457174
rect 455782 456938 455866 457174
rect 456102 456938 456134 457174
rect 455514 456854 456134 456938
rect 455514 456618 455546 456854
rect 455782 456618 455866 456854
rect 456102 456618 456134 456854
rect 455514 421174 456134 456618
rect 455514 420938 455546 421174
rect 455782 420938 455866 421174
rect 456102 420938 456134 421174
rect 455514 420854 456134 420938
rect 455514 420618 455546 420854
rect 455782 420618 455866 420854
rect 456102 420618 456134 420854
rect 455514 385174 456134 420618
rect 455514 384938 455546 385174
rect 455782 384938 455866 385174
rect 456102 384938 456134 385174
rect 455514 384854 456134 384938
rect 455514 384618 455546 384854
rect 455782 384618 455866 384854
rect 456102 384618 456134 384854
rect 455514 349174 456134 384618
rect 455514 348938 455546 349174
rect 455782 348938 455866 349174
rect 456102 348938 456134 349174
rect 455514 348854 456134 348938
rect 455514 348618 455546 348854
rect 455782 348618 455866 348854
rect 456102 348618 456134 348854
rect 455514 313174 456134 348618
rect 455514 312938 455546 313174
rect 455782 312938 455866 313174
rect 456102 312938 456134 313174
rect 455514 312854 456134 312938
rect 455514 312618 455546 312854
rect 455782 312618 455866 312854
rect 456102 312618 456134 312854
rect 455514 277174 456134 312618
rect 455514 276938 455546 277174
rect 455782 276938 455866 277174
rect 456102 276938 456134 277174
rect 455514 276854 456134 276938
rect 455514 276618 455546 276854
rect 455782 276618 455866 276854
rect 456102 276618 456134 276854
rect 455514 241174 456134 276618
rect 455514 240938 455546 241174
rect 455782 240938 455866 241174
rect 456102 240938 456134 241174
rect 455514 240854 456134 240938
rect 455514 240618 455546 240854
rect 455782 240618 455866 240854
rect 456102 240618 456134 240854
rect 455514 205174 456134 240618
rect 455514 204938 455546 205174
rect 455782 204938 455866 205174
rect 456102 204938 456134 205174
rect 455514 204854 456134 204938
rect 455514 204618 455546 204854
rect 455782 204618 455866 204854
rect 456102 204618 456134 204854
rect 455514 169174 456134 204618
rect 455514 168938 455546 169174
rect 455782 168938 455866 169174
rect 456102 168938 456134 169174
rect 455514 168854 456134 168938
rect 455514 168618 455546 168854
rect 455782 168618 455866 168854
rect 456102 168618 456134 168854
rect 455514 133174 456134 168618
rect 455514 132938 455546 133174
rect 455782 132938 455866 133174
rect 456102 132938 456134 133174
rect 455514 132854 456134 132938
rect 455514 132618 455546 132854
rect 455782 132618 455866 132854
rect 456102 132618 456134 132854
rect 455514 97174 456134 132618
rect 455514 96938 455546 97174
rect 455782 96938 455866 97174
rect 456102 96938 456134 97174
rect 455514 96854 456134 96938
rect 455514 96618 455546 96854
rect 455782 96618 455866 96854
rect 456102 96618 456134 96854
rect 455514 61174 456134 96618
rect 455514 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 456134 61174
rect 455514 60854 456134 60938
rect 455514 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 456134 60854
rect 455514 25174 456134 60618
rect 455514 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 456134 25174
rect 455514 24854 456134 24938
rect 455514 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 456134 24854
rect 455514 -3226 456134 24618
rect 455514 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 456134 -3226
rect 455514 -3546 456134 -3462
rect 455514 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 456134 -3546
rect 455514 -3814 456134 -3782
rect 459234 676894 459854 709082
rect 459234 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 459854 676894
rect 459234 676574 459854 676658
rect 459234 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 459854 676574
rect 459234 640894 459854 676338
rect 459234 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 459854 640894
rect 459234 640574 459854 640658
rect 459234 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 459854 640574
rect 459234 604894 459854 640338
rect 459234 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 459854 604894
rect 459234 604574 459854 604658
rect 459234 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 459854 604574
rect 459234 568894 459854 604338
rect 459234 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 459854 568894
rect 459234 568574 459854 568658
rect 459234 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 459854 568574
rect 459234 532894 459854 568338
rect 459234 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 459854 532894
rect 459234 532574 459854 532658
rect 459234 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 459854 532574
rect 459234 496894 459854 532338
rect 459234 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 459854 496894
rect 459234 496574 459854 496658
rect 459234 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 459854 496574
rect 459234 460894 459854 496338
rect 459234 460658 459266 460894
rect 459502 460658 459586 460894
rect 459822 460658 459854 460894
rect 459234 460574 459854 460658
rect 459234 460338 459266 460574
rect 459502 460338 459586 460574
rect 459822 460338 459854 460574
rect 459234 424894 459854 460338
rect 459234 424658 459266 424894
rect 459502 424658 459586 424894
rect 459822 424658 459854 424894
rect 459234 424574 459854 424658
rect 459234 424338 459266 424574
rect 459502 424338 459586 424574
rect 459822 424338 459854 424574
rect 459234 388894 459854 424338
rect 459234 388658 459266 388894
rect 459502 388658 459586 388894
rect 459822 388658 459854 388894
rect 459234 388574 459854 388658
rect 459234 388338 459266 388574
rect 459502 388338 459586 388574
rect 459822 388338 459854 388574
rect 459234 352894 459854 388338
rect 459234 352658 459266 352894
rect 459502 352658 459586 352894
rect 459822 352658 459854 352894
rect 459234 352574 459854 352658
rect 459234 352338 459266 352574
rect 459502 352338 459586 352574
rect 459822 352338 459854 352574
rect 459234 316894 459854 352338
rect 459234 316658 459266 316894
rect 459502 316658 459586 316894
rect 459822 316658 459854 316894
rect 459234 316574 459854 316658
rect 459234 316338 459266 316574
rect 459502 316338 459586 316574
rect 459822 316338 459854 316574
rect 459234 280894 459854 316338
rect 459234 280658 459266 280894
rect 459502 280658 459586 280894
rect 459822 280658 459854 280894
rect 459234 280574 459854 280658
rect 459234 280338 459266 280574
rect 459502 280338 459586 280574
rect 459822 280338 459854 280574
rect 459234 244894 459854 280338
rect 459234 244658 459266 244894
rect 459502 244658 459586 244894
rect 459822 244658 459854 244894
rect 459234 244574 459854 244658
rect 459234 244338 459266 244574
rect 459502 244338 459586 244574
rect 459822 244338 459854 244574
rect 459234 208894 459854 244338
rect 459234 208658 459266 208894
rect 459502 208658 459586 208894
rect 459822 208658 459854 208894
rect 459234 208574 459854 208658
rect 459234 208338 459266 208574
rect 459502 208338 459586 208574
rect 459822 208338 459854 208574
rect 459234 172894 459854 208338
rect 459234 172658 459266 172894
rect 459502 172658 459586 172894
rect 459822 172658 459854 172894
rect 459234 172574 459854 172658
rect 459234 172338 459266 172574
rect 459502 172338 459586 172574
rect 459822 172338 459854 172574
rect 459234 136894 459854 172338
rect 459234 136658 459266 136894
rect 459502 136658 459586 136894
rect 459822 136658 459854 136894
rect 459234 136574 459854 136658
rect 459234 136338 459266 136574
rect 459502 136338 459586 136574
rect 459822 136338 459854 136574
rect 459234 100894 459854 136338
rect 459234 100658 459266 100894
rect 459502 100658 459586 100894
rect 459822 100658 459854 100894
rect 459234 100574 459854 100658
rect 459234 100338 459266 100574
rect 459502 100338 459586 100574
rect 459822 100338 459854 100574
rect 459234 64894 459854 100338
rect 459234 64658 459266 64894
rect 459502 64658 459586 64894
rect 459822 64658 459854 64894
rect 459234 64574 459854 64658
rect 459234 64338 459266 64574
rect 459502 64338 459586 64574
rect 459822 64338 459854 64574
rect 459234 28894 459854 64338
rect 459234 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 459854 28894
rect 459234 28574 459854 28658
rect 459234 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 459854 28574
rect 459234 -5146 459854 28338
rect 459234 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 459854 -5146
rect 459234 -5466 459854 -5382
rect 459234 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 459854 -5466
rect 459234 -5734 459854 -5702
rect 462954 680614 463574 711002
rect 480954 710598 481574 711590
rect 480954 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 481574 710598
rect 480954 710278 481574 710362
rect 480954 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 481574 710278
rect 477234 708678 477854 709670
rect 477234 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 477854 708678
rect 477234 708358 477854 708442
rect 477234 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 477854 708358
rect 473514 706758 474134 707750
rect 473514 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 474134 706758
rect 473514 706438 474134 706522
rect 473514 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 474134 706438
rect 462954 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 463574 680614
rect 462954 680294 463574 680378
rect 462954 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 463574 680294
rect 462954 644614 463574 680058
rect 462954 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 463574 644614
rect 462954 644294 463574 644378
rect 462954 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 463574 644294
rect 462954 608614 463574 644058
rect 462954 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 463574 608614
rect 462954 608294 463574 608378
rect 462954 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 463574 608294
rect 462954 572614 463574 608058
rect 462954 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 463574 572614
rect 462954 572294 463574 572378
rect 462954 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 463574 572294
rect 462954 536614 463574 572058
rect 462954 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 463574 536614
rect 462954 536294 463574 536378
rect 462954 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 463574 536294
rect 462954 500614 463574 536058
rect 462954 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 463574 500614
rect 462954 500294 463574 500378
rect 462954 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 463574 500294
rect 462954 464614 463574 500058
rect 462954 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 463574 464614
rect 462954 464294 463574 464378
rect 462954 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 463574 464294
rect 462954 428614 463574 464058
rect 462954 428378 462986 428614
rect 463222 428378 463306 428614
rect 463542 428378 463574 428614
rect 462954 428294 463574 428378
rect 462954 428058 462986 428294
rect 463222 428058 463306 428294
rect 463542 428058 463574 428294
rect 462954 392614 463574 428058
rect 462954 392378 462986 392614
rect 463222 392378 463306 392614
rect 463542 392378 463574 392614
rect 462954 392294 463574 392378
rect 462954 392058 462986 392294
rect 463222 392058 463306 392294
rect 463542 392058 463574 392294
rect 462954 356614 463574 392058
rect 462954 356378 462986 356614
rect 463222 356378 463306 356614
rect 463542 356378 463574 356614
rect 462954 356294 463574 356378
rect 462954 356058 462986 356294
rect 463222 356058 463306 356294
rect 463542 356058 463574 356294
rect 462954 320614 463574 356058
rect 462954 320378 462986 320614
rect 463222 320378 463306 320614
rect 463542 320378 463574 320614
rect 462954 320294 463574 320378
rect 462954 320058 462986 320294
rect 463222 320058 463306 320294
rect 463542 320058 463574 320294
rect 462954 284614 463574 320058
rect 462954 284378 462986 284614
rect 463222 284378 463306 284614
rect 463542 284378 463574 284614
rect 462954 284294 463574 284378
rect 462954 284058 462986 284294
rect 463222 284058 463306 284294
rect 463542 284058 463574 284294
rect 462954 248614 463574 284058
rect 462954 248378 462986 248614
rect 463222 248378 463306 248614
rect 463542 248378 463574 248614
rect 462954 248294 463574 248378
rect 462954 248058 462986 248294
rect 463222 248058 463306 248294
rect 463542 248058 463574 248294
rect 462954 212614 463574 248058
rect 462954 212378 462986 212614
rect 463222 212378 463306 212614
rect 463542 212378 463574 212614
rect 462954 212294 463574 212378
rect 462954 212058 462986 212294
rect 463222 212058 463306 212294
rect 463542 212058 463574 212294
rect 462954 176614 463574 212058
rect 462954 176378 462986 176614
rect 463222 176378 463306 176614
rect 463542 176378 463574 176614
rect 462954 176294 463574 176378
rect 462954 176058 462986 176294
rect 463222 176058 463306 176294
rect 463542 176058 463574 176294
rect 462954 140614 463574 176058
rect 462954 140378 462986 140614
rect 463222 140378 463306 140614
rect 463542 140378 463574 140614
rect 462954 140294 463574 140378
rect 462954 140058 462986 140294
rect 463222 140058 463306 140294
rect 463542 140058 463574 140294
rect 462954 104614 463574 140058
rect 462954 104378 462986 104614
rect 463222 104378 463306 104614
rect 463542 104378 463574 104614
rect 462954 104294 463574 104378
rect 462954 104058 462986 104294
rect 463222 104058 463306 104294
rect 463542 104058 463574 104294
rect 462954 68614 463574 104058
rect 462954 68378 462986 68614
rect 463222 68378 463306 68614
rect 463542 68378 463574 68614
rect 462954 68294 463574 68378
rect 462954 68058 462986 68294
rect 463222 68058 463306 68294
rect 463542 68058 463574 68294
rect 462954 32614 463574 68058
rect 462954 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 463574 32614
rect 462954 32294 463574 32378
rect 462954 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 463574 32294
rect 444954 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 445574 -6106
rect 444954 -6426 445574 -6342
rect 444954 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 445574 -6426
rect 444954 -7654 445574 -6662
rect 462954 -7066 463574 32058
rect 469794 704838 470414 705830
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 363454 470414 398898
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 291454 470414 326898
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -1894 470414 -902
rect 473514 691174 474134 706202
rect 473514 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 474134 691174
rect 473514 690854 474134 690938
rect 473514 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 474134 690854
rect 473514 655174 474134 690618
rect 473514 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 474134 655174
rect 473514 654854 474134 654938
rect 473514 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 474134 654854
rect 473514 619174 474134 654618
rect 473514 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 474134 619174
rect 473514 618854 474134 618938
rect 473514 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 474134 618854
rect 473514 583174 474134 618618
rect 473514 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 474134 583174
rect 473514 582854 474134 582938
rect 473514 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 474134 582854
rect 473514 547174 474134 582618
rect 473514 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 474134 547174
rect 473514 546854 474134 546938
rect 473514 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 474134 546854
rect 473514 511174 474134 546618
rect 473514 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 474134 511174
rect 473514 510854 474134 510938
rect 473514 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 474134 510854
rect 473514 475174 474134 510618
rect 473514 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 474134 475174
rect 473514 474854 474134 474938
rect 473514 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 474134 474854
rect 473514 439174 474134 474618
rect 473514 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 474134 439174
rect 473514 438854 474134 438938
rect 473514 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 474134 438854
rect 473514 403174 474134 438618
rect 473514 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 474134 403174
rect 473514 402854 474134 402938
rect 473514 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 474134 402854
rect 473514 367174 474134 402618
rect 473514 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 474134 367174
rect 473514 366854 474134 366938
rect 473514 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 474134 366854
rect 473514 331174 474134 366618
rect 473514 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 474134 331174
rect 473514 330854 474134 330938
rect 473514 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 474134 330854
rect 473514 295174 474134 330618
rect 473514 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 474134 295174
rect 473514 294854 474134 294938
rect 473514 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 474134 294854
rect 473514 259174 474134 294618
rect 473514 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 474134 259174
rect 473514 258854 474134 258938
rect 473514 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 474134 258854
rect 473514 223174 474134 258618
rect 473514 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 474134 223174
rect 473514 222854 474134 222938
rect 473514 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 474134 222854
rect 473514 187174 474134 222618
rect 473514 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 474134 187174
rect 473514 186854 474134 186938
rect 473514 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 474134 186854
rect 473514 151174 474134 186618
rect 473514 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 474134 151174
rect 473514 150854 474134 150938
rect 473514 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 474134 150854
rect 473514 115174 474134 150618
rect 473514 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 474134 115174
rect 473514 114854 474134 114938
rect 473514 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 474134 114854
rect 473514 79174 474134 114618
rect 473514 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 474134 79174
rect 473514 78854 474134 78938
rect 473514 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 474134 78854
rect 473514 43174 474134 78618
rect 473514 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 474134 43174
rect 473514 42854 474134 42938
rect 473514 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 474134 42854
rect 473514 7174 474134 42618
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -2266 474134 6618
rect 473514 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 474134 -2266
rect 473514 -2586 474134 -2502
rect 473514 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 474134 -2586
rect 473514 -3814 474134 -2822
rect 477234 694894 477854 708122
rect 477234 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 477854 694894
rect 477234 694574 477854 694658
rect 477234 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 477854 694574
rect 477234 658894 477854 694338
rect 477234 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 477854 658894
rect 477234 658574 477854 658658
rect 477234 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 477854 658574
rect 477234 622894 477854 658338
rect 477234 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 477854 622894
rect 477234 622574 477854 622658
rect 477234 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 477854 622574
rect 477234 586894 477854 622338
rect 477234 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 477854 586894
rect 477234 586574 477854 586658
rect 477234 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 477854 586574
rect 477234 550894 477854 586338
rect 477234 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 477854 550894
rect 477234 550574 477854 550658
rect 477234 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 477854 550574
rect 477234 514894 477854 550338
rect 477234 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 477854 514894
rect 477234 514574 477854 514658
rect 477234 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 477854 514574
rect 477234 478894 477854 514338
rect 477234 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 477854 478894
rect 477234 478574 477854 478658
rect 477234 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 477854 478574
rect 477234 442894 477854 478338
rect 477234 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 477854 442894
rect 477234 442574 477854 442658
rect 477234 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 477854 442574
rect 477234 406894 477854 442338
rect 477234 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 477854 406894
rect 477234 406574 477854 406658
rect 477234 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 477854 406574
rect 477234 370894 477854 406338
rect 477234 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 477854 370894
rect 477234 370574 477854 370658
rect 477234 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 477854 370574
rect 477234 334894 477854 370338
rect 477234 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 477854 334894
rect 477234 334574 477854 334658
rect 477234 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 477854 334574
rect 477234 298894 477854 334338
rect 477234 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 477854 298894
rect 477234 298574 477854 298658
rect 477234 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 477854 298574
rect 477234 262894 477854 298338
rect 477234 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 477854 262894
rect 477234 262574 477854 262658
rect 477234 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 477854 262574
rect 477234 226894 477854 262338
rect 477234 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 477854 226894
rect 477234 226574 477854 226658
rect 477234 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 477854 226574
rect 477234 190894 477854 226338
rect 477234 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 477854 190894
rect 477234 190574 477854 190658
rect 477234 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 477854 190574
rect 477234 154894 477854 190338
rect 477234 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 477854 154894
rect 477234 154574 477854 154658
rect 477234 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 477854 154574
rect 477234 118894 477854 154338
rect 477234 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 477854 118894
rect 477234 118574 477854 118658
rect 477234 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 477854 118574
rect 477234 82894 477854 118338
rect 477234 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 477854 82894
rect 477234 82574 477854 82658
rect 477234 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 477854 82574
rect 477234 46894 477854 82338
rect 477234 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 477854 46894
rect 477234 46574 477854 46658
rect 477234 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 477854 46574
rect 477234 10894 477854 46338
rect 477234 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 477854 10894
rect 477234 10574 477854 10658
rect 477234 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 477854 10574
rect 477234 -4186 477854 10338
rect 477234 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 477854 -4186
rect 477234 -4506 477854 -4422
rect 477234 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 477854 -4506
rect 477234 -5734 477854 -4742
rect 480954 698614 481574 710042
rect 498954 711558 499574 711590
rect 498954 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 499574 711558
rect 498954 711238 499574 711322
rect 498954 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 499574 711238
rect 495234 709638 495854 709670
rect 495234 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 495854 709638
rect 495234 709318 495854 709402
rect 495234 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 495854 709318
rect 491514 707718 492134 707750
rect 491514 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 492134 707718
rect 491514 707398 492134 707482
rect 491514 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 492134 707398
rect 480954 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 481574 698614
rect 480954 698294 481574 698378
rect 480954 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 481574 698294
rect 480954 662614 481574 698058
rect 480954 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 481574 662614
rect 480954 662294 481574 662378
rect 480954 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 481574 662294
rect 480954 626614 481574 662058
rect 480954 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 481574 626614
rect 480954 626294 481574 626378
rect 480954 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 481574 626294
rect 480954 590614 481574 626058
rect 480954 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 481574 590614
rect 480954 590294 481574 590378
rect 480954 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 481574 590294
rect 480954 554614 481574 590058
rect 480954 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 481574 554614
rect 480954 554294 481574 554378
rect 480954 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 481574 554294
rect 480954 518614 481574 554058
rect 480954 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 481574 518614
rect 480954 518294 481574 518378
rect 480954 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 481574 518294
rect 480954 482614 481574 518058
rect 480954 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 481574 482614
rect 480954 482294 481574 482378
rect 480954 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 481574 482294
rect 480954 446614 481574 482058
rect 480954 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 481574 446614
rect 480954 446294 481574 446378
rect 480954 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 481574 446294
rect 480954 410614 481574 446058
rect 480954 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 481574 410614
rect 480954 410294 481574 410378
rect 480954 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 481574 410294
rect 480954 374614 481574 410058
rect 480954 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 481574 374614
rect 480954 374294 481574 374378
rect 480954 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 481574 374294
rect 480954 338614 481574 374058
rect 480954 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 481574 338614
rect 480954 338294 481574 338378
rect 480954 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 481574 338294
rect 480954 302614 481574 338058
rect 480954 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 481574 302614
rect 480954 302294 481574 302378
rect 480954 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 481574 302294
rect 480954 266614 481574 302058
rect 480954 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 481574 266614
rect 480954 266294 481574 266378
rect 480954 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 481574 266294
rect 480954 230614 481574 266058
rect 480954 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 481574 230614
rect 480954 230294 481574 230378
rect 480954 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 481574 230294
rect 480954 194614 481574 230058
rect 480954 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 481574 194614
rect 480954 194294 481574 194378
rect 480954 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 481574 194294
rect 480954 158614 481574 194058
rect 480954 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 481574 158614
rect 480954 158294 481574 158378
rect 480954 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 481574 158294
rect 480954 122614 481574 158058
rect 480954 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 481574 122614
rect 480954 122294 481574 122378
rect 480954 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 481574 122294
rect 480954 86614 481574 122058
rect 480954 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 481574 86614
rect 480954 86294 481574 86378
rect 480954 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 481574 86294
rect 480954 50614 481574 86058
rect 480954 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 481574 50614
rect 480954 50294 481574 50378
rect 480954 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 481574 50294
rect 480954 14614 481574 50058
rect 480954 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 481574 14614
rect 480954 14294 481574 14378
rect 480954 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 481574 14294
rect 462954 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 463574 -7066
rect 462954 -7386 463574 -7302
rect 462954 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 463574 -7386
rect 462954 -7654 463574 -7622
rect 480954 -6106 481574 14058
rect 487794 705798 488414 705830
rect 487794 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 488414 705798
rect 487794 705478 488414 705562
rect 487794 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 488414 705478
rect 487794 669454 488414 705242
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597454 488414 632898
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 561454 488414 596898
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 453454 488414 488898
rect 487794 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 488414 453454
rect 487794 453134 488414 453218
rect 487794 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 488414 453134
rect 487794 417454 488414 452898
rect 487794 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 488414 417454
rect 487794 417134 488414 417218
rect 487794 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 488414 417134
rect 487794 381454 488414 416898
rect 487794 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 488414 381454
rect 487794 381134 488414 381218
rect 487794 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 488414 381134
rect 487794 345454 488414 380898
rect 487794 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 488414 345454
rect 487794 345134 488414 345218
rect 487794 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 488414 345134
rect 487794 309454 488414 344898
rect 487794 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 488414 309454
rect 487794 309134 488414 309218
rect 487794 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 488414 309134
rect 487794 273454 488414 308898
rect 487794 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 488414 273454
rect 487794 273134 488414 273218
rect 487794 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 488414 273134
rect 487794 237454 488414 272898
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 487794 201454 488414 236898
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 165454 488414 200898
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 129454 488414 164898
rect 487794 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 488414 129454
rect 487794 129134 488414 129218
rect 487794 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 488414 129134
rect 487794 93454 488414 128898
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -1306 488414 20898
rect 487794 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 488414 -1306
rect 487794 -1626 488414 -1542
rect 487794 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 488414 -1626
rect 487794 -1894 488414 -1862
rect 491514 673174 492134 707162
rect 491514 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 492134 673174
rect 491514 672854 492134 672938
rect 491514 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 492134 672854
rect 491514 637174 492134 672618
rect 491514 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 492134 637174
rect 491514 636854 492134 636938
rect 491514 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 492134 636854
rect 491514 601174 492134 636618
rect 491514 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 492134 601174
rect 491514 600854 492134 600938
rect 491514 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 492134 600854
rect 491514 565174 492134 600618
rect 491514 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 492134 565174
rect 491514 564854 492134 564938
rect 491514 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 492134 564854
rect 491514 529174 492134 564618
rect 491514 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 492134 529174
rect 491514 528854 492134 528938
rect 491514 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 492134 528854
rect 491514 493174 492134 528618
rect 491514 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 492134 493174
rect 491514 492854 492134 492938
rect 491514 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 492134 492854
rect 491514 457174 492134 492618
rect 491514 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 492134 457174
rect 491514 456854 492134 456938
rect 491514 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 492134 456854
rect 491514 421174 492134 456618
rect 491514 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 492134 421174
rect 491514 420854 492134 420938
rect 491514 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 492134 420854
rect 491514 385174 492134 420618
rect 491514 384938 491546 385174
rect 491782 384938 491866 385174
rect 492102 384938 492134 385174
rect 491514 384854 492134 384938
rect 491514 384618 491546 384854
rect 491782 384618 491866 384854
rect 492102 384618 492134 384854
rect 491514 349174 492134 384618
rect 491514 348938 491546 349174
rect 491782 348938 491866 349174
rect 492102 348938 492134 349174
rect 491514 348854 492134 348938
rect 491514 348618 491546 348854
rect 491782 348618 491866 348854
rect 492102 348618 492134 348854
rect 491514 313174 492134 348618
rect 491514 312938 491546 313174
rect 491782 312938 491866 313174
rect 492102 312938 492134 313174
rect 491514 312854 492134 312938
rect 491514 312618 491546 312854
rect 491782 312618 491866 312854
rect 492102 312618 492134 312854
rect 491514 277174 492134 312618
rect 491514 276938 491546 277174
rect 491782 276938 491866 277174
rect 492102 276938 492134 277174
rect 491514 276854 492134 276938
rect 491514 276618 491546 276854
rect 491782 276618 491866 276854
rect 492102 276618 492134 276854
rect 491514 241174 492134 276618
rect 491514 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 492134 241174
rect 491514 240854 492134 240938
rect 491514 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 492134 240854
rect 491514 205174 492134 240618
rect 491514 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 492134 205174
rect 491514 204854 492134 204938
rect 491514 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 492134 204854
rect 491514 169174 492134 204618
rect 491514 168938 491546 169174
rect 491782 168938 491866 169174
rect 492102 168938 492134 169174
rect 491514 168854 492134 168938
rect 491514 168618 491546 168854
rect 491782 168618 491866 168854
rect 492102 168618 492134 168854
rect 491514 133174 492134 168618
rect 491514 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 492134 133174
rect 491514 132854 492134 132938
rect 491514 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 492134 132854
rect 491514 97174 492134 132618
rect 491514 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 492134 97174
rect 491514 96854 492134 96938
rect 491514 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 492134 96854
rect 491514 61174 492134 96618
rect 491514 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 492134 61174
rect 491514 60854 492134 60938
rect 491514 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 492134 60854
rect 491514 25174 492134 60618
rect 491514 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 492134 25174
rect 491514 24854 492134 24938
rect 491514 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 492134 24854
rect 491514 -3226 492134 24618
rect 491514 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 492134 -3226
rect 491514 -3546 492134 -3462
rect 491514 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 492134 -3546
rect 491514 -3814 492134 -3782
rect 495234 676894 495854 709082
rect 495234 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 495854 676894
rect 495234 676574 495854 676658
rect 495234 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 495854 676574
rect 495234 640894 495854 676338
rect 495234 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 495854 640894
rect 495234 640574 495854 640658
rect 495234 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 495854 640574
rect 495234 604894 495854 640338
rect 495234 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 495854 604894
rect 495234 604574 495854 604658
rect 495234 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 495854 604574
rect 495234 568894 495854 604338
rect 495234 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 495854 568894
rect 495234 568574 495854 568658
rect 495234 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 495854 568574
rect 495234 532894 495854 568338
rect 495234 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 495854 532894
rect 495234 532574 495854 532658
rect 495234 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 495854 532574
rect 495234 496894 495854 532338
rect 495234 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 495854 496894
rect 495234 496574 495854 496658
rect 495234 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 495854 496574
rect 495234 460894 495854 496338
rect 495234 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 495854 460894
rect 495234 460574 495854 460658
rect 495234 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 495854 460574
rect 495234 424894 495854 460338
rect 495234 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 495854 424894
rect 495234 424574 495854 424658
rect 495234 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 495854 424574
rect 495234 388894 495854 424338
rect 495234 388658 495266 388894
rect 495502 388658 495586 388894
rect 495822 388658 495854 388894
rect 495234 388574 495854 388658
rect 495234 388338 495266 388574
rect 495502 388338 495586 388574
rect 495822 388338 495854 388574
rect 495234 352894 495854 388338
rect 495234 352658 495266 352894
rect 495502 352658 495586 352894
rect 495822 352658 495854 352894
rect 495234 352574 495854 352658
rect 495234 352338 495266 352574
rect 495502 352338 495586 352574
rect 495822 352338 495854 352574
rect 495234 316894 495854 352338
rect 495234 316658 495266 316894
rect 495502 316658 495586 316894
rect 495822 316658 495854 316894
rect 495234 316574 495854 316658
rect 495234 316338 495266 316574
rect 495502 316338 495586 316574
rect 495822 316338 495854 316574
rect 495234 280894 495854 316338
rect 495234 280658 495266 280894
rect 495502 280658 495586 280894
rect 495822 280658 495854 280894
rect 495234 280574 495854 280658
rect 495234 280338 495266 280574
rect 495502 280338 495586 280574
rect 495822 280338 495854 280574
rect 495234 244894 495854 280338
rect 495234 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 495854 244894
rect 495234 244574 495854 244658
rect 495234 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 495854 244574
rect 495234 208894 495854 244338
rect 495234 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 495854 208894
rect 495234 208574 495854 208658
rect 495234 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 495854 208574
rect 495234 172894 495854 208338
rect 495234 172658 495266 172894
rect 495502 172658 495586 172894
rect 495822 172658 495854 172894
rect 495234 172574 495854 172658
rect 495234 172338 495266 172574
rect 495502 172338 495586 172574
rect 495822 172338 495854 172574
rect 495234 136894 495854 172338
rect 495234 136658 495266 136894
rect 495502 136658 495586 136894
rect 495822 136658 495854 136894
rect 495234 136574 495854 136658
rect 495234 136338 495266 136574
rect 495502 136338 495586 136574
rect 495822 136338 495854 136574
rect 495234 100894 495854 136338
rect 495234 100658 495266 100894
rect 495502 100658 495586 100894
rect 495822 100658 495854 100894
rect 495234 100574 495854 100658
rect 495234 100338 495266 100574
rect 495502 100338 495586 100574
rect 495822 100338 495854 100574
rect 495234 64894 495854 100338
rect 495234 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 495854 64894
rect 495234 64574 495854 64658
rect 495234 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 495854 64574
rect 495234 28894 495854 64338
rect 495234 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 495854 28894
rect 495234 28574 495854 28658
rect 495234 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 495854 28574
rect 495234 -5146 495854 28338
rect 495234 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 495854 -5146
rect 495234 -5466 495854 -5382
rect 495234 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 495854 -5466
rect 495234 -5734 495854 -5702
rect 498954 680614 499574 711002
rect 516954 710598 517574 711590
rect 516954 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 517574 710598
rect 516954 710278 517574 710362
rect 516954 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 517574 710278
rect 513234 708678 513854 709670
rect 513234 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 513854 708678
rect 513234 708358 513854 708442
rect 513234 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 513854 708358
rect 509514 706758 510134 707750
rect 509514 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 510134 706758
rect 509514 706438 510134 706522
rect 509514 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 510134 706438
rect 498954 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 499574 680614
rect 498954 680294 499574 680378
rect 498954 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 499574 680294
rect 498954 644614 499574 680058
rect 498954 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 499574 644614
rect 498954 644294 499574 644378
rect 498954 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 499574 644294
rect 498954 608614 499574 644058
rect 498954 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 499574 608614
rect 498954 608294 499574 608378
rect 498954 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 499574 608294
rect 498954 572614 499574 608058
rect 498954 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 499574 572614
rect 498954 572294 499574 572378
rect 498954 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 499574 572294
rect 498954 536614 499574 572058
rect 498954 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 499574 536614
rect 498954 536294 499574 536378
rect 498954 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 499574 536294
rect 498954 500614 499574 536058
rect 498954 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 499574 500614
rect 498954 500294 499574 500378
rect 498954 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 499574 500294
rect 498954 464614 499574 500058
rect 498954 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 499574 464614
rect 498954 464294 499574 464378
rect 498954 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 499574 464294
rect 498954 428614 499574 464058
rect 498954 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 499574 428614
rect 498954 428294 499574 428378
rect 498954 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 499574 428294
rect 498954 392614 499574 428058
rect 498954 392378 498986 392614
rect 499222 392378 499306 392614
rect 499542 392378 499574 392614
rect 498954 392294 499574 392378
rect 498954 392058 498986 392294
rect 499222 392058 499306 392294
rect 499542 392058 499574 392294
rect 498954 356614 499574 392058
rect 498954 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 499574 356614
rect 498954 356294 499574 356378
rect 498954 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 499574 356294
rect 498954 320614 499574 356058
rect 498954 320378 498986 320614
rect 499222 320378 499306 320614
rect 499542 320378 499574 320614
rect 498954 320294 499574 320378
rect 498954 320058 498986 320294
rect 499222 320058 499306 320294
rect 499542 320058 499574 320294
rect 498954 284614 499574 320058
rect 498954 284378 498986 284614
rect 499222 284378 499306 284614
rect 499542 284378 499574 284614
rect 498954 284294 499574 284378
rect 498954 284058 498986 284294
rect 499222 284058 499306 284294
rect 499542 284058 499574 284294
rect 498954 248614 499574 284058
rect 498954 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 499574 248614
rect 498954 248294 499574 248378
rect 498954 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 499574 248294
rect 498954 212614 499574 248058
rect 498954 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 499574 212614
rect 498954 212294 499574 212378
rect 498954 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 499574 212294
rect 498954 176614 499574 212058
rect 498954 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 499574 176614
rect 498954 176294 499574 176378
rect 498954 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 499574 176294
rect 498954 140614 499574 176058
rect 498954 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 499574 140614
rect 498954 140294 499574 140378
rect 498954 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 499574 140294
rect 498954 104614 499574 140058
rect 498954 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 499574 104614
rect 498954 104294 499574 104378
rect 498954 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 499574 104294
rect 498954 68614 499574 104058
rect 498954 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 499574 68614
rect 498954 68294 499574 68378
rect 498954 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 499574 68294
rect 498954 32614 499574 68058
rect 498954 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 499574 32614
rect 498954 32294 499574 32378
rect 498954 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 499574 32294
rect 480954 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 481574 -6106
rect 480954 -6426 481574 -6342
rect 480954 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 481574 -6426
rect 480954 -7654 481574 -6662
rect 498954 -7066 499574 32058
rect 505794 704838 506414 705830
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -1894 506414 -902
rect 509514 691174 510134 706202
rect 509514 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 510134 691174
rect 509514 690854 510134 690938
rect 509514 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 510134 690854
rect 509514 655174 510134 690618
rect 509514 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 510134 655174
rect 509514 654854 510134 654938
rect 509514 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 510134 654854
rect 509514 619174 510134 654618
rect 509514 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 510134 619174
rect 509514 618854 510134 618938
rect 509514 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 510134 618854
rect 509514 583174 510134 618618
rect 509514 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 510134 583174
rect 509514 582854 510134 582938
rect 509514 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 510134 582854
rect 509514 547174 510134 582618
rect 509514 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 510134 547174
rect 509514 546854 510134 546938
rect 509514 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 510134 546854
rect 509514 511174 510134 546618
rect 509514 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 510134 511174
rect 509514 510854 510134 510938
rect 509514 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 510134 510854
rect 509514 475174 510134 510618
rect 509514 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 510134 475174
rect 509514 474854 510134 474938
rect 509514 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 510134 474854
rect 509514 439174 510134 474618
rect 509514 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 510134 439174
rect 509514 438854 510134 438938
rect 509514 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 510134 438854
rect 509514 403174 510134 438618
rect 509514 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 510134 403174
rect 509514 402854 510134 402938
rect 509514 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 510134 402854
rect 509514 367174 510134 402618
rect 509514 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 510134 367174
rect 509514 366854 510134 366938
rect 509514 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 510134 366854
rect 509514 331174 510134 366618
rect 509514 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 510134 331174
rect 509514 330854 510134 330938
rect 509514 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 510134 330854
rect 509514 295174 510134 330618
rect 509514 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 510134 295174
rect 509514 294854 510134 294938
rect 509514 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 510134 294854
rect 509514 259174 510134 294618
rect 509514 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 510134 259174
rect 509514 258854 510134 258938
rect 509514 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 510134 258854
rect 509514 223174 510134 258618
rect 509514 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 510134 223174
rect 509514 222854 510134 222938
rect 509514 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 510134 222854
rect 509514 187174 510134 222618
rect 509514 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 510134 187174
rect 509514 186854 510134 186938
rect 509514 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 510134 186854
rect 509514 151174 510134 186618
rect 509514 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 510134 151174
rect 509514 150854 510134 150938
rect 509514 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 510134 150854
rect 509514 115174 510134 150618
rect 509514 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 510134 115174
rect 509514 114854 510134 114938
rect 509514 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 510134 114854
rect 509514 79174 510134 114618
rect 509514 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 510134 79174
rect 509514 78854 510134 78938
rect 509514 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 510134 78854
rect 509514 43174 510134 78618
rect 509514 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 510134 43174
rect 509514 42854 510134 42938
rect 509514 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 510134 42854
rect 509514 7174 510134 42618
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -2266 510134 6618
rect 509514 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 510134 -2266
rect 509514 -2586 510134 -2502
rect 509514 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 510134 -2586
rect 509514 -3814 510134 -2822
rect 513234 694894 513854 708122
rect 513234 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 513854 694894
rect 513234 694574 513854 694658
rect 513234 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 513854 694574
rect 513234 658894 513854 694338
rect 513234 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 513854 658894
rect 513234 658574 513854 658658
rect 513234 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 513854 658574
rect 513234 622894 513854 658338
rect 513234 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 513854 622894
rect 513234 622574 513854 622658
rect 513234 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 513854 622574
rect 513234 586894 513854 622338
rect 513234 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 513854 586894
rect 513234 586574 513854 586658
rect 513234 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 513854 586574
rect 513234 550894 513854 586338
rect 513234 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 513854 550894
rect 513234 550574 513854 550658
rect 513234 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 513854 550574
rect 513234 514894 513854 550338
rect 513234 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 513854 514894
rect 513234 514574 513854 514658
rect 513234 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 513854 514574
rect 513234 478894 513854 514338
rect 513234 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 513854 478894
rect 513234 478574 513854 478658
rect 513234 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 513854 478574
rect 513234 442894 513854 478338
rect 513234 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 513854 442894
rect 513234 442574 513854 442658
rect 513234 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 513854 442574
rect 513234 406894 513854 442338
rect 513234 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 513854 406894
rect 513234 406574 513854 406658
rect 513234 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 513854 406574
rect 513234 370894 513854 406338
rect 513234 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 513854 370894
rect 513234 370574 513854 370658
rect 513234 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 513854 370574
rect 513234 334894 513854 370338
rect 513234 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 513854 334894
rect 513234 334574 513854 334658
rect 513234 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 513854 334574
rect 513234 298894 513854 334338
rect 513234 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 513854 298894
rect 513234 298574 513854 298658
rect 513234 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 513854 298574
rect 513234 262894 513854 298338
rect 513234 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 513854 262894
rect 513234 262574 513854 262658
rect 513234 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 513854 262574
rect 513234 226894 513854 262338
rect 513234 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 513854 226894
rect 513234 226574 513854 226658
rect 513234 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 513854 226574
rect 513234 190894 513854 226338
rect 513234 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 513854 190894
rect 513234 190574 513854 190658
rect 513234 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 513854 190574
rect 513234 154894 513854 190338
rect 513234 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 513854 154894
rect 513234 154574 513854 154658
rect 513234 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 513854 154574
rect 513234 118894 513854 154338
rect 513234 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 513854 118894
rect 513234 118574 513854 118658
rect 513234 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 513854 118574
rect 513234 82894 513854 118338
rect 513234 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 513854 82894
rect 513234 82574 513854 82658
rect 513234 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 513854 82574
rect 513234 46894 513854 82338
rect 513234 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 513854 46894
rect 513234 46574 513854 46658
rect 513234 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 513854 46574
rect 513234 10894 513854 46338
rect 513234 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 513854 10894
rect 513234 10574 513854 10658
rect 513234 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 513854 10574
rect 513234 -4186 513854 10338
rect 513234 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 513854 -4186
rect 513234 -4506 513854 -4422
rect 513234 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 513854 -4506
rect 513234 -5734 513854 -4742
rect 516954 698614 517574 710042
rect 534954 711558 535574 711590
rect 534954 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 535574 711558
rect 534954 711238 535574 711322
rect 534954 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 535574 711238
rect 531234 709638 531854 709670
rect 531234 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 531854 709638
rect 531234 709318 531854 709402
rect 531234 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 531854 709318
rect 527514 707718 528134 707750
rect 527514 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 528134 707718
rect 527514 707398 528134 707482
rect 527514 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 528134 707398
rect 516954 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 517574 698614
rect 516954 698294 517574 698378
rect 516954 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 517574 698294
rect 516954 662614 517574 698058
rect 516954 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 517574 662614
rect 516954 662294 517574 662378
rect 516954 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 517574 662294
rect 516954 626614 517574 662058
rect 516954 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 517574 626614
rect 516954 626294 517574 626378
rect 516954 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 517574 626294
rect 516954 590614 517574 626058
rect 516954 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 517574 590614
rect 516954 590294 517574 590378
rect 516954 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 517574 590294
rect 516954 554614 517574 590058
rect 516954 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 517574 554614
rect 516954 554294 517574 554378
rect 516954 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 517574 554294
rect 516954 518614 517574 554058
rect 516954 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 517574 518614
rect 516954 518294 517574 518378
rect 516954 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 517574 518294
rect 516954 482614 517574 518058
rect 516954 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 517574 482614
rect 516954 482294 517574 482378
rect 516954 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 517574 482294
rect 516954 446614 517574 482058
rect 516954 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 517574 446614
rect 516954 446294 517574 446378
rect 516954 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 517574 446294
rect 516954 410614 517574 446058
rect 516954 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 517574 410614
rect 516954 410294 517574 410378
rect 516954 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 517574 410294
rect 516954 374614 517574 410058
rect 516954 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 517574 374614
rect 516954 374294 517574 374378
rect 516954 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 517574 374294
rect 516954 338614 517574 374058
rect 516954 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 517574 338614
rect 516954 338294 517574 338378
rect 516954 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 517574 338294
rect 516954 302614 517574 338058
rect 516954 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 517574 302614
rect 516954 302294 517574 302378
rect 516954 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 517574 302294
rect 516954 266614 517574 302058
rect 516954 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 517574 266614
rect 516954 266294 517574 266378
rect 516954 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 517574 266294
rect 516954 230614 517574 266058
rect 516954 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 517574 230614
rect 516954 230294 517574 230378
rect 516954 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 517574 230294
rect 516954 194614 517574 230058
rect 516954 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 517574 194614
rect 516954 194294 517574 194378
rect 516954 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 517574 194294
rect 516954 158614 517574 194058
rect 516954 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 517574 158614
rect 516954 158294 517574 158378
rect 516954 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 517574 158294
rect 516954 122614 517574 158058
rect 516954 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 517574 122614
rect 516954 122294 517574 122378
rect 516954 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 517574 122294
rect 516954 86614 517574 122058
rect 516954 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 517574 86614
rect 516954 86294 517574 86378
rect 516954 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 517574 86294
rect 516954 50614 517574 86058
rect 516954 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 517574 50614
rect 516954 50294 517574 50378
rect 516954 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 517574 50294
rect 516954 14614 517574 50058
rect 516954 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 517574 14614
rect 516954 14294 517574 14378
rect 516954 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 517574 14294
rect 498954 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 499574 -7066
rect 498954 -7386 499574 -7302
rect 498954 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 499574 -7386
rect 498954 -7654 499574 -7622
rect 516954 -6106 517574 14058
rect 523794 705798 524414 705830
rect 523794 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 524414 705798
rect 523794 705478 524414 705562
rect 523794 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 524414 705478
rect 523794 669454 524414 705242
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -1306 524414 20898
rect 523794 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 524414 -1306
rect 523794 -1626 524414 -1542
rect 523794 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 524414 -1626
rect 523794 -1894 524414 -1862
rect 527514 673174 528134 707162
rect 527514 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 528134 673174
rect 527514 672854 528134 672938
rect 527514 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 528134 672854
rect 527514 637174 528134 672618
rect 527514 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 528134 637174
rect 527514 636854 528134 636938
rect 527514 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 528134 636854
rect 527514 601174 528134 636618
rect 527514 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 528134 601174
rect 527514 600854 528134 600938
rect 527514 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 528134 600854
rect 527514 565174 528134 600618
rect 527514 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 528134 565174
rect 527514 564854 528134 564938
rect 527514 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 528134 564854
rect 527514 529174 528134 564618
rect 527514 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 528134 529174
rect 527514 528854 528134 528938
rect 527514 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 528134 528854
rect 527514 493174 528134 528618
rect 527514 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 528134 493174
rect 527514 492854 528134 492938
rect 527514 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 528134 492854
rect 527514 457174 528134 492618
rect 527514 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 528134 457174
rect 527514 456854 528134 456938
rect 527514 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 528134 456854
rect 527514 421174 528134 456618
rect 527514 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 528134 421174
rect 527514 420854 528134 420938
rect 527514 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 528134 420854
rect 527514 385174 528134 420618
rect 527514 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 528134 385174
rect 527514 384854 528134 384938
rect 527514 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 528134 384854
rect 527514 349174 528134 384618
rect 527514 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 528134 349174
rect 527514 348854 528134 348938
rect 527514 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 528134 348854
rect 527514 313174 528134 348618
rect 527514 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 528134 313174
rect 527514 312854 528134 312938
rect 527514 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 528134 312854
rect 527514 277174 528134 312618
rect 527514 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 528134 277174
rect 527514 276854 528134 276938
rect 527514 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 528134 276854
rect 527514 241174 528134 276618
rect 527514 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 528134 241174
rect 527514 240854 528134 240938
rect 527514 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 528134 240854
rect 527514 205174 528134 240618
rect 527514 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 528134 205174
rect 527514 204854 528134 204938
rect 527514 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 528134 204854
rect 527514 169174 528134 204618
rect 527514 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 528134 169174
rect 527514 168854 528134 168938
rect 527514 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 528134 168854
rect 527514 133174 528134 168618
rect 527514 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 528134 133174
rect 527514 132854 528134 132938
rect 527514 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 528134 132854
rect 527514 97174 528134 132618
rect 527514 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 528134 97174
rect 527514 96854 528134 96938
rect 527514 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 528134 96854
rect 527514 61174 528134 96618
rect 527514 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 528134 61174
rect 527514 60854 528134 60938
rect 527514 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 528134 60854
rect 527514 25174 528134 60618
rect 527514 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 528134 25174
rect 527514 24854 528134 24938
rect 527514 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 528134 24854
rect 527514 -3226 528134 24618
rect 527514 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 528134 -3226
rect 527514 -3546 528134 -3462
rect 527514 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 528134 -3546
rect 527514 -3814 528134 -3782
rect 531234 676894 531854 709082
rect 531234 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 531854 676894
rect 531234 676574 531854 676658
rect 531234 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 531854 676574
rect 531234 640894 531854 676338
rect 531234 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 531854 640894
rect 531234 640574 531854 640658
rect 531234 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 531854 640574
rect 531234 604894 531854 640338
rect 531234 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 531854 604894
rect 531234 604574 531854 604658
rect 531234 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 531854 604574
rect 531234 568894 531854 604338
rect 531234 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 531854 568894
rect 531234 568574 531854 568658
rect 531234 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 531854 568574
rect 531234 532894 531854 568338
rect 531234 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 531854 532894
rect 531234 532574 531854 532658
rect 531234 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 531854 532574
rect 531234 496894 531854 532338
rect 531234 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 531854 496894
rect 531234 496574 531854 496658
rect 531234 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 531854 496574
rect 531234 460894 531854 496338
rect 531234 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 531854 460894
rect 531234 460574 531854 460658
rect 531234 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 531854 460574
rect 531234 424894 531854 460338
rect 531234 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 531854 424894
rect 531234 424574 531854 424658
rect 531234 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 531854 424574
rect 531234 388894 531854 424338
rect 531234 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 531854 388894
rect 531234 388574 531854 388658
rect 531234 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 531854 388574
rect 531234 352894 531854 388338
rect 531234 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 531854 352894
rect 531234 352574 531854 352658
rect 531234 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 531854 352574
rect 531234 316894 531854 352338
rect 531234 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 531854 316894
rect 531234 316574 531854 316658
rect 531234 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 531854 316574
rect 531234 280894 531854 316338
rect 531234 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 531854 280894
rect 531234 280574 531854 280658
rect 531234 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 531854 280574
rect 531234 244894 531854 280338
rect 531234 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 531854 244894
rect 531234 244574 531854 244658
rect 531234 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 531854 244574
rect 531234 208894 531854 244338
rect 531234 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 531854 208894
rect 531234 208574 531854 208658
rect 531234 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 531854 208574
rect 531234 172894 531854 208338
rect 531234 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 531854 172894
rect 531234 172574 531854 172658
rect 531234 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 531854 172574
rect 531234 136894 531854 172338
rect 531234 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 531854 136894
rect 531234 136574 531854 136658
rect 531234 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 531854 136574
rect 531234 100894 531854 136338
rect 531234 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 531854 100894
rect 531234 100574 531854 100658
rect 531234 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 531854 100574
rect 531234 64894 531854 100338
rect 531234 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 531854 64894
rect 531234 64574 531854 64658
rect 531234 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 531854 64574
rect 531234 28894 531854 64338
rect 531234 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 531854 28894
rect 531234 28574 531854 28658
rect 531234 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 531854 28574
rect 531234 -5146 531854 28338
rect 531234 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 531854 -5146
rect 531234 -5466 531854 -5382
rect 531234 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 531854 -5466
rect 531234 -5734 531854 -5702
rect 534954 680614 535574 711002
rect 552954 710598 553574 711590
rect 552954 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 553574 710598
rect 552954 710278 553574 710362
rect 552954 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 553574 710278
rect 549234 708678 549854 709670
rect 549234 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 549854 708678
rect 549234 708358 549854 708442
rect 549234 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 549854 708358
rect 545514 706758 546134 707750
rect 545514 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 546134 706758
rect 545514 706438 546134 706522
rect 545514 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 546134 706438
rect 534954 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 535574 680614
rect 534954 680294 535574 680378
rect 534954 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 535574 680294
rect 534954 644614 535574 680058
rect 534954 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 535574 644614
rect 534954 644294 535574 644378
rect 534954 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 535574 644294
rect 534954 608614 535574 644058
rect 534954 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 535574 608614
rect 534954 608294 535574 608378
rect 534954 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 535574 608294
rect 534954 572614 535574 608058
rect 534954 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 535574 572614
rect 534954 572294 535574 572378
rect 534954 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 535574 572294
rect 534954 536614 535574 572058
rect 534954 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 535574 536614
rect 534954 536294 535574 536378
rect 534954 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 535574 536294
rect 534954 500614 535574 536058
rect 534954 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 535574 500614
rect 534954 500294 535574 500378
rect 534954 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 535574 500294
rect 534954 464614 535574 500058
rect 534954 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 535574 464614
rect 534954 464294 535574 464378
rect 534954 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 535574 464294
rect 534954 428614 535574 464058
rect 534954 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 535574 428614
rect 534954 428294 535574 428378
rect 534954 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 535574 428294
rect 534954 392614 535574 428058
rect 534954 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 535574 392614
rect 534954 392294 535574 392378
rect 534954 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 535574 392294
rect 534954 356614 535574 392058
rect 534954 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 535574 356614
rect 534954 356294 535574 356378
rect 534954 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 535574 356294
rect 534954 320614 535574 356058
rect 534954 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 535574 320614
rect 534954 320294 535574 320378
rect 534954 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 535574 320294
rect 534954 284614 535574 320058
rect 534954 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 535574 284614
rect 534954 284294 535574 284378
rect 534954 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 535574 284294
rect 534954 248614 535574 284058
rect 534954 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 535574 248614
rect 534954 248294 535574 248378
rect 534954 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 535574 248294
rect 534954 212614 535574 248058
rect 534954 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 535574 212614
rect 534954 212294 535574 212378
rect 534954 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 535574 212294
rect 534954 176614 535574 212058
rect 534954 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 535574 176614
rect 534954 176294 535574 176378
rect 534954 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 535574 176294
rect 534954 140614 535574 176058
rect 534954 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 535574 140614
rect 534954 140294 535574 140378
rect 534954 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 535574 140294
rect 534954 104614 535574 140058
rect 534954 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 535574 104614
rect 534954 104294 535574 104378
rect 534954 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 535574 104294
rect 534954 68614 535574 104058
rect 534954 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 535574 68614
rect 534954 68294 535574 68378
rect 534954 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 535574 68294
rect 534954 32614 535574 68058
rect 534954 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 535574 32614
rect 534954 32294 535574 32378
rect 534954 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 535574 32294
rect 516954 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 517574 -6106
rect 516954 -6426 517574 -6342
rect 516954 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 517574 -6426
rect 516954 -7654 517574 -6662
rect 534954 -7066 535574 32058
rect 541794 704838 542414 705830
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -1894 542414 -902
rect 545514 691174 546134 706202
rect 545514 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 546134 691174
rect 545514 690854 546134 690938
rect 545514 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 546134 690854
rect 545514 655174 546134 690618
rect 545514 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 546134 655174
rect 545514 654854 546134 654938
rect 545514 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 546134 654854
rect 545514 619174 546134 654618
rect 545514 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 546134 619174
rect 545514 618854 546134 618938
rect 545514 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 546134 618854
rect 545514 583174 546134 618618
rect 545514 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 546134 583174
rect 545514 582854 546134 582938
rect 545514 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 546134 582854
rect 545514 547174 546134 582618
rect 545514 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 546134 547174
rect 545514 546854 546134 546938
rect 545514 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 546134 546854
rect 545514 511174 546134 546618
rect 545514 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 546134 511174
rect 545514 510854 546134 510938
rect 545514 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 546134 510854
rect 545514 475174 546134 510618
rect 545514 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 546134 475174
rect 545514 474854 546134 474938
rect 545514 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 546134 474854
rect 545514 439174 546134 474618
rect 545514 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 546134 439174
rect 545514 438854 546134 438938
rect 545514 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 546134 438854
rect 545514 403174 546134 438618
rect 545514 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 546134 403174
rect 545514 402854 546134 402938
rect 545514 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 546134 402854
rect 545514 367174 546134 402618
rect 545514 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 546134 367174
rect 545514 366854 546134 366938
rect 545514 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 546134 366854
rect 545514 331174 546134 366618
rect 545514 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 546134 331174
rect 545514 330854 546134 330938
rect 545514 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 546134 330854
rect 545514 295174 546134 330618
rect 545514 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 546134 295174
rect 545514 294854 546134 294938
rect 545514 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 546134 294854
rect 545514 259174 546134 294618
rect 545514 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 546134 259174
rect 545514 258854 546134 258938
rect 545514 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 546134 258854
rect 545514 223174 546134 258618
rect 545514 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 546134 223174
rect 545514 222854 546134 222938
rect 545514 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 546134 222854
rect 545514 187174 546134 222618
rect 545514 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 546134 187174
rect 545514 186854 546134 186938
rect 545514 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 546134 186854
rect 545514 151174 546134 186618
rect 545514 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 546134 151174
rect 545514 150854 546134 150938
rect 545514 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 546134 150854
rect 545514 115174 546134 150618
rect 545514 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 546134 115174
rect 545514 114854 546134 114938
rect 545514 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 546134 114854
rect 545514 79174 546134 114618
rect 545514 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 546134 79174
rect 545514 78854 546134 78938
rect 545514 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 546134 78854
rect 545514 43174 546134 78618
rect 545514 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 546134 43174
rect 545514 42854 546134 42938
rect 545514 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 546134 42854
rect 545514 7174 546134 42618
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -2266 546134 6618
rect 545514 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 546134 -2266
rect 545514 -2586 546134 -2502
rect 545514 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 546134 -2586
rect 545514 -3814 546134 -2822
rect 549234 694894 549854 708122
rect 549234 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 549854 694894
rect 549234 694574 549854 694658
rect 549234 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 549854 694574
rect 549234 658894 549854 694338
rect 549234 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 549854 658894
rect 549234 658574 549854 658658
rect 549234 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 549854 658574
rect 549234 622894 549854 658338
rect 549234 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 549854 622894
rect 549234 622574 549854 622658
rect 549234 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 549854 622574
rect 549234 586894 549854 622338
rect 549234 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 549854 586894
rect 549234 586574 549854 586658
rect 549234 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 549854 586574
rect 549234 550894 549854 586338
rect 549234 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 549854 550894
rect 549234 550574 549854 550658
rect 549234 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 549854 550574
rect 549234 514894 549854 550338
rect 549234 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 549854 514894
rect 549234 514574 549854 514658
rect 549234 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 549854 514574
rect 549234 478894 549854 514338
rect 549234 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 549854 478894
rect 549234 478574 549854 478658
rect 549234 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 549854 478574
rect 549234 442894 549854 478338
rect 549234 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 549854 442894
rect 549234 442574 549854 442658
rect 549234 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 549854 442574
rect 549234 406894 549854 442338
rect 549234 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 549854 406894
rect 549234 406574 549854 406658
rect 549234 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 549854 406574
rect 549234 370894 549854 406338
rect 549234 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 549854 370894
rect 549234 370574 549854 370658
rect 549234 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 549854 370574
rect 549234 334894 549854 370338
rect 549234 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 549854 334894
rect 549234 334574 549854 334658
rect 549234 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 549854 334574
rect 549234 298894 549854 334338
rect 549234 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 549854 298894
rect 549234 298574 549854 298658
rect 549234 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 549854 298574
rect 549234 262894 549854 298338
rect 549234 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 549854 262894
rect 549234 262574 549854 262658
rect 549234 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 549854 262574
rect 549234 226894 549854 262338
rect 549234 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 549854 226894
rect 549234 226574 549854 226658
rect 549234 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 549854 226574
rect 549234 190894 549854 226338
rect 549234 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 549854 190894
rect 549234 190574 549854 190658
rect 549234 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 549854 190574
rect 549234 154894 549854 190338
rect 549234 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 549854 154894
rect 549234 154574 549854 154658
rect 549234 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 549854 154574
rect 549234 118894 549854 154338
rect 549234 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 549854 118894
rect 549234 118574 549854 118658
rect 549234 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 549854 118574
rect 549234 82894 549854 118338
rect 549234 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 549854 82894
rect 549234 82574 549854 82658
rect 549234 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 549854 82574
rect 549234 46894 549854 82338
rect 549234 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 549854 46894
rect 549234 46574 549854 46658
rect 549234 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 549854 46574
rect 549234 10894 549854 46338
rect 549234 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 549854 10894
rect 549234 10574 549854 10658
rect 549234 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 549854 10574
rect 549234 -4186 549854 10338
rect 549234 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 549854 -4186
rect 549234 -4506 549854 -4422
rect 549234 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 549854 -4506
rect 549234 -5734 549854 -4742
rect 552954 698614 553574 710042
rect 570954 711558 571574 711590
rect 570954 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 571574 711558
rect 570954 711238 571574 711322
rect 570954 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 571574 711238
rect 567234 709638 567854 709670
rect 567234 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 567854 709638
rect 567234 709318 567854 709402
rect 567234 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 567854 709318
rect 563514 707718 564134 707750
rect 563514 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 564134 707718
rect 563514 707398 564134 707482
rect 563514 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 564134 707398
rect 552954 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 553574 698614
rect 552954 698294 553574 698378
rect 552954 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 553574 698294
rect 552954 662614 553574 698058
rect 552954 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 553574 662614
rect 552954 662294 553574 662378
rect 552954 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 553574 662294
rect 552954 626614 553574 662058
rect 552954 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 553574 626614
rect 552954 626294 553574 626378
rect 552954 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 553574 626294
rect 552954 590614 553574 626058
rect 552954 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 553574 590614
rect 552954 590294 553574 590378
rect 552954 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 553574 590294
rect 552954 554614 553574 590058
rect 552954 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 553574 554614
rect 552954 554294 553574 554378
rect 552954 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 553574 554294
rect 552954 518614 553574 554058
rect 552954 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 553574 518614
rect 552954 518294 553574 518378
rect 552954 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 553574 518294
rect 552954 482614 553574 518058
rect 552954 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 553574 482614
rect 552954 482294 553574 482378
rect 552954 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 553574 482294
rect 552954 446614 553574 482058
rect 552954 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 553574 446614
rect 552954 446294 553574 446378
rect 552954 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 553574 446294
rect 552954 410614 553574 446058
rect 552954 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 553574 410614
rect 552954 410294 553574 410378
rect 552954 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 553574 410294
rect 552954 374614 553574 410058
rect 552954 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 553574 374614
rect 552954 374294 553574 374378
rect 552954 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 553574 374294
rect 552954 338614 553574 374058
rect 552954 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 553574 338614
rect 552954 338294 553574 338378
rect 552954 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 553574 338294
rect 552954 302614 553574 338058
rect 552954 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 553574 302614
rect 552954 302294 553574 302378
rect 552954 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 553574 302294
rect 552954 266614 553574 302058
rect 552954 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 553574 266614
rect 552954 266294 553574 266378
rect 552954 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 553574 266294
rect 552954 230614 553574 266058
rect 552954 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 553574 230614
rect 552954 230294 553574 230378
rect 552954 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 553574 230294
rect 552954 194614 553574 230058
rect 552954 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 553574 194614
rect 552954 194294 553574 194378
rect 552954 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 553574 194294
rect 552954 158614 553574 194058
rect 552954 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 553574 158614
rect 552954 158294 553574 158378
rect 552954 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 553574 158294
rect 552954 122614 553574 158058
rect 552954 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 553574 122614
rect 552954 122294 553574 122378
rect 552954 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 553574 122294
rect 552954 86614 553574 122058
rect 552954 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 553574 86614
rect 552954 86294 553574 86378
rect 552954 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 553574 86294
rect 552954 50614 553574 86058
rect 552954 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 553574 50614
rect 552954 50294 553574 50378
rect 552954 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 553574 50294
rect 552954 14614 553574 50058
rect 552954 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 553574 14614
rect 552954 14294 553574 14378
rect 552954 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 553574 14294
rect 534954 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 535574 -7066
rect 534954 -7386 535574 -7302
rect 534954 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 535574 -7386
rect 534954 -7654 535574 -7622
rect 552954 -6106 553574 14058
rect 559794 705798 560414 705830
rect 559794 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 560414 705798
rect 559794 705478 560414 705562
rect 559794 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 560414 705478
rect 559794 669454 560414 705242
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -1306 560414 20898
rect 559794 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 560414 -1306
rect 559794 -1626 560414 -1542
rect 559794 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 560414 -1626
rect 559794 -1894 560414 -1862
rect 563514 673174 564134 707162
rect 563514 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 564134 673174
rect 563514 672854 564134 672938
rect 563514 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 564134 672854
rect 563514 637174 564134 672618
rect 563514 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 564134 637174
rect 563514 636854 564134 636938
rect 563514 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 564134 636854
rect 563514 601174 564134 636618
rect 563514 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 564134 601174
rect 563514 600854 564134 600938
rect 563514 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 564134 600854
rect 563514 565174 564134 600618
rect 563514 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 564134 565174
rect 563514 564854 564134 564938
rect 563514 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 564134 564854
rect 563514 529174 564134 564618
rect 563514 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 564134 529174
rect 563514 528854 564134 528938
rect 563514 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 564134 528854
rect 563514 493174 564134 528618
rect 563514 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 564134 493174
rect 563514 492854 564134 492938
rect 563514 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 564134 492854
rect 563514 457174 564134 492618
rect 563514 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 564134 457174
rect 563514 456854 564134 456938
rect 563514 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 564134 456854
rect 563514 421174 564134 456618
rect 563514 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 564134 421174
rect 563514 420854 564134 420938
rect 563514 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 564134 420854
rect 563514 385174 564134 420618
rect 563514 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 564134 385174
rect 563514 384854 564134 384938
rect 563514 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 564134 384854
rect 563514 349174 564134 384618
rect 563514 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 564134 349174
rect 563514 348854 564134 348938
rect 563514 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 564134 348854
rect 563514 313174 564134 348618
rect 563514 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 564134 313174
rect 563514 312854 564134 312938
rect 563514 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 564134 312854
rect 563514 277174 564134 312618
rect 563514 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 564134 277174
rect 563514 276854 564134 276938
rect 563514 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 564134 276854
rect 563514 241174 564134 276618
rect 563514 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 564134 241174
rect 563514 240854 564134 240938
rect 563514 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 564134 240854
rect 563514 205174 564134 240618
rect 563514 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 564134 205174
rect 563514 204854 564134 204938
rect 563514 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 564134 204854
rect 563514 169174 564134 204618
rect 563514 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 564134 169174
rect 563514 168854 564134 168938
rect 563514 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 564134 168854
rect 563514 133174 564134 168618
rect 563514 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 564134 133174
rect 563514 132854 564134 132938
rect 563514 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 564134 132854
rect 563514 97174 564134 132618
rect 563514 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 564134 97174
rect 563514 96854 564134 96938
rect 563514 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 564134 96854
rect 563514 61174 564134 96618
rect 563514 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 564134 61174
rect 563514 60854 564134 60938
rect 563514 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 564134 60854
rect 563514 25174 564134 60618
rect 563514 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 564134 25174
rect 563514 24854 564134 24938
rect 563514 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 564134 24854
rect 563514 -3226 564134 24618
rect 563514 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 564134 -3226
rect 563514 -3546 564134 -3462
rect 563514 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 564134 -3546
rect 563514 -3814 564134 -3782
rect 567234 676894 567854 709082
rect 567234 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 567854 676894
rect 567234 676574 567854 676658
rect 567234 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 567854 676574
rect 567234 640894 567854 676338
rect 567234 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 567854 640894
rect 567234 640574 567854 640658
rect 567234 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 567854 640574
rect 567234 604894 567854 640338
rect 567234 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 567854 604894
rect 567234 604574 567854 604658
rect 567234 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 567854 604574
rect 567234 568894 567854 604338
rect 567234 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 567854 568894
rect 567234 568574 567854 568658
rect 567234 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 567854 568574
rect 567234 532894 567854 568338
rect 567234 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 567854 532894
rect 567234 532574 567854 532658
rect 567234 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 567854 532574
rect 567234 496894 567854 532338
rect 567234 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 567854 496894
rect 567234 496574 567854 496658
rect 567234 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 567854 496574
rect 567234 460894 567854 496338
rect 567234 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 567854 460894
rect 567234 460574 567854 460658
rect 567234 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 567854 460574
rect 567234 424894 567854 460338
rect 567234 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 567854 424894
rect 567234 424574 567854 424658
rect 567234 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 567854 424574
rect 567234 388894 567854 424338
rect 567234 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 567854 388894
rect 567234 388574 567854 388658
rect 567234 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 567854 388574
rect 567234 352894 567854 388338
rect 567234 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 567854 352894
rect 567234 352574 567854 352658
rect 567234 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 567854 352574
rect 567234 316894 567854 352338
rect 567234 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 567854 316894
rect 567234 316574 567854 316658
rect 567234 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 567854 316574
rect 567234 280894 567854 316338
rect 567234 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 567854 280894
rect 567234 280574 567854 280658
rect 567234 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 567854 280574
rect 567234 244894 567854 280338
rect 567234 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 567854 244894
rect 567234 244574 567854 244658
rect 567234 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 567854 244574
rect 567234 208894 567854 244338
rect 567234 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 567854 208894
rect 567234 208574 567854 208658
rect 567234 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 567854 208574
rect 567234 172894 567854 208338
rect 567234 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 567854 172894
rect 567234 172574 567854 172658
rect 567234 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 567854 172574
rect 567234 136894 567854 172338
rect 567234 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 567854 136894
rect 567234 136574 567854 136658
rect 567234 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 567854 136574
rect 567234 100894 567854 136338
rect 567234 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 567854 100894
rect 567234 100574 567854 100658
rect 567234 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 567854 100574
rect 567234 64894 567854 100338
rect 567234 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 567854 64894
rect 567234 64574 567854 64658
rect 567234 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 567854 64574
rect 567234 28894 567854 64338
rect 567234 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 567854 28894
rect 567234 28574 567854 28658
rect 567234 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 567854 28574
rect 567234 -5146 567854 28338
rect 567234 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 567854 -5146
rect 567234 -5466 567854 -5382
rect 567234 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 567854 -5466
rect 567234 -5734 567854 -5702
rect 570954 680614 571574 711002
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 581514 706758 582134 707750
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 581514 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 582134 706758
rect 581514 706438 582134 706522
rect 581514 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 582134 706438
rect 570954 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 571574 680614
rect 570954 680294 571574 680378
rect 570954 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 571574 680294
rect 570954 644614 571574 680058
rect 570954 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 571574 644614
rect 570954 644294 571574 644378
rect 570954 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 571574 644294
rect 570954 608614 571574 644058
rect 570954 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 571574 608614
rect 570954 608294 571574 608378
rect 570954 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 571574 608294
rect 570954 572614 571574 608058
rect 570954 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 571574 572614
rect 570954 572294 571574 572378
rect 570954 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 571574 572294
rect 570954 536614 571574 572058
rect 570954 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 571574 536614
rect 570954 536294 571574 536378
rect 570954 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 571574 536294
rect 570954 500614 571574 536058
rect 570954 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 571574 500614
rect 570954 500294 571574 500378
rect 570954 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 571574 500294
rect 570954 464614 571574 500058
rect 570954 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 571574 464614
rect 570954 464294 571574 464378
rect 570954 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 571574 464294
rect 570954 428614 571574 464058
rect 570954 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 571574 428614
rect 570954 428294 571574 428378
rect 570954 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 571574 428294
rect 570954 392614 571574 428058
rect 570954 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 571574 392614
rect 570954 392294 571574 392378
rect 570954 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 571574 392294
rect 570954 356614 571574 392058
rect 570954 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 571574 356614
rect 570954 356294 571574 356378
rect 570954 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 571574 356294
rect 570954 320614 571574 356058
rect 570954 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 571574 320614
rect 570954 320294 571574 320378
rect 570954 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 571574 320294
rect 570954 284614 571574 320058
rect 570954 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 571574 284614
rect 570954 284294 571574 284378
rect 570954 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 571574 284294
rect 570954 248614 571574 284058
rect 570954 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 571574 248614
rect 570954 248294 571574 248378
rect 570954 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 571574 248294
rect 570954 212614 571574 248058
rect 570954 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 571574 212614
rect 570954 212294 571574 212378
rect 570954 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 571574 212294
rect 570954 176614 571574 212058
rect 570954 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 571574 176614
rect 570954 176294 571574 176378
rect 570954 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 571574 176294
rect 570954 140614 571574 176058
rect 570954 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 571574 140614
rect 570954 140294 571574 140378
rect 570954 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 571574 140294
rect 570954 104614 571574 140058
rect 570954 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 571574 104614
rect 570954 104294 571574 104378
rect 570954 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 571574 104294
rect 570954 68614 571574 104058
rect 570954 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 571574 68614
rect 570954 68294 571574 68378
rect 570954 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 571574 68294
rect 570954 32614 571574 68058
rect 570954 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 571574 32614
rect 570954 32294 571574 32378
rect 570954 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 571574 32294
rect 552954 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 553574 -6106
rect 552954 -6426 553574 -6342
rect 552954 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 553574 -6426
rect 552954 -7654 553574 -6662
rect 570954 -7066 571574 32058
rect 577794 704838 578414 705830
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -1894 578414 -902
rect 581514 691174 582134 706202
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -2266 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 669454 586890 705242
rect 586270 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect 586270 669134 586890 669218
rect 586270 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect 586270 633454 586890 668898
rect 586270 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect 586270 633134 586890 633218
rect 586270 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect 586270 597454 586890 632898
rect 586270 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect 586270 597134 586890 597218
rect 586270 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect 586270 561454 586890 596898
rect 586270 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect 586270 561134 586890 561218
rect 586270 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect 586270 525454 586890 560898
rect 586270 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect 586270 525134 586890 525218
rect 586270 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect 586270 489454 586890 524898
rect 586270 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect 586270 489134 586890 489218
rect 586270 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect 586270 453454 586890 488898
rect 586270 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect 586270 453134 586890 453218
rect 586270 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect 586270 417454 586890 452898
rect 586270 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect 586270 417134 586890 417218
rect 586270 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect 586270 381454 586890 416898
rect 586270 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect 586270 381134 586890 381218
rect 586270 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect 586270 345454 586890 380898
rect 586270 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect 586270 345134 586890 345218
rect 586270 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect 586270 309454 586890 344898
rect 586270 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect 586270 309134 586890 309218
rect 586270 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect 586270 273454 586890 308898
rect 586270 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect 586270 273134 586890 273218
rect 586270 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect 586270 237454 586890 272898
rect 586270 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect 586270 237134 586890 237218
rect 586270 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect 586270 201454 586890 236898
rect 586270 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect 586270 201134 586890 201218
rect 586270 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect 586270 165454 586890 200898
rect 586270 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect 586270 165134 586890 165218
rect 586270 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect 586270 129454 586890 164898
rect 586270 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect 586270 129134 586890 129218
rect 586270 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect 586270 93454 586890 128898
rect 586270 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect 586270 93134 586890 93218
rect 586270 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect 586270 57454 586890 92898
rect 586270 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect 586270 57134 586890 57218
rect 586270 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect 586270 21454 586890 56898
rect 586270 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect 586270 21134 586890 21218
rect 586270 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect 586270 -1306 586890 20898
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 691174 587850 706202
rect 587230 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 587850 691174
rect 587230 690854 587850 690938
rect 587230 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 587850 690854
rect 587230 655174 587850 690618
rect 587230 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 587850 655174
rect 587230 654854 587850 654938
rect 587230 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 587850 654854
rect 587230 619174 587850 654618
rect 587230 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 587850 619174
rect 587230 618854 587850 618938
rect 587230 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 587850 618854
rect 587230 583174 587850 618618
rect 587230 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 587850 583174
rect 587230 582854 587850 582938
rect 587230 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 587850 582854
rect 587230 547174 587850 582618
rect 587230 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 587850 547174
rect 587230 546854 587850 546938
rect 587230 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 587850 546854
rect 587230 511174 587850 546618
rect 587230 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 587850 511174
rect 587230 510854 587850 510938
rect 587230 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 587850 510854
rect 587230 475174 587850 510618
rect 587230 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 587850 475174
rect 587230 474854 587850 474938
rect 587230 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 587850 474854
rect 587230 439174 587850 474618
rect 587230 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 587850 439174
rect 587230 438854 587850 438938
rect 587230 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 587850 438854
rect 587230 403174 587850 438618
rect 587230 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 587850 403174
rect 587230 402854 587850 402938
rect 587230 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 587850 402854
rect 587230 367174 587850 402618
rect 587230 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 587850 367174
rect 587230 366854 587850 366938
rect 587230 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 587850 366854
rect 587230 331174 587850 366618
rect 587230 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 587850 331174
rect 587230 330854 587850 330938
rect 587230 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 587850 330854
rect 587230 295174 587850 330618
rect 587230 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 587850 295174
rect 587230 294854 587850 294938
rect 587230 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 587850 294854
rect 587230 259174 587850 294618
rect 587230 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 587850 259174
rect 587230 258854 587850 258938
rect 587230 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 587850 258854
rect 587230 223174 587850 258618
rect 587230 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 587850 223174
rect 587230 222854 587850 222938
rect 587230 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 587850 222854
rect 587230 187174 587850 222618
rect 587230 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 587850 187174
rect 587230 186854 587850 186938
rect 587230 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 587850 186854
rect 587230 151174 587850 186618
rect 587230 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 587850 151174
rect 587230 150854 587850 150938
rect 587230 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 587850 150854
rect 587230 115174 587850 150618
rect 587230 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 587850 115174
rect 587230 114854 587850 114938
rect 587230 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 587850 114854
rect 587230 79174 587850 114618
rect 587230 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 587850 79174
rect 587230 78854 587850 78938
rect 587230 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 587850 78854
rect 587230 43174 587850 78618
rect 587230 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 587850 43174
rect 587230 42854 587850 42938
rect 587230 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 587850 42854
rect 587230 7174 587850 42618
rect 587230 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 587850 7174
rect 587230 6854 587850 6938
rect 587230 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 587850 6854
rect 581514 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 582134 -2266
rect 581514 -2586 582134 -2502
rect 581514 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 582134 -2586
rect 581514 -3814 582134 -2822
rect 587230 -2266 587850 6618
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 673174 588810 707162
rect 588190 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect 588190 672854 588810 672938
rect 588190 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect 588190 637174 588810 672618
rect 588190 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect 588190 636854 588810 636938
rect 588190 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect 588190 601174 588810 636618
rect 588190 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect 588190 600854 588810 600938
rect 588190 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect 588190 565174 588810 600618
rect 588190 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect 588190 564854 588810 564938
rect 588190 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect 588190 529174 588810 564618
rect 588190 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect 588190 528854 588810 528938
rect 588190 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect 588190 493174 588810 528618
rect 588190 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect 588190 492854 588810 492938
rect 588190 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect 588190 457174 588810 492618
rect 588190 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect 588190 456854 588810 456938
rect 588190 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect 588190 421174 588810 456618
rect 588190 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect 588190 420854 588810 420938
rect 588190 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect 588190 385174 588810 420618
rect 588190 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect 588190 384854 588810 384938
rect 588190 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect 588190 349174 588810 384618
rect 588190 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect 588190 348854 588810 348938
rect 588190 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect 588190 313174 588810 348618
rect 588190 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect 588190 312854 588810 312938
rect 588190 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect 588190 277174 588810 312618
rect 588190 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect 588190 276854 588810 276938
rect 588190 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect 588190 241174 588810 276618
rect 588190 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect 588190 240854 588810 240938
rect 588190 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect 588190 205174 588810 240618
rect 588190 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect 588190 204854 588810 204938
rect 588190 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect 588190 169174 588810 204618
rect 588190 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect 588190 168854 588810 168938
rect 588190 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect 588190 133174 588810 168618
rect 588190 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect 588190 132854 588810 132938
rect 588190 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect 588190 97174 588810 132618
rect 588190 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect 588190 96854 588810 96938
rect 588190 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect 588190 61174 588810 96618
rect 588190 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect 588190 60854 588810 60938
rect 588190 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect 588190 25174 588810 60618
rect 588190 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect 588190 24854 588810 24938
rect 588190 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect 588190 -3226 588810 24618
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 694894 589770 708122
rect 589150 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 589770 694894
rect 589150 694574 589770 694658
rect 589150 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 589770 694574
rect 589150 658894 589770 694338
rect 589150 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 589770 658894
rect 589150 658574 589770 658658
rect 589150 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 589770 658574
rect 589150 622894 589770 658338
rect 589150 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 589770 622894
rect 589150 622574 589770 622658
rect 589150 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 589770 622574
rect 589150 586894 589770 622338
rect 589150 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 589770 586894
rect 589150 586574 589770 586658
rect 589150 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 589770 586574
rect 589150 550894 589770 586338
rect 589150 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 589770 550894
rect 589150 550574 589770 550658
rect 589150 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 589770 550574
rect 589150 514894 589770 550338
rect 589150 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 589770 514894
rect 589150 514574 589770 514658
rect 589150 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 589770 514574
rect 589150 478894 589770 514338
rect 589150 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 589770 478894
rect 589150 478574 589770 478658
rect 589150 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 589770 478574
rect 589150 442894 589770 478338
rect 589150 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 589770 442894
rect 589150 442574 589770 442658
rect 589150 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 589770 442574
rect 589150 406894 589770 442338
rect 589150 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 589770 406894
rect 589150 406574 589770 406658
rect 589150 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 589770 406574
rect 589150 370894 589770 406338
rect 589150 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 589770 370894
rect 589150 370574 589770 370658
rect 589150 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 589770 370574
rect 589150 334894 589770 370338
rect 589150 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 589770 334894
rect 589150 334574 589770 334658
rect 589150 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 589770 334574
rect 589150 298894 589770 334338
rect 589150 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 589770 298894
rect 589150 298574 589770 298658
rect 589150 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 589770 298574
rect 589150 262894 589770 298338
rect 589150 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 589770 262894
rect 589150 262574 589770 262658
rect 589150 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 589770 262574
rect 589150 226894 589770 262338
rect 589150 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 589770 226894
rect 589150 226574 589770 226658
rect 589150 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 589770 226574
rect 589150 190894 589770 226338
rect 589150 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 589770 190894
rect 589150 190574 589770 190658
rect 589150 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 589770 190574
rect 589150 154894 589770 190338
rect 589150 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 589770 154894
rect 589150 154574 589770 154658
rect 589150 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 589770 154574
rect 589150 118894 589770 154338
rect 589150 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 589770 118894
rect 589150 118574 589770 118658
rect 589150 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 589770 118574
rect 589150 82894 589770 118338
rect 589150 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 589770 82894
rect 589150 82574 589770 82658
rect 589150 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 589770 82574
rect 589150 46894 589770 82338
rect 589150 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 589770 46894
rect 589150 46574 589770 46658
rect 589150 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 589770 46574
rect 589150 10894 589770 46338
rect 589150 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 589770 10894
rect 589150 10574 589770 10658
rect 589150 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 589770 10574
rect 589150 -4186 589770 10338
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 676894 590730 709082
rect 590110 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect 590110 676574 590730 676658
rect 590110 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect 590110 640894 590730 676338
rect 590110 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect 590110 640574 590730 640658
rect 590110 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect 590110 604894 590730 640338
rect 590110 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect 590110 604574 590730 604658
rect 590110 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect 590110 568894 590730 604338
rect 590110 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect 590110 568574 590730 568658
rect 590110 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect 590110 532894 590730 568338
rect 590110 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect 590110 532574 590730 532658
rect 590110 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect 590110 496894 590730 532338
rect 590110 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect 590110 496574 590730 496658
rect 590110 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect 590110 460894 590730 496338
rect 590110 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect 590110 460574 590730 460658
rect 590110 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect 590110 424894 590730 460338
rect 590110 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect 590110 424574 590730 424658
rect 590110 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect 590110 388894 590730 424338
rect 590110 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect 590110 388574 590730 388658
rect 590110 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect 590110 352894 590730 388338
rect 590110 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect 590110 352574 590730 352658
rect 590110 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect 590110 316894 590730 352338
rect 590110 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect 590110 316574 590730 316658
rect 590110 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect 590110 280894 590730 316338
rect 590110 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect 590110 280574 590730 280658
rect 590110 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect 590110 244894 590730 280338
rect 590110 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect 590110 244574 590730 244658
rect 590110 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect 590110 208894 590730 244338
rect 590110 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect 590110 208574 590730 208658
rect 590110 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect 590110 172894 590730 208338
rect 590110 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect 590110 172574 590730 172658
rect 590110 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect 590110 136894 590730 172338
rect 590110 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect 590110 136574 590730 136658
rect 590110 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect 590110 100894 590730 136338
rect 590110 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect 590110 100574 590730 100658
rect 590110 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect 590110 64894 590730 100338
rect 590110 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect 590110 64574 590730 64658
rect 590110 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect 590110 28894 590730 64338
rect 590110 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect 590110 28574 590730 28658
rect 590110 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect 590110 -5146 590730 28338
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 698614 591690 710042
rect 591070 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 591690 698614
rect 591070 698294 591690 698378
rect 591070 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 591690 698294
rect 591070 662614 591690 698058
rect 591070 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 591690 662614
rect 591070 662294 591690 662378
rect 591070 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 591690 662294
rect 591070 626614 591690 662058
rect 591070 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 591690 626614
rect 591070 626294 591690 626378
rect 591070 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 591690 626294
rect 591070 590614 591690 626058
rect 591070 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 591690 590614
rect 591070 590294 591690 590378
rect 591070 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 591690 590294
rect 591070 554614 591690 590058
rect 591070 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 591690 554614
rect 591070 554294 591690 554378
rect 591070 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 591690 554294
rect 591070 518614 591690 554058
rect 591070 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 591690 518614
rect 591070 518294 591690 518378
rect 591070 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 591690 518294
rect 591070 482614 591690 518058
rect 591070 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 591690 482614
rect 591070 482294 591690 482378
rect 591070 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 591690 482294
rect 591070 446614 591690 482058
rect 591070 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 591690 446614
rect 591070 446294 591690 446378
rect 591070 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 591690 446294
rect 591070 410614 591690 446058
rect 591070 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 591690 410614
rect 591070 410294 591690 410378
rect 591070 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 591690 410294
rect 591070 374614 591690 410058
rect 591070 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 591690 374614
rect 591070 374294 591690 374378
rect 591070 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 591690 374294
rect 591070 338614 591690 374058
rect 591070 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 591690 338614
rect 591070 338294 591690 338378
rect 591070 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 591690 338294
rect 591070 302614 591690 338058
rect 591070 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 591690 302614
rect 591070 302294 591690 302378
rect 591070 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 591690 302294
rect 591070 266614 591690 302058
rect 591070 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 591690 266614
rect 591070 266294 591690 266378
rect 591070 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 591690 266294
rect 591070 230614 591690 266058
rect 591070 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 591690 230614
rect 591070 230294 591690 230378
rect 591070 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 591690 230294
rect 591070 194614 591690 230058
rect 591070 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 591690 194614
rect 591070 194294 591690 194378
rect 591070 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 591690 194294
rect 591070 158614 591690 194058
rect 591070 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 591690 158614
rect 591070 158294 591690 158378
rect 591070 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 591690 158294
rect 591070 122614 591690 158058
rect 591070 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 591690 122614
rect 591070 122294 591690 122378
rect 591070 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 591690 122294
rect 591070 86614 591690 122058
rect 591070 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 591690 86614
rect 591070 86294 591690 86378
rect 591070 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 591690 86294
rect 591070 50614 591690 86058
rect 591070 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 591690 50614
rect 591070 50294 591690 50378
rect 591070 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 591690 50294
rect 591070 14614 591690 50058
rect 591070 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 591690 14614
rect 591070 14294 591690 14378
rect 591070 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 591690 14294
rect 591070 -6106 591690 14058
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 680614 592650 711002
rect 592030 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect 592030 680294 592650 680378
rect 592030 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect 592030 644614 592650 680058
rect 592030 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect 592030 644294 592650 644378
rect 592030 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect 592030 608614 592650 644058
rect 592030 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect 592030 608294 592650 608378
rect 592030 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect 592030 572614 592650 608058
rect 592030 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect 592030 572294 592650 572378
rect 592030 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect 592030 536614 592650 572058
rect 592030 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect 592030 536294 592650 536378
rect 592030 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect 592030 500614 592650 536058
rect 592030 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect 592030 500294 592650 500378
rect 592030 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect 592030 464614 592650 500058
rect 592030 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect 592030 464294 592650 464378
rect 592030 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect 592030 428614 592650 464058
rect 592030 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect 592030 428294 592650 428378
rect 592030 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect 592030 392614 592650 428058
rect 592030 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect 592030 392294 592650 392378
rect 592030 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect 592030 356614 592650 392058
rect 592030 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect 592030 356294 592650 356378
rect 592030 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect 592030 320614 592650 356058
rect 592030 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect 592030 320294 592650 320378
rect 592030 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect 592030 284614 592650 320058
rect 592030 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect 592030 284294 592650 284378
rect 592030 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect 592030 248614 592650 284058
rect 592030 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect 592030 248294 592650 248378
rect 592030 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect 592030 212614 592650 248058
rect 592030 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect 592030 212294 592650 212378
rect 592030 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect 592030 176614 592650 212058
rect 592030 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect 592030 176294 592650 176378
rect 592030 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect 592030 140614 592650 176058
rect 592030 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect 592030 140294 592650 140378
rect 592030 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect 592030 104614 592650 140058
rect 592030 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect 592030 104294 592650 104378
rect 592030 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect 592030 68614 592650 104058
rect 592030 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect 592030 68294 592650 68378
rect 592030 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect 592030 32614 592650 68058
rect 592030 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect 592030 32294 592650 32378
rect 592030 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect 570954 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 571574 -7066
rect 570954 -7386 571574 -7302
rect 570954 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 571574 -7386
rect 570954 -7654 571574 -7622
rect 592030 -7066 592650 32058
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 680378 -8458 680614
rect -8374 680378 -8138 680614
rect -8694 680058 -8458 680294
rect -8374 680058 -8138 680294
rect -8694 644378 -8458 644614
rect -8374 644378 -8138 644614
rect -8694 644058 -8458 644294
rect -8374 644058 -8138 644294
rect -8694 608378 -8458 608614
rect -8374 608378 -8138 608614
rect -8694 608058 -8458 608294
rect -8374 608058 -8138 608294
rect -8694 572378 -8458 572614
rect -8374 572378 -8138 572614
rect -8694 572058 -8458 572294
rect -8374 572058 -8138 572294
rect -8694 536378 -8458 536614
rect -8374 536378 -8138 536614
rect -8694 536058 -8458 536294
rect -8374 536058 -8138 536294
rect -8694 500378 -8458 500614
rect -8374 500378 -8138 500614
rect -8694 500058 -8458 500294
rect -8374 500058 -8138 500294
rect -8694 464378 -8458 464614
rect -8374 464378 -8138 464614
rect -8694 464058 -8458 464294
rect -8374 464058 -8138 464294
rect -8694 428378 -8458 428614
rect -8374 428378 -8138 428614
rect -8694 428058 -8458 428294
rect -8374 428058 -8138 428294
rect -8694 392378 -8458 392614
rect -8374 392378 -8138 392614
rect -8694 392058 -8458 392294
rect -8374 392058 -8138 392294
rect -8694 356378 -8458 356614
rect -8374 356378 -8138 356614
rect -8694 356058 -8458 356294
rect -8374 356058 -8138 356294
rect -8694 320378 -8458 320614
rect -8374 320378 -8138 320614
rect -8694 320058 -8458 320294
rect -8374 320058 -8138 320294
rect -8694 284378 -8458 284614
rect -8374 284378 -8138 284614
rect -8694 284058 -8458 284294
rect -8374 284058 -8138 284294
rect -8694 248378 -8458 248614
rect -8374 248378 -8138 248614
rect -8694 248058 -8458 248294
rect -8374 248058 -8138 248294
rect -8694 212378 -8458 212614
rect -8374 212378 -8138 212614
rect -8694 212058 -8458 212294
rect -8374 212058 -8138 212294
rect -8694 176378 -8458 176614
rect -8374 176378 -8138 176614
rect -8694 176058 -8458 176294
rect -8374 176058 -8138 176294
rect -8694 140378 -8458 140614
rect -8374 140378 -8138 140614
rect -8694 140058 -8458 140294
rect -8374 140058 -8138 140294
rect -8694 104378 -8458 104614
rect -8374 104378 -8138 104614
rect -8694 104058 -8458 104294
rect -8374 104058 -8138 104294
rect -8694 68378 -8458 68614
rect -8374 68378 -8138 68614
rect -8694 68058 -8458 68294
rect -8374 68058 -8138 68294
rect -8694 32378 -8458 32614
rect -8374 32378 -8138 32614
rect -8694 32058 -8458 32294
rect -8374 32058 -8138 32294
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect 12986 710362 13222 710598
rect 13306 710362 13542 710598
rect 12986 710042 13222 710278
rect 13306 710042 13542 710278
rect -7734 698378 -7498 698614
rect -7414 698378 -7178 698614
rect -7734 698058 -7498 698294
rect -7414 698058 -7178 698294
rect -7734 662378 -7498 662614
rect -7414 662378 -7178 662614
rect -7734 662058 -7498 662294
rect -7414 662058 -7178 662294
rect -7734 626378 -7498 626614
rect -7414 626378 -7178 626614
rect -7734 626058 -7498 626294
rect -7414 626058 -7178 626294
rect -7734 590378 -7498 590614
rect -7414 590378 -7178 590614
rect -7734 590058 -7498 590294
rect -7414 590058 -7178 590294
rect -7734 554378 -7498 554614
rect -7414 554378 -7178 554614
rect -7734 554058 -7498 554294
rect -7414 554058 -7178 554294
rect -7734 518378 -7498 518614
rect -7414 518378 -7178 518614
rect -7734 518058 -7498 518294
rect -7414 518058 -7178 518294
rect -7734 482378 -7498 482614
rect -7414 482378 -7178 482614
rect -7734 482058 -7498 482294
rect -7414 482058 -7178 482294
rect -7734 446378 -7498 446614
rect -7414 446378 -7178 446614
rect -7734 446058 -7498 446294
rect -7414 446058 -7178 446294
rect -7734 410378 -7498 410614
rect -7414 410378 -7178 410614
rect -7734 410058 -7498 410294
rect -7414 410058 -7178 410294
rect -7734 374378 -7498 374614
rect -7414 374378 -7178 374614
rect -7734 374058 -7498 374294
rect -7414 374058 -7178 374294
rect -7734 338378 -7498 338614
rect -7414 338378 -7178 338614
rect -7734 338058 -7498 338294
rect -7414 338058 -7178 338294
rect -7734 302378 -7498 302614
rect -7414 302378 -7178 302614
rect -7734 302058 -7498 302294
rect -7414 302058 -7178 302294
rect -7734 266378 -7498 266614
rect -7414 266378 -7178 266614
rect -7734 266058 -7498 266294
rect -7414 266058 -7178 266294
rect -7734 230378 -7498 230614
rect -7414 230378 -7178 230614
rect -7734 230058 -7498 230294
rect -7414 230058 -7178 230294
rect -7734 194378 -7498 194614
rect -7414 194378 -7178 194614
rect -7734 194058 -7498 194294
rect -7414 194058 -7178 194294
rect -7734 158378 -7498 158614
rect -7414 158378 -7178 158614
rect -7734 158058 -7498 158294
rect -7414 158058 -7178 158294
rect -7734 122378 -7498 122614
rect -7414 122378 -7178 122614
rect -7734 122058 -7498 122294
rect -7414 122058 -7178 122294
rect -7734 86378 -7498 86614
rect -7414 86378 -7178 86614
rect -7734 86058 -7498 86294
rect -7414 86058 -7178 86294
rect -7734 50378 -7498 50614
rect -7414 50378 -7178 50614
rect -7734 50058 -7498 50294
rect -7414 50058 -7178 50294
rect -7734 14378 -7498 14614
rect -7414 14378 -7178 14614
rect -7734 14058 -7498 14294
rect -7414 14058 -7178 14294
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 676658 -6538 676894
rect -6454 676658 -6218 676894
rect -6774 676338 -6538 676574
rect -6454 676338 -6218 676574
rect -6774 640658 -6538 640894
rect -6454 640658 -6218 640894
rect -6774 640338 -6538 640574
rect -6454 640338 -6218 640574
rect -6774 604658 -6538 604894
rect -6454 604658 -6218 604894
rect -6774 604338 -6538 604574
rect -6454 604338 -6218 604574
rect -6774 568658 -6538 568894
rect -6454 568658 -6218 568894
rect -6774 568338 -6538 568574
rect -6454 568338 -6218 568574
rect -6774 532658 -6538 532894
rect -6454 532658 -6218 532894
rect -6774 532338 -6538 532574
rect -6454 532338 -6218 532574
rect -6774 496658 -6538 496894
rect -6454 496658 -6218 496894
rect -6774 496338 -6538 496574
rect -6454 496338 -6218 496574
rect -6774 460658 -6538 460894
rect -6454 460658 -6218 460894
rect -6774 460338 -6538 460574
rect -6454 460338 -6218 460574
rect -6774 424658 -6538 424894
rect -6454 424658 -6218 424894
rect -6774 424338 -6538 424574
rect -6454 424338 -6218 424574
rect -6774 388658 -6538 388894
rect -6454 388658 -6218 388894
rect -6774 388338 -6538 388574
rect -6454 388338 -6218 388574
rect -6774 352658 -6538 352894
rect -6454 352658 -6218 352894
rect -6774 352338 -6538 352574
rect -6454 352338 -6218 352574
rect -6774 316658 -6538 316894
rect -6454 316658 -6218 316894
rect -6774 316338 -6538 316574
rect -6454 316338 -6218 316574
rect -6774 280658 -6538 280894
rect -6454 280658 -6218 280894
rect -6774 280338 -6538 280574
rect -6454 280338 -6218 280574
rect -6774 244658 -6538 244894
rect -6454 244658 -6218 244894
rect -6774 244338 -6538 244574
rect -6454 244338 -6218 244574
rect -6774 208658 -6538 208894
rect -6454 208658 -6218 208894
rect -6774 208338 -6538 208574
rect -6454 208338 -6218 208574
rect -6774 172658 -6538 172894
rect -6454 172658 -6218 172894
rect -6774 172338 -6538 172574
rect -6454 172338 -6218 172574
rect -6774 136658 -6538 136894
rect -6454 136658 -6218 136894
rect -6774 136338 -6538 136574
rect -6454 136338 -6218 136574
rect -6774 100658 -6538 100894
rect -6454 100658 -6218 100894
rect -6774 100338 -6538 100574
rect -6454 100338 -6218 100574
rect -6774 64658 -6538 64894
rect -6454 64658 -6218 64894
rect -6774 64338 -6538 64574
rect -6454 64338 -6218 64574
rect -6774 28658 -6538 28894
rect -6454 28658 -6218 28894
rect -6774 28338 -6538 28574
rect -6454 28338 -6218 28574
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect 9266 708442 9502 708678
rect 9586 708442 9822 708678
rect 9266 708122 9502 708358
rect 9586 708122 9822 708358
rect -5814 694658 -5578 694894
rect -5494 694658 -5258 694894
rect -5814 694338 -5578 694574
rect -5494 694338 -5258 694574
rect -5814 658658 -5578 658894
rect -5494 658658 -5258 658894
rect -5814 658338 -5578 658574
rect -5494 658338 -5258 658574
rect -5814 622658 -5578 622894
rect -5494 622658 -5258 622894
rect -5814 622338 -5578 622574
rect -5494 622338 -5258 622574
rect -5814 586658 -5578 586894
rect -5494 586658 -5258 586894
rect -5814 586338 -5578 586574
rect -5494 586338 -5258 586574
rect -5814 550658 -5578 550894
rect -5494 550658 -5258 550894
rect -5814 550338 -5578 550574
rect -5494 550338 -5258 550574
rect -5814 514658 -5578 514894
rect -5494 514658 -5258 514894
rect -5814 514338 -5578 514574
rect -5494 514338 -5258 514574
rect -5814 478658 -5578 478894
rect -5494 478658 -5258 478894
rect -5814 478338 -5578 478574
rect -5494 478338 -5258 478574
rect -5814 442658 -5578 442894
rect -5494 442658 -5258 442894
rect -5814 442338 -5578 442574
rect -5494 442338 -5258 442574
rect -5814 406658 -5578 406894
rect -5494 406658 -5258 406894
rect -5814 406338 -5578 406574
rect -5494 406338 -5258 406574
rect -5814 370658 -5578 370894
rect -5494 370658 -5258 370894
rect -5814 370338 -5578 370574
rect -5494 370338 -5258 370574
rect -5814 334658 -5578 334894
rect -5494 334658 -5258 334894
rect -5814 334338 -5578 334574
rect -5494 334338 -5258 334574
rect -5814 298658 -5578 298894
rect -5494 298658 -5258 298894
rect -5814 298338 -5578 298574
rect -5494 298338 -5258 298574
rect -5814 262658 -5578 262894
rect -5494 262658 -5258 262894
rect -5814 262338 -5578 262574
rect -5494 262338 -5258 262574
rect -5814 226658 -5578 226894
rect -5494 226658 -5258 226894
rect -5814 226338 -5578 226574
rect -5494 226338 -5258 226574
rect -5814 190658 -5578 190894
rect -5494 190658 -5258 190894
rect -5814 190338 -5578 190574
rect -5494 190338 -5258 190574
rect -5814 154658 -5578 154894
rect -5494 154658 -5258 154894
rect -5814 154338 -5578 154574
rect -5494 154338 -5258 154574
rect -5814 118658 -5578 118894
rect -5494 118658 -5258 118894
rect -5814 118338 -5578 118574
rect -5494 118338 -5258 118574
rect -5814 82658 -5578 82894
rect -5494 82658 -5258 82894
rect -5814 82338 -5578 82574
rect -5494 82338 -5258 82574
rect -5814 46658 -5578 46894
rect -5494 46658 -5258 46894
rect -5814 46338 -5578 46574
rect -5494 46338 -5258 46574
rect -5814 10658 -5578 10894
rect -5494 10658 -5258 10894
rect -5814 10338 -5578 10574
rect -5494 10338 -5258 10574
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 672938 -4618 673174
rect -4534 672938 -4298 673174
rect -4854 672618 -4618 672854
rect -4534 672618 -4298 672854
rect -4854 636938 -4618 637174
rect -4534 636938 -4298 637174
rect -4854 636618 -4618 636854
rect -4534 636618 -4298 636854
rect -4854 600938 -4618 601174
rect -4534 600938 -4298 601174
rect -4854 600618 -4618 600854
rect -4534 600618 -4298 600854
rect -4854 564938 -4618 565174
rect -4534 564938 -4298 565174
rect -4854 564618 -4618 564854
rect -4534 564618 -4298 564854
rect -4854 528938 -4618 529174
rect -4534 528938 -4298 529174
rect -4854 528618 -4618 528854
rect -4534 528618 -4298 528854
rect -4854 492938 -4618 493174
rect -4534 492938 -4298 493174
rect -4854 492618 -4618 492854
rect -4534 492618 -4298 492854
rect -4854 456938 -4618 457174
rect -4534 456938 -4298 457174
rect -4854 456618 -4618 456854
rect -4534 456618 -4298 456854
rect -4854 420938 -4618 421174
rect -4534 420938 -4298 421174
rect -4854 420618 -4618 420854
rect -4534 420618 -4298 420854
rect -4854 384938 -4618 385174
rect -4534 384938 -4298 385174
rect -4854 384618 -4618 384854
rect -4534 384618 -4298 384854
rect -4854 348938 -4618 349174
rect -4534 348938 -4298 349174
rect -4854 348618 -4618 348854
rect -4534 348618 -4298 348854
rect -4854 312938 -4618 313174
rect -4534 312938 -4298 313174
rect -4854 312618 -4618 312854
rect -4534 312618 -4298 312854
rect -4854 276938 -4618 277174
rect -4534 276938 -4298 277174
rect -4854 276618 -4618 276854
rect -4534 276618 -4298 276854
rect -4854 240938 -4618 241174
rect -4534 240938 -4298 241174
rect -4854 240618 -4618 240854
rect -4534 240618 -4298 240854
rect -4854 204938 -4618 205174
rect -4534 204938 -4298 205174
rect -4854 204618 -4618 204854
rect -4534 204618 -4298 204854
rect -4854 168938 -4618 169174
rect -4534 168938 -4298 169174
rect -4854 168618 -4618 168854
rect -4534 168618 -4298 168854
rect -4854 132938 -4618 133174
rect -4534 132938 -4298 133174
rect -4854 132618 -4618 132854
rect -4534 132618 -4298 132854
rect -4854 96938 -4618 97174
rect -4534 96938 -4298 97174
rect -4854 96618 -4618 96854
rect -4534 96618 -4298 96854
rect -4854 60938 -4618 61174
rect -4534 60938 -4298 61174
rect -4854 60618 -4618 60854
rect -4534 60618 -4298 60854
rect -4854 24938 -4618 25174
rect -4534 24938 -4298 25174
rect -4854 24618 -4618 24854
rect -4534 24618 -4298 24854
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect 5546 706522 5782 706758
rect 5866 706522 6102 706758
rect 5546 706202 5782 706438
rect 5866 706202 6102 706438
rect -3894 690938 -3658 691174
rect -3574 690938 -3338 691174
rect -3894 690618 -3658 690854
rect -3574 690618 -3338 690854
rect -3894 654938 -3658 655174
rect -3574 654938 -3338 655174
rect -3894 654618 -3658 654854
rect -3574 654618 -3338 654854
rect -3894 618938 -3658 619174
rect -3574 618938 -3338 619174
rect -3894 618618 -3658 618854
rect -3574 618618 -3338 618854
rect -3894 582938 -3658 583174
rect -3574 582938 -3338 583174
rect -3894 582618 -3658 582854
rect -3574 582618 -3338 582854
rect -3894 546938 -3658 547174
rect -3574 546938 -3338 547174
rect -3894 546618 -3658 546854
rect -3574 546618 -3338 546854
rect -3894 510938 -3658 511174
rect -3574 510938 -3338 511174
rect -3894 510618 -3658 510854
rect -3574 510618 -3338 510854
rect -3894 474938 -3658 475174
rect -3574 474938 -3338 475174
rect -3894 474618 -3658 474854
rect -3574 474618 -3338 474854
rect -3894 438938 -3658 439174
rect -3574 438938 -3338 439174
rect -3894 438618 -3658 438854
rect -3574 438618 -3338 438854
rect -3894 402938 -3658 403174
rect -3574 402938 -3338 403174
rect -3894 402618 -3658 402854
rect -3574 402618 -3338 402854
rect -3894 366938 -3658 367174
rect -3574 366938 -3338 367174
rect -3894 366618 -3658 366854
rect -3574 366618 -3338 366854
rect -3894 330938 -3658 331174
rect -3574 330938 -3338 331174
rect -3894 330618 -3658 330854
rect -3574 330618 -3338 330854
rect -3894 294938 -3658 295174
rect -3574 294938 -3338 295174
rect -3894 294618 -3658 294854
rect -3574 294618 -3338 294854
rect -3894 258938 -3658 259174
rect -3574 258938 -3338 259174
rect -3894 258618 -3658 258854
rect -3574 258618 -3338 258854
rect -3894 222938 -3658 223174
rect -3574 222938 -3338 223174
rect -3894 222618 -3658 222854
rect -3574 222618 -3338 222854
rect -3894 186938 -3658 187174
rect -3574 186938 -3338 187174
rect -3894 186618 -3658 186854
rect -3574 186618 -3338 186854
rect -3894 150938 -3658 151174
rect -3574 150938 -3338 151174
rect -3894 150618 -3658 150854
rect -3574 150618 -3338 150854
rect -3894 114938 -3658 115174
rect -3574 114938 -3338 115174
rect -3894 114618 -3658 114854
rect -3574 114618 -3338 114854
rect -3894 78938 -3658 79174
rect -3574 78938 -3338 79174
rect -3894 78618 -3658 78854
rect -3574 78618 -3338 78854
rect -3894 42938 -3658 43174
rect -3574 42938 -3338 43174
rect -3894 42618 -3658 42854
rect -3574 42618 -3338 42854
rect -3894 6938 -3658 7174
rect -3574 6938 -3338 7174
rect -3894 6618 -3658 6854
rect -3574 6618 -3338 6854
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 669218 -2698 669454
rect -2614 669218 -2378 669454
rect -2934 668898 -2698 669134
rect -2614 668898 -2378 669134
rect -2934 633218 -2698 633454
rect -2614 633218 -2378 633454
rect -2934 632898 -2698 633134
rect -2614 632898 -2378 633134
rect -2934 597218 -2698 597454
rect -2614 597218 -2378 597454
rect -2934 596898 -2698 597134
rect -2614 596898 -2378 597134
rect -2934 561218 -2698 561454
rect -2614 561218 -2378 561454
rect -2934 560898 -2698 561134
rect -2614 560898 -2378 561134
rect -2934 525218 -2698 525454
rect -2614 525218 -2378 525454
rect -2934 524898 -2698 525134
rect -2614 524898 -2378 525134
rect -2934 489218 -2698 489454
rect -2614 489218 -2378 489454
rect -2934 488898 -2698 489134
rect -2614 488898 -2378 489134
rect -2934 453218 -2698 453454
rect -2614 453218 -2378 453454
rect -2934 452898 -2698 453134
rect -2614 452898 -2378 453134
rect -2934 417218 -2698 417454
rect -2614 417218 -2378 417454
rect -2934 416898 -2698 417134
rect -2614 416898 -2378 417134
rect -2934 381218 -2698 381454
rect -2614 381218 -2378 381454
rect -2934 380898 -2698 381134
rect -2614 380898 -2378 381134
rect -2934 345218 -2698 345454
rect -2614 345218 -2378 345454
rect -2934 344898 -2698 345134
rect -2614 344898 -2378 345134
rect -2934 309218 -2698 309454
rect -2614 309218 -2378 309454
rect -2934 308898 -2698 309134
rect -2614 308898 -2378 309134
rect -2934 273218 -2698 273454
rect -2614 273218 -2378 273454
rect -2934 272898 -2698 273134
rect -2614 272898 -2378 273134
rect -2934 237218 -2698 237454
rect -2614 237218 -2378 237454
rect -2934 236898 -2698 237134
rect -2614 236898 -2378 237134
rect -2934 201218 -2698 201454
rect -2614 201218 -2378 201454
rect -2934 200898 -2698 201134
rect -2614 200898 -2378 201134
rect -2934 165218 -2698 165454
rect -2614 165218 -2378 165454
rect -2934 164898 -2698 165134
rect -2614 164898 -2378 165134
rect -2934 129218 -2698 129454
rect -2614 129218 -2378 129454
rect -2934 128898 -2698 129134
rect -2614 128898 -2378 129134
rect -2934 93218 -2698 93454
rect -2614 93218 -2378 93454
rect -2934 92898 -2698 93134
rect -2614 92898 -2378 93134
rect -2934 57218 -2698 57454
rect -2614 57218 -2378 57454
rect -2934 56898 -2698 57134
rect -2614 56898 -2378 57134
rect -2934 21218 -2698 21454
rect -2614 21218 -2378 21454
rect -2934 20898 -2698 21134
rect -2614 20898 -2378 21134
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect 5546 -2502 5782 -2266
rect 5866 -2502 6102 -2266
rect 5546 -2822 5782 -2586
rect 5866 -2822 6102 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect 9266 694658 9502 694894
rect 9586 694658 9822 694894
rect 9266 694338 9502 694574
rect 9586 694338 9822 694574
rect 9266 658658 9502 658894
rect 9586 658658 9822 658894
rect 9266 658338 9502 658574
rect 9586 658338 9822 658574
rect 9266 622658 9502 622894
rect 9586 622658 9822 622894
rect 9266 622338 9502 622574
rect 9586 622338 9822 622574
rect 9266 586658 9502 586894
rect 9586 586658 9822 586894
rect 9266 586338 9502 586574
rect 9586 586338 9822 586574
rect 9266 550658 9502 550894
rect 9586 550658 9822 550894
rect 9266 550338 9502 550574
rect 9586 550338 9822 550574
rect 9266 514658 9502 514894
rect 9586 514658 9822 514894
rect 9266 514338 9502 514574
rect 9586 514338 9822 514574
rect 9266 478658 9502 478894
rect 9586 478658 9822 478894
rect 9266 478338 9502 478574
rect 9586 478338 9822 478574
rect 9266 442658 9502 442894
rect 9586 442658 9822 442894
rect 9266 442338 9502 442574
rect 9586 442338 9822 442574
rect 9266 406658 9502 406894
rect 9586 406658 9822 406894
rect 9266 406338 9502 406574
rect 9586 406338 9822 406574
rect 9266 370658 9502 370894
rect 9586 370658 9822 370894
rect 9266 370338 9502 370574
rect 9586 370338 9822 370574
rect 9266 334658 9502 334894
rect 9586 334658 9822 334894
rect 9266 334338 9502 334574
rect 9586 334338 9822 334574
rect 9266 298658 9502 298894
rect 9586 298658 9822 298894
rect 9266 298338 9502 298574
rect 9586 298338 9822 298574
rect 9266 262658 9502 262894
rect 9586 262658 9822 262894
rect 9266 262338 9502 262574
rect 9586 262338 9822 262574
rect 9266 226658 9502 226894
rect 9586 226658 9822 226894
rect 9266 226338 9502 226574
rect 9586 226338 9822 226574
rect 9266 190658 9502 190894
rect 9586 190658 9822 190894
rect 9266 190338 9502 190574
rect 9586 190338 9822 190574
rect 9266 154658 9502 154894
rect 9586 154658 9822 154894
rect 9266 154338 9502 154574
rect 9586 154338 9822 154574
rect 9266 118658 9502 118894
rect 9586 118658 9822 118894
rect 9266 118338 9502 118574
rect 9586 118338 9822 118574
rect 9266 82658 9502 82894
rect 9586 82658 9822 82894
rect 9266 82338 9502 82574
rect 9586 82338 9822 82574
rect 9266 46658 9502 46894
rect 9586 46658 9822 46894
rect 9266 46338 9502 46574
rect 9586 46338 9822 46574
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect 9266 -4422 9502 -4186
rect 9586 -4422 9822 -4186
rect 9266 -4742 9502 -4506
rect 9586 -4742 9822 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect 30986 711322 31222 711558
rect 31306 711322 31542 711558
rect 30986 711002 31222 711238
rect 31306 711002 31542 711238
rect 27266 709402 27502 709638
rect 27586 709402 27822 709638
rect 27266 709082 27502 709318
rect 27586 709082 27822 709318
rect 23546 707482 23782 707718
rect 23866 707482 24102 707718
rect 23546 707162 23782 707398
rect 23866 707162 24102 707398
rect 12986 698378 13222 698614
rect 13306 698378 13542 698614
rect 12986 698058 13222 698294
rect 13306 698058 13542 698294
rect 12986 662378 13222 662614
rect 13306 662378 13542 662614
rect 12986 662058 13222 662294
rect 13306 662058 13542 662294
rect 12986 626378 13222 626614
rect 13306 626378 13542 626614
rect 12986 626058 13222 626294
rect 13306 626058 13542 626294
rect 12986 590378 13222 590614
rect 13306 590378 13542 590614
rect 12986 590058 13222 590294
rect 13306 590058 13542 590294
rect 12986 554378 13222 554614
rect 13306 554378 13542 554614
rect 12986 554058 13222 554294
rect 13306 554058 13542 554294
rect 12986 518378 13222 518614
rect 13306 518378 13542 518614
rect 12986 518058 13222 518294
rect 13306 518058 13542 518294
rect 12986 482378 13222 482614
rect 13306 482378 13542 482614
rect 12986 482058 13222 482294
rect 13306 482058 13542 482294
rect 12986 446378 13222 446614
rect 13306 446378 13542 446614
rect 12986 446058 13222 446294
rect 13306 446058 13542 446294
rect 12986 410378 13222 410614
rect 13306 410378 13542 410614
rect 12986 410058 13222 410294
rect 13306 410058 13542 410294
rect 12986 374378 13222 374614
rect 13306 374378 13542 374614
rect 12986 374058 13222 374294
rect 13306 374058 13542 374294
rect 12986 338378 13222 338614
rect 13306 338378 13542 338614
rect 12986 338058 13222 338294
rect 13306 338058 13542 338294
rect 12986 302378 13222 302614
rect 13306 302378 13542 302614
rect 12986 302058 13222 302294
rect 13306 302058 13542 302294
rect 12986 266378 13222 266614
rect 13306 266378 13542 266614
rect 12986 266058 13222 266294
rect 13306 266058 13542 266294
rect 12986 230378 13222 230614
rect 13306 230378 13542 230614
rect 12986 230058 13222 230294
rect 13306 230058 13542 230294
rect 12986 194378 13222 194614
rect 13306 194378 13542 194614
rect 12986 194058 13222 194294
rect 13306 194058 13542 194294
rect 12986 158378 13222 158614
rect 13306 158378 13542 158614
rect 12986 158058 13222 158294
rect 13306 158058 13542 158294
rect 12986 122378 13222 122614
rect 13306 122378 13542 122614
rect 12986 122058 13222 122294
rect 13306 122058 13542 122294
rect 12986 86378 13222 86614
rect 13306 86378 13542 86614
rect 12986 86058 13222 86294
rect 13306 86058 13542 86294
rect 12986 50378 13222 50614
rect 13306 50378 13542 50614
rect 12986 50058 13222 50294
rect 13306 50058 13542 50294
rect 12986 14378 13222 14614
rect 13306 14378 13542 14614
rect 12986 14058 13222 14294
rect 13306 14058 13542 14294
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect 19826 705562 20062 705798
rect 20146 705562 20382 705798
rect 19826 705242 20062 705478
rect 20146 705242 20382 705478
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -1542 20062 -1306
rect 20146 -1542 20382 -1306
rect 19826 -1862 20062 -1626
rect 20146 -1862 20382 -1626
rect 23546 672938 23782 673174
rect 23866 672938 24102 673174
rect 23546 672618 23782 672854
rect 23866 672618 24102 672854
rect 23546 636938 23782 637174
rect 23866 636938 24102 637174
rect 23546 636618 23782 636854
rect 23866 636618 24102 636854
rect 23546 600938 23782 601174
rect 23866 600938 24102 601174
rect 23546 600618 23782 600854
rect 23866 600618 24102 600854
rect 23546 564938 23782 565174
rect 23866 564938 24102 565174
rect 23546 564618 23782 564854
rect 23866 564618 24102 564854
rect 23546 528938 23782 529174
rect 23866 528938 24102 529174
rect 23546 528618 23782 528854
rect 23866 528618 24102 528854
rect 23546 492938 23782 493174
rect 23866 492938 24102 493174
rect 23546 492618 23782 492854
rect 23866 492618 24102 492854
rect 23546 456938 23782 457174
rect 23866 456938 24102 457174
rect 23546 456618 23782 456854
rect 23866 456618 24102 456854
rect 23546 420938 23782 421174
rect 23866 420938 24102 421174
rect 23546 420618 23782 420854
rect 23866 420618 24102 420854
rect 23546 384938 23782 385174
rect 23866 384938 24102 385174
rect 23546 384618 23782 384854
rect 23866 384618 24102 384854
rect 23546 348938 23782 349174
rect 23866 348938 24102 349174
rect 23546 348618 23782 348854
rect 23866 348618 24102 348854
rect 23546 312938 23782 313174
rect 23866 312938 24102 313174
rect 23546 312618 23782 312854
rect 23866 312618 24102 312854
rect 23546 276938 23782 277174
rect 23866 276938 24102 277174
rect 23546 276618 23782 276854
rect 23866 276618 24102 276854
rect 23546 240938 23782 241174
rect 23866 240938 24102 241174
rect 23546 240618 23782 240854
rect 23866 240618 24102 240854
rect 23546 204938 23782 205174
rect 23866 204938 24102 205174
rect 23546 204618 23782 204854
rect 23866 204618 24102 204854
rect 23546 168938 23782 169174
rect 23866 168938 24102 169174
rect 23546 168618 23782 168854
rect 23866 168618 24102 168854
rect 23546 132938 23782 133174
rect 23866 132938 24102 133174
rect 23546 132618 23782 132854
rect 23866 132618 24102 132854
rect 23546 96938 23782 97174
rect 23866 96938 24102 97174
rect 23546 96618 23782 96854
rect 23866 96618 24102 96854
rect 23546 60938 23782 61174
rect 23866 60938 24102 61174
rect 23546 60618 23782 60854
rect 23866 60618 24102 60854
rect 23546 24938 23782 25174
rect 23866 24938 24102 25174
rect 23546 24618 23782 24854
rect 23866 24618 24102 24854
rect 23546 -3462 23782 -3226
rect 23866 -3462 24102 -3226
rect 23546 -3782 23782 -3546
rect 23866 -3782 24102 -3546
rect 27266 676658 27502 676894
rect 27586 676658 27822 676894
rect 27266 676338 27502 676574
rect 27586 676338 27822 676574
rect 27266 640658 27502 640894
rect 27586 640658 27822 640894
rect 27266 640338 27502 640574
rect 27586 640338 27822 640574
rect 27266 604658 27502 604894
rect 27586 604658 27822 604894
rect 27266 604338 27502 604574
rect 27586 604338 27822 604574
rect 27266 568658 27502 568894
rect 27586 568658 27822 568894
rect 27266 568338 27502 568574
rect 27586 568338 27822 568574
rect 27266 532658 27502 532894
rect 27586 532658 27822 532894
rect 27266 532338 27502 532574
rect 27586 532338 27822 532574
rect 27266 496658 27502 496894
rect 27586 496658 27822 496894
rect 27266 496338 27502 496574
rect 27586 496338 27822 496574
rect 27266 460658 27502 460894
rect 27586 460658 27822 460894
rect 27266 460338 27502 460574
rect 27586 460338 27822 460574
rect 27266 424658 27502 424894
rect 27586 424658 27822 424894
rect 27266 424338 27502 424574
rect 27586 424338 27822 424574
rect 27266 388658 27502 388894
rect 27586 388658 27822 388894
rect 27266 388338 27502 388574
rect 27586 388338 27822 388574
rect 27266 352658 27502 352894
rect 27586 352658 27822 352894
rect 27266 352338 27502 352574
rect 27586 352338 27822 352574
rect 27266 316658 27502 316894
rect 27586 316658 27822 316894
rect 27266 316338 27502 316574
rect 27586 316338 27822 316574
rect 27266 280658 27502 280894
rect 27586 280658 27822 280894
rect 27266 280338 27502 280574
rect 27586 280338 27822 280574
rect 27266 244658 27502 244894
rect 27586 244658 27822 244894
rect 27266 244338 27502 244574
rect 27586 244338 27822 244574
rect 27266 208658 27502 208894
rect 27586 208658 27822 208894
rect 27266 208338 27502 208574
rect 27586 208338 27822 208574
rect 27266 172658 27502 172894
rect 27586 172658 27822 172894
rect 27266 172338 27502 172574
rect 27586 172338 27822 172574
rect 27266 136658 27502 136894
rect 27586 136658 27822 136894
rect 27266 136338 27502 136574
rect 27586 136338 27822 136574
rect 27266 100658 27502 100894
rect 27586 100658 27822 100894
rect 27266 100338 27502 100574
rect 27586 100338 27822 100574
rect 27266 64658 27502 64894
rect 27586 64658 27822 64894
rect 27266 64338 27502 64574
rect 27586 64338 27822 64574
rect 27266 28658 27502 28894
rect 27586 28658 27822 28894
rect 27266 28338 27502 28574
rect 27586 28338 27822 28574
rect 27266 -5382 27502 -5146
rect 27586 -5382 27822 -5146
rect 27266 -5702 27502 -5466
rect 27586 -5702 27822 -5466
rect 48986 710362 49222 710598
rect 49306 710362 49542 710598
rect 48986 710042 49222 710278
rect 49306 710042 49542 710278
rect 45266 708442 45502 708678
rect 45586 708442 45822 708678
rect 45266 708122 45502 708358
rect 45586 708122 45822 708358
rect 41546 706522 41782 706758
rect 41866 706522 42102 706758
rect 41546 706202 41782 706438
rect 41866 706202 42102 706438
rect 30986 680378 31222 680614
rect 31306 680378 31542 680614
rect 30986 680058 31222 680294
rect 31306 680058 31542 680294
rect 30986 644378 31222 644614
rect 31306 644378 31542 644614
rect 30986 644058 31222 644294
rect 31306 644058 31542 644294
rect 30986 608378 31222 608614
rect 31306 608378 31542 608614
rect 30986 608058 31222 608294
rect 31306 608058 31542 608294
rect 30986 572378 31222 572614
rect 31306 572378 31542 572614
rect 30986 572058 31222 572294
rect 31306 572058 31542 572294
rect 30986 536378 31222 536614
rect 31306 536378 31542 536614
rect 30986 536058 31222 536294
rect 31306 536058 31542 536294
rect 30986 500378 31222 500614
rect 31306 500378 31542 500614
rect 30986 500058 31222 500294
rect 31306 500058 31542 500294
rect 30986 464378 31222 464614
rect 31306 464378 31542 464614
rect 30986 464058 31222 464294
rect 31306 464058 31542 464294
rect 30986 428378 31222 428614
rect 31306 428378 31542 428614
rect 30986 428058 31222 428294
rect 31306 428058 31542 428294
rect 30986 392378 31222 392614
rect 31306 392378 31542 392614
rect 30986 392058 31222 392294
rect 31306 392058 31542 392294
rect 30986 356378 31222 356614
rect 31306 356378 31542 356614
rect 30986 356058 31222 356294
rect 31306 356058 31542 356294
rect 30986 320378 31222 320614
rect 31306 320378 31542 320614
rect 30986 320058 31222 320294
rect 31306 320058 31542 320294
rect 30986 284378 31222 284614
rect 31306 284378 31542 284614
rect 30986 284058 31222 284294
rect 31306 284058 31542 284294
rect 30986 248378 31222 248614
rect 31306 248378 31542 248614
rect 30986 248058 31222 248294
rect 31306 248058 31542 248294
rect 30986 212378 31222 212614
rect 31306 212378 31542 212614
rect 30986 212058 31222 212294
rect 31306 212058 31542 212294
rect 30986 176378 31222 176614
rect 31306 176378 31542 176614
rect 30986 176058 31222 176294
rect 31306 176058 31542 176294
rect 30986 140378 31222 140614
rect 31306 140378 31542 140614
rect 30986 140058 31222 140294
rect 31306 140058 31542 140294
rect 30986 104378 31222 104614
rect 31306 104378 31542 104614
rect 30986 104058 31222 104294
rect 31306 104058 31542 104294
rect 30986 68378 31222 68614
rect 31306 68378 31542 68614
rect 30986 68058 31222 68294
rect 31306 68058 31542 68294
rect 30986 32378 31222 32614
rect 31306 32378 31542 32614
rect 30986 32058 31222 32294
rect 31306 32058 31542 32294
rect 12986 -6342 13222 -6106
rect 13306 -6342 13542 -6106
rect 12986 -6662 13222 -6426
rect 13306 -6662 13542 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 41546 654938 41782 655174
rect 41866 654938 42102 655174
rect 41546 654618 41782 654854
rect 41866 654618 42102 654854
rect 41546 618938 41782 619174
rect 41866 618938 42102 619174
rect 41546 618618 41782 618854
rect 41866 618618 42102 618854
rect 41546 582938 41782 583174
rect 41866 582938 42102 583174
rect 41546 582618 41782 582854
rect 41866 582618 42102 582854
rect 41546 546938 41782 547174
rect 41866 546938 42102 547174
rect 41546 546618 41782 546854
rect 41866 546618 42102 546854
rect 41546 510938 41782 511174
rect 41866 510938 42102 511174
rect 41546 510618 41782 510854
rect 41866 510618 42102 510854
rect 41546 474938 41782 475174
rect 41866 474938 42102 475174
rect 41546 474618 41782 474854
rect 41866 474618 42102 474854
rect 41546 438938 41782 439174
rect 41866 438938 42102 439174
rect 41546 438618 41782 438854
rect 41866 438618 42102 438854
rect 41546 402938 41782 403174
rect 41866 402938 42102 403174
rect 41546 402618 41782 402854
rect 41866 402618 42102 402854
rect 41546 366938 41782 367174
rect 41866 366938 42102 367174
rect 41546 366618 41782 366854
rect 41866 366618 42102 366854
rect 41546 330938 41782 331174
rect 41866 330938 42102 331174
rect 41546 330618 41782 330854
rect 41866 330618 42102 330854
rect 41546 294938 41782 295174
rect 41866 294938 42102 295174
rect 41546 294618 41782 294854
rect 41866 294618 42102 294854
rect 41546 258938 41782 259174
rect 41866 258938 42102 259174
rect 41546 258618 41782 258854
rect 41866 258618 42102 258854
rect 41546 222938 41782 223174
rect 41866 222938 42102 223174
rect 41546 222618 41782 222854
rect 41866 222618 42102 222854
rect 41546 186938 41782 187174
rect 41866 186938 42102 187174
rect 41546 186618 41782 186854
rect 41866 186618 42102 186854
rect 41546 150938 41782 151174
rect 41866 150938 42102 151174
rect 41546 150618 41782 150854
rect 41866 150618 42102 150854
rect 41546 114938 41782 115174
rect 41866 114938 42102 115174
rect 41546 114618 41782 114854
rect 41866 114618 42102 114854
rect 41546 78938 41782 79174
rect 41866 78938 42102 79174
rect 41546 78618 41782 78854
rect 41866 78618 42102 78854
rect 41546 42938 41782 43174
rect 41866 42938 42102 43174
rect 41546 42618 41782 42854
rect 41866 42618 42102 42854
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 41546 -2502 41782 -2266
rect 41866 -2502 42102 -2266
rect 41546 -2822 41782 -2586
rect 41866 -2822 42102 -2586
rect 45266 694658 45502 694894
rect 45586 694658 45822 694894
rect 45266 694338 45502 694574
rect 45586 694338 45822 694574
rect 45266 658658 45502 658894
rect 45586 658658 45822 658894
rect 45266 658338 45502 658574
rect 45586 658338 45822 658574
rect 45266 622658 45502 622894
rect 45586 622658 45822 622894
rect 45266 622338 45502 622574
rect 45586 622338 45822 622574
rect 45266 586658 45502 586894
rect 45586 586658 45822 586894
rect 45266 586338 45502 586574
rect 45586 586338 45822 586574
rect 45266 550658 45502 550894
rect 45586 550658 45822 550894
rect 45266 550338 45502 550574
rect 45586 550338 45822 550574
rect 45266 514658 45502 514894
rect 45586 514658 45822 514894
rect 45266 514338 45502 514574
rect 45586 514338 45822 514574
rect 45266 478658 45502 478894
rect 45586 478658 45822 478894
rect 45266 478338 45502 478574
rect 45586 478338 45822 478574
rect 45266 442658 45502 442894
rect 45586 442658 45822 442894
rect 45266 442338 45502 442574
rect 45586 442338 45822 442574
rect 45266 406658 45502 406894
rect 45586 406658 45822 406894
rect 45266 406338 45502 406574
rect 45586 406338 45822 406574
rect 45266 370658 45502 370894
rect 45586 370658 45822 370894
rect 45266 370338 45502 370574
rect 45586 370338 45822 370574
rect 45266 334658 45502 334894
rect 45586 334658 45822 334894
rect 45266 334338 45502 334574
rect 45586 334338 45822 334574
rect 45266 298658 45502 298894
rect 45586 298658 45822 298894
rect 45266 298338 45502 298574
rect 45586 298338 45822 298574
rect 45266 262658 45502 262894
rect 45586 262658 45822 262894
rect 45266 262338 45502 262574
rect 45586 262338 45822 262574
rect 45266 226658 45502 226894
rect 45586 226658 45822 226894
rect 45266 226338 45502 226574
rect 45586 226338 45822 226574
rect 45266 190658 45502 190894
rect 45586 190658 45822 190894
rect 45266 190338 45502 190574
rect 45586 190338 45822 190574
rect 45266 154658 45502 154894
rect 45586 154658 45822 154894
rect 45266 154338 45502 154574
rect 45586 154338 45822 154574
rect 45266 118658 45502 118894
rect 45586 118658 45822 118894
rect 45266 118338 45502 118574
rect 45586 118338 45822 118574
rect 45266 82658 45502 82894
rect 45586 82658 45822 82894
rect 45266 82338 45502 82574
rect 45586 82338 45822 82574
rect 45266 46658 45502 46894
rect 45586 46658 45822 46894
rect 45266 46338 45502 46574
rect 45586 46338 45822 46574
rect 45266 10658 45502 10894
rect 45586 10658 45822 10894
rect 45266 10338 45502 10574
rect 45586 10338 45822 10574
rect 45266 -4422 45502 -4186
rect 45586 -4422 45822 -4186
rect 45266 -4742 45502 -4506
rect 45586 -4742 45822 -4506
rect 66986 711322 67222 711558
rect 67306 711322 67542 711558
rect 66986 711002 67222 711238
rect 67306 711002 67542 711238
rect 63266 709402 63502 709638
rect 63586 709402 63822 709638
rect 63266 709082 63502 709318
rect 63586 709082 63822 709318
rect 59546 707482 59782 707718
rect 59866 707482 60102 707718
rect 59546 707162 59782 707398
rect 59866 707162 60102 707398
rect 48986 698378 49222 698614
rect 49306 698378 49542 698614
rect 48986 698058 49222 698294
rect 49306 698058 49542 698294
rect 48986 662378 49222 662614
rect 49306 662378 49542 662614
rect 48986 662058 49222 662294
rect 49306 662058 49542 662294
rect 48986 626378 49222 626614
rect 49306 626378 49542 626614
rect 48986 626058 49222 626294
rect 49306 626058 49542 626294
rect 48986 590378 49222 590614
rect 49306 590378 49542 590614
rect 48986 590058 49222 590294
rect 49306 590058 49542 590294
rect 48986 554378 49222 554614
rect 49306 554378 49542 554614
rect 48986 554058 49222 554294
rect 49306 554058 49542 554294
rect 48986 518378 49222 518614
rect 49306 518378 49542 518614
rect 48986 518058 49222 518294
rect 49306 518058 49542 518294
rect 48986 482378 49222 482614
rect 49306 482378 49542 482614
rect 48986 482058 49222 482294
rect 49306 482058 49542 482294
rect 48986 446378 49222 446614
rect 49306 446378 49542 446614
rect 48986 446058 49222 446294
rect 49306 446058 49542 446294
rect 48986 410378 49222 410614
rect 49306 410378 49542 410614
rect 48986 410058 49222 410294
rect 49306 410058 49542 410294
rect 48986 374378 49222 374614
rect 49306 374378 49542 374614
rect 48986 374058 49222 374294
rect 49306 374058 49542 374294
rect 48986 338378 49222 338614
rect 49306 338378 49542 338614
rect 48986 338058 49222 338294
rect 49306 338058 49542 338294
rect 48986 302378 49222 302614
rect 49306 302378 49542 302614
rect 48986 302058 49222 302294
rect 49306 302058 49542 302294
rect 48986 266378 49222 266614
rect 49306 266378 49542 266614
rect 48986 266058 49222 266294
rect 49306 266058 49542 266294
rect 48986 230378 49222 230614
rect 49306 230378 49542 230614
rect 48986 230058 49222 230294
rect 49306 230058 49542 230294
rect 48986 194378 49222 194614
rect 49306 194378 49542 194614
rect 48986 194058 49222 194294
rect 49306 194058 49542 194294
rect 48986 158378 49222 158614
rect 49306 158378 49542 158614
rect 48986 158058 49222 158294
rect 49306 158058 49542 158294
rect 48986 122378 49222 122614
rect 49306 122378 49542 122614
rect 48986 122058 49222 122294
rect 49306 122058 49542 122294
rect 48986 86378 49222 86614
rect 49306 86378 49542 86614
rect 48986 86058 49222 86294
rect 49306 86058 49542 86294
rect 48986 50378 49222 50614
rect 49306 50378 49542 50614
rect 48986 50058 49222 50294
rect 49306 50058 49542 50294
rect 48986 14378 49222 14614
rect 49306 14378 49542 14614
rect 48986 14058 49222 14294
rect 49306 14058 49542 14294
rect 30986 -7302 31222 -7066
rect 31306 -7302 31542 -7066
rect 30986 -7622 31222 -7386
rect 31306 -7622 31542 -7386
rect 55826 705562 56062 705798
rect 56146 705562 56382 705798
rect 55826 705242 56062 705478
rect 56146 705242 56382 705478
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -1542 56062 -1306
rect 56146 -1542 56382 -1306
rect 55826 -1862 56062 -1626
rect 56146 -1862 56382 -1626
rect 59546 672938 59782 673174
rect 59866 672938 60102 673174
rect 59546 672618 59782 672854
rect 59866 672618 60102 672854
rect 59546 636938 59782 637174
rect 59866 636938 60102 637174
rect 59546 636618 59782 636854
rect 59866 636618 60102 636854
rect 59546 600938 59782 601174
rect 59866 600938 60102 601174
rect 59546 600618 59782 600854
rect 59866 600618 60102 600854
rect 59546 564938 59782 565174
rect 59866 564938 60102 565174
rect 59546 564618 59782 564854
rect 59866 564618 60102 564854
rect 59546 528938 59782 529174
rect 59866 528938 60102 529174
rect 59546 528618 59782 528854
rect 59866 528618 60102 528854
rect 59546 492938 59782 493174
rect 59866 492938 60102 493174
rect 59546 492618 59782 492854
rect 59866 492618 60102 492854
rect 59546 456938 59782 457174
rect 59866 456938 60102 457174
rect 59546 456618 59782 456854
rect 59866 456618 60102 456854
rect 59546 420938 59782 421174
rect 59866 420938 60102 421174
rect 59546 420618 59782 420854
rect 59866 420618 60102 420854
rect 59546 384938 59782 385174
rect 59866 384938 60102 385174
rect 59546 384618 59782 384854
rect 59866 384618 60102 384854
rect 59546 348938 59782 349174
rect 59866 348938 60102 349174
rect 59546 348618 59782 348854
rect 59866 348618 60102 348854
rect 59546 312938 59782 313174
rect 59866 312938 60102 313174
rect 59546 312618 59782 312854
rect 59866 312618 60102 312854
rect 59546 276938 59782 277174
rect 59866 276938 60102 277174
rect 59546 276618 59782 276854
rect 59866 276618 60102 276854
rect 59546 240938 59782 241174
rect 59866 240938 60102 241174
rect 59546 240618 59782 240854
rect 59866 240618 60102 240854
rect 59546 204938 59782 205174
rect 59866 204938 60102 205174
rect 59546 204618 59782 204854
rect 59866 204618 60102 204854
rect 59546 168938 59782 169174
rect 59866 168938 60102 169174
rect 59546 168618 59782 168854
rect 59866 168618 60102 168854
rect 59546 132938 59782 133174
rect 59866 132938 60102 133174
rect 59546 132618 59782 132854
rect 59866 132618 60102 132854
rect 59546 96938 59782 97174
rect 59866 96938 60102 97174
rect 59546 96618 59782 96854
rect 59866 96618 60102 96854
rect 59546 60938 59782 61174
rect 59866 60938 60102 61174
rect 59546 60618 59782 60854
rect 59866 60618 60102 60854
rect 59546 24938 59782 25174
rect 59866 24938 60102 25174
rect 59546 24618 59782 24854
rect 59866 24618 60102 24854
rect 59546 -3462 59782 -3226
rect 59866 -3462 60102 -3226
rect 59546 -3782 59782 -3546
rect 59866 -3782 60102 -3546
rect 63266 676658 63502 676894
rect 63586 676658 63822 676894
rect 63266 676338 63502 676574
rect 63586 676338 63822 676574
rect 63266 640658 63502 640894
rect 63586 640658 63822 640894
rect 63266 640338 63502 640574
rect 63586 640338 63822 640574
rect 63266 604658 63502 604894
rect 63586 604658 63822 604894
rect 63266 604338 63502 604574
rect 63586 604338 63822 604574
rect 63266 568658 63502 568894
rect 63586 568658 63822 568894
rect 63266 568338 63502 568574
rect 63586 568338 63822 568574
rect 63266 532658 63502 532894
rect 63586 532658 63822 532894
rect 63266 532338 63502 532574
rect 63586 532338 63822 532574
rect 63266 496658 63502 496894
rect 63586 496658 63822 496894
rect 63266 496338 63502 496574
rect 63586 496338 63822 496574
rect 63266 460658 63502 460894
rect 63586 460658 63822 460894
rect 63266 460338 63502 460574
rect 63586 460338 63822 460574
rect 63266 424658 63502 424894
rect 63586 424658 63822 424894
rect 63266 424338 63502 424574
rect 63586 424338 63822 424574
rect 63266 388658 63502 388894
rect 63586 388658 63822 388894
rect 63266 388338 63502 388574
rect 63586 388338 63822 388574
rect 63266 352658 63502 352894
rect 63586 352658 63822 352894
rect 63266 352338 63502 352574
rect 63586 352338 63822 352574
rect 63266 316658 63502 316894
rect 63586 316658 63822 316894
rect 63266 316338 63502 316574
rect 63586 316338 63822 316574
rect 63266 280658 63502 280894
rect 63586 280658 63822 280894
rect 63266 280338 63502 280574
rect 63586 280338 63822 280574
rect 63266 244658 63502 244894
rect 63586 244658 63822 244894
rect 63266 244338 63502 244574
rect 63586 244338 63822 244574
rect 63266 208658 63502 208894
rect 63586 208658 63822 208894
rect 63266 208338 63502 208574
rect 63586 208338 63822 208574
rect 63266 172658 63502 172894
rect 63586 172658 63822 172894
rect 63266 172338 63502 172574
rect 63586 172338 63822 172574
rect 63266 136658 63502 136894
rect 63586 136658 63822 136894
rect 63266 136338 63502 136574
rect 63586 136338 63822 136574
rect 63266 100658 63502 100894
rect 63586 100658 63822 100894
rect 63266 100338 63502 100574
rect 63586 100338 63822 100574
rect 63266 64658 63502 64894
rect 63586 64658 63822 64894
rect 63266 64338 63502 64574
rect 63586 64338 63822 64574
rect 63266 28658 63502 28894
rect 63586 28658 63822 28894
rect 63266 28338 63502 28574
rect 63586 28338 63822 28574
rect 63266 -5382 63502 -5146
rect 63586 -5382 63822 -5146
rect 63266 -5702 63502 -5466
rect 63586 -5702 63822 -5466
rect 84986 710362 85222 710598
rect 85306 710362 85542 710598
rect 84986 710042 85222 710278
rect 85306 710042 85542 710278
rect 81266 708442 81502 708678
rect 81586 708442 81822 708678
rect 81266 708122 81502 708358
rect 81586 708122 81822 708358
rect 77546 706522 77782 706758
rect 77866 706522 78102 706758
rect 77546 706202 77782 706438
rect 77866 706202 78102 706438
rect 66986 680378 67222 680614
rect 67306 680378 67542 680614
rect 66986 680058 67222 680294
rect 67306 680058 67542 680294
rect 66986 644378 67222 644614
rect 67306 644378 67542 644614
rect 66986 644058 67222 644294
rect 67306 644058 67542 644294
rect 66986 608378 67222 608614
rect 67306 608378 67542 608614
rect 66986 608058 67222 608294
rect 67306 608058 67542 608294
rect 66986 572378 67222 572614
rect 67306 572378 67542 572614
rect 66986 572058 67222 572294
rect 67306 572058 67542 572294
rect 66986 536378 67222 536614
rect 67306 536378 67542 536614
rect 66986 536058 67222 536294
rect 67306 536058 67542 536294
rect 66986 500378 67222 500614
rect 67306 500378 67542 500614
rect 66986 500058 67222 500294
rect 67306 500058 67542 500294
rect 66986 464378 67222 464614
rect 67306 464378 67542 464614
rect 66986 464058 67222 464294
rect 67306 464058 67542 464294
rect 66986 428378 67222 428614
rect 67306 428378 67542 428614
rect 66986 428058 67222 428294
rect 67306 428058 67542 428294
rect 66986 392378 67222 392614
rect 67306 392378 67542 392614
rect 66986 392058 67222 392294
rect 67306 392058 67542 392294
rect 66986 356378 67222 356614
rect 67306 356378 67542 356614
rect 66986 356058 67222 356294
rect 67306 356058 67542 356294
rect 66986 320378 67222 320614
rect 67306 320378 67542 320614
rect 66986 320058 67222 320294
rect 67306 320058 67542 320294
rect 66986 284378 67222 284614
rect 67306 284378 67542 284614
rect 66986 284058 67222 284294
rect 67306 284058 67542 284294
rect 66986 248378 67222 248614
rect 67306 248378 67542 248614
rect 66986 248058 67222 248294
rect 67306 248058 67542 248294
rect 66986 212378 67222 212614
rect 67306 212378 67542 212614
rect 66986 212058 67222 212294
rect 67306 212058 67542 212294
rect 66986 176378 67222 176614
rect 67306 176378 67542 176614
rect 66986 176058 67222 176294
rect 67306 176058 67542 176294
rect 66986 140378 67222 140614
rect 67306 140378 67542 140614
rect 66986 140058 67222 140294
rect 67306 140058 67542 140294
rect 66986 104378 67222 104614
rect 67306 104378 67542 104614
rect 66986 104058 67222 104294
rect 67306 104058 67542 104294
rect 66986 68378 67222 68614
rect 67306 68378 67542 68614
rect 66986 68058 67222 68294
rect 67306 68058 67542 68294
rect 66986 32378 67222 32614
rect 67306 32378 67542 32614
rect 66986 32058 67222 32294
rect 67306 32058 67542 32294
rect 48986 -6342 49222 -6106
rect 49306 -6342 49542 -6106
rect 48986 -6662 49222 -6426
rect 49306 -6662 49542 -6426
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 73826 579218 74062 579454
rect 74146 579218 74382 579454
rect 73826 578898 74062 579134
rect 74146 578898 74382 579134
rect 73826 543218 74062 543454
rect 74146 543218 74382 543454
rect 73826 542898 74062 543134
rect 74146 542898 74382 543134
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 73826 435218 74062 435454
rect 74146 435218 74382 435454
rect 73826 434898 74062 435134
rect 74146 434898 74382 435134
rect 73826 399218 74062 399454
rect 74146 399218 74382 399454
rect 73826 398898 74062 399134
rect 74146 398898 74382 399134
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 73826 327218 74062 327454
rect 74146 327218 74382 327454
rect 73826 326898 74062 327134
rect 74146 326898 74382 327134
rect 73826 291218 74062 291454
rect 74146 291218 74382 291454
rect 73826 290898 74062 291134
rect 74146 290898 74382 291134
rect 73826 255218 74062 255454
rect 74146 255218 74382 255454
rect 73826 254898 74062 255134
rect 74146 254898 74382 255134
rect 73826 219218 74062 219454
rect 74146 219218 74382 219454
rect 73826 218898 74062 219134
rect 74146 218898 74382 219134
rect 73826 183218 74062 183454
rect 74146 183218 74382 183454
rect 73826 182898 74062 183134
rect 74146 182898 74382 183134
rect 73826 147218 74062 147454
rect 74146 147218 74382 147454
rect 73826 146898 74062 147134
rect 74146 146898 74382 147134
rect 73826 111218 74062 111454
rect 74146 111218 74382 111454
rect 73826 110898 74062 111134
rect 74146 110898 74382 111134
rect 73826 75218 74062 75454
rect 74146 75218 74382 75454
rect 73826 74898 74062 75134
rect 74146 74898 74382 75134
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 77546 654938 77782 655174
rect 77866 654938 78102 655174
rect 77546 654618 77782 654854
rect 77866 654618 78102 654854
rect 77546 618938 77782 619174
rect 77866 618938 78102 619174
rect 77546 618618 77782 618854
rect 77866 618618 78102 618854
rect 77546 582938 77782 583174
rect 77866 582938 78102 583174
rect 77546 582618 77782 582854
rect 77866 582618 78102 582854
rect 77546 546938 77782 547174
rect 77866 546938 78102 547174
rect 77546 546618 77782 546854
rect 77866 546618 78102 546854
rect 77546 510938 77782 511174
rect 77866 510938 78102 511174
rect 77546 510618 77782 510854
rect 77866 510618 78102 510854
rect 77546 474938 77782 475174
rect 77866 474938 78102 475174
rect 77546 474618 77782 474854
rect 77866 474618 78102 474854
rect 77546 438938 77782 439174
rect 77866 438938 78102 439174
rect 77546 438618 77782 438854
rect 77866 438618 78102 438854
rect 77546 402938 77782 403174
rect 77866 402938 78102 403174
rect 77546 402618 77782 402854
rect 77866 402618 78102 402854
rect 77546 366938 77782 367174
rect 77866 366938 78102 367174
rect 77546 366618 77782 366854
rect 77866 366618 78102 366854
rect 77546 330938 77782 331174
rect 77866 330938 78102 331174
rect 77546 330618 77782 330854
rect 77866 330618 78102 330854
rect 77546 294938 77782 295174
rect 77866 294938 78102 295174
rect 77546 294618 77782 294854
rect 77866 294618 78102 294854
rect 77546 258938 77782 259174
rect 77866 258938 78102 259174
rect 77546 258618 77782 258854
rect 77866 258618 78102 258854
rect 77546 222938 77782 223174
rect 77866 222938 78102 223174
rect 77546 222618 77782 222854
rect 77866 222618 78102 222854
rect 77546 186938 77782 187174
rect 77866 186938 78102 187174
rect 77546 186618 77782 186854
rect 77866 186618 78102 186854
rect 77546 150938 77782 151174
rect 77866 150938 78102 151174
rect 77546 150618 77782 150854
rect 77866 150618 78102 150854
rect 77546 114938 77782 115174
rect 77866 114938 78102 115174
rect 77546 114618 77782 114854
rect 77866 114618 78102 114854
rect 77546 78938 77782 79174
rect 77866 78938 78102 79174
rect 77546 78618 77782 78854
rect 77866 78618 78102 78854
rect 77546 42938 77782 43174
rect 77866 42938 78102 43174
rect 77546 42618 77782 42854
rect 77866 42618 78102 42854
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 77546 -2502 77782 -2266
rect 77866 -2502 78102 -2266
rect 77546 -2822 77782 -2586
rect 77866 -2822 78102 -2586
rect 81266 694658 81502 694894
rect 81586 694658 81822 694894
rect 81266 694338 81502 694574
rect 81586 694338 81822 694574
rect 81266 658658 81502 658894
rect 81586 658658 81822 658894
rect 81266 658338 81502 658574
rect 81586 658338 81822 658574
rect 81266 622658 81502 622894
rect 81586 622658 81822 622894
rect 81266 622338 81502 622574
rect 81586 622338 81822 622574
rect 81266 586658 81502 586894
rect 81586 586658 81822 586894
rect 81266 586338 81502 586574
rect 81586 586338 81822 586574
rect 81266 550658 81502 550894
rect 81586 550658 81822 550894
rect 81266 550338 81502 550574
rect 81586 550338 81822 550574
rect 81266 514658 81502 514894
rect 81586 514658 81822 514894
rect 81266 514338 81502 514574
rect 81586 514338 81822 514574
rect 81266 478658 81502 478894
rect 81586 478658 81822 478894
rect 81266 478338 81502 478574
rect 81586 478338 81822 478574
rect 81266 442658 81502 442894
rect 81586 442658 81822 442894
rect 81266 442338 81502 442574
rect 81586 442338 81822 442574
rect 81266 406658 81502 406894
rect 81586 406658 81822 406894
rect 81266 406338 81502 406574
rect 81586 406338 81822 406574
rect 81266 370658 81502 370894
rect 81586 370658 81822 370894
rect 81266 370338 81502 370574
rect 81586 370338 81822 370574
rect 81266 334658 81502 334894
rect 81586 334658 81822 334894
rect 81266 334338 81502 334574
rect 81586 334338 81822 334574
rect 81266 298658 81502 298894
rect 81586 298658 81822 298894
rect 81266 298338 81502 298574
rect 81586 298338 81822 298574
rect 81266 262658 81502 262894
rect 81586 262658 81822 262894
rect 81266 262338 81502 262574
rect 81586 262338 81822 262574
rect 81266 226658 81502 226894
rect 81586 226658 81822 226894
rect 81266 226338 81502 226574
rect 81586 226338 81822 226574
rect 81266 190658 81502 190894
rect 81586 190658 81822 190894
rect 81266 190338 81502 190574
rect 81586 190338 81822 190574
rect 81266 154658 81502 154894
rect 81586 154658 81822 154894
rect 81266 154338 81502 154574
rect 81586 154338 81822 154574
rect 81266 118658 81502 118894
rect 81586 118658 81822 118894
rect 81266 118338 81502 118574
rect 81586 118338 81822 118574
rect 81266 82658 81502 82894
rect 81586 82658 81822 82894
rect 81266 82338 81502 82574
rect 81586 82338 81822 82574
rect 81266 46658 81502 46894
rect 81586 46658 81822 46894
rect 81266 46338 81502 46574
rect 81586 46338 81822 46574
rect 81266 10658 81502 10894
rect 81586 10658 81822 10894
rect 81266 10338 81502 10574
rect 81586 10338 81822 10574
rect 81266 -4422 81502 -4186
rect 81586 -4422 81822 -4186
rect 81266 -4742 81502 -4506
rect 81586 -4742 81822 -4506
rect 102986 711322 103222 711558
rect 103306 711322 103542 711558
rect 102986 711002 103222 711238
rect 103306 711002 103542 711238
rect 99266 709402 99502 709638
rect 99586 709402 99822 709638
rect 99266 709082 99502 709318
rect 99586 709082 99822 709318
rect 95546 707482 95782 707718
rect 95866 707482 96102 707718
rect 95546 707162 95782 707398
rect 95866 707162 96102 707398
rect 84986 698378 85222 698614
rect 85306 698378 85542 698614
rect 84986 698058 85222 698294
rect 85306 698058 85542 698294
rect 84986 662378 85222 662614
rect 85306 662378 85542 662614
rect 84986 662058 85222 662294
rect 85306 662058 85542 662294
rect 84986 626378 85222 626614
rect 85306 626378 85542 626614
rect 84986 626058 85222 626294
rect 85306 626058 85542 626294
rect 84986 590378 85222 590614
rect 85306 590378 85542 590614
rect 84986 590058 85222 590294
rect 85306 590058 85542 590294
rect 84986 554378 85222 554614
rect 85306 554378 85542 554614
rect 84986 554058 85222 554294
rect 85306 554058 85542 554294
rect 84986 518378 85222 518614
rect 85306 518378 85542 518614
rect 84986 518058 85222 518294
rect 85306 518058 85542 518294
rect 84986 482378 85222 482614
rect 85306 482378 85542 482614
rect 84986 482058 85222 482294
rect 85306 482058 85542 482294
rect 84986 446378 85222 446614
rect 85306 446378 85542 446614
rect 84986 446058 85222 446294
rect 85306 446058 85542 446294
rect 84986 410378 85222 410614
rect 85306 410378 85542 410614
rect 84986 410058 85222 410294
rect 85306 410058 85542 410294
rect 84986 374378 85222 374614
rect 85306 374378 85542 374614
rect 84986 374058 85222 374294
rect 85306 374058 85542 374294
rect 84986 338378 85222 338614
rect 85306 338378 85542 338614
rect 84986 338058 85222 338294
rect 85306 338058 85542 338294
rect 84986 302378 85222 302614
rect 85306 302378 85542 302614
rect 84986 302058 85222 302294
rect 85306 302058 85542 302294
rect 84986 266378 85222 266614
rect 85306 266378 85542 266614
rect 84986 266058 85222 266294
rect 85306 266058 85542 266294
rect 84986 230378 85222 230614
rect 85306 230378 85542 230614
rect 84986 230058 85222 230294
rect 85306 230058 85542 230294
rect 84986 194378 85222 194614
rect 85306 194378 85542 194614
rect 84986 194058 85222 194294
rect 85306 194058 85542 194294
rect 84986 158378 85222 158614
rect 85306 158378 85542 158614
rect 84986 158058 85222 158294
rect 85306 158058 85542 158294
rect 84986 122378 85222 122614
rect 85306 122378 85542 122614
rect 84986 122058 85222 122294
rect 85306 122058 85542 122294
rect 84986 86378 85222 86614
rect 85306 86378 85542 86614
rect 84986 86058 85222 86294
rect 85306 86058 85542 86294
rect 84986 50378 85222 50614
rect 85306 50378 85542 50614
rect 84986 50058 85222 50294
rect 85306 50058 85542 50294
rect 84986 14378 85222 14614
rect 85306 14378 85542 14614
rect 84986 14058 85222 14294
rect 85306 14058 85542 14294
rect 66986 -7302 67222 -7066
rect 67306 -7302 67542 -7066
rect 66986 -7622 67222 -7386
rect 67306 -7622 67542 -7386
rect 91826 705562 92062 705798
rect 92146 705562 92382 705798
rect 91826 705242 92062 705478
rect 92146 705242 92382 705478
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 91826 561218 92062 561454
rect 92146 561218 92382 561454
rect 91826 560898 92062 561134
rect 92146 560898 92382 561134
rect 91826 525218 92062 525454
rect 92146 525218 92382 525454
rect 91826 524898 92062 525134
rect 92146 524898 92382 525134
rect 91826 489218 92062 489454
rect 92146 489218 92382 489454
rect 91826 488898 92062 489134
rect 92146 488898 92382 489134
rect 91826 453218 92062 453454
rect 92146 453218 92382 453454
rect 91826 452898 92062 453134
rect 92146 452898 92382 453134
rect 91826 417218 92062 417454
rect 92146 417218 92382 417454
rect 91826 416898 92062 417134
rect 92146 416898 92382 417134
rect 91826 381218 92062 381454
rect 92146 381218 92382 381454
rect 91826 380898 92062 381134
rect 92146 380898 92382 381134
rect 91826 345218 92062 345454
rect 92146 345218 92382 345454
rect 91826 344898 92062 345134
rect 92146 344898 92382 345134
rect 91826 309218 92062 309454
rect 92146 309218 92382 309454
rect 91826 308898 92062 309134
rect 92146 308898 92382 309134
rect 91826 273218 92062 273454
rect 92146 273218 92382 273454
rect 91826 272898 92062 273134
rect 92146 272898 92382 273134
rect 91826 237218 92062 237454
rect 92146 237218 92382 237454
rect 91826 236898 92062 237134
rect 92146 236898 92382 237134
rect 91826 201218 92062 201454
rect 92146 201218 92382 201454
rect 91826 200898 92062 201134
rect 92146 200898 92382 201134
rect 91826 165218 92062 165454
rect 92146 165218 92382 165454
rect 91826 164898 92062 165134
rect 92146 164898 92382 165134
rect 91826 129218 92062 129454
rect 92146 129218 92382 129454
rect 91826 128898 92062 129134
rect 92146 128898 92382 129134
rect 91826 93218 92062 93454
rect 92146 93218 92382 93454
rect 91826 92898 92062 93134
rect 92146 92898 92382 93134
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -1542 92062 -1306
rect 92146 -1542 92382 -1306
rect 91826 -1862 92062 -1626
rect 92146 -1862 92382 -1626
rect 95546 672938 95782 673174
rect 95866 672938 96102 673174
rect 95546 672618 95782 672854
rect 95866 672618 96102 672854
rect 95546 636938 95782 637174
rect 95866 636938 96102 637174
rect 95546 636618 95782 636854
rect 95866 636618 96102 636854
rect 95546 600938 95782 601174
rect 95866 600938 96102 601174
rect 95546 600618 95782 600854
rect 95866 600618 96102 600854
rect 95546 564938 95782 565174
rect 95866 564938 96102 565174
rect 95546 564618 95782 564854
rect 95866 564618 96102 564854
rect 95546 528938 95782 529174
rect 95866 528938 96102 529174
rect 95546 528618 95782 528854
rect 95866 528618 96102 528854
rect 95546 492938 95782 493174
rect 95866 492938 96102 493174
rect 95546 492618 95782 492854
rect 95866 492618 96102 492854
rect 95546 456938 95782 457174
rect 95866 456938 96102 457174
rect 95546 456618 95782 456854
rect 95866 456618 96102 456854
rect 95546 420938 95782 421174
rect 95866 420938 96102 421174
rect 95546 420618 95782 420854
rect 95866 420618 96102 420854
rect 95546 384938 95782 385174
rect 95866 384938 96102 385174
rect 95546 384618 95782 384854
rect 95866 384618 96102 384854
rect 95546 348938 95782 349174
rect 95866 348938 96102 349174
rect 95546 348618 95782 348854
rect 95866 348618 96102 348854
rect 95546 312938 95782 313174
rect 95866 312938 96102 313174
rect 95546 312618 95782 312854
rect 95866 312618 96102 312854
rect 95546 276938 95782 277174
rect 95866 276938 96102 277174
rect 95546 276618 95782 276854
rect 95866 276618 96102 276854
rect 95546 240938 95782 241174
rect 95866 240938 96102 241174
rect 95546 240618 95782 240854
rect 95866 240618 96102 240854
rect 95546 204938 95782 205174
rect 95866 204938 96102 205174
rect 95546 204618 95782 204854
rect 95866 204618 96102 204854
rect 95546 168938 95782 169174
rect 95866 168938 96102 169174
rect 95546 168618 95782 168854
rect 95866 168618 96102 168854
rect 95546 132938 95782 133174
rect 95866 132938 96102 133174
rect 95546 132618 95782 132854
rect 95866 132618 96102 132854
rect 95546 96938 95782 97174
rect 95866 96938 96102 97174
rect 95546 96618 95782 96854
rect 95866 96618 96102 96854
rect 95546 60938 95782 61174
rect 95866 60938 96102 61174
rect 95546 60618 95782 60854
rect 95866 60618 96102 60854
rect 95546 24938 95782 25174
rect 95866 24938 96102 25174
rect 95546 24618 95782 24854
rect 95866 24618 96102 24854
rect 95546 -3462 95782 -3226
rect 95866 -3462 96102 -3226
rect 95546 -3782 95782 -3546
rect 95866 -3782 96102 -3546
rect 99266 676658 99502 676894
rect 99586 676658 99822 676894
rect 99266 676338 99502 676574
rect 99586 676338 99822 676574
rect 99266 640658 99502 640894
rect 99586 640658 99822 640894
rect 99266 640338 99502 640574
rect 99586 640338 99822 640574
rect 99266 604658 99502 604894
rect 99586 604658 99822 604894
rect 99266 604338 99502 604574
rect 99586 604338 99822 604574
rect 99266 568658 99502 568894
rect 99586 568658 99822 568894
rect 99266 568338 99502 568574
rect 99586 568338 99822 568574
rect 99266 532658 99502 532894
rect 99586 532658 99822 532894
rect 99266 532338 99502 532574
rect 99586 532338 99822 532574
rect 99266 496658 99502 496894
rect 99586 496658 99822 496894
rect 99266 496338 99502 496574
rect 99586 496338 99822 496574
rect 99266 460658 99502 460894
rect 99586 460658 99822 460894
rect 99266 460338 99502 460574
rect 99586 460338 99822 460574
rect 99266 424658 99502 424894
rect 99586 424658 99822 424894
rect 99266 424338 99502 424574
rect 99586 424338 99822 424574
rect 99266 388658 99502 388894
rect 99586 388658 99822 388894
rect 99266 388338 99502 388574
rect 99586 388338 99822 388574
rect 99266 352658 99502 352894
rect 99586 352658 99822 352894
rect 99266 352338 99502 352574
rect 99586 352338 99822 352574
rect 99266 316658 99502 316894
rect 99586 316658 99822 316894
rect 99266 316338 99502 316574
rect 99586 316338 99822 316574
rect 99266 280658 99502 280894
rect 99586 280658 99822 280894
rect 99266 280338 99502 280574
rect 99586 280338 99822 280574
rect 99266 244658 99502 244894
rect 99586 244658 99822 244894
rect 99266 244338 99502 244574
rect 99586 244338 99822 244574
rect 99266 208658 99502 208894
rect 99586 208658 99822 208894
rect 99266 208338 99502 208574
rect 99586 208338 99822 208574
rect 99266 172658 99502 172894
rect 99586 172658 99822 172894
rect 99266 172338 99502 172574
rect 99586 172338 99822 172574
rect 99266 136658 99502 136894
rect 99586 136658 99822 136894
rect 99266 136338 99502 136574
rect 99586 136338 99822 136574
rect 99266 100658 99502 100894
rect 99586 100658 99822 100894
rect 99266 100338 99502 100574
rect 99586 100338 99822 100574
rect 99266 64658 99502 64894
rect 99586 64658 99822 64894
rect 99266 64338 99502 64574
rect 99586 64338 99822 64574
rect 99266 28658 99502 28894
rect 99586 28658 99822 28894
rect 99266 28338 99502 28574
rect 99586 28338 99822 28574
rect 99266 -5382 99502 -5146
rect 99586 -5382 99822 -5146
rect 99266 -5702 99502 -5466
rect 99586 -5702 99822 -5466
rect 120986 710362 121222 710598
rect 121306 710362 121542 710598
rect 120986 710042 121222 710278
rect 121306 710042 121542 710278
rect 117266 708442 117502 708678
rect 117586 708442 117822 708678
rect 117266 708122 117502 708358
rect 117586 708122 117822 708358
rect 113546 706522 113782 706758
rect 113866 706522 114102 706758
rect 113546 706202 113782 706438
rect 113866 706202 114102 706438
rect 102986 680378 103222 680614
rect 103306 680378 103542 680614
rect 102986 680058 103222 680294
rect 103306 680058 103542 680294
rect 102986 644378 103222 644614
rect 103306 644378 103542 644614
rect 102986 644058 103222 644294
rect 103306 644058 103542 644294
rect 102986 608378 103222 608614
rect 103306 608378 103542 608614
rect 102986 608058 103222 608294
rect 103306 608058 103542 608294
rect 102986 572378 103222 572614
rect 103306 572378 103542 572614
rect 102986 572058 103222 572294
rect 103306 572058 103542 572294
rect 102986 536378 103222 536614
rect 103306 536378 103542 536614
rect 102986 536058 103222 536294
rect 103306 536058 103542 536294
rect 102986 500378 103222 500614
rect 103306 500378 103542 500614
rect 102986 500058 103222 500294
rect 103306 500058 103542 500294
rect 102986 464378 103222 464614
rect 103306 464378 103542 464614
rect 102986 464058 103222 464294
rect 103306 464058 103542 464294
rect 102986 428378 103222 428614
rect 103306 428378 103542 428614
rect 102986 428058 103222 428294
rect 103306 428058 103542 428294
rect 102986 392378 103222 392614
rect 103306 392378 103542 392614
rect 102986 392058 103222 392294
rect 103306 392058 103542 392294
rect 102986 356378 103222 356614
rect 103306 356378 103542 356614
rect 102986 356058 103222 356294
rect 103306 356058 103542 356294
rect 102986 320378 103222 320614
rect 103306 320378 103542 320614
rect 102986 320058 103222 320294
rect 103306 320058 103542 320294
rect 102986 284378 103222 284614
rect 103306 284378 103542 284614
rect 102986 284058 103222 284294
rect 103306 284058 103542 284294
rect 102986 248378 103222 248614
rect 103306 248378 103542 248614
rect 102986 248058 103222 248294
rect 103306 248058 103542 248294
rect 102986 212378 103222 212614
rect 103306 212378 103542 212614
rect 102986 212058 103222 212294
rect 103306 212058 103542 212294
rect 102986 176378 103222 176614
rect 103306 176378 103542 176614
rect 102986 176058 103222 176294
rect 103306 176058 103542 176294
rect 102986 140378 103222 140614
rect 103306 140378 103542 140614
rect 102986 140058 103222 140294
rect 103306 140058 103542 140294
rect 102986 104378 103222 104614
rect 103306 104378 103542 104614
rect 102986 104058 103222 104294
rect 103306 104058 103542 104294
rect 102986 68378 103222 68614
rect 103306 68378 103542 68614
rect 102986 68058 103222 68294
rect 103306 68058 103542 68294
rect 102986 32378 103222 32614
rect 103306 32378 103542 32614
rect 102986 32058 103222 32294
rect 103306 32058 103542 32294
rect 84986 -6342 85222 -6106
rect 85306 -6342 85542 -6106
rect 84986 -6662 85222 -6426
rect 85306 -6662 85542 -6426
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 109826 507218 110062 507454
rect 110146 507218 110382 507454
rect 109826 506898 110062 507134
rect 110146 506898 110382 507134
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 109826 435218 110062 435454
rect 110146 435218 110382 435454
rect 109826 434898 110062 435134
rect 110146 434898 110382 435134
rect 109826 399218 110062 399454
rect 110146 399218 110382 399454
rect 109826 398898 110062 399134
rect 110146 398898 110382 399134
rect 109826 363218 110062 363454
rect 110146 363218 110382 363454
rect 109826 362898 110062 363134
rect 110146 362898 110382 363134
rect 109826 327218 110062 327454
rect 110146 327218 110382 327454
rect 109826 326898 110062 327134
rect 110146 326898 110382 327134
rect 109826 291218 110062 291454
rect 110146 291218 110382 291454
rect 109826 290898 110062 291134
rect 110146 290898 110382 291134
rect 109826 255218 110062 255454
rect 110146 255218 110382 255454
rect 109826 254898 110062 255134
rect 110146 254898 110382 255134
rect 109826 219218 110062 219454
rect 110146 219218 110382 219454
rect 109826 218898 110062 219134
rect 110146 218898 110382 219134
rect 109826 183218 110062 183454
rect 110146 183218 110382 183454
rect 109826 182898 110062 183134
rect 110146 182898 110382 183134
rect 109826 147218 110062 147454
rect 110146 147218 110382 147454
rect 109826 146898 110062 147134
rect 110146 146898 110382 147134
rect 109826 111218 110062 111454
rect 110146 111218 110382 111454
rect 109826 110898 110062 111134
rect 110146 110898 110382 111134
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 690938 113782 691174
rect 113866 690938 114102 691174
rect 113546 690618 113782 690854
rect 113866 690618 114102 690854
rect 113546 654938 113782 655174
rect 113866 654938 114102 655174
rect 113546 654618 113782 654854
rect 113866 654618 114102 654854
rect 113546 618938 113782 619174
rect 113866 618938 114102 619174
rect 113546 618618 113782 618854
rect 113866 618618 114102 618854
rect 113546 582938 113782 583174
rect 113866 582938 114102 583174
rect 113546 582618 113782 582854
rect 113866 582618 114102 582854
rect 113546 546938 113782 547174
rect 113866 546938 114102 547174
rect 113546 546618 113782 546854
rect 113866 546618 114102 546854
rect 113546 510938 113782 511174
rect 113866 510938 114102 511174
rect 113546 510618 113782 510854
rect 113866 510618 114102 510854
rect 113546 474938 113782 475174
rect 113866 474938 114102 475174
rect 113546 474618 113782 474854
rect 113866 474618 114102 474854
rect 113546 438938 113782 439174
rect 113866 438938 114102 439174
rect 113546 438618 113782 438854
rect 113866 438618 114102 438854
rect 113546 402938 113782 403174
rect 113866 402938 114102 403174
rect 113546 402618 113782 402854
rect 113866 402618 114102 402854
rect 113546 366938 113782 367174
rect 113866 366938 114102 367174
rect 113546 366618 113782 366854
rect 113866 366618 114102 366854
rect 113546 330938 113782 331174
rect 113866 330938 114102 331174
rect 113546 330618 113782 330854
rect 113866 330618 114102 330854
rect 113546 294938 113782 295174
rect 113866 294938 114102 295174
rect 113546 294618 113782 294854
rect 113866 294618 114102 294854
rect 113546 258938 113782 259174
rect 113866 258938 114102 259174
rect 113546 258618 113782 258854
rect 113866 258618 114102 258854
rect 113546 222938 113782 223174
rect 113866 222938 114102 223174
rect 113546 222618 113782 222854
rect 113866 222618 114102 222854
rect 113546 186938 113782 187174
rect 113866 186938 114102 187174
rect 113546 186618 113782 186854
rect 113866 186618 114102 186854
rect 113546 150938 113782 151174
rect 113866 150938 114102 151174
rect 113546 150618 113782 150854
rect 113866 150618 114102 150854
rect 113546 114938 113782 115174
rect 113866 114938 114102 115174
rect 113546 114618 113782 114854
rect 113866 114618 114102 114854
rect 113546 78938 113782 79174
rect 113866 78938 114102 79174
rect 113546 78618 113782 78854
rect 113866 78618 114102 78854
rect 113546 42938 113782 43174
rect 113866 42938 114102 43174
rect 113546 42618 113782 42854
rect 113866 42618 114102 42854
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 113546 -2502 113782 -2266
rect 113866 -2502 114102 -2266
rect 113546 -2822 113782 -2586
rect 113866 -2822 114102 -2586
rect 117266 694658 117502 694894
rect 117586 694658 117822 694894
rect 117266 694338 117502 694574
rect 117586 694338 117822 694574
rect 117266 658658 117502 658894
rect 117586 658658 117822 658894
rect 117266 658338 117502 658574
rect 117586 658338 117822 658574
rect 117266 622658 117502 622894
rect 117586 622658 117822 622894
rect 117266 622338 117502 622574
rect 117586 622338 117822 622574
rect 117266 586658 117502 586894
rect 117586 586658 117822 586894
rect 117266 586338 117502 586574
rect 117586 586338 117822 586574
rect 117266 550658 117502 550894
rect 117586 550658 117822 550894
rect 117266 550338 117502 550574
rect 117586 550338 117822 550574
rect 117266 514658 117502 514894
rect 117586 514658 117822 514894
rect 117266 514338 117502 514574
rect 117586 514338 117822 514574
rect 117266 478658 117502 478894
rect 117586 478658 117822 478894
rect 117266 478338 117502 478574
rect 117586 478338 117822 478574
rect 117266 442658 117502 442894
rect 117586 442658 117822 442894
rect 117266 442338 117502 442574
rect 117586 442338 117822 442574
rect 117266 406658 117502 406894
rect 117586 406658 117822 406894
rect 117266 406338 117502 406574
rect 117586 406338 117822 406574
rect 117266 370658 117502 370894
rect 117586 370658 117822 370894
rect 117266 370338 117502 370574
rect 117586 370338 117822 370574
rect 117266 334658 117502 334894
rect 117586 334658 117822 334894
rect 117266 334338 117502 334574
rect 117586 334338 117822 334574
rect 117266 298658 117502 298894
rect 117586 298658 117822 298894
rect 117266 298338 117502 298574
rect 117586 298338 117822 298574
rect 117266 262658 117502 262894
rect 117586 262658 117822 262894
rect 117266 262338 117502 262574
rect 117586 262338 117822 262574
rect 117266 226658 117502 226894
rect 117586 226658 117822 226894
rect 117266 226338 117502 226574
rect 117586 226338 117822 226574
rect 117266 190658 117502 190894
rect 117586 190658 117822 190894
rect 117266 190338 117502 190574
rect 117586 190338 117822 190574
rect 117266 154658 117502 154894
rect 117586 154658 117822 154894
rect 117266 154338 117502 154574
rect 117586 154338 117822 154574
rect 117266 118658 117502 118894
rect 117586 118658 117822 118894
rect 117266 118338 117502 118574
rect 117586 118338 117822 118574
rect 117266 82658 117502 82894
rect 117586 82658 117822 82894
rect 117266 82338 117502 82574
rect 117586 82338 117822 82574
rect 117266 46658 117502 46894
rect 117586 46658 117822 46894
rect 117266 46338 117502 46574
rect 117586 46338 117822 46574
rect 117266 10658 117502 10894
rect 117586 10658 117822 10894
rect 117266 10338 117502 10574
rect 117586 10338 117822 10574
rect 117266 -4422 117502 -4186
rect 117586 -4422 117822 -4186
rect 117266 -4742 117502 -4506
rect 117586 -4742 117822 -4506
rect 138986 711322 139222 711558
rect 139306 711322 139542 711558
rect 138986 711002 139222 711238
rect 139306 711002 139542 711238
rect 135266 709402 135502 709638
rect 135586 709402 135822 709638
rect 135266 709082 135502 709318
rect 135586 709082 135822 709318
rect 131546 707482 131782 707718
rect 131866 707482 132102 707718
rect 131546 707162 131782 707398
rect 131866 707162 132102 707398
rect 120986 698378 121222 698614
rect 121306 698378 121542 698614
rect 120986 698058 121222 698294
rect 121306 698058 121542 698294
rect 120986 662378 121222 662614
rect 121306 662378 121542 662614
rect 120986 662058 121222 662294
rect 121306 662058 121542 662294
rect 120986 626378 121222 626614
rect 121306 626378 121542 626614
rect 120986 626058 121222 626294
rect 121306 626058 121542 626294
rect 120986 590378 121222 590614
rect 121306 590378 121542 590614
rect 120986 590058 121222 590294
rect 121306 590058 121542 590294
rect 120986 554378 121222 554614
rect 121306 554378 121542 554614
rect 120986 554058 121222 554294
rect 121306 554058 121542 554294
rect 120986 518378 121222 518614
rect 121306 518378 121542 518614
rect 120986 518058 121222 518294
rect 121306 518058 121542 518294
rect 120986 482378 121222 482614
rect 121306 482378 121542 482614
rect 120986 482058 121222 482294
rect 121306 482058 121542 482294
rect 120986 446378 121222 446614
rect 121306 446378 121542 446614
rect 120986 446058 121222 446294
rect 121306 446058 121542 446294
rect 120986 410378 121222 410614
rect 121306 410378 121542 410614
rect 120986 410058 121222 410294
rect 121306 410058 121542 410294
rect 120986 374378 121222 374614
rect 121306 374378 121542 374614
rect 120986 374058 121222 374294
rect 121306 374058 121542 374294
rect 120986 338378 121222 338614
rect 121306 338378 121542 338614
rect 120986 338058 121222 338294
rect 121306 338058 121542 338294
rect 120986 302378 121222 302614
rect 121306 302378 121542 302614
rect 120986 302058 121222 302294
rect 121306 302058 121542 302294
rect 120986 266378 121222 266614
rect 121306 266378 121542 266614
rect 120986 266058 121222 266294
rect 121306 266058 121542 266294
rect 120986 230378 121222 230614
rect 121306 230378 121542 230614
rect 120986 230058 121222 230294
rect 121306 230058 121542 230294
rect 120986 194378 121222 194614
rect 121306 194378 121542 194614
rect 120986 194058 121222 194294
rect 121306 194058 121542 194294
rect 120986 158378 121222 158614
rect 121306 158378 121542 158614
rect 120986 158058 121222 158294
rect 121306 158058 121542 158294
rect 120986 122378 121222 122614
rect 121306 122378 121542 122614
rect 120986 122058 121222 122294
rect 121306 122058 121542 122294
rect 120986 86378 121222 86614
rect 121306 86378 121542 86614
rect 120986 86058 121222 86294
rect 121306 86058 121542 86294
rect 120986 50378 121222 50614
rect 121306 50378 121542 50614
rect 120986 50058 121222 50294
rect 121306 50058 121542 50294
rect 120986 14378 121222 14614
rect 121306 14378 121542 14614
rect 120986 14058 121222 14294
rect 121306 14058 121542 14294
rect 102986 -7302 103222 -7066
rect 103306 -7302 103542 -7066
rect 102986 -7622 103222 -7386
rect 103306 -7622 103542 -7386
rect 127826 705562 128062 705798
rect 128146 705562 128382 705798
rect 127826 705242 128062 705478
rect 128146 705242 128382 705478
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 127826 561218 128062 561454
rect 128146 561218 128382 561454
rect 127826 560898 128062 561134
rect 128146 560898 128382 561134
rect 127826 525218 128062 525454
rect 128146 525218 128382 525454
rect 127826 524898 128062 525134
rect 128146 524898 128382 525134
rect 127826 489218 128062 489454
rect 128146 489218 128382 489454
rect 127826 488898 128062 489134
rect 128146 488898 128382 489134
rect 127826 453218 128062 453454
rect 128146 453218 128382 453454
rect 127826 452898 128062 453134
rect 128146 452898 128382 453134
rect 127826 417218 128062 417454
rect 128146 417218 128382 417454
rect 127826 416898 128062 417134
rect 128146 416898 128382 417134
rect 127826 381218 128062 381454
rect 128146 381218 128382 381454
rect 127826 380898 128062 381134
rect 128146 380898 128382 381134
rect 127826 345218 128062 345454
rect 128146 345218 128382 345454
rect 127826 344898 128062 345134
rect 128146 344898 128382 345134
rect 127826 309218 128062 309454
rect 128146 309218 128382 309454
rect 127826 308898 128062 309134
rect 128146 308898 128382 309134
rect 127826 273218 128062 273454
rect 128146 273218 128382 273454
rect 127826 272898 128062 273134
rect 128146 272898 128382 273134
rect 127826 237218 128062 237454
rect 128146 237218 128382 237454
rect 127826 236898 128062 237134
rect 128146 236898 128382 237134
rect 127826 201218 128062 201454
rect 128146 201218 128382 201454
rect 127826 200898 128062 201134
rect 128146 200898 128382 201134
rect 127826 165218 128062 165454
rect 128146 165218 128382 165454
rect 127826 164898 128062 165134
rect 128146 164898 128382 165134
rect 127826 129218 128062 129454
rect 128146 129218 128382 129454
rect 127826 128898 128062 129134
rect 128146 128898 128382 129134
rect 127826 93218 128062 93454
rect 128146 93218 128382 93454
rect 127826 92898 128062 93134
rect 128146 92898 128382 93134
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -1542 128062 -1306
rect 128146 -1542 128382 -1306
rect 127826 -1862 128062 -1626
rect 128146 -1862 128382 -1626
rect 131546 672938 131782 673174
rect 131866 672938 132102 673174
rect 131546 672618 131782 672854
rect 131866 672618 132102 672854
rect 131546 636938 131782 637174
rect 131866 636938 132102 637174
rect 131546 636618 131782 636854
rect 131866 636618 132102 636854
rect 131546 600938 131782 601174
rect 131866 600938 132102 601174
rect 131546 600618 131782 600854
rect 131866 600618 132102 600854
rect 131546 564938 131782 565174
rect 131866 564938 132102 565174
rect 131546 564618 131782 564854
rect 131866 564618 132102 564854
rect 131546 528938 131782 529174
rect 131866 528938 132102 529174
rect 131546 528618 131782 528854
rect 131866 528618 132102 528854
rect 131546 492938 131782 493174
rect 131866 492938 132102 493174
rect 131546 492618 131782 492854
rect 131866 492618 132102 492854
rect 131546 456938 131782 457174
rect 131866 456938 132102 457174
rect 131546 456618 131782 456854
rect 131866 456618 132102 456854
rect 131546 420938 131782 421174
rect 131866 420938 132102 421174
rect 131546 420618 131782 420854
rect 131866 420618 132102 420854
rect 131546 384938 131782 385174
rect 131866 384938 132102 385174
rect 131546 384618 131782 384854
rect 131866 384618 132102 384854
rect 131546 348938 131782 349174
rect 131866 348938 132102 349174
rect 131546 348618 131782 348854
rect 131866 348618 132102 348854
rect 131546 312938 131782 313174
rect 131866 312938 132102 313174
rect 131546 312618 131782 312854
rect 131866 312618 132102 312854
rect 131546 276938 131782 277174
rect 131866 276938 132102 277174
rect 131546 276618 131782 276854
rect 131866 276618 132102 276854
rect 131546 240938 131782 241174
rect 131866 240938 132102 241174
rect 131546 240618 131782 240854
rect 131866 240618 132102 240854
rect 131546 204938 131782 205174
rect 131866 204938 132102 205174
rect 131546 204618 131782 204854
rect 131866 204618 132102 204854
rect 131546 168938 131782 169174
rect 131866 168938 132102 169174
rect 131546 168618 131782 168854
rect 131866 168618 132102 168854
rect 131546 132938 131782 133174
rect 131866 132938 132102 133174
rect 131546 132618 131782 132854
rect 131866 132618 132102 132854
rect 131546 96938 131782 97174
rect 131866 96938 132102 97174
rect 131546 96618 131782 96854
rect 131866 96618 132102 96854
rect 131546 60938 131782 61174
rect 131866 60938 132102 61174
rect 131546 60618 131782 60854
rect 131866 60618 132102 60854
rect 131546 24938 131782 25174
rect 131866 24938 132102 25174
rect 131546 24618 131782 24854
rect 131866 24618 132102 24854
rect 131546 -3462 131782 -3226
rect 131866 -3462 132102 -3226
rect 131546 -3782 131782 -3546
rect 131866 -3782 132102 -3546
rect 135266 676658 135502 676894
rect 135586 676658 135822 676894
rect 135266 676338 135502 676574
rect 135586 676338 135822 676574
rect 135266 640658 135502 640894
rect 135586 640658 135822 640894
rect 135266 640338 135502 640574
rect 135586 640338 135822 640574
rect 135266 604658 135502 604894
rect 135586 604658 135822 604894
rect 135266 604338 135502 604574
rect 135586 604338 135822 604574
rect 135266 568658 135502 568894
rect 135586 568658 135822 568894
rect 135266 568338 135502 568574
rect 135586 568338 135822 568574
rect 135266 532658 135502 532894
rect 135586 532658 135822 532894
rect 135266 532338 135502 532574
rect 135586 532338 135822 532574
rect 135266 496658 135502 496894
rect 135586 496658 135822 496894
rect 135266 496338 135502 496574
rect 135586 496338 135822 496574
rect 135266 460658 135502 460894
rect 135586 460658 135822 460894
rect 135266 460338 135502 460574
rect 135586 460338 135822 460574
rect 135266 424658 135502 424894
rect 135586 424658 135822 424894
rect 135266 424338 135502 424574
rect 135586 424338 135822 424574
rect 135266 388658 135502 388894
rect 135586 388658 135822 388894
rect 135266 388338 135502 388574
rect 135586 388338 135822 388574
rect 135266 352658 135502 352894
rect 135586 352658 135822 352894
rect 135266 352338 135502 352574
rect 135586 352338 135822 352574
rect 135266 316658 135502 316894
rect 135586 316658 135822 316894
rect 135266 316338 135502 316574
rect 135586 316338 135822 316574
rect 135266 280658 135502 280894
rect 135586 280658 135822 280894
rect 135266 280338 135502 280574
rect 135586 280338 135822 280574
rect 135266 244658 135502 244894
rect 135586 244658 135822 244894
rect 135266 244338 135502 244574
rect 135586 244338 135822 244574
rect 135266 208658 135502 208894
rect 135586 208658 135822 208894
rect 135266 208338 135502 208574
rect 135586 208338 135822 208574
rect 135266 172658 135502 172894
rect 135586 172658 135822 172894
rect 135266 172338 135502 172574
rect 135586 172338 135822 172574
rect 135266 136658 135502 136894
rect 135586 136658 135822 136894
rect 135266 136338 135502 136574
rect 135586 136338 135822 136574
rect 135266 100658 135502 100894
rect 135586 100658 135822 100894
rect 135266 100338 135502 100574
rect 135586 100338 135822 100574
rect 135266 64658 135502 64894
rect 135586 64658 135822 64894
rect 135266 64338 135502 64574
rect 135586 64338 135822 64574
rect 135266 28658 135502 28894
rect 135586 28658 135822 28894
rect 135266 28338 135502 28574
rect 135586 28338 135822 28574
rect 135266 -5382 135502 -5146
rect 135586 -5382 135822 -5146
rect 135266 -5702 135502 -5466
rect 135586 -5702 135822 -5466
rect 156986 710362 157222 710598
rect 157306 710362 157542 710598
rect 156986 710042 157222 710278
rect 157306 710042 157542 710278
rect 153266 708442 153502 708678
rect 153586 708442 153822 708678
rect 153266 708122 153502 708358
rect 153586 708122 153822 708358
rect 149546 706522 149782 706758
rect 149866 706522 150102 706758
rect 149546 706202 149782 706438
rect 149866 706202 150102 706438
rect 138986 680378 139222 680614
rect 139306 680378 139542 680614
rect 138986 680058 139222 680294
rect 139306 680058 139542 680294
rect 138986 644378 139222 644614
rect 139306 644378 139542 644614
rect 138986 644058 139222 644294
rect 139306 644058 139542 644294
rect 138986 608378 139222 608614
rect 139306 608378 139542 608614
rect 138986 608058 139222 608294
rect 139306 608058 139542 608294
rect 138986 572378 139222 572614
rect 139306 572378 139542 572614
rect 138986 572058 139222 572294
rect 139306 572058 139542 572294
rect 138986 536378 139222 536614
rect 139306 536378 139542 536614
rect 138986 536058 139222 536294
rect 139306 536058 139542 536294
rect 138986 500378 139222 500614
rect 139306 500378 139542 500614
rect 138986 500058 139222 500294
rect 139306 500058 139542 500294
rect 138986 464378 139222 464614
rect 139306 464378 139542 464614
rect 138986 464058 139222 464294
rect 139306 464058 139542 464294
rect 138986 428378 139222 428614
rect 139306 428378 139542 428614
rect 138986 428058 139222 428294
rect 139306 428058 139542 428294
rect 138986 392378 139222 392614
rect 139306 392378 139542 392614
rect 138986 392058 139222 392294
rect 139306 392058 139542 392294
rect 138986 356378 139222 356614
rect 139306 356378 139542 356614
rect 138986 356058 139222 356294
rect 139306 356058 139542 356294
rect 138986 320378 139222 320614
rect 139306 320378 139542 320614
rect 138986 320058 139222 320294
rect 139306 320058 139542 320294
rect 138986 284378 139222 284614
rect 139306 284378 139542 284614
rect 138986 284058 139222 284294
rect 139306 284058 139542 284294
rect 138986 248378 139222 248614
rect 139306 248378 139542 248614
rect 138986 248058 139222 248294
rect 139306 248058 139542 248294
rect 138986 212378 139222 212614
rect 139306 212378 139542 212614
rect 138986 212058 139222 212294
rect 139306 212058 139542 212294
rect 138986 176378 139222 176614
rect 139306 176378 139542 176614
rect 138986 176058 139222 176294
rect 139306 176058 139542 176294
rect 138986 140378 139222 140614
rect 139306 140378 139542 140614
rect 138986 140058 139222 140294
rect 139306 140058 139542 140294
rect 138986 104378 139222 104614
rect 139306 104378 139542 104614
rect 138986 104058 139222 104294
rect 139306 104058 139542 104294
rect 138986 68378 139222 68614
rect 139306 68378 139542 68614
rect 138986 68058 139222 68294
rect 139306 68058 139542 68294
rect 138986 32378 139222 32614
rect 139306 32378 139542 32614
rect 138986 32058 139222 32294
rect 139306 32058 139542 32294
rect 120986 -6342 121222 -6106
rect 121306 -6342 121542 -6106
rect 120986 -6662 121222 -6426
rect 121306 -6662 121542 -6426
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 145826 507218 146062 507454
rect 146146 507218 146382 507454
rect 145826 506898 146062 507134
rect 146146 506898 146382 507134
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 145826 435218 146062 435454
rect 146146 435218 146382 435454
rect 145826 434898 146062 435134
rect 146146 434898 146382 435134
rect 145826 399218 146062 399454
rect 146146 399218 146382 399454
rect 145826 398898 146062 399134
rect 146146 398898 146382 399134
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 145826 327218 146062 327454
rect 146146 327218 146382 327454
rect 145826 326898 146062 327134
rect 146146 326898 146382 327134
rect 145826 291218 146062 291454
rect 146146 291218 146382 291454
rect 145826 290898 146062 291134
rect 146146 290898 146382 291134
rect 145826 255218 146062 255454
rect 146146 255218 146382 255454
rect 145826 254898 146062 255134
rect 146146 254898 146382 255134
rect 145826 219218 146062 219454
rect 146146 219218 146382 219454
rect 145826 218898 146062 219134
rect 146146 218898 146382 219134
rect 145826 183218 146062 183454
rect 146146 183218 146382 183454
rect 145826 182898 146062 183134
rect 146146 182898 146382 183134
rect 145826 147218 146062 147454
rect 146146 147218 146382 147454
rect 145826 146898 146062 147134
rect 146146 146898 146382 147134
rect 145826 111218 146062 111454
rect 146146 111218 146382 111454
rect 145826 110898 146062 111134
rect 146146 110898 146382 111134
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 149546 654938 149782 655174
rect 149866 654938 150102 655174
rect 149546 654618 149782 654854
rect 149866 654618 150102 654854
rect 149546 618938 149782 619174
rect 149866 618938 150102 619174
rect 149546 618618 149782 618854
rect 149866 618618 150102 618854
rect 149546 582938 149782 583174
rect 149866 582938 150102 583174
rect 149546 582618 149782 582854
rect 149866 582618 150102 582854
rect 149546 546938 149782 547174
rect 149866 546938 150102 547174
rect 149546 546618 149782 546854
rect 149866 546618 150102 546854
rect 149546 510938 149782 511174
rect 149866 510938 150102 511174
rect 149546 510618 149782 510854
rect 149866 510618 150102 510854
rect 149546 474938 149782 475174
rect 149866 474938 150102 475174
rect 149546 474618 149782 474854
rect 149866 474618 150102 474854
rect 149546 438938 149782 439174
rect 149866 438938 150102 439174
rect 149546 438618 149782 438854
rect 149866 438618 150102 438854
rect 149546 402938 149782 403174
rect 149866 402938 150102 403174
rect 149546 402618 149782 402854
rect 149866 402618 150102 402854
rect 149546 366938 149782 367174
rect 149866 366938 150102 367174
rect 149546 366618 149782 366854
rect 149866 366618 150102 366854
rect 149546 330938 149782 331174
rect 149866 330938 150102 331174
rect 149546 330618 149782 330854
rect 149866 330618 150102 330854
rect 149546 294938 149782 295174
rect 149866 294938 150102 295174
rect 149546 294618 149782 294854
rect 149866 294618 150102 294854
rect 149546 258938 149782 259174
rect 149866 258938 150102 259174
rect 149546 258618 149782 258854
rect 149866 258618 150102 258854
rect 149546 222938 149782 223174
rect 149866 222938 150102 223174
rect 149546 222618 149782 222854
rect 149866 222618 150102 222854
rect 149546 186938 149782 187174
rect 149866 186938 150102 187174
rect 149546 186618 149782 186854
rect 149866 186618 150102 186854
rect 149546 150938 149782 151174
rect 149866 150938 150102 151174
rect 149546 150618 149782 150854
rect 149866 150618 150102 150854
rect 149546 114938 149782 115174
rect 149866 114938 150102 115174
rect 149546 114618 149782 114854
rect 149866 114618 150102 114854
rect 149546 78938 149782 79174
rect 149866 78938 150102 79174
rect 149546 78618 149782 78854
rect 149866 78618 150102 78854
rect 149546 42938 149782 43174
rect 149866 42938 150102 43174
rect 149546 42618 149782 42854
rect 149866 42618 150102 42854
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 149546 -2502 149782 -2266
rect 149866 -2502 150102 -2266
rect 149546 -2822 149782 -2586
rect 149866 -2822 150102 -2586
rect 153266 694658 153502 694894
rect 153586 694658 153822 694894
rect 153266 694338 153502 694574
rect 153586 694338 153822 694574
rect 153266 658658 153502 658894
rect 153586 658658 153822 658894
rect 153266 658338 153502 658574
rect 153586 658338 153822 658574
rect 153266 622658 153502 622894
rect 153586 622658 153822 622894
rect 153266 622338 153502 622574
rect 153586 622338 153822 622574
rect 153266 586658 153502 586894
rect 153586 586658 153822 586894
rect 153266 586338 153502 586574
rect 153586 586338 153822 586574
rect 153266 550658 153502 550894
rect 153586 550658 153822 550894
rect 153266 550338 153502 550574
rect 153586 550338 153822 550574
rect 153266 514658 153502 514894
rect 153586 514658 153822 514894
rect 153266 514338 153502 514574
rect 153586 514338 153822 514574
rect 153266 478658 153502 478894
rect 153586 478658 153822 478894
rect 153266 478338 153502 478574
rect 153586 478338 153822 478574
rect 153266 442658 153502 442894
rect 153586 442658 153822 442894
rect 153266 442338 153502 442574
rect 153586 442338 153822 442574
rect 153266 406658 153502 406894
rect 153586 406658 153822 406894
rect 153266 406338 153502 406574
rect 153586 406338 153822 406574
rect 153266 370658 153502 370894
rect 153586 370658 153822 370894
rect 153266 370338 153502 370574
rect 153586 370338 153822 370574
rect 153266 334658 153502 334894
rect 153586 334658 153822 334894
rect 153266 334338 153502 334574
rect 153586 334338 153822 334574
rect 153266 298658 153502 298894
rect 153586 298658 153822 298894
rect 153266 298338 153502 298574
rect 153586 298338 153822 298574
rect 153266 262658 153502 262894
rect 153586 262658 153822 262894
rect 153266 262338 153502 262574
rect 153586 262338 153822 262574
rect 153266 226658 153502 226894
rect 153586 226658 153822 226894
rect 153266 226338 153502 226574
rect 153586 226338 153822 226574
rect 153266 190658 153502 190894
rect 153586 190658 153822 190894
rect 153266 190338 153502 190574
rect 153586 190338 153822 190574
rect 153266 154658 153502 154894
rect 153586 154658 153822 154894
rect 153266 154338 153502 154574
rect 153586 154338 153822 154574
rect 153266 118658 153502 118894
rect 153586 118658 153822 118894
rect 153266 118338 153502 118574
rect 153586 118338 153822 118574
rect 153266 82658 153502 82894
rect 153586 82658 153822 82894
rect 153266 82338 153502 82574
rect 153586 82338 153822 82574
rect 153266 46658 153502 46894
rect 153586 46658 153822 46894
rect 153266 46338 153502 46574
rect 153586 46338 153822 46574
rect 153266 10658 153502 10894
rect 153586 10658 153822 10894
rect 153266 10338 153502 10574
rect 153586 10338 153822 10574
rect 153266 -4422 153502 -4186
rect 153586 -4422 153822 -4186
rect 153266 -4742 153502 -4506
rect 153586 -4742 153822 -4506
rect 174986 711322 175222 711558
rect 175306 711322 175542 711558
rect 174986 711002 175222 711238
rect 175306 711002 175542 711238
rect 171266 709402 171502 709638
rect 171586 709402 171822 709638
rect 171266 709082 171502 709318
rect 171586 709082 171822 709318
rect 167546 707482 167782 707718
rect 167866 707482 168102 707718
rect 167546 707162 167782 707398
rect 167866 707162 168102 707398
rect 156986 698378 157222 698614
rect 157306 698378 157542 698614
rect 156986 698058 157222 698294
rect 157306 698058 157542 698294
rect 156986 662378 157222 662614
rect 157306 662378 157542 662614
rect 156986 662058 157222 662294
rect 157306 662058 157542 662294
rect 156986 626378 157222 626614
rect 157306 626378 157542 626614
rect 156986 626058 157222 626294
rect 157306 626058 157542 626294
rect 156986 590378 157222 590614
rect 157306 590378 157542 590614
rect 156986 590058 157222 590294
rect 157306 590058 157542 590294
rect 156986 554378 157222 554614
rect 157306 554378 157542 554614
rect 156986 554058 157222 554294
rect 157306 554058 157542 554294
rect 156986 518378 157222 518614
rect 157306 518378 157542 518614
rect 156986 518058 157222 518294
rect 157306 518058 157542 518294
rect 156986 482378 157222 482614
rect 157306 482378 157542 482614
rect 156986 482058 157222 482294
rect 157306 482058 157542 482294
rect 156986 446378 157222 446614
rect 157306 446378 157542 446614
rect 156986 446058 157222 446294
rect 157306 446058 157542 446294
rect 156986 410378 157222 410614
rect 157306 410378 157542 410614
rect 156986 410058 157222 410294
rect 157306 410058 157542 410294
rect 156986 374378 157222 374614
rect 157306 374378 157542 374614
rect 156986 374058 157222 374294
rect 157306 374058 157542 374294
rect 156986 338378 157222 338614
rect 157306 338378 157542 338614
rect 156986 338058 157222 338294
rect 157306 338058 157542 338294
rect 156986 302378 157222 302614
rect 157306 302378 157542 302614
rect 156986 302058 157222 302294
rect 157306 302058 157542 302294
rect 156986 266378 157222 266614
rect 157306 266378 157542 266614
rect 156986 266058 157222 266294
rect 157306 266058 157542 266294
rect 156986 230378 157222 230614
rect 157306 230378 157542 230614
rect 156986 230058 157222 230294
rect 157306 230058 157542 230294
rect 156986 194378 157222 194614
rect 157306 194378 157542 194614
rect 156986 194058 157222 194294
rect 157306 194058 157542 194294
rect 163826 705562 164062 705798
rect 164146 705562 164382 705798
rect 163826 705242 164062 705478
rect 164146 705242 164382 705478
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 163826 561218 164062 561454
rect 164146 561218 164382 561454
rect 163826 560898 164062 561134
rect 164146 560898 164382 561134
rect 163826 525218 164062 525454
rect 164146 525218 164382 525454
rect 163826 524898 164062 525134
rect 164146 524898 164382 525134
rect 163826 489218 164062 489454
rect 164146 489218 164382 489454
rect 163826 488898 164062 489134
rect 164146 488898 164382 489134
rect 163826 453218 164062 453454
rect 164146 453218 164382 453454
rect 163826 452898 164062 453134
rect 164146 452898 164382 453134
rect 163826 417218 164062 417454
rect 164146 417218 164382 417454
rect 163826 416898 164062 417134
rect 164146 416898 164382 417134
rect 163826 381218 164062 381454
rect 164146 381218 164382 381454
rect 163826 380898 164062 381134
rect 164146 380898 164382 381134
rect 163826 345218 164062 345454
rect 164146 345218 164382 345454
rect 163826 344898 164062 345134
rect 164146 344898 164382 345134
rect 163826 309218 164062 309454
rect 164146 309218 164382 309454
rect 163826 308898 164062 309134
rect 164146 308898 164382 309134
rect 163826 273218 164062 273454
rect 164146 273218 164382 273454
rect 163826 272898 164062 273134
rect 164146 272898 164382 273134
rect 163826 237218 164062 237454
rect 164146 237218 164382 237454
rect 163826 236898 164062 237134
rect 164146 236898 164382 237134
rect 163826 201218 164062 201454
rect 164146 201218 164382 201454
rect 163826 200898 164062 201134
rect 164146 200898 164382 201134
rect 167546 672938 167782 673174
rect 167866 672938 168102 673174
rect 167546 672618 167782 672854
rect 167866 672618 168102 672854
rect 167546 636938 167782 637174
rect 167866 636938 168102 637174
rect 167546 636618 167782 636854
rect 167866 636618 168102 636854
rect 167546 600938 167782 601174
rect 167866 600938 168102 601174
rect 167546 600618 167782 600854
rect 167866 600618 168102 600854
rect 167546 564938 167782 565174
rect 167866 564938 168102 565174
rect 167546 564618 167782 564854
rect 167866 564618 168102 564854
rect 167546 528938 167782 529174
rect 167866 528938 168102 529174
rect 167546 528618 167782 528854
rect 167866 528618 168102 528854
rect 167546 492938 167782 493174
rect 167866 492938 168102 493174
rect 167546 492618 167782 492854
rect 167866 492618 168102 492854
rect 167546 456938 167782 457174
rect 167866 456938 168102 457174
rect 167546 456618 167782 456854
rect 167866 456618 168102 456854
rect 167546 420938 167782 421174
rect 167866 420938 168102 421174
rect 167546 420618 167782 420854
rect 167866 420618 168102 420854
rect 167546 384938 167782 385174
rect 167866 384938 168102 385174
rect 167546 384618 167782 384854
rect 167866 384618 168102 384854
rect 167546 348938 167782 349174
rect 167866 348938 168102 349174
rect 167546 348618 167782 348854
rect 167866 348618 168102 348854
rect 167546 312938 167782 313174
rect 167866 312938 168102 313174
rect 167546 312618 167782 312854
rect 167866 312618 168102 312854
rect 167546 276938 167782 277174
rect 167866 276938 168102 277174
rect 167546 276618 167782 276854
rect 167866 276618 168102 276854
rect 167546 240938 167782 241174
rect 167866 240938 168102 241174
rect 167546 240618 167782 240854
rect 167866 240618 168102 240854
rect 167546 204938 167782 205174
rect 167866 204938 168102 205174
rect 167546 204618 167782 204854
rect 167866 204618 168102 204854
rect 171266 676658 171502 676894
rect 171586 676658 171822 676894
rect 171266 676338 171502 676574
rect 171586 676338 171822 676574
rect 171266 640658 171502 640894
rect 171586 640658 171822 640894
rect 171266 640338 171502 640574
rect 171586 640338 171822 640574
rect 171266 604658 171502 604894
rect 171586 604658 171822 604894
rect 171266 604338 171502 604574
rect 171586 604338 171822 604574
rect 171266 568658 171502 568894
rect 171586 568658 171822 568894
rect 171266 568338 171502 568574
rect 171586 568338 171822 568574
rect 171266 532658 171502 532894
rect 171586 532658 171822 532894
rect 171266 532338 171502 532574
rect 171586 532338 171822 532574
rect 171266 496658 171502 496894
rect 171586 496658 171822 496894
rect 171266 496338 171502 496574
rect 171586 496338 171822 496574
rect 171266 460658 171502 460894
rect 171586 460658 171822 460894
rect 171266 460338 171502 460574
rect 171586 460338 171822 460574
rect 171266 424658 171502 424894
rect 171586 424658 171822 424894
rect 171266 424338 171502 424574
rect 171586 424338 171822 424574
rect 171266 388658 171502 388894
rect 171586 388658 171822 388894
rect 171266 388338 171502 388574
rect 171586 388338 171822 388574
rect 171266 352658 171502 352894
rect 171586 352658 171822 352894
rect 171266 352338 171502 352574
rect 171586 352338 171822 352574
rect 171266 316658 171502 316894
rect 171586 316658 171822 316894
rect 171266 316338 171502 316574
rect 171586 316338 171822 316574
rect 171266 280658 171502 280894
rect 171586 280658 171822 280894
rect 171266 280338 171502 280574
rect 171586 280338 171822 280574
rect 171266 244658 171502 244894
rect 171586 244658 171822 244894
rect 171266 244338 171502 244574
rect 171586 244338 171822 244574
rect 171266 208658 171502 208894
rect 171586 208658 171822 208894
rect 171266 208338 171502 208574
rect 171586 208338 171822 208574
rect 192986 710362 193222 710598
rect 193306 710362 193542 710598
rect 192986 710042 193222 710278
rect 193306 710042 193542 710278
rect 189266 708442 189502 708678
rect 189586 708442 189822 708678
rect 189266 708122 189502 708358
rect 189586 708122 189822 708358
rect 185546 706522 185782 706758
rect 185866 706522 186102 706758
rect 185546 706202 185782 706438
rect 185866 706202 186102 706438
rect 174986 680378 175222 680614
rect 175306 680378 175542 680614
rect 174986 680058 175222 680294
rect 175306 680058 175542 680294
rect 174986 644378 175222 644614
rect 175306 644378 175542 644614
rect 174986 644058 175222 644294
rect 175306 644058 175542 644294
rect 174986 608378 175222 608614
rect 175306 608378 175542 608614
rect 174986 608058 175222 608294
rect 175306 608058 175542 608294
rect 174986 572378 175222 572614
rect 175306 572378 175542 572614
rect 174986 572058 175222 572294
rect 175306 572058 175542 572294
rect 174986 536378 175222 536614
rect 175306 536378 175542 536614
rect 174986 536058 175222 536294
rect 175306 536058 175542 536294
rect 174986 500378 175222 500614
rect 175306 500378 175542 500614
rect 174986 500058 175222 500294
rect 175306 500058 175542 500294
rect 174986 464378 175222 464614
rect 175306 464378 175542 464614
rect 174986 464058 175222 464294
rect 175306 464058 175542 464294
rect 174986 428378 175222 428614
rect 175306 428378 175542 428614
rect 174986 428058 175222 428294
rect 175306 428058 175542 428294
rect 174986 392378 175222 392614
rect 175306 392378 175542 392614
rect 174986 392058 175222 392294
rect 175306 392058 175542 392294
rect 174986 356378 175222 356614
rect 175306 356378 175542 356614
rect 174986 356058 175222 356294
rect 175306 356058 175542 356294
rect 174986 320378 175222 320614
rect 175306 320378 175542 320614
rect 174986 320058 175222 320294
rect 175306 320058 175542 320294
rect 174986 284378 175222 284614
rect 175306 284378 175542 284614
rect 174986 284058 175222 284294
rect 175306 284058 175542 284294
rect 174986 248378 175222 248614
rect 175306 248378 175542 248614
rect 174986 248058 175222 248294
rect 175306 248058 175542 248294
rect 174986 212378 175222 212614
rect 175306 212378 175542 212614
rect 174986 212058 175222 212294
rect 175306 212058 175542 212294
rect 162285 183218 162521 183454
rect 162285 182898 162521 183134
rect 164882 183218 165118 183454
rect 164882 182898 165118 183134
rect 167479 183218 167715 183454
rect 167479 182898 167715 183134
rect 174986 176378 175222 176614
rect 175306 176378 175542 176614
rect 174986 176058 175222 176294
rect 175306 176058 175542 176294
rect 163583 165218 163819 165454
rect 163583 164898 163819 165134
rect 166180 165218 166416 165454
rect 166180 164898 166416 165134
rect 156986 158378 157222 158614
rect 157306 158378 157542 158614
rect 156986 158058 157222 158294
rect 157306 158058 157542 158294
rect 162285 147218 162521 147454
rect 162285 146898 162521 147134
rect 164882 147218 165118 147454
rect 164882 146898 165118 147134
rect 167479 147218 167715 147454
rect 167479 146898 167715 147134
rect 174986 140378 175222 140614
rect 175306 140378 175542 140614
rect 174986 140058 175222 140294
rect 175306 140058 175542 140294
rect 163583 129218 163819 129454
rect 163583 128898 163819 129134
rect 166180 129218 166416 129454
rect 166180 128898 166416 129134
rect 156986 122378 157222 122614
rect 157306 122378 157542 122614
rect 156986 122058 157222 122294
rect 157306 122058 157542 122294
rect 156986 86378 157222 86614
rect 157306 86378 157542 86614
rect 156986 86058 157222 86294
rect 157306 86058 157542 86294
rect 156986 50378 157222 50614
rect 157306 50378 157542 50614
rect 156986 50058 157222 50294
rect 157306 50058 157542 50294
rect 156986 14378 157222 14614
rect 157306 14378 157542 14614
rect 156986 14058 157222 14294
rect 157306 14058 157542 14294
rect 138986 -7302 139222 -7066
rect 139306 -7302 139542 -7066
rect 138986 -7622 139222 -7386
rect 139306 -7622 139542 -7386
rect 163826 93218 164062 93454
rect 164146 93218 164382 93454
rect 163826 92898 164062 93134
rect 164146 92898 164382 93134
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -1542 164062 -1306
rect 164146 -1542 164382 -1306
rect 163826 -1862 164062 -1626
rect 164146 -1862 164382 -1626
rect 167546 96938 167782 97174
rect 167866 96938 168102 97174
rect 167546 96618 167782 96854
rect 167866 96618 168102 96854
rect 167546 60938 167782 61174
rect 167866 60938 168102 61174
rect 167546 60618 167782 60854
rect 167866 60618 168102 60854
rect 167546 24938 167782 25174
rect 167866 24938 168102 25174
rect 167546 24618 167782 24854
rect 167866 24618 168102 24854
rect 167546 -3462 167782 -3226
rect 167866 -3462 168102 -3226
rect 167546 -3782 167782 -3546
rect 167866 -3782 168102 -3546
rect 171266 100658 171502 100894
rect 171586 100658 171822 100894
rect 171266 100338 171502 100574
rect 171586 100338 171822 100574
rect 171266 64658 171502 64894
rect 171586 64658 171822 64894
rect 171266 64338 171502 64574
rect 171586 64338 171822 64574
rect 171266 28658 171502 28894
rect 171586 28658 171822 28894
rect 171266 28338 171502 28574
rect 171586 28338 171822 28574
rect 171266 -5382 171502 -5146
rect 171586 -5382 171822 -5146
rect 171266 -5702 171502 -5466
rect 171586 -5702 171822 -5466
rect 174986 104378 175222 104614
rect 175306 104378 175542 104614
rect 174986 104058 175222 104294
rect 175306 104058 175542 104294
rect 174986 68378 175222 68614
rect 175306 68378 175542 68614
rect 174986 68058 175222 68294
rect 175306 68058 175542 68294
rect 174986 32378 175222 32614
rect 175306 32378 175542 32614
rect 174986 32058 175222 32294
rect 175306 32058 175542 32294
rect 156986 -6342 157222 -6106
rect 157306 -6342 157542 -6106
rect 156986 -6662 157222 -6426
rect 157306 -6662 157542 -6426
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 181826 435218 182062 435454
rect 182146 435218 182382 435454
rect 181826 434898 182062 435134
rect 182146 434898 182382 435134
rect 181826 399218 182062 399454
rect 182146 399218 182382 399454
rect 181826 398898 182062 399134
rect 182146 398898 182382 399134
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 181826 327218 182062 327454
rect 182146 327218 182382 327454
rect 181826 326898 182062 327134
rect 182146 326898 182382 327134
rect 181826 291218 182062 291454
rect 182146 291218 182382 291454
rect 181826 290898 182062 291134
rect 182146 290898 182382 291134
rect 181826 255218 182062 255454
rect 182146 255218 182382 255454
rect 181826 254898 182062 255134
rect 182146 254898 182382 255134
rect 181826 219218 182062 219454
rect 182146 219218 182382 219454
rect 181826 218898 182062 219134
rect 182146 218898 182382 219134
rect 181826 183218 182062 183454
rect 182146 183218 182382 183454
rect 181826 182898 182062 183134
rect 182146 182898 182382 183134
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 181826 111218 182062 111454
rect 182146 111218 182382 111454
rect 181826 110898 182062 111134
rect 182146 110898 182382 111134
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 185546 690938 185782 691174
rect 185866 690938 186102 691174
rect 185546 690618 185782 690854
rect 185866 690618 186102 690854
rect 185546 654938 185782 655174
rect 185866 654938 186102 655174
rect 185546 654618 185782 654854
rect 185866 654618 186102 654854
rect 185546 618938 185782 619174
rect 185866 618938 186102 619174
rect 185546 618618 185782 618854
rect 185866 618618 186102 618854
rect 185546 582938 185782 583174
rect 185866 582938 186102 583174
rect 185546 582618 185782 582854
rect 185866 582618 186102 582854
rect 185546 546938 185782 547174
rect 185866 546938 186102 547174
rect 185546 546618 185782 546854
rect 185866 546618 186102 546854
rect 185546 510938 185782 511174
rect 185866 510938 186102 511174
rect 185546 510618 185782 510854
rect 185866 510618 186102 510854
rect 185546 474938 185782 475174
rect 185866 474938 186102 475174
rect 185546 474618 185782 474854
rect 185866 474618 186102 474854
rect 185546 438938 185782 439174
rect 185866 438938 186102 439174
rect 185546 438618 185782 438854
rect 185866 438618 186102 438854
rect 185546 402938 185782 403174
rect 185866 402938 186102 403174
rect 185546 402618 185782 402854
rect 185866 402618 186102 402854
rect 185546 366938 185782 367174
rect 185866 366938 186102 367174
rect 185546 366618 185782 366854
rect 185866 366618 186102 366854
rect 185546 330938 185782 331174
rect 185866 330938 186102 331174
rect 185546 330618 185782 330854
rect 185866 330618 186102 330854
rect 185546 294938 185782 295174
rect 185866 294938 186102 295174
rect 185546 294618 185782 294854
rect 185866 294618 186102 294854
rect 185546 258938 185782 259174
rect 185866 258938 186102 259174
rect 185546 258618 185782 258854
rect 185866 258618 186102 258854
rect 185546 222938 185782 223174
rect 185866 222938 186102 223174
rect 185546 222618 185782 222854
rect 185866 222618 186102 222854
rect 185546 186938 185782 187174
rect 185866 186938 186102 187174
rect 185546 186618 185782 186854
rect 185866 186618 186102 186854
rect 185546 150938 185782 151174
rect 185866 150938 186102 151174
rect 185546 150618 185782 150854
rect 185866 150618 186102 150854
rect 185546 114938 185782 115174
rect 185866 114938 186102 115174
rect 185546 114618 185782 114854
rect 185866 114618 186102 114854
rect 185546 78938 185782 79174
rect 185866 78938 186102 79174
rect 185546 78618 185782 78854
rect 185866 78618 186102 78854
rect 185546 42938 185782 43174
rect 185866 42938 186102 43174
rect 185546 42618 185782 42854
rect 185866 42618 186102 42854
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 185546 -2502 185782 -2266
rect 185866 -2502 186102 -2266
rect 185546 -2822 185782 -2586
rect 185866 -2822 186102 -2586
rect 189266 694658 189502 694894
rect 189586 694658 189822 694894
rect 189266 694338 189502 694574
rect 189586 694338 189822 694574
rect 189266 658658 189502 658894
rect 189586 658658 189822 658894
rect 189266 658338 189502 658574
rect 189586 658338 189822 658574
rect 189266 622658 189502 622894
rect 189586 622658 189822 622894
rect 189266 622338 189502 622574
rect 189586 622338 189822 622574
rect 189266 586658 189502 586894
rect 189586 586658 189822 586894
rect 189266 586338 189502 586574
rect 189586 586338 189822 586574
rect 189266 550658 189502 550894
rect 189586 550658 189822 550894
rect 189266 550338 189502 550574
rect 189586 550338 189822 550574
rect 189266 514658 189502 514894
rect 189586 514658 189822 514894
rect 189266 514338 189502 514574
rect 189586 514338 189822 514574
rect 189266 478658 189502 478894
rect 189586 478658 189822 478894
rect 189266 478338 189502 478574
rect 189586 478338 189822 478574
rect 189266 442658 189502 442894
rect 189586 442658 189822 442894
rect 189266 442338 189502 442574
rect 189586 442338 189822 442574
rect 189266 406658 189502 406894
rect 189586 406658 189822 406894
rect 189266 406338 189502 406574
rect 189586 406338 189822 406574
rect 189266 370658 189502 370894
rect 189586 370658 189822 370894
rect 189266 370338 189502 370574
rect 189586 370338 189822 370574
rect 189266 334658 189502 334894
rect 189586 334658 189822 334894
rect 189266 334338 189502 334574
rect 189586 334338 189822 334574
rect 189266 298658 189502 298894
rect 189586 298658 189822 298894
rect 189266 298338 189502 298574
rect 189586 298338 189822 298574
rect 189266 262658 189502 262894
rect 189586 262658 189822 262894
rect 189266 262338 189502 262574
rect 189586 262338 189822 262574
rect 189266 226658 189502 226894
rect 189586 226658 189822 226894
rect 189266 226338 189502 226574
rect 189586 226338 189822 226574
rect 189266 190658 189502 190894
rect 189586 190658 189822 190894
rect 189266 190338 189502 190574
rect 189586 190338 189822 190574
rect 189266 154658 189502 154894
rect 189586 154658 189822 154894
rect 189266 154338 189502 154574
rect 189586 154338 189822 154574
rect 189266 118658 189502 118894
rect 189586 118658 189822 118894
rect 189266 118338 189502 118574
rect 189586 118338 189822 118574
rect 189266 82658 189502 82894
rect 189586 82658 189822 82894
rect 189266 82338 189502 82574
rect 189586 82338 189822 82574
rect 189266 46658 189502 46894
rect 189586 46658 189822 46894
rect 189266 46338 189502 46574
rect 189586 46338 189822 46574
rect 189266 10658 189502 10894
rect 189586 10658 189822 10894
rect 189266 10338 189502 10574
rect 189586 10338 189822 10574
rect 189266 -4422 189502 -4186
rect 189586 -4422 189822 -4186
rect 189266 -4742 189502 -4506
rect 189586 -4742 189822 -4506
rect 210986 711322 211222 711558
rect 211306 711322 211542 711558
rect 210986 711002 211222 711238
rect 211306 711002 211542 711238
rect 207266 709402 207502 709638
rect 207586 709402 207822 709638
rect 207266 709082 207502 709318
rect 207586 709082 207822 709318
rect 203546 707482 203782 707718
rect 203866 707482 204102 707718
rect 203546 707162 203782 707398
rect 203866 707162 204102 707398
rect 192986 698378 193222 698614
rect 193306 698378 193542 698614
rect 192986 698058 193222 698294
rect 193306 698058 193542 698294
rect 192986 662378 193222 662614
rect 193306 662378 193542 662614
rect 192986 662058 193222 662294
rect 193306 662058 193542 662294
rect 192986 626378 193222 626614
rect 193306 626378 193542 626614
rect 192986 626058 193222 626294
rect 193306 626058 193542 626294
rect 192986 590378 193222 590614
rect 193306 590378 193542 590614
rect 192986 590058 193222 590294
rect 193306 590058 193542 590294
rect 192986 554378 193222 554614
rect 193306 554378 193542 554614
rect 192986 554058 193222 554294
rect 193306 554058 193542 554294
rect 192986 518378 193222 518614
rect 193306 518378 193542 518614
rect 192986 518058 193222 518294
rect 193306 518058 193542 518294
rect 192986 482378 193222 482614
rect 193306 482378 193542 482614
rect 192986 482058 193222 482294
rect 193306 482058 193542 482294
rect 192986 446378 193222 446614
rect 193306 446378 193542 446614
rect 192986 446058 193222 446294
rect 193306 446058 193542 446294
rect 192986 410378 193222 410614
rect 193306 410378 193542 410614
rect 192986 410058 193222 410294
rect 193306 410058 193542 410294
rect 192986 374378 193222 374614
rect 193306 374378 193542 374614
rect 192986 374058 193222 374294
rect 193306 374058 193542 374294
rect 192986 338378 193222 338614
rect 193306 338378 193542 338614
rect 192986 338058 193222 338294
rect 193306 338058 193542 338294
rect 192986 302378 193222 302614
rect 193306 302378 193542 302614
rect 192986 302058 193222 302294
rect 193306 302058 193542 302294
rect 192986 266378 193222 266614
rect 193306 266378 193542 266614
rect 192986 266058 193222 266294
rect 193306 266058 193542 266294
rect 192986 230378 193222 230614
rect 193306 230378 193542 230614
rect 192986 230058 193222 230294
rect 193306 230058 193542 230294
rect 199826 705562 200062 705798
rect 200146 705562 200382 705798
rect 199826 705242 200062 705478
rect 200146 705242 200382 705478
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 199826 561218 200062 561454
rect 200146 561218 200382 561454
rect 199826 560898 200062 561134
rect 200146 560898 200382 561134
rect 199826 525218 200062 525454
rect 200146 525218 200382 525454
rect 199826 524898 200062 525134
rect 200146 524898 200382 525134
rect 199826 489218 200062 489454
rect 200146 489218 200382 489454
rect 199826 488898 200062 489134
rect 200146 488898 200382 489134
rect 199826 453218 200062 453454
rect 200146 453218 200382 453454
rect 199826 452898 200062 453134
rect 200146 452898 200382 453134
rect 199826 417218 200062 417454
rect 200146 417218 200382 417454
rect 199826 416898 200062 417134
rect 200146 416898 200382 417134
rect 199826 381218 200062 381454
rect 200146 381218 200382 381454
rect 199826 380898 200062 381134
rect 200146 380898 200382 381134
rect 199826 345218 200062 345454
rect 200146 345218 200382 345454
rect 199826 344898 200062 345134
rect 200146 344898 200382 345134
rect 199826 309218 200062 309454
rect 200146 309218 200382 309454
rect 199826 308898 200062 309134
rect 200146 308898 200382 309134
rect 199826 273218 200062 273454
rect 200146 273218 200382 273454
rect 199826 272898 200062 273134
rect 200146 272898 200382 273134
rect 199826 237218 200062 237454
rect 200146 237218 200382 237454
rect 199826 236898 200062 237134
rect 200146 236898 200382 237134
rect 203546 672938 203782 673174
rect 203866 672938 204102 673174
rect 203546 672618 203782 672854
rect 203866 672618 204102 672854
rect 203546 636938 203782 637174
rect 203866 636938 204102 637174
rect 203546 636618 203782 636854
rect 203866 636618 204102 636854
rect 203546 600938 203782 601174
rect 203866 600938 204102 601174
rect 203546 600618 203782 600854
rect 203866 600618 204102 600854
rect 203546 564938 203782 565174
rect 203866 564938 204102 565174
rect 203546 564618 203782 564854
rect 203866 564618 204102 564854
rect 203546 528938 203782 529174
rect 203866 528938 204102 529174
rect 203546 528618 203782 528854
rect 203866 528618 204102 528854
rect 203546 492938 203782 493174
rect 203866 492938 204102 493174
rect 203546 492618 203782 492854
rect 203866 492618 204102 492854
rect 203546 456938 203782 457174
rect 203866 456938 204102 457174
rect 203546 456618 203782 456854
rect 203866 456618 204102 456854
rect 203546 420938 203782 421174
rect 203866 420938 204102 421174
rect 203546 420618 203782 420854
rect 203866 420618 204102 420854
rect 203546 384938 203782 385174
rect 203866 384938 204102 385174
rect 203546 384618 203782 384854
rect 203866 384618 204102 384854
rect 203546 348938 203782 349174
rect 203866 348938 204102 349174
rect 203546 348618 203782 348854
rect 203866 348618 204102 348854
rect 203546 312938 203782 313174
rect 203866 312938 204102 313174
rect 203546 312618 203782 312854
rect 203866 312618 204102 312854
rect 203546 276938 203782 277174
rect 203866 276938 204102 277174
rect 203546 276618 203782 276854
rect 203866 276618 204102 276854
rect 203546 240938 203782 241174
rect 203866 240938 204102 241174
rect 203546 240618 203782 240854
rect 203866 240618 204102 240854
rect 203546 204938 203782 205174
rect 203866 204938 204102 205174
rect 203546 204618 203782 204854
rect 203866 204618 204102 204854
rect 207266 676658 207502 676894
rect 207586 676658 207822 676894
rect 207266 676338 207502 676574
rect 207586 676338 207822 676574
rect 207266 640658 207502 640894
rect 207586 640658 207822 640894
rect 207266 640338 207502 640574
rect 207586 640338 207822 640574
rect 207266 604658 207502 604894
rect 207586 604658 207822 604894
rect 207266 604338 207502 604574
rect 207586 604338 207822 604574
rect 207266 568658 207502 568894
rect 207586 568658 207822 568894
rect 207266 568338 207502 568574
rect 207586 568338 207822 568574
rect 207266 532658 207502 532894
rect 207586 532658 207822 532894
rect 207266 532338 207502 532574
rect 207586 532338 207822 532574
rect 207266 496658 207502 496894
rect 207586 496658 207822 496894
rect 207266 496338 207502 496574
rect 207586 496338 207822 496574
rect 207266 460658 207502 460894
rect 207586 460658 207822 460894
rect 207266 460338 207502 460574
rect 207586 460338 207822 460574
rect 207266 424658 207502 424894
rect 207586 424658 207822 424894
rect 207266 424338 207502 424574
rect 207586 424338 207822 424574
rect 207266 388658 207502 388894
rect 207586 388658 207822 388894
rect 207266 388338 207502 388574
rect 207586 388338 207822 388574
rect 207266 352658 207502 352894
rect 207586 352658 207822 352894
rect 207266 352338 207502 352574
rect 207586 352338 207822 352574
rect 207266 316658 207502 316894
rect 207586 316658 207822 316894
rect 207266 316338 207502 316574
rect 207586 316338 207822 316574
rect 207266 280658 207502 280894
rect 207586 280658 207822 280894
rect 207266 280338 207502 280574
rect 207586 280338 207822 280574
rect 207266 244658 207502 244894
rect 207586 244658 207822 244894
rect 207266 244338 207502 244574
rect 207586 244338 207822 244574
rect 207266 208658 207502 208894
rect 207586 208658 207822 208894
rect 207266 208338 207502 208574
rect 207586 208338 207822 208574
rect 228986 710362 229222 710598
rect 229306 710362 229542 710598
rect 228986 710042 229222 710278
rect 229306 710042 229542 710278
rect 225266 708442 225502 708678
rect 225586 708442 225822 708678
rect 225266 708122 225502 708358
rect 225586 708122 225822 708358
rect 221546 706522 221782 706758
rect 221866 706522 222102 706758
rect 221546 706202 221782 706438
rect 221866 706202 222102 706438
rect 210986 680378 211222 680614
rect 211306 680378 211542 680614
rect 210986 680058 211222 680294
rect 211306 680058 211542 680294
rect 210986 644378 211222 644614
rect 211306 644378 211542 644614
rect 210986 644058 211222 644294
rect 211306 644058 211542 644294
rect 210986 608378 211222 608614
rect 211306 608378 211542 608614
rect 210986 608058 211222 608294
rect 211306 608058 211542 608294
rect 210986 572378 211222 572614
rect 211306 572378 211542 572614
rect 210986 572058 211222 572294
rect 211306 572058 211542 572294
rect 210986 536378 211222 536614
rect 211306 536378 211542 536614
rect 210986 536058 211222 536294
rect 211306 536058 211542 536294
rect 210986 500378 211222 500614
rect 211306 500378 211542 500614
rect 210986 500058 211222 500294
rect 211306 500058 211542 500294
rect 210986 464378 211222 464614
rect 211306 464378 211542 464614
rect 210986 464058 211222 464294
rect 211306 464058 211542 464294
rect 210986 428378 211222 428614
rect 211306 428378 211542 428614
rect 210986 428058 211222 428294
rect 211306 428058 211542 428294
rect 210986 392378 211222 392614
rect 211306 392378 211542 392614
rect 210986 392058 211222 392294
rect 211306 392058 211542 392294
rect 210986 356378 211222 356614
rect 211306 356378 211542 356614
rect 210986 356058 211222 356294
rect 211306 356058 211542 356294
rect 210986 320378 211222 320614
rect 211306 320378 211542 320614
rect 210986 320058 211222 320294
rect 211306 320058 211542 320294
rect 210986 284378 211222 284614
rect 211306 284378 211542 284614
rect 210986 284058 211222 284294
rect 211306 284058 211542 284294
rect 210986 248378 211222 248614
rect 211306 248378 211542 248614
rect 210986 248058 211222 248294
rect 211306 248058 211542 248294
rect 210986 212378 211222 212614
rect 211306 212378 211542 212614
rect 210986 212058 211222 212294
rect 211306 212058 211542 212294
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 217826 543218 218062 543454
rect 218146 543218 218382 543454
rect 217826 542898 218062 543134
rect 218146 542898 218382 543134
rect 217826 507218 218062 507454
rect 218146 507218 218382 507454
rect 217826 506898 218062 507134
rect 218146 506898 218382 507134
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 217826 435218 218062 435454
rect 218146 435218 218382 435454
rect 217826 434898 218062 435134
rect 218146 434898 218382 435134
rect 217826 399218 218062 399454
rect 218146 399218 218382 399454
rect 217826 398898 218062 399134
rect 218146 398898 218382 399134
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 217826 327218 218062 327454
rect 218146 327218 218382 327454
rect 217826 326898 218062 327134
rect 218146 326898 218382 327134
rect 217826 291218 218062 291454
rect 218146 291218 218382 291454
rect 217826 290898 218062 291134
rect 218146 290898 218382 291134
rect 217826 255218 218062 255454
rect 218146 255218 218382 255454
rect 217826 254898 218062 255134
rect 218146 254898 218382 255134
rect 217826 219218 218062 219454
rect 218146 219218 218382 219454
rect 217826 218898 218062 219134
rect 218146 218898 218382 219134
rect 221546 690938 221782 691174
rect 221866 690938 222102 691174
rect 221546 690618 221782 690854
rect 221866 690618 222102 690854
rect 221546 654938 221782 655174
rect 221866 654938 222102 655174
rect 221546 654618 221782 654854
rect 221866 654618 222102 654854
rect 221546 618938 221782 619174
rect 221866 618938 222102 619174
rect 221546 618618 221782 618854
rect 221866 618618 222102 618854
rect 221546 582938 221782 583174
rect 221866 582938 222102 583174
rect 221546 582618 221782 582854
rect 221866 582618 222102 582854
rect 221546 546938 221782 547174
rect 221866 546938 222102 547174
rect 221546 546618 221782 546854
rect 221866 546618 222102 546854
rect 221546 510938 221782 511174
rect 221866 510938 222102 511174
rect 221546 510618 221782 510854
rect 221866 510618 222102 510854
rect 221546 474938 221782 475174
rect 221866 474938 222102 475174
rect 221546 474618 221782 474854
rect 221866 474618 222102 474854
rect 221546 438938 221782 439174
rect 221866 438938 222102 439174
rect 221546 438618 221782 438854
rect 221866 438618 222102 438854
rect 221546 402938 221782 403174
rect 221866 402938 222102 403174
rect 221546 402618 221782 402854
rect 221866 402618 222102 402854
rect 221546 366938 221782 367174
rect 221866 366938 222102 367174
rect 221546 366618 221782 366854
rect 221866 366618 222102 366854
rect 221546 330938 221782 331174
rect 221866 330938 222102 331174
rect 221546 330618 221782 330854
rect 221866 330618 222102 330854
rect 221546 294938 221782 295174
rect 221866 294938 222102 295174
rect 221546 294618 221782 294854
rect 221866 294618 222102 294854
rect 221546 258938 221782 259174
rect 221866 258938 222102 259174
rect 221546 258618 221782 258854
rect 221866 258618 222102 258854
rect 221546 222938 221782 223174
rect 221866 222938 222102 223174
rect 221546 222618 221782 222854
rect 221866 222618 222102 222854
rect 225266 694658 225502 694894
rect 225586 694658 225822 694894
rect 225266 694338 225502 694574
rect 225586 694338 225822 694574
rect 225266 658658 225502 658894
rect 225586 658658 225822 658894
rect 225266 658338 225502 658574
rect 225586 658338 225822 658574
rect 225266 622658 225502 622894
rect 225586 622658 225822 622894
rect 225266 622338 225502 622574
rect 225586 622338 225822 622574
rect 225266 586658 225502 586894
rect 225586 586658 225822 586894
rect 225266 586338 225502 586574
rect 225586 586338 225822 586574
rect 225266 550658 225502 550894
rect 225586 550658 225822 550894
rect 225266 550338 225502 550574
rect 225586 550338 225822 550574
rect 225266 514658 225502 514894
rect 225586 514658 225822 514894
rect 225266 514338 225502 514574
rect 225586 514338 225822 514574
rect 225266 478658 225502 478894
rect 225586 478658 225822 478894
rect 225266 478338 225502 478574
rect 225586 478338 225822 478574
rect 225266 442658 225502 442894
rect 225586 442658 225822 442894
rect 225266 442338 225502 442574
rect 225586 442338 225822 442574
rect 225266 406658 225502 406894
rect 225586 406658 225822 406894
rect 225266 406338 225502 406574
rect 225586 406338 225822 406574
rect 225266 370658 225502 370894
rect 225586 370658 225822 370894
rect 225266 370338 225502 370574
rect 225586 370338 225822 370574
rect 225266 334658 225502 334894
rect 225586 334658 225822 334894
rect 225266 334338 225502 334574
rect 225586 334338 225822 334574
rect 225266 298658 225502 298894
rect 225586 298658 225822 298894
rect 225266 298338 225502 298574
rect 225586 298338 225822 298574
rect 225266 262658 225502 262894
rect 225586 262658 225822 262894
rect 225266 262338 225502 262574
rect 225586 262338 225822 262574
rect 225266 226658 225502 226894
rect 225586 226658 225822 226894
rect 225266 226338 225502 226574
rect 225586 226338 225822 226574
rect 246986 711322 247222 711558
rect 247306 711322 247542 711558
rect 246986 711002 247222 711238
rect 247306 711002 247542 711238
rect 243266 709402 243502 709638
rect 243586 709402 243822 709638
rect 243266 709082 243502 709318
rect 243586 709082 243822 709318
rect 239546 707482 239782 707718
rect 239866 707482 240102 707718
rect 239546 707162 239782 707398
rect 239866 707162 240102 707398
rect 228986 698378 229222 698614
rect 229306 698378 229542 698614
rect 228986 698058 229222 698294
rect 229306 698058 229542 698294
rect 228986 662378 229222 662614
rect 229306 662378 229542 662614
rect 228986 662058 229222 662294
rect 229306 662058 229542 662294
rect 228986 626378 229222 626614
rect 229306 626378 229542 626614
rect 228986 626058 229222 626294
rect 229306 626058 229542 626294
rect 228986 590378 229222 590614
rect 229306 590378 229542 590614
rect 228986 590058 229222 590294
rect 229306 590058 229542 590294
rect 228986 554378 229222 554614
rect 229306 554378 229542 554614
rect 228986 554058 229222 554294
rect 229306 554058 229542 554294
rect 228986 518378 229222 518614
rect 229306 518378 229542 518614
rect 228986 518058 229222 518294
rect 229306 518058 229542 518294
rect 228986 482378 229222 482614
rect 229306 482378 229542 482614
rect 228986 482058 229222 482294
rect 229306 482058 229542 482294
rect 228986 446378 229222 446614
rect 229306 446378 229542 446614
rect 228986 446058 229222 446294
rect 229306 446058 229542 446294
rect 228986 410378 229222 410614
rect 229306 410378 229542 410614
rect 228986 410058 229222 410294
rect 229306 410058 229542 410294
rect 228986 374378 229222 374614
rect 229306 374378 229542 374614
rect 228986 374058 229222 374294
rect 229306 374058 229542 374294
rect 228986 338378 229222 338614
rect 229306 338378 229542 338614
rect 228986 338058 229222 338294
rect 229306 338058 229542 338294
rect 228986 302378 229222 302614
rect 229306 302378 229542 302614
rect 228986 302058 229222 302294
rect 229306 302058 229542 302294
rect 228986 266378 229222 266614
rect 229306 266378 229542 266614
rect 228986 266058 229222 266294
rect 229306 266058 229542 266294
rect 228986 230378 229222 230614
rect 229306 230378 229542 230614
rect 228986 230058 229222 230294
rect 229306 230058 229542 230294
rect 235826 705562 236062 705798
rect 236146 705562 236382 705798
rect 235826 705242 236062 705478
rect 236146 705242 236382 705478
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 235826 561218 236062 561454
rect 236146 561218 236382 561454
rect 235826 560898 236062 561134
rect 236146 560898 236382 561134
rect 235826 525218 236062 525454
rect 236146 525218 236382 525454
rect 235826 524898 236062 525134
rect 236146 524898 236382 525134
rect 235826 489218 236062 489454
rect 236146 489218 236382 489454
rect 235826 488898 236062 489134
rect 236146 488898 236382 489134
rect 235826 453218 236062 453454
rect 236146 453218 236382 453454
rect 235826 452898 236062 453134
rect 236146 452898 236382 453134
rect 235826 417218 236062 417454
rect 236146 417218 236382 417454
rect 235826 416898 236062 417134
rect 236146 416898 236382 417134
rect 235826 381218 236062 381454
rect 236146 381218 236382 381454
rect 235826 380898 236062 381134
rect 236146 380898 236382 381134
rect 235826 345218 236062 345454
rect 236146 345218 236382 345454
rect 235826 344898 236062 345134
rect 236146 344898 236382 345134
rect 235826 309218 236062 309454
rect 236146 309218 236382 309454
rect 235826 308898 236062 309134
rect 236146 308898 236382 309134
rect 235826 273218 236062 273454
rect 236146 273218 236382 273454
rect 235826 272898 236062 273134
rect 236146 272898 236382 273134
rect 235826 237218 236062 237454
rect 236146 237218 236382 237454
rect 235826 236898 236062 237134
rect 236146 236898 236382 237134
rect 239546 672938 239782 673174
rect 239866 672938 240102 673174
rect 239546 672618 239782 672854
rect 239866 672618 240102 672854
rect 239546 636938 239782 637174
rect 239866 636938 240102 637174
rect 239546 636618 239782 636854
rect 239866 636618 240102 636854
rect 239546 600938 239782 601174
rect 239866 600938 240102 601174
rect 239546 600618 239782 600854
rect 239866 600618 240102 600854
rect 239546 564938 239782 565174
rect 239866 564938 240102 565174
rect 239546 564618 239782 564854
rect 239866 564618 240102 564854
rect 239546 528938 239782 529174
rect 239866 528938 240102 529174
rect 239546 528618 239782 528854
rect 239866 528618 240102 528854
rect 239546 492938 239782 493174
rect 239866 492938 240102 493174
rect 239546 492618 239782 492854
rect 239866 492618 240102 492854
rect 239546 456938 239782 457174
rect 239866 456938 240102 457174
rect 239546 456618 239782 456854
rect 239866 456618 240102 456854
rect 239546 420938 239782 421174
rect 239866 420938 240102 421174
rect 239546 420618 239782 420854
rect 239866 420618 240102 420854
rect 239546 384938 239782 385174
rect 239866 384938 240102 385174
rect 239546 384618 239782 384854
rect 239866 384618 240102 384854
rect 239546 348938 239782 349174
rect 239866 348938 240102 349174
rect 239546 348618 239782 348854
rect 239866 348618 240102 348854
rect 239546 312938 239782 313174
rect 239866 312938 240102 313174
rect 239546 312618 239782 312854
rect 239866 312618 240102 312854
rect 239546 276938 239782 277174
rect 239866 276938 240102 277174
rect 239546 276618 239782 276854
rect 239866 276618 240102 276854
rect 239546 240938 239782 241174
rect 239866 240938 240102 241174
rect 239546 240618 239782 240854
rect 239866 240618 240102 240854
rect 239546 204938 239782 205174
rect 239866 204938 240102 205174
rect 239546 204618 239782 204854
rect 239866 204618 240102 204854
rect 243266 676658 243502 676894
rect 243586 676658 243822 676894
rect 243266 676338 243502 676574
rect 243586 676338 243822 676574
rect 243266 640658 243502 640894
rect 243586 640658 243822 640894
rect 243266 640338 243502 640574
rect 243586 640338 243822 640574
rect 243266 604658 243502 604894
rect 243586 604658 243822 604894
rect 243266 604338 243502 604574
rect 243586 604338 243822 604574
rect 243266 568658 243502 568894
rect 243586 568658 243822 568894
rect 243266 568338 243502 568574
rect 243586 568338 243822 568574
rect 243266 532658 243502 532894
rect 243586 532658 243822 532894
rect 243266 532338 243502 532574
rect 243586 532338 243822 532574
rect 243266 496658 243502 496894
rect 243586 496658 243822 496894
rect 243266 496338 243502 496574
rect 243586 496338 243822 496574
rect 243266 460658 243502 460894
rect 243586 460658 243822 460894
rect 243266 460338 243502 460574
rect 243586 460338 243822 460574
rect 243266 424658 243502 424894
rect 243586 424658 243822 424894
rect 243266 424338 243502 424574
rect 243586 424338 243822 424574
rect 243266 388658 243502 388894
rect 243586 388658 243822 388894
rect 243266 388338 243502 388574
rect 243586 388338 243822 388574
rect 243266 352658 243502 352894
rect 243586 352658 243822 352894
rect 243266 352338 243502 352574
rect 243586 352338 243822 352574
rect 243266 316658 243502 316894
rect 243586 316658 243822 316894
rect 243266 316338 243502 316574
rect 243586 316338 243822 316574
rect 243266 280658 243502 280894
rect 243586 280658 243822 280894
rect 243266 280338 243502 280574
rect 243586 280338 243822 280574
rect 243266 244658 243502 244894
rect 243586 244658 243822 244894
rect 243266 244338 243502 244574
rect 243586 244338 243822 244574
rect 243266 208658 243502 208894
rect 243586 208658 243822 208894
rect 243266 208338 243502 208574
rect 243586 208338 243822 208574
rect 264986 710362 265222 710598
rect 265306 710362 265542 710598
rect 264986 710042 265222 710278
rect 265306 710042 265542 710278
rect 261266 708442 261502 708678
rect 261586 708442 261822 708678
rect 261266 708122 261502 708358
rect 261586 708122 261822 708358
rect 257546 706522 257782 706758
rect 257866 706522 258102 706758
rect 257546 706202 257782 706438
rect 257866 706202 258102 706438
rect 246986 680378 247222 680614
rect 247306 680378 247542 680614
rect 246986 680058 247222 680294
rect 247306 680058 247542 680294
rect 246986 644378 247222 644614
rect 247306 644378 247542 644614
rect 246986 644058 247222 644294
rect 247306 644058 247542 644294
rect 246986 608378 247222 608614
rect 247306 608378 247542 608614
rect 246986 608058 247222 608294
rect 247306 608058 247542 608294
rect 246986 572378 247222 572614
rect 247306 572378 247542 572614
rect 246986 572058 247222 572294
rect 247306 572058 247542 572294
rect 246986 536378 247222 536614
rect 247306 536378 247542 536614
rect 246986 536058 247222 536294
rect 247306 536058 247542 536294
rect 246986 500378 247222 500614
rect 247306 500378 247542 500614
rect 246986 500058 247222 500294
rect 247306 500058 247542 500294
rect 246986 464378 247222 464614
rect 247306 464378 247542 464614
rect 246986 464058 247222 464294
rect 247306 464058 247542 464294
rect 246986 428378 247222 428614
rect 247306 428378 247542 428614
rect 246986 428058 247222 428294
rect 247306 428058 247542 428294
rect 246986 392378 247222 392614
rect 247306 392378 247542 392614
rect 246986 392058 247222 392294
rect 247306 392058 247542 392294
rect 246986 356378 247222 356614
rect 247306 356378 247542 356614
rect 246986 356058 247222 356294
rect 247306 356058 247542 356294
rect 246986 320378 247222 320614
rect 247306 320378 247542 320614
rect 246986 320058 247222 320294
rect 247306 320058 247542 320294
rect 246986 284378 247222 284614
rect 247306 284378 247542 284614
rect 246986 284058 247222 284294
rect 247306 284058 247542 284294
rect 246986 248378 247222 248614
rect 247306 248378 247542 248614
rect 246986 248058 247222 248294
rect 247306 248058 247542 248294
rect 246986 212378 247222 212614
rect 247306 212378 247542 212614
rect 246986 212058 247222 212294
rect 247306 212058 247542 212294
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 253826 543218 254062 543454
rect 254146 543218 254382 543454
rect 253826 542898 254062 543134
rect 254146 542898 254382 543134
rect 253826 507218 254062 507454
rect 254146 507218 254382 507454
rect 253826 506898 254062 507134
rect 254146 506898 254382 507134
rect 253826 471218 254062 471454
rect 254146 471218 254382 471454
rect 253826 470898 254062 471134
rect 254146 470898 254382 471134
rect 253826 435218 254062 435454
rect 254146 435218 254382 435454
rect 253826 434898 254062 435134
rect 254146 434898 254382 435134
rect 253826 399218 254062 399454
rect 254146 399218 254382 399454
rect 253826 398898 254062 399134
rect 254146 398898 254382 399134
rect 253826 363218 254062 363454
rect 254146 363218 254382 363454
rect 253826 362898 254062 363134
rect 254146 362898 254382 363134
rect 253826 327218 254062 327454
rect 254146 327218 254382 327454
rect 253826 326898 254062 327134
rect 254146 326898 254382 327134
rect 253826 291218 254062 291454
rect 254146 291218 254382 291454
rect 253826 290898 254062 291134
rect 254146 290898 254382 291134
rect 253826 255218 254062 255454
rect 254146 255218 254382 255454
rect 253826 254898 254062 255134
rect 254146 254898 254382 255134
rect 253826 219218 254062 219454
rect 254146 219218 254382 219454
rect 253826 218898 254062 219134
rect 254146 218898 254382 219134
rect 257546 690938 257782 691174
rect 257866 690938 258102 691174
rect 257546 690618 257782 690854
rect 257866 690618 258102 690854
rect 257546 654938 257782 655174
rect 257866 654938 258102 655174
rect 257546 654618 257782 654854
rect 257866 654618 258102 654854
rect 257546 618938 257782 619174
rect 257866 618938 258102 619174
rect 257546 618618 257782 618854
rect 257866 618618 258102 618854
rect 257546 582938 257782 583174
rect 257866 582938 258102 583174
rect 257546 582618 257782 582854
rect 257866 582618 258102 582854
rect 257546 546938 257782 547174
rect 257866 546938 258102 547174
rect 257546 546618 257782 546854
rect 257866 546618 258102 546854
rect 257546 510938 257782 511174
rect 257866 510938 258102 511174
rect 257546 510618 257782 510854
rect 257866 510618 258102 510854
rect 257546 474938 257782 475174
rect 257866 474938 258102 475174
rect 257546 474618 257782 474854
rect 257866 474618 258102 474854
rect 257546 438938 257782 439174
rect 257866 438938 258102 439174
rect 257546 438618 257782 438854
rect 257866 438618 258102 438854
rect 257546 402938 257782 403174
rect 257866 402938 258102 403174
rect 257546 402618 257782 402854
rect 257866 402618 258102 402854
rect 257546 366938 257782 367174
rect 257866 366938 258102 367174
rect 257546 366618 257782 366854
rect 257866 366618 258102 366854
rect 257546 330938 257782 331174
rect 257866 330938 258102 331174
rect 257546 330618 257782 330854
rect 257866 330618 258102 330854
rect 257546 294938 257782 295174
rect 257866 294938 258102 295174
rect 257546 294618 257782 294854
rect 257866 294618 258102 294854
rect 257546 258938 257782 259174
rect 257866 258938 258102 259174
rect 257546 258618 257782 258854
rect 257866 258618 258102 258854
rect 257546 222938 257782 223174
rect 257866 222938 258102 223174
rect 257546 222618 257782 222854
rect 257866 222618 258102 222854
rect 261266 694658 261502 694894
rect 261586 694658 261822 694894
rect 261266 694338 261502 694574
rect 261586 694338 261822 694574
rect 261266 658658 261502 658894
rect 261586 658658 261822 658894
rect 261266 658338 261502 658574
rect 261586 658338 261822 658574
rect 261266 622658 261502 622894
rect 261586 622658 261822 622894
rect 261266 622338 261502 622574
rect 261586 622338 261822 622574
rect 261266 586658 261502 586894
rect 261586 586658 261822 586894
rect 261266 586338 261502 586574
rect 261586 586338 261822 586574
rect 261266 550658 261502 550894
rect 261586 550658 261822 550894
rect 261266 550338 261502 550574
rect 261586 550338 261822 550574
rect 261266 514658 261502 514894
rect 261586 514658 261822 514894
rect 261266 514338 261502 514574
rect 261586 514338 261822 514574
rect 261266 478658 261502 478894
rect 261586 478658 261822 478894
rect 261266 478338 261502 478574
rect 261586 478338 261822 478574
rect 261266 442658 261502 442894
rect 261586 442658 261822 442894
rect 261266 442338 261502 442574
rect 261586 442338 261822 442574
rect 261266 406658 261502 406894
rect 261586 406658 261822 406894
rect 261266 406338 261502 406574
rect 261586 406338 261822 406574
rect 261266 370658 261502 370894
rect 261586 370658 261822 370894
rect 261266 370338 261502 370574
rect 261586 370338 261822 370574
rect 261266 334658 261502 334894
rect 261586 334658 261822 334894
rect 261266 334338 261502 334574
rect 261586 334338 261822 334574
rect 261266 298658 261502 298894
rect 261586 298658 261822 298894
rect 261266 298338 261502 298574
rect 261586 298338 261822 298574
rect 261266 262658 261502 262894
rect 261586 262658 261822 262894
rect 261266 262338 261502 262574
rect 261586 262338 261822 262574
rect 261266 226658 261502 226894
rect 261586 226658 261822 226894
rect 261266 226338 261502 226574
rect 261586 226338 261822 226574
rect 282986 711322 283222 711558
rect 283306 711322 283542 711558
rect 282986 711002 283222 711238
rect 283306 711002 283542 711238
rect 279266 709402 279502 709638
rect 279586 709402 279822 709638
rect 279266 709082 279502 709318
rect 279586 709082 279822 709318
rect 275546 707482 275782 707718
rect 275866 707482 276102 707718
rect 275546 707162 275782 707398
rect 275866 707162 276102 707398
rect 264986 698378 265222 698614
rect 265306 698378 265542 698614
rect 264986 698058 265222 698294
rect 265306 698058 265542 698294
rect 264986 662378 265222 662614
rect 265306 662378 265542 662614
rect 264986 662058 265222 662294
rect 265306 662058 265542 662294
rect 264986 626378 265222 626614
rect 265306 626378 265542 626614
rect 264986 626058 265222 626294
rect 265306 626058 265542 626294
rect 264986 590378 265222 590614
rect 265306 590378 265542 590614
rect 264986 590058 265222 590294
rect 265306 590058 265542 590294
rect 264986 554378 265222 554614
rect 265306 554378 265542 554614
rect 264986 554058 265222 554294
rect 265306 554058 265542 554294
rect 264986 518378 265222 518614
rect 265306 518378 265542 518614
rect 264986 518058 265222 518294
rect 265306 518058 265542 518294
rect 264986 482378 265222 482614
rect 265306 482378 265542 482614
rect 264986 482058 265222 482294
rect 265306 482058 265542 482294
rect 264986 446378 265222 446614
rect 265306 446378 265542 446614
rect 264986 446058 265222 446294
rect 265306 446058 265542 446294
rect 264986 410378 265222 410614
rect 265306 410378 265542 410614
rect 264986 410058 265222 410294
rect 265306 410058 265542 410294
rect 264986 374378 265222 374614
rect 265306 374378 265542 374614
rect 264986 374058 265222 374294
rect 265306 374058 265542 374294
rect 264986 338378 265222 338614
rect 265306 338378 265542 338614
rect 264986 338058 265222 338294
rect 265306 338058 265542 338294
rect 264986 302378 265222 302614
rect 265306 302378 265542 302614
rect 264986 302058 265222 302294
rect 265306 302058 265542 302294
rect 264986 266378 265222 266614
rect 265306 266378 265542 266614
rect 264986 266058 265222 266294
rect 265306 266058 265542 266294
rect 264986 230378 265222 230614
rect 265306 230378 265542 230614
rect 264986 230058 265222 230294
rect 265306 230058 265542 230294
rect 271826 705562 272062 705798
rect 272146 705562 272382 705798
rect 271826 705242 272062 705478
rect 272146 705242 272382 705478
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 271826 561218 272062 561454
rect 272146 561218 272382 561454
rect 271826 560898 272062 561134
rect 272146 560898 272382 561134
rect 271826 525218 272062 525454
rect 272146 525218 272382 525454
rect 271826 524898 272062 525134
rect 272146 524898 272382 525134
rect 271826 489218 272062 489454
rect 272146 489218 272382 489454
rect 271826 488898 272062 489134
rect 272146 488898 272382 489134
rect 271826 453218 272062 453454
rect 272146 453218 272382 453454
rect 271826 452898 272062 453134
rect 272146 452898 272382 453134
rect 271826 417218 272062 417454
rect 272146 417218 272382 417454
rect 271826 416898 272062 417134
rect 272146 416898 272382 417134
rect 271826 381218 272062 381454
rect 272146 381218 272382 381454
rect 271826 380898 272062 381134
rect 272146 380898 272382 381134
rect 271826 345218 272062 345454
rect 272146 345218 272382 345454
rect 271826 344898 272062 345134
rect 272146 344898 272382 345134
rect 271826 309218 272062 309454
rect 272146 309218 272382 309454
rect 271826 308898 272062 309134
rect 272146 308898 272382 309134
rect 271826 273218 272062 273454
rect 272146 273218 272382 273454
rect 271826 272898 272062 273134
rect 272146 272898 272382 273134
rect 271826 237218 272062 237454
rect 272146 237218 272382 237454
rect 271826 236898 272062 237134
rect 272146 236898 272382 237134
rect 275546 672938 275782 673174
rect 275866 672938 276102 673174
rect 275546 672618 275782 672854
rect 275866 672618 276102 672854
rect 275546 636938 275782 637174
rect 275866 636938 276102 637174
rect 275546 636618 275782 636854
rect 275866 636618 276102 636854
rect 275546 600938 275782 601174
rect 275866 600938 276102 601174
rect 275546 600618 275782 600854
rect 275866 600618 276102 600854
rect 275546 564938 275782 565174
rect 275866 564938 276102 565174
rect 275546 564618 275782 564854
rect 275866 564618 276102 564854
rect 275546 528938 275782 529174
rect 275866 528938 276102 529174
rect 275546 528618 275782 528854
rect 275866 528618 276102 528854
rect 275546 492938 275782 493174
rect 275866 492938 276102 493174
rect 275546 492618 275782 492854
rect 275866 492618 276102 492854
rect 275546 456938 275782 457174
rect 275866 456938 276102 457174
rect 275546 456618 275782 456854
rect 275866 456618 276102 456854
rect 275546 420938 275782 421174
rect 275866 420938 276102 421174
rect 275546 420618 275782 420854
rect 275866 420618 276102 420854
rect 275546 384938 275782 385174
rect 275866 384938 276102 385174
rect 275546 384618 275782 384854
rect 275866 384618 276102 384854
rect 275546 348938 275782 349174
rect 275866 348938 276102 349174
rect 275546 348618 275782 348854
rect 275866 348618 276102 348854
rect 275546 312938 275782 313174
rect 275866 312938 276102 313174
rect 275546 312618 275782 312854
rect 275866 312618 276102 312854
rect 275546 276938 275782 277174
rect 275866 276938 276102 277174
rect 275546 276618 275782 276854
rect 275866 276618 276102 276854
rect 275546 240938 275782 241174
rect 275866 240938 276102 241174
rect 275546 240618 275782 240854
rect 275866 240618 276102 240854
rect 275546 204938 275782 205174
rect 275866 204938 276102 205174
rect 275546 204618 275782 204854
rect 275866 204618 276102 204854
rect 279266 676658 279502 676894
rect 279586 676658 279822 676894
rect 279266 676338 279502 676574
rect 279586 676338 279822 676574
rect 279266 640658 279502 640894
rect 279586 640658 279822 640894
rect 279266 640338 279502 640574
rect 279586 640338 279822 640574
rect 279266 604658 279502 604894
rect 279586 604658 279822 604894
rect 279266 604338 279502 604574
rect 279586 604338 279822 604574
rect 279266 568658 279502 568894
rect 279586 568658 279822 568894
rect 279266 568338 279502 568574
rect 279586 568338 279822 568574
rect 279266 532658 279502 532894
rect 279586 532658 279822 532894
rect 279266 532338 279502 532574
rect 279586 532338 279822 532574
rect 279266 496658 279502 496894
rect 279586 496658 279822 496894
rect 279266 496338 279502 496574
rect 279586 496338 279822 496574
rect 279266 460658 279502 460894
rect 279586 460658 279822 460894
rect 279266 460338 279502 460574
rect 279586 460338 279822 460574
rect 279266 424658 279502 424894
rect 279586 424658 279822 424894
rect 279266 424338 279502 424574
rect 279586 424338 279822 424574
rect 279266 388658 279502 388894
rect 279586 388658 279822 388894
rect 279266 388338 279502 388574
rect 279586 388338 279822 388574
rect 279266 352658 279502 352894
rect 279586 352658 279822 352894
rect 279266 352338 279502 352574
rect 279586 352338 279822 352574
rect 279266 316658 279502 316894
rect 279586 316658 279822 316894
rect 279266 316338 279502 316574
rect 279586 316338 279822 316574
rect 279266 280658 279502 280894
rect 279586 280658 279822 280894
rect 279266 280338 279502 280574
rect 279586 280338 279822 280574
rect 279266 244658 279502 244894
rect 279586 244658 279822 244894
rect 279266 244338 279502 244574
rect 279586 244338 279822 244574
rect 279266 208658 279502 208894
rect 279586 208658 279822 208894
rect 279266 208338 279502 208574
rect 279586 208338 279822 208574
rect 300986 710362 301222 710598
rect 301306 710362 301542 710598
rect 300986 710042 301222 710278
rect 301306 710042 301542 710278
rect 297266 708442 297502 708678
rect 297586 708442 297822 708678
rect 297266 708122 297502 708358
rect 297586 708122 297822 708358
rect 293546 706522 293782 706758
rect 293866 706522 294102 706758
rect 293546 706202 293782 706438
rect 293866 706202 294102 706438
rect 282986 680378 283222 680614
rect 283306 680378 283542 680614
rect 282986 680058 283222 680294
rect 283306 680058 283542 680294
rect 282986 644378 283222 644614
rect 283306 644378 283542 644614
rect 282986 644058 283222 644294
rect 283306 644058 283542 644294
rect 282986 608378 283222 608614
rect 283306 608378 283542 608614
rect 282986 608058 283222 608294
rect 283306 608058 283542 608294
rect 282986 572378 283222 572614
rect 283306 572378 283542 572614
rect 282986 572058 283222 572294
rect 283306 572058 283542 572294
rect 282986 536378 283222 536614
rect 283306 536378 283542 536614
rect 282986 536058 283222 536294
rect 283306 536058 283542 536294
rect 282986 500378 283222 500614
rect 283306 500378 283542 500614
rect 282986 500058 283222 500294
rect 283306 500058 283542 500294
rect 282986 464378 283222 464614
rect 283306 464378 283542 464614
rect 282986 464058 283222 464294
rect 283306 464058 283542 464294
rect 282986 428378 283222 428614
rect 283306 428378 283542 428614
rect 282986 428058 283222 428294
rect 283306 428058 283542 428294
rect 282986 392378 283222 392614
rect 283306 392378 283542 392614
rect 282986 392058 283222 392294
rect 283306 392058 283542 392294
rect 282986 356378 283222 356614
rect 283306 356378 283542 356614
rect 282986 356058 283222 356294
rect 283306 356058 283542 356294
rect 282986 320378 283222 320614
rect 283306 320378 283542 320614
rect 282986 320058 283222 320294
rect 283306 320058 283542 320294
rect 282986 284378 283222 284614
rect 283306 284378 283542 284614
rect 282986 284058 283222 284294
rect 283306 284058 283542 284294
rect 282986 248378 283222 248614
rect 283306 248378 283542 248614
rect 282986 248058 283222 248294
rect 283306 248058 283542 248294
rect 282986 212378 283222 212614
rect 283306 212378 283542 212614
rect 282986 212058 283222 212294
rect 283306 212058 283542 212294
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 289826 507218 290062 507454
rect 290146 507218 290382 507454
rect 289826 506898 290062 507134
rect 290146 506898 290382 507134
rect 289826 471218 290062 471454
rect 290146 471218 290382 471454
rect 289826 470898 290062 471134
rect 290146 470898 290382 471134
rect 289826 435218 290062 435454
rect 290146 435218 290382 435454
rect 289826 434898 290062 435134
rect 290146 434898 290382 435134
rect 289826 399218 290062 399454
rect 290146 399218 290382 399454
rect 289826 398898 290062 399134
rect 290146 398898 290382 399134
rect 289826 363218 290062 363454
rect 290146 363218 290382 363454
rect 289826 362898 290062 363134
rect 290146 362898 290382 363134
rect 289826 327218 290062 327454
rect 290146 327218 290382 327454
rect 289826 326898 290062 327134
rect 290146 326898 290382 327134
rect 289826 291218 290062 291454
rect 290146 291218 290382 291454
rect 289826 290898 290062 291134
rect 290146 290898 290382 291134
rect 289826 255218 290062 255454
rect 290146 255218 290382 255454
rect 289826 254898 290062 255134
rect 290146 254898 290382 255134
rect 289826 219218 290062 219454
rect 290146 219218 290382 219454
rect 289826 218898 290062 219134
rect 290146 218898 290382 219134
rect 293546 690938 293782 691174
rect 293866 690938 294102 691174
rect 293546 690618 293782 690854
rect 293866 690618 294102 690854
rect 293546 654938 293782 655174
rect 293866 654938 294102 655174
rect 293546 654618 293782 654854
rect 293866 654618 294102 654854
rect 293546 618938 293782 619174
rect 293866 618938 294102 619174
rect 293546 618618 293782 618854
rect 293866 618618 294102 618854
rect 293546 582938 293782 583174
rect 293866 582938 294102 583174
rect 293546 582618 293782 582854
rect 293866 582618 294102 582854
rect 293546 546938 293782 547174
rect 293866 546938 294102 547174
rect 293546 546618 293782 546854
rect 293866 546618 294102 546854
rect 293546 510938 293782 511174
rect 293866 510938 294102 511174
rect 293546 510618 293782 510854
rect 293866 510618 294102 510854
rect 293546 474938 293782 475174
rect 293866 474938 294102 475174
rect 293546 474618 293782 474854
rect 293866 474618 294102 474854
rect 293546 438938 293782 439174
rect 293866 438938 294102 439174
rect 293546 438618 293782 438854
rect 293866 438618 294102 438854
rect 293546 402938 293782 403174
rect 293866 402938 294102 403174
rect 293546 402618 293782 402854
rect 293866 402618 294102 402854
rect 293546 366938 293782 367174
rect 293866 366938 294102 367174
rect 293546 366618 293782 366854
rect 293866 366618 294102 366854
rect 293546 330938 293782 331174
rect 293866 330938 294102 331174
rect 293546 330618 293782 330854
rect 293866 330618 294102 330854
rect 293546 294938 293782 295174
rect 293866 294938 294102 295174
rect 293546 294618 293782 294854
rect 293866 294618 294102 294854
rect 293546 258938 293782 259174
rect 293866 258938 294102 259174
rect 293546 258618 293782 258854
rect 293866 258618 294102 258854
rect 293546 222938 293782 223174
rect 293866 222938 294102 223174
rect 293546 222618 293782 222854
rect 293866 222618 294102 222854
rect 297266 694658 297502 694894
rect 297586 694658 297822 694894
rect 297266 694338 297502 694574
rect 297586 694338 297822 694574
rect 297266 658658 297502 658894
rect 297586 658658 297822 658894
rect 297266 658338 297502 658574
rect 297586 658338 297822 658574
rect 297266 622658 297502 622894
rect 297586 622658 297822 622894
rect 297266 622338 297502 622574
rect 297586 622338 297822 622574
rect 297266 586658 297502 586894
rect 297586 586658 297822 586894
rect 297266 586338 297502 586574
rect 297586 586338 297822 586574
rect 297266 550658 297502 550894
rect 297586 550658 297822 550894
rect 297266 550338 297502 550574
rect 297586 550338 297822 550574
rect 297266 514658 297502 514894
rect 297586 514658 297822 514894
rect 297266 514338 297502 514574
rect 297586 514338 297822 514574
rect 297266 478658 297502 478894
rect 297586 478658 297822 478894
rect 297266 478338 297502 478574
rect 297586 478338 297822 478574
rect 297266 442658 297502 442894
rect 297586 442658 297822 442894
rect 297266 442338 297502 442574
rect 297586 442338 297822 442574
rect 297266 406658 297502 406894
rect 297586 406658 297822 406894
rect 297266 406338 297502 406574
rect 297586 406338 297822 406574
rect 297266 370658 297502 370894
rect 297586 370658 297822 370894
rect 297266 370338 297502 370574
rect 297586 370338 297822 370574
rect 297266 334658 297502 334894
rect 297586 334658 297822 334894
rect 297266 334338 297502 334574
rect 297586 334338 297822 334574
rect 297266 298658 297502 298894
rect 297586 298658 297822 298894
rect 297266 298338 297502 298574
rect 297586 298338 297822 298574
rect 297266 262658 297502 262894
rect 297586 262658 297822 262894
rect 297266 262338 297502 262574
rect 297586 262338 297822 262574
rect 297266 226658 297502 226894
rect 297586 226658 297822 226894
rect 297266 226338 297502 226574
rect 297586 226338 297822 226574
rect 318986 711322 319222 711558
rect 319306 711322 319542 711558
rect 318986 711002 319222 711238
rect 319306 711002 319542 711238
rect 315266 709402 315502 709638
rect 315586 709402 315822 709638
rect 315266 709082 315502 709318
rect 315586 709082 315822 709318
rect 311546 707482 311782 707718
rect 311866 707482 312102 707718
rect 311546 707162 311782 707398
rect 311866 707162 312102 707398
rect 300986 698378 301222 698614
rect 301306 698378 301542 698614
rect 300986 698058 301222 698294
rect 301306 698058 301542 698294
rect 300986 662378 301222 662614
rect 301306 662378 301542 662614
rect 300986 662058 301222 662294
rect 301306 662058 301542 662294
rect 300986 626378 301222 626614
rect 301306 626378 301542 626614
rect 300986 626058 301222 626294
rect 301306 626058 301542 626294
rect 300986 590378 301222 590614
rect 301306 590378 301542 590614
rect 300986 590058 301222 590294
rect 301306 590058 301542 590294
rect 300986 554378 301222 554614
rect 301306 554378 301542 554614
rect 300986 554058 301222 554294
rect 301306 554058 301542 554294
rect 300986 518378 301222 518614
rect 301306 518378 301542 518614
rect 300986 518058 301222 518294
rect 301306 518058 301542 518294
rect 300986 482378 301222 482614
rect 301306 482378 301542 482614
rect 300986 482058 301222 482294
rect 301306 482058 301542 482294
rect 300986 446378 301222 446614
rect 301306 446378 301542 446614
rect 300986 446058 301222 446294
rect 301306 446058 301542 446294
rect 300986 410378 301222 410614
rect 301306 410378 301542 410614
rect 300986 410058 301222 410294
rect 301306 410058 301542 410294
rect 300986 374378 301222 374614
rect 301306 374378 301542 374614
rect 300986 374058 301222 374294
rect 301306 374058 301542 374294
rect 300986 338378 301222 338614
rect 301306 338378 301542 338614
rect 300986 338058 301222 338294
rect 301306 338058 301542 338294
rect 300986 302378 301222 302614
rect 301306 302378 301542 302614
rect 300986 302058 301222 302294
rect 301306 302058 301542 302294
rect 300986 266378 301222 266614
rect 301306 266378 301542 266614
rect 300986 266058 301222 266294
rect 301306 266058 301542 266294
rect 300986 230378 301222 230614
rect 301306 230378 301542 230614
rect 300986 230058 301222 230294
rect 301306 230058 301542 230294
rect 307826 705562 308062 705798
rect 308146 705562 308382 705798
rect 307826 705242 308062 705478
rect 308146 705242 308382 705478
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 307826 561218 308062 561454
rect 308146 561218 308382 561454
rect 307826 560898 308062 561134
rect 308146 560898 308382 561134
rect 307826 525218 308062 525454
rect 308146 525218 308382 525454
rect 307826 524898 308062 525134
rect 308146 524898 308382 525134
rect 307826 489218 308062 489454
rect 308146 489218 308382 489454
rect 307826 488898 308062 489134
rect 308146 488898 308382 489134
rect 307826 453218 308062 453454
rect 308146 453218 308382 453454
rect 307826 452898 308062 453134
rect 308146 452898 308382 453134
rect 307826 417218 308062 417454
rect 308146 417218 308382 417454
rect 307826 416898 308062 417134
rect 308146 416898 308382 417134
rect 307826 381218 308062 381454
rect 308146 381218 308382 381454
rect 307826 380898 308062 381134
rect 308146 380898 308382 381134
rect 307826 345218 308062 345454
rect 308146 345218 308382 345454
rect 307826 344898 308062 345134
rect 308146 344898 308382 345134
rect 307826 309218 308062 309454
rect 308146 309218 308382 309454
rect 307826 308898 308062 309134
rect 308146 308898 308382 309134
rect 307826 273218 308062 273454
rect 308146 273218 308382 273454
rect 307826 272898 308062 273134
rect 308146 272898 308382 273134
rect 307826 237218 308062 237454
rect 308146 237218 308382 237454
rect 307826 236898 308062 237134
rect 308146 236898 308382 237134
rect 192986 194378 193222 194614
rect 193306 194378 193542 194614
rect 192986 194058 193222 194294
rect 193306 194058 193542 194294
rect 307826 201218 308062 201454
rect 308146 201218 308382 201454
rect 307826 200898 308062 201134
rect 308146 200898 308382 201134
rect 204250 183218 204486 183454
rect 204250 182898 204486 183134
rect 234970 183218 235206 183454
rect 234970 182898 235206 183134
rect 265690 183218 265926 183454
rect 265690 182898 265926 183134
rect 296410 183218 296646 183454
rect 296410 182898 296646 183134
rect 219610 165218 219846 165454
rect 219610 164898 219846 165134
rect 250330 165218 250566 165454
rect 250330 164898 250566 165134
rect 281050 165218 281286 165454
rect 281050 164898 281286 165134
rect 307826 165218 308062 165454
rect 308146 165218 308382 165454
rect 307826 164898 308062 165134
rect 308146 164898 308382 165134
rect 192986 158378 193222 158614
rect 193306 158378 193542 158614
rect 192986 158058 193222 158294
rect 193306 158058 193542 158294
rect 204250 147218 204486 147454
rect 204250 146898 204486 147134
rect 234970 147218 235206 147454
rect 234970 146898 235206 147134
rect 265690 147218 265926 147454
rect 265690 146898 265926 147134
rect 296410 147218 296646 147454
rect 296410 146898 296646 147134
rect 219610 129218 219846 129454
rect 219610 128898 219846 129134
rect 250330 129218 250566 129454
rect 250330 128898 250566 129134
rect 281050 129218 281286 129454
rect 281050 128898 281286 129134
rect 307826 129218 308062 129454
rect 308146 129218 308382 129454
rect 307826 128898 308062 129134
rect 308146 128898 308382 129134
rect 192986 122378 193222 122614
rect 193306 122378 193542 122614
rect 192986 122058 193222 122294
rect 193306 122058 193542 122294
rect 204250 111218 204486 111454
rect 204250 110898 204486 111134
rect 234970 111218 235206 111454
rect 234970 110898 235206 111134
rect 265690 111218 265926 111454
rect 265690 110898 265926 111134
rect 296410 111218 296646 111454
rect 296410 110898 296646 111134
rect 192986 86378 193222 86614
rect 193306 86378 193542 86614
rect 192986 86058 193222 86294
rect 193306 86058 193542 86294
rect 192986 50378 193222 50614
rect 193306 50378 193542 50614
rect 192986 50058 193222 50294
rect 193306 50058 193542 50294
rect 192986 14378 193222 14614
rect 193306 14378 193542 14614
rect 192986 14058 193222 14294
rect 193306 14058 193542 14294
rect 174986 -7302 175222 -7066
rect 175306 -7302 175542 -7066
rect 174986 -7622 175222 -7386
rect 175306 -7622 175542 -7386
rect 203546 96938 203782 97174
rect 203866 96938 204102 97174
rect 199826 93218 200062 93454
rect 200146 93218 200382 93454
rect 199826 92898 200062 93134
rect 200146 92898 200382 93134
rect 203546 96618 203782 96854
rect 203866 96618 204102 96854
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -1542 200062 -1306
rect 200146 -1542 200382 -1306
rect 199826 -1862 200062 -1626
rect 200146 -1862 200382 -1626
rect 203546 60938 203782 61174
rect 203866 60938 204102 61174
rect 203546 60618 203782 60854
rect 203866 60618 204102 60854
rect 203546 24938 203782 25174
rect 203866 24938 204102 25174
rect 203546 24618 203782 24854
rect 203866 24618 204102 24854
rect 203546 -3462 203782 -3226
rect 203866 -3462 204102 -3226
rect 203546 -3782 203782 -3546
rect 203866 -3782 204102 -3546
rect 207266 64658 207502 64894
rect 207586 64658 207822 64894
rect 207266 64338 207502 64574
rect 207586 64338 207822 64574
rect 207266 28658 207502 28894
rect 207586 28658 207822 28894
rect 207266 28338 207502 28574
rect 207586 28338 207822 28574
rect 207266 -5382 207502 -5146
rect 207586 -5382 207822 -5146
rect 207266 -5702 207502 -5466
rect 207586 -5702 207822 -5466
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 210986 68378 211222 68614
rect 211306 68378 211542 68614
rect 210986 68058 211222 68294
rect 211306 68058 211542 68294
rect 210986 32378 211222 32614
rect 211306 32378 211542 32614
rect 210986 32058 211222 32294
rect 211306 32058 211542 32294
rect 192986 -6342 193222 -6106
rect 193306 -6342 193542 -6106
rect 192986 -6662 193222 -6426
rect 193306 -6662 193542 -6426
rect 221546 78938 221782 79174
rect 221866 78938 222102 79174
rect 221546 78618 221782 78854
rect 221866 78618 222102 78854
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 221546 42938 221782 43174
rect 221866 42938 222102 43174
rect 221546 42618 221782 42854
rect 221866 42618 222102 42854
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 221546 -2502 221782 -2266
rect 221866 -2502 222102 -2266
rect 221546 -2822 221782 -2586
rect 221866 -2822 222102 -2586
rect 225266 82658 225502 82894
rect 225586 82658 225822 82894
rect 225266 82338 225502 82574
rect 225586 82338 225822 82574
rect 225266 46658 225502 46894
rect 225586 46658 225822 46894
rect 225266 46338 225502 46574
rect 225586 46338 225822 46574
rect 225266 10658 225502 10894
rect 225586 10658 225822 10894
rect 225266 10338 225502 10574
rect 225586 10338 225822 10574
rect 225266 -4422 225502 -4186
rect 225586 -4422 225822 -4186
rect 225266 -4742 225502 -4506
rect 225586 -4742 225822 -4506
rect 228986 86378 229222 86614
rect 229306 86378 229542 86614
rect 228986 86058 229222 86294
rect 229306 86058 229542 86294
rect 239546 96938 239782 97174
rect 239866 96938 240102 97174
rect 235826 93218 236062 93454
rect 236146 93218 236382 93454
rect 235826 92898 236062 93134
rect 236146 92898 236382 93134
rect 228986 50378 229222 50614
rect 229306 50378 229542 50614
rect 228986 50058 229222 50294
rect 229306 50058 229542 50294
rect 228986 14378 229222 14614
rect 229306 14378 229542 14614
rect 228986 14058 229222 14294
rect 229306 14058 229542 14294
rect 210986 -7302 211222 -7066
rect 211306 -7302 211542 -7066
rect 210986 -7622 211222 -7386
rect 211306 -7622 211542 -7386
rect 239546 96618 239782 96854
rect 239866 96618 240102 96854
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -1542 236062 -1306
rect 236146 -1542 236382 -1306
rect 235826 -1862 236062 -1626
rect 236146 -1862 236382 -1626
rect 239546 60938 239782 61174
rect 239866 60938 240102 61174
rect 239546 60618 239782 60854
rect 239866 60618 240102 60854
rect 239546 24938 239782 25174
rect 239866 24938 240102 25174
rect 239546 24618 239782 24854
rect 239866 24618 240102 24854
rect 239546 -3462 239782 -3226
rect 239866 -3462 240102 -3226
rect 239546 -3782 239782 -3546
rect 239866 -3782 240102 -3546
rect 243266 64658 243502 64894
rect 243586 64658 243822 64894
rect 243266 64338 243502 64574
rect 243586 64338 243822 64574
rect 243266 28658 243502 28894
rect 243586 28658 243822 28894
rect 243266 28338 243502 28574
rect 243586 28338 243822 28574
rect 246986 68378 247222 68614
rect 247306 68378 247542 68614
rect 246986 68058 247222 68294
rect 247306 68058 247542 68294
rect 246986 32378 247222 32614
rect 247306 32378 247542 32614
rect 246986 32058 247222 32294
rect 247306 32058 247542 32294
rect 243266 -5382 243502 -5146
rect 243586 -5382 243822 -5146
rect 243266 -5702 243502 -5466
rect 243586 -5702 243822 -5466
rect 228986 -6342 229222 -6106
rect 229306 -6342 229542 -6106
rect 228986 -6662 229222 -6426
rect 229306 -6662 229542 -6426
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 257546 78938 257782 79174
rect 257866 78938 258102 79174
rect 257546 78618 257782 78854
rect 257866 78618 258102 78854
rect 261266 82658 261502 82894
rect 261586 82658 261822 82894
rect 261266 82338 261502 82574
rect 261586 82338 261822 82574
rect 257546 42938 257782 43174
rect 257866 42938 258102 43174
rect 257546 42618 257782 42854
rect 257866 42618 258102 42854
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 257546 -2502 257782 -2266
rect 257866 -2502 258102 -2266
rect 257546 -2822 257782 -2586
rect 257866 -2822 258102 -2586
rect 261266 46658 261502 46894
rect 261586 46658 261822 46894
rect 261266 46338 261502 46574
rect 261586 46338 261822 46574
rect 264986 86378 265222 86614
rect 265306 86378 265542 86614
rect 264986 86058 265222 86294
rect 265306 86058 265542 86294
rect 271826 93218 272062 93454
rect 272146 93218 272382 93454
rect 271826 92898 272062 93134
rect 272146 92898 272382 93134
rect 264986 50378 265222 50614
rect 265306 50378 265542 50614
rect 264986 50058 265222 50294
rect 265306 50058 265542 50294
rect 261266 10658 261502 10894
rect 261586 10658 261822 10894
rect 261266 10338 261502 10574
rect 261586 10338 261822 10574
rect 261266 -4422 261502 -4186
rect 261586 -4422 261822 -4186
rect 261266 -4742 261502 -4506
rect 261586 -4742 261822 -4506
rect 264986 14378 265222 14614
rect 265306 14378 265542 14614
rect 264986 14058 265222 14294
rect 265306 14058 265542 14294
rect 246986 -7302 247222 -7066
rect 247306 -7302 247542 -7066
rect 246986 -7622 247222 -7386
rect 247306 -7622 247542 -7386
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 275546 96938 275782 97174
rect 275866 96938 276102 97174
rect 275546 96618 275782 96854
rect 275866 96618 276102 96854
rect 275546 60938 275782 61174
rect 275866 60938 276102 61174
rect 275546 60618 275782 60854
rect 275866 60618 276102 60854
rect 275546 24938 275782 25174
rect 275866 24938 276102 25174
rect 275546 24618 275782 24854
rect 275866 24618 276102 24854
rect 271826 -1542 272062 -1306
rect 272146 -1542 272382 -1306
rect 271826 -1862 272062 -1626
rect 272146 -1862 272382 -1626
rect 275546 -3462 275782 -3226
rect 275866 -3462 276102 -3226
rect 275546 -3782 275782 -3546
rect 275866 -3782 276102 -3546
rect 279266 64658 279502 64894
rect 279586 64658 279822 64894
rect 279266 64338 279502 64574
rect 279586 64338 279822 64574
rect 279266 28658 279502 28894
rect 279586 28658 279822 28894
rect 279266 28338 279502 28574
rect 279586 28338 279822 28574
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 282986 68378 283222 68614
rect 283306 68378 283542 68614
rect 282986 68058 283222 68294
rect 283306 68058 283542 68294
rect 282986 32378 283222 32614
rect 283306 32378 283542 32614
rect 282986 32058 283222 32294
rect 283306 32058 283542 32294
rect 279266 -5382 279502 -5146
rect 279586 -5382 279822 -5146
rect 279266 -5702 279502 -5466
rect 279586 -5702 279822 -5466
rect 264986 -6342 265222 -6106
rect 265306 -6342 265542 -6106
rect 264986 -6662 265222 -6426
rect 265306 -6662 265542 -6426
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 293546 78938 293782 79174
rect 293866 78938 294102 79174
rect 293546 78618 293782 78854
rect 293866 78618 294102 78854
rect 293546 42938 293782 43174
rect 293866 42938 294102 43174
rect 293546 42618 293782 42854
rect 293866 42618 294102 42854
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 293546 -2502 293782 -2266
rect 293866 -2502 294102 -2266
rect 293546 -2822 293782 -2586
rect 293866 -2822 294102 -2586
rect 297266 82658 297502 82894
rect 297586 82658 297822 82894
rect 297266 82338 297502 82574
rect 297586 82338 297822 82574
rect 300986 86378 301222 86614
rect 301306 86378 301542 86614
rect 300986 86058 301222 86294
rect 301306 86058 301542 86294
rect 300986 50378 301222 50614
rect 301306 50378 301542 50614
rect 297266 46658 297502 46894
rect 297586 46658 297822 46894
rect 297266 46338 297502 46574
rect 297586 46338 297822 46574
rect 297266 10658 297502 10894
rect 297586 10658 297822 10894
rect 297266 10338 297502 10574
rect 297586 10338 297822 10574
rect 297266 -4422 297502 -4186
rect 297586 -4422 297822 -4186
rect 297266 -4742 297502 -4506
rect 297586 -4742 297822 -4506
rect 300986 50058 301222 50294
rect 301306 50058 301542 50294
rect 300986 14378 301222 14614
rect 301306 14378 301542 14614
rect 300986 14058 301222 14294
rect 301306 14058 301542 14294
rect 282986 -7302 283222 -7066
rect 283306 -7302 283542 -7066
rect 282986 -7622 283222 -7386
rect 283306 -7622 283542 -7386
rect 307826 93218 308062 93454
rect 308146 93218 308382 93454
rect 307826 92898 308062 93134
rect 308146 92898 308382 93134
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -1542 308062 -1306
rect 308146 -1542 308382 -1306
rect 307826 -1862 308062 -1626
rect 308146 -1862 308382 -1626
rect 311546 672938 311782 673174
rect 311866 672938 312102 673174
rect 311546 672618 311782 672854
rect 311866 672618 312102 672854
rect 311546 636938 311782 637174
rect 311866 636938 312102 637174
rect 311546 636618 311782 636854
rect 311866 636618 312102 636854
rect 311546 600938 311782 601174
rect 311866 600938 312102 601174
rect 311546 600618 311782 600854
rect 311866 600618 312102 600854
rect 311546 564938 311782 565174
rect 311866 564938 312102 565174
rect 311546 564618 311782 564854
rect 311866 564618 312102 564854
rect 311546 528938 311782 529174
rect 311866 528938 312102 529174
rect 311546 528618 311782 528854
rect 311866 528618 312102 528854
rect 311546 492938 311782 493174
rect 311866 492938 312102 493174
rect 311546 492618 311782 492854
rect 311866 492618 312102 492854
rect 311546 456938 311782 457174
rect 311866 456938 312102 457174
rect 311546 456618 311782 456854
rect 311866 456618 312102 456854
rect 311546 420938 311782 421174
rect 311866 420938 312102 421174
rect 311546 420618 311782 420854
rect 311866 420618 312102 420854
rect 311546 384938 311782 385174
rect 311866 384938 312102 385174
rect 311546 384618 311782 384854
rect 311866 384618 312102 384854
rect 311546 348938 311782 349174
rect 311866 348938 312102 349174
rect 311546 348618 311782 348854
rect 311866 348618 312102 348854
rect 311546 312938 311782 313174
rect 311866 312938 312102 313174
rect 311546 312618 311782 312854
rect 311866 312618 312102 312854
rect 311546 276938 311782 277174
rect 311866 276938 312102 277174
rect 311546 276618 311782 276854
rect 311866 276618 312102 276854
rect 311546 240938 311782 241174
rect 311866 240938 312102 241174
rect 311546 240618 311782 240854
rect 311866 240618 312102 240854
rect 311546 204938 311782 205174
rect 311866 204938 312102 205174
rect 311546 204618 311782 204854
rect 311866 204618 312102 204854
rect 311546 168938 311782 169174
rect 311866 168938 312102 169174
rect 311546 168618 311782 168854
rect 311866 168618 312102 168854
rect 311546 132938 311782 133174
rect 311866 132938 312102 133174
rect 311546 132618 311782 132854
rect 311866 132618 312102 132854
rect 311546 96938 311782 97174
rect 311866 96938 312102 97174
rect 311546 96618 311782 96854
rect 311866 96618 312102 96854
rect 311546 60938 311782 61174
rect 311866 60938 312102 61174
rect 311546 60618 311782 60854
rect 311866 60618 312102 60854
rect 311546 24938 311782 25174
rect 311866 24938 312102 25174
rect 311546 24618 311782 24854
rect 311866 24618 312102 24854
rect 311546 -3462 311782 -3226
rect 311866 -3462 312102 -3226
rect 311546 -3782 311782 -3546
rect 311866 -3782 312102 -3546
rect 315266 676658 315502 676894
rect 315586 676658 315822 676894
rect 315266 676338 315502 676574
rect 315586 676338 315822 676574
rect 315266 640658 315502 640894
rect 315586 640658 315822 640894
rect 315266 640338 315502 640574
rect 315586 640338 315822 640574
rect 315266 604658 315502 604894
rect 315586 604658 315822 604894
rect 315266 604338 315502 604574
rect 315586 604338 315822 604574
rect 315266 568658 315502 568894
rect 315586 568658 315822 568894
rect 315266 568338 315502 568574
rect 315586 568338 315822 568574
rect 315266 532658 315502 532894
rect 315586 532658 315822 532894
rect 315266 532338 315502 532574
rect 315586 532338 315822 532574
rect 315266 496658 315502 496894
rect 315586 496658 315822 496894
rect 315266 496338 315502 496574
rect 315586 496338 315822 496574
rect 315266 460658 315502 460894
rect 315586 460658 315822 460894
rect 315266 460338 315502 460574
rect 315586 460338 315822 460574
rect 315266 424658 315502 424894
rect 315586 424658 315822 424894
rect 315266 424338 315502 424574
rect 315586 424338 315822 424574
rect 315266 388658 315502 388894
rect 315586 388658 315822 388894
rect 315266 388338 315502 388574
rect 315586 388338 315822 388574
rect 315266 352658 315502 352894
rect 315586 352658 315822 352894
rect 315266 352338 315502 352574
rect 315586 352338 315822 352574
rect 315266 316658 315502 316894
rect 315586 316658 315822 316894
rect 315266 316338 315502 316574
rect 315586 316338 315822 316574
rect 315266 280658 315502 280894
rect 315586 280658 315822 280894
rect 315266 280338 315502 280574
rect 315586 280338 315822 280574
rect 315266 244658 315502 244894
rect 315586 244658 315822 244894
rect 315266 244338 315502 244574
rect 315586 244338 315822 244574
rect 315266 208658 315502 208894
rect 315586 208658 315822 208894
rect 315266 208338 315502 208574
rect 315586 208338 315822 208574
rect 315266 172658 315502 172894
rect 315586 172658 315822 172894
rect 315266 172338 315502 172574
rect 315586 172338 315822 172574
rect 315266 136658 315502 136894
rect 315586 136658 315822 136894
rect 315266 136338 315502 136574
rect 315586 136338 315822 136574
rect 315266 100658 315502 100894
rect 315586 100658 315822 100894
rect 315266 100338 315502 100574
rect 315586 100338 315822 100574
rect 315266 64658 315502 64894
rect 315586 64658 315822 64894
rect 315266 64338 315502 64574
rect 315586 64338 315822 64574
rect 315266 28658 315502 28894
rect 315586 28658 315822 28894
rect 315266 28338 315502 28574
rect 315586 28338 315822 28574
rect 315266 -5382 315502 -5146
rect 315586 -5382 315822 -5146
rect 315266 -5702 315502 -5466
rect 315586 -5702 315822 -5466
rect 336986 710362 337222 710598
rect 337306 710362 337542 710598
rect 336986 710042 337222 710278
rect 337306 710042 337542 710278
rect 333266 708442 333502 708678
rect 333586 708442 333822 708678
rect 333266 708122 333502 708358
rect 333586 708122 333822 708358
rect 329546 706522 329782 706758
rect 329866 706522 330102 706758
rect 329546 706202 329782 706438
rect 329866 706202 330102 706438
rect 318986 680378 319222 680614
rect 319306 680378 319542 680614
rect 318986 680058 319222 680294
rect 319306 680058 319542 680294
rect 318986 644378 319222 644614
rect 319306 644378 319542 644614
rect 318986 644058 319222 644294
rect 319306 644058 319542 644294
rect 318986 608378 319222 608614
rect 319306 608378 319542 608614
rect 318986 608058 319222 608294
rect 319306 608058 319542 608294
rect 318986 572378 319222 572614
rect 319306 572378 319542 572614
rect 318986 572058 319222 572294
rect 319306 572058 319542 572294
rect 318986 536378 319222 536614
rect 319306 536378 319542 536614
rect 318986 536058 319222 536294
rect 319306 536058 319542 536294
rect 318986 500378 319222 500614
rect 319306 500378 319542 500614
rect 318986 500058 319222 500294
rect 319306 500058 319542 500294
rect 318986 464378 319222 464614
rect 319306 464378 319542 464614
rect 318986 464058 319222 464294
rect 319306 464058 319542 464294
rect 318986 428378 319222 428614
rect 319306 428378 319542 428614
rect 318986 428058 319222 428294
rect 319306 428058 319542 428294
rect 318986 392378 319222 392614
rect 319306 392378 319542 392614
rect 318986 392058 319222 392294
rect 319306 392058 319542 392294
rect 318986 356378 319222 356614
rect 319306 356378 319542 356614
rect 318986 356058 319222 356294
rect 319306 356058 319542 356294
rect 318986 320378 319222 320614
rect 319306 320378 319542 320614
rect 318986 320058 319222 320294
rect 319306 320058 319542 320294
rect 318986 284378 319222 284614
rect 319306 284378 319542 284614
rect 318986 284058 319222 284294
rect 319306 284058 319542 284294
rect 318986 248378 319222 248614
rect 319306 248378 319542 248614
rect 318986 248058 319222 248294
rect 319306 248058 319542 248294
rect 318986 212378 319222 212614
rect 319306 212378 319542 212614
rect 318986 212058 319222 212294
rect 319306 212058 319542 212294
rect 318986 176378 319222 176614
rect 319306 176378 319542 176614
rect 318986 176058 319222 176294
rect 319306 176058 319542 176294
rect 318986 140378 319222 140614
rect 319306 140378 319542 140614
rect 318986 140058 319222 140294
rect 319306 140058 319542 140294
rect 318986 104378 319222 104614
rect 319306 104378 319542 104614
rect 318986 104058 319222 104294
rect 319306 104058 319542 104294
rect 318986 68378 319222 68614
rect 319306 68378 319542 68614
rect 318986 68058 319222 68294
rect 319306 68058 319542 68294
rect 318986 32378 319222 32614
rect 319306 32378 319542 32614
rect 318986 32058 319222 32294
rect 319306 32058 319542 32294
rect 300986 -6342 301222 -6106
rect 301306 -6342 301542 -6106
rect 300986 -6662 301222 -6426
rect 301306 -6662 301542 -6426
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 325826 543218 326062 543454
rect 326146 543218 326382 543454
rect 325826 542898 326062 543134
rect 326146 542898 326382 543134
rect 325826 507218 326062 507454
rect 326146 507218 326382 507454
rect 325826 506898 326062 507134
rect 326146 506898 326382 507134
rect 325826 471218 326062 471454
rect 326146 471218 326382 471454
rect 325826 470898 326062 471134
rect 326146 470898 326382 471134
rect 325826 435218 326062 435454
rect 326146 435218 326382 435454
rect 325826 434898 326062 435134
rect 326146 434898 326382 435134
rect 325826 399218 326062 399454
rect 326146 399218 326382 399454
rect 325826 398898 326062 399134
rect 326146 398898 326382 399134
rect 325826 363218 326062 363454
rect 326146 363218 326382 363454
rect 325826 362898 326062 363134
rect 326146 362898 326382 363134
rect 325826 327218 326062 327454
rect 326146 327218 326382 327454
rect 325826 326898 326062 327134
rect 326146 326898 326382 327134
rect 325826 291218 326062 291454
rect 326146 291218 326382 291454
rect 325826 290898 326062 291134
rect 326146 290898 326382 291134
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 325826 219218 326062 219454
rect 326146 219218 326382 219454
rect 325826 218898 326062 219134
rect 326146 218898 326382 219134
rect 325826 183218 326062 183454
rect 326146 183218 326382 183454
rect 325826 182898 326062 183134
rect 326146 182898 326382 183134
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 325826 111218 326062 111454
rect 326146 111218 326382 111454
rect 325826 110898 326062 111134
rect 326146 110898 326382 111134
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 690938 329782 691174
rect 329866 690938 330102 691174
rect 329546 690618 329782 690854
rect 329866 690618 330102 690854
rect 329546 654938 329782 655174
rect 329866 654938 330102 655174
rect 329546 654618 329782 654854
rect 329866 654618 330102 654854
rect 329546 618938 329782 619174
rect 329866 618938 330102 619174
rect 329546 618618 329782 618854
rect 329866 618618 330102 618854
rect 329546 582938 329782 583174
rect 329866 582938 330102 583174
rect 329546 582618 329782 582854
rect 329866 582618 330102 582854
rect 329546 546938 329782 547174
rect 329866 546938 330102 547174
rect 329546 546618 329782 546854
rect 329866 546618 330102 546854
rect 329546 510938 329782 511174
rect 329866 510938 330102 511174
rect 329546 510618 329782 510854
rect 329866 510618 330102 510854
rect 329546 474938 329782 475174
rect 329866 474938 330102 475174
rect 329546 474618 329782 474854
rect 329866 474618 330102 474854
rect 329546 438938 329782 439174
rect 329866 438938 330102 439174
rect 329546 438618 329782 438854
rect 329866 438618 330102 438854
rect 329546 402938 329782 403174
rect 329866 402938 330102 403174
rect 329546 402618 329782 402854
rect 329866 402618 330102 402854
rect 329546 366938 329782 367174
rect 329866 366938 330102 367174
rect 329546 366618 329782 366854
rect 329866 366618 330102 366854
rect 329546 330938 329782 331174
rect 329866 330938 330102 331174
rect 329546 330618 329782 330854
rect 329866 330618 330102 330854
rect 329546 294938 329782 295174
rect 329866 294938 330102 295174
rect 329546 294618 329782 294854
rect 329866 294618 330102 294854
rect 329546 258938 329782 259174
rect 329866 258938 330102 259174
rect 329546 258618 329782 258854
rect 329866 258618 330102 258854
rect 329546 222938 329782 223174
rect 329866 222938 330102 223174
rect 329546 222618 329782 222854
rect 329866 222618 330102 222854
rect 329546 186938 329782 187174
rect 329866 186938 330102 187174
rect 329546 186618 329782 186854
rect 329866 186618 330102 186854
rect 329546 150938 329782 151174
rect 329866 150938 330102 151174
rect 329546 150618 329782 150854
rect 329866 150618 330102 150854
rect 329546 114938 329782 115174
rect 329866 114938 330102 115174
rect 329546 114618 329782 114854
rect 329866 114618 330102 114854
rect 329546 78938 329782 79174
rect 329866 78938 330102 79174
rect 329546 78618 329782 78854
rect 329866 78618 330102 78854
rect 329546 42938 329782 43174
rect 329866 42938 330102 43174
rect 329546 42618 329782 42854
rect 329866 42618 330102 42854
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 329546 -2502 329782 -2266
rect 329866 -2502 330102 -2266
rect 329546 -2822 329782 -2586
rect 329866 -2822 330102 -2586
rect 333266 694658 333502 694894
rect 333586 694658 333822 694894
rect 333266 694338 333502 694574
rect 333586 694338 333822 694574
rect 333266 658658 333502 658894
rect 333586 658658 333822 658894
rect 333266 658338 333502 658574
rect 333586 658338 333822 658574
rect 333266 622658 333502 622894
rect 333586 622658 333822 622894
rect 333266 622338 333502 622574
rect 333586 622338 333822 622574
rect 333266 586658 333502 586894
rect 333586 586658 333822 586894
rect 333266 586338 333502 586574
rect 333586 586338 333822 586574
rect 333266 550658 333502 550894
rect 333586 550658 333822 550894
rect 333266 550338 333502 550574
rect 333586 550338 333822 550574
rect 333266 514658 333502 514894
rect 333586 514658 333822 514894
rect 333266 514338 333502 514574
rect 333586 514338 333822 514574
rect 333266 478658 333502 478894
rect 333586 478658 333822 478894
rect 333266 478338 333502 478574
rect 333586 478338 333822 478574
rect 333266 442658 333502 442894
rect 333586 442658 333822 442894
rect 333266 442338 333502 442574
rect 333586 442338 333822 442574
rect 333266 406658 333502 406894
rect 333586 406658 333822 406894
rect 333266 406338 333502 406574
rect 333586 406338 333822 406574
rect 333266 370658 333502 370894
rect 333586 370658 333822 370894
rect 333266 370338 333502 370574
rect 333586 370338 333822 370574
rect 333266 334658 333502 334894
rect 333586 334658 333822 334894
rect 333266 334338 333502 334574
rect 333586 334338 333822 334574
rect 333266 298658 333502 298894
rect 333586 298658 333822 298894
rect 333266 298338 333502 298574
rect 333586 298338 333822 298574
rect 333266 262658 333502 262894
rect 333586 262658 333822 262894
rect 333266 262338 333502 262574
rect 333586 262338 333822 262574
rect 333266 226658 333502 226894
rect 333586 226658 333822 226894
rect 333266 226338 333502 226574
rect 333586 226338 333822 226574
rect 333266 190658 333502 190894
rect 333586 190658 333822 190894
rect 333266 190338 333502 190574
rect 333586 190338 333822 190574
rect 333266 154658 333502 154894
rect 333586 154658 333822 154894
rect 333266 154338 333502 154574
rect 333586 154338 333822 154574
rect 333266 118658 333502 118894
rect 333586 118658 333822 118894
rect 333266 118338 333502 118574
rect 333586 118338 333822 118574
rect 333266 82658 333502 82894
rect 333586 82658 333822 82894
rect 333266 82338 333502 82574
rect 333586 82338 333822 82574
rect 333266 46658 333502 46894
rect 333586 46658 333822 46894
rect 333266 46338 333502 46574
rect 333586 46338 333822 46574
rect 333266 10658 333502 10894
rect 333586 10658 333822 10894
rect 333266 10338 333502 10574
rect 333586 10338 333822 10574
rect 333266 -4422 333502 -4186
rect 333586 -4422 333822 -4186
rect 333266 -4742 333502 -4506
rect 333586 -4742 333822 -4506
rect 354986 711322 355222 711558
rect 355306 711322 355542 711558
rect 354986 711002 355222 711238
rect 355306 711002 355542 711238
rect 351266 709402 351502 709638
rect 351586 709402 351822 709638
rect 351266 709082 351502 709318
rect 351586 709082 351822 709318
rect 347546 707482 347782 707718
rect 347866 707482 348102 707718
rect 347546 707162 347782 707398
rect 347866 707162 348102 707398
rect 336986 698378 337222 698614
rect 337306 698378 337542 698614
rect 336986 698058 337222 698294
rect 337306 698058 337542 698294
rect 336986 662378 337222 662614
rect 337306 662378 337542 662614
rect 336986 662058 337222 662294
rect 337306 662058 337542 662294
rect 336986 626378 337222 626614
rect 337306 626378 337542 626614
rect 336986 626058 337222 626294
rect 337306 626058 337542 626294
rect 336986 590378 337222 590614
rect 337306 590378 337542 590614
rect 336986 590058 337222 590294
rect 337306 590058 337542 590294
rect 336986 554378 337222 554614
rect 337306 554378 337542 554614
rect 336986 554058 337222 554294
rect 337306 554058 337542 554294
rect 336986 518378 337222 518614
rect 337306 518378 337542 518614
rect 336986 518058 337222 518294
rect 337306 518058 337542 518294
rect 336986 482378 337222 482614
rect 337306 482378 337542 482614
rect 336986 482058 337222 482294
rect 337306 482058 337542 482294
rect 336986 446378 337222 446614
rect 337306 446378 337542 446614
rect 336986 446058 337222 446294
rect 337306 446058 337542 446294
rect 336986 410378 337222 410614
rect 337306 410378 337542 410614
rect 336986 410058 337222 410294
rect 337306 410058 337542 410294
rect 336986 374378 337222 374614
rect 337306 374378 337542 374614
rect 336986 374058 337222 374294
rect 337306 374058 337542 374294
rect 336986 338378 337222 338614
rect 337306 338378 337542 338614
rect 336986 338058 337222 338294
rect 337306 338058 337542 338294
rect 336986 302378 337222 302614
rect 337306 302378 337542 302614
rect 336986 302058 337222 302294
rect 337306 302058 337542 302294
rect 336986 266378 337222 266614
rect 337306 266378 337542 266614
rect 336986 266058 337222 266294
rect 337306 266058 337542 266294
rect 336986 230378 337222 230614
rect 337306 230378 337542 230614
rect 336986 230058 337222 230294
rect 337306 230058 337542 230294
rect 336986 194378 337222 194614
rect 337306 194378 337542 194614
rect 336986 194058 337222 194294
rect 337306 194058 337542 194294
rect 336986 158378 337222 158614
rect 337306 158378 337542 158614
rect 336986 158058 337222 158294
rect 337306 158058 337542 158294
rect 336986 122378 337222 122614
rect 337306 122378 337542 122614
rect 336986 122058 337222 122294
rect 337306 122058 337542 122294
rect 336986 86378 337222 86614
rect 337306 86378 337542 86614
rect 336986 86058 337222 86294
rect 337306 86058 337542 86294
rect 336986 50378 337222 50614
rect 337306 50378 337542 50614
rect 336986 50058 337222 50294
rect 337306 50058 337542 50294
rect 336986 14378 337222 14614
rect 337306 14378 337542 14614
rect 336986 14058 337222 14294
rect 337306 14058 337542 14294
rect 318986 -7302 319222 -7066
rect 319306 -7302 319542 -7066
rect 318986 -7622 319222 -7386
rect 319306 -7622 319542 -7386
rect 343826 705562 344062 705798
rect 344146 705562 344382 705798
rect 343826 705242 344062 705478
rect 344146 705242 344382 705478
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 343826 561218 344062 561454
rect 344146 561218 344382 561454
rect 343826 560898 344062 561134
rect 344146 560898 344382 561134
rect 343826 525218 344062 525454
rect 344146 525218 344382 525454
rect 343826 524898 344062 525134
rect 344146 524898 344382 525134
rect 343826 489218 344062 489454
rect 344146 489218 344382 489454
rect 343826 488898 344062 489134
rect 344146 488898 344382 489134
rect 343826 453218 344062 453454
rect 344146 453218 344382 453454
rect 343826 452898 344062 453134
rect 344146 452898 344382 453134
rect 343826 417218 344062 417454
rect 344146 417218 344382 417454
rect 343826 416898 344062 417134
rect 344146 416898 344382 417134
rect 343826 381218 344062 381454
rect 344146 381218 344382 381454
rect 343826 380898 344062 381134
rect 344146 380898 344382 381134
rect 343826 345218 344062 345454
rect 344146 345218 344382 345454
rect 343826 344898 344062 345134
rect 344146 344898 344382 345134
rect 343826 309218 344062 309454
rect 344146 309218 344382 309454
rect 343826 308898 344062 309134
rect 344146 308898 344382 309134
rect 343826 273218 344062 273454
rect 344146 273218 344382 273454
rect 343826 272898 344062 273134
rect 344146 272898 344382 273134
rect 343826 237218 344062 237454
rect 344146 237218 344382 237454
rect 343826 236898 344062 237134
rect 344146 236898 344382 237134
rect 343826 201218 344062 201454
rect 344146 201218 344382 201454
rect 343826 200898 344062 201134
rect 344146 200898 344382 201134
rect 343826 165218 344062 165454
rect 344146 165218 344382 165454
rect 343826 164898 344062 165134
rect 344146 164898 344382 165134
rect 343826 129218 344062 129454
rect 344146 129218 344382 129454
rect 343826 128898 344062 129134
rect 344146 128898 344382 129134
rect 343826 93218 344062 93454
rect 344146 93218 344382 93454
rect 343826 92898 344062 93134
rect 344146 92898 344382 93134
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -1542 344062 -1306
rect 344146 -1542 344382 -1306
rect 343826 -1862 344062 -1626
rect 344146 -1862 344382 -1626
rect 347546 672938 347782 673174
rect 347866 672938 348102 673174
rect 347546 672618 347782 672854
rect 347866 672618 348102 672854
rect 347546 636938 347782 637174
rect 347866 636938 348102 637174
rect 347546 636618 347782 636854
rect 347866 636618 348102 636854
rect 347546 600938 347782 601174
rect 347866 600938 348102 601174
rect 347546 600618 347782 600854
rect 347866 600618 348102 600854
rect 347546 564938 347782 565174
rect 347866 564938 348102 565174
rect 347546 564618 347782 564854
rect 347866 564618 348102 564854
rect 347546 528938 347782 529174
rect 347866 528938 348102 529174
rect 347546 528618 347782 528854
rect 347866 528618 348102 528854
rect 347546 492938 347782 493174
rect 347866 492938 348102 493174
rect 347546 492618 347782 492854
rect 347866 492618 348102 492854
rect 347546 456938 347782 457174
rect 347866 456938 348102 457174
rect 347546 456618 347782 456854
rect 347866 456618 348102 456854
rect 347546 420938 347782 421174
rect 347866 420938 348102 421174
rect 347546 420618 347782 420854
rect 347866 420618 348102 420854
rect 347546 384938 347782 385174
rect 347866 384938 348102 385174
rect 347546 384618 347782 384854
rect 347866 384618 348102 384854
rect 347546 348938 347782 349174
rect 347866 348938 348102 349174
rect 347546 348618 347782 348854
rect 347866 348618 348102 348854
rect 347546 312938 347782 313174
rect 347866 312938 348102 313174
rect 347546 312618 347782 312854
rect 347866 312618 348102 312854
rect 347546 276938 347782 277174
rect 347866 276938 348102 277174
rect 347546 276618 347782 276854
rect 347866 276618 348102 276854
rect 347546 240938 347782 241174
rect 347866 240938 348102 241174
rect 347546 240618 347782 240854
rect 347866 240618 348102 240854
rect 347546 204938 347782 205174
rect 347866 204938 348102 205174
rect 347546 204618 347782 204854
rect 347866 204618 348102 204854
rect 347546 168938 347782 169174
rect 347866 168938 348102 169174
rect 347546 168618 347782 168854
rect 347866 168618 348102 168854
rect 347546 132938 347782 133174
rect 347866 132938 348102 133174
rect 347546 132618 347782 132854
rect 347866 132618 348102 132854
rect 347546 96938 347782 97174
rect 347866 96938 348102 97174
rect 347546 96618 347782 96854
rect 347866 96618 348102 96854
rect 347546 60938 347782 61174
rect 347866 60938 348102 61174
rect 347546 60618 347782 60854
rect 347866 60618 348102 60854
rect 347546 24938 347782 25174
rect 347866 24938 348102 25174
rect 347546 24618 347782 24854
rect 347866 24618 348102 24854
rect 347546 -3462 347782 -3226
rect 347866 -3462 348102 -3226
rect 347546 -3782 347782 -3546
rect 347866 -3782 348102 -3546
rect 351266 676658 351502 676894
rect 351586 676658 351822 676894
rect 351266 676338 351502 676574
rect 351586 676338 351822 676574
rect 351266 640658 351502 640894
rect 351586 640658 351822 640894
rect 351266 640338 351502 640574
rect 351586 640338 351822 640574
rect 351266 604658 351502 604894
rect 351586 604658 351822 604894
rect 351266 604338 351502 604574
rect 351586 604338 351822 604574
rect 351266 568658 351502 568894
rect 351586 568658 351822 568894
rect 351266 568338 351502 568574
rect 351586 568338 351822 568574
rect 351266 532658 351502 532894
rect 351586 532658 351822 532894
rect 351266 532338 351502 532574
rect 351586 532338 351822 532574
rect 351266 496658 351502 496894
rect 351586 496658 351822 496894
rect 351266 496338 351502 496574
rect 351586 496338 351822 496574
rect 351266 460658 351502 460894
rect 351586 460658 351822 460894
rect 351266 460338 351502 460574
rect 351586 460338 351822 460574
rect 351266 424658 351502 424894
rect 351586 424658 351822 424894
rect 351266 424338 351502 424574
rect 351586 424338 351822 424574
rect 351266 388658 351502 388894
rect 351586 388658 351822 388894
rect 351266 388338 351502 388574
rect 351586 388338 351822 388574
rect 351266 352658 351502 352894
rect 351586 352658 351822 352894
rect 351266 352338 351502 352574
rect 351586 352338 351822 352574
rect 351266 316658 351502 316894
rect 351586 316658 351822 316894
rect 351266 316338 351502 316574
rect 351586 316338 351822 316574
rect 351266 280658 351502 280894
rect 351586 280658 351822 280894
rect 351266 280338 351502 280574
rect 351586 280338 351822 280574
rect 351266 244658 351502 244894
rect 351586 244658 351822 244894
rect 351266 244338 351502 244574
rect 351586 244338 351822 244574
rect 351266 208658 351502 208894
rect 351586 208658 351822 208894
rect 351266 208338 351502 208574
rect 351586 208338 351822 208574
rect 351266 172658 351502 172894
rect 351586 172658 351822 172894
rect 351266 172338 351502 172574
rect 351586 172338 351822 172574
rect 351266 136658 351502 136894
rect 351586 136658 351822 136894
rect 351266 136338 351502 136574
rect 351586 136338 351822 136574
rect 351266 100658 351502 100894
rect 351586 100658 351822 100894
rect 351266 100338 351502 100574
rect 351586 100338 351822 100574
rect 351266 64658 351502 64894
rect 351586 64658 351822 64894
rect 351266 64338 351502 64574
rect 351586 64338 351822 64574
rect 351266 28658 351502 28894
rect 351586 28658 351822 28894
rect 351266 28338 351502 28574
rect 351586 28338 351822 28574
rect 351266 -5382 351502 -5146
rect 351586 -5382 351822 -5146
rect 351266 -5702 351502 -5466
rect 351586 -5702 351822 -5466
rect 372986 710362 373222 710598
rect 373306 710362 373542 710598
rect 372986 710042 373222 710278
rect 373306 710042 373542 710278
rect 369266 708442 369502 708678
rect 369586 708442 369822 708678
rect 369266 708122 369502 708358
rect 369586 708122 369822 708358
rect 365546 706522 365782 706758
rect 365866 706522 366102 706758
rect 365546 706202 365782 706438
rect 365866 706202 366102 706438
rect 354986 680378 355222 680614
rect 355306 680378 355542 680614
rect 354986 680058 355222 680294
rect 355306 680058 355542 680294
rect 354986 644378 355222 644614
rect 355306 644378 355542 644614
rect 354986 644058 355222 644294
rect 355306 644058 355542 644294
rect 354986 608378 355222 608614
rect 355306 608378 355542 608614
rect 354986 608058 355222 608294
rect 355306 608058 355542 608294
rect 354986 572378 355222 572614
rect 355306 572378 355542 572614
rect 354986 572058 355222 572294
rect 355306 572058 355542 572294
rect 354986 536378 355222 536614
rect 355306 536378 355542 536614
rect 354986 536058 355222 536294
rect 355306 536058 355542 536294
rect 354986 500378 355222 500614
rect 355306 500378 355542 500614
rect 354986 500058 355222 500294
rect 355306 500058 355542 500294
rect 354986 464378 355222 464614
rect 355306 464378 355542 464614
rect 354986 464058 355222 464294
rect 355306 464058 355542 464294
rect 354986 428378 355222 428614
rect 355306 428378 355542 428614
rect 354986 428058 355222 428294
rect 355306 428058 355542 428294
rect 354986 392378 355222 392614
rect 355306 392378 355542 392614
rect 354986 392058 355222 392294
rect 355306 392058 355542 392294
rect 354986 356378 355222 356614
rect 355306 356378 355542 356614
rect 354986 356058 355222 356294
rect 355306 356058 355542 356294
rect 354986 320378 355222 320614
rect 355306 320378 355542 320614
rect 354986 320058 355222 320294
rect 355306 320058 355542 320294
rect 354986 284378 355222 284614
rect 355306 284378 355542 284614
rect 354986 284058 355222 284294
rect 355306 284058 355542 284294
rect 354986 248378 355222 248614
rect 355306 248378 355542 248614
rect 354986 248058 355222 248294
rect 355306 248058 355542 248294
rect 354986 212378 355222 212614
rect 355306 212378 355542 212614
rect 354986 212058 355222 212294
rect 355306 212058 355542 212294
rect 354986 176378 355222 176614
rect 355306 176378 355542 176614
rect 354986 176058 355222 176294
rect 355306 176058 355542 176294
rect 354986 140378 355222 140614
rect 355306 140378 355542 140614
rect 354986 140058 355222 140294
rect 355306 140058 355542 140294
rect 354986 104378 355222 104614
rect 355306 104378 355542 104614
rect 354986 104058 355222 104294
rect 355306 104058 355542 104294
rect 354986 68378 355222 68614
rect 355306 68378 355542 68614
rect 354986 68058 355222 68294
rect 355306 68058 355542 68294
rect 354986 32378 355222 32614
rect 355306 32378 355542 32614
rect 354986 32058 355222 32294
rect 355306 32058 355542 32294
rect 336986 -6342 337222 -6106
rect 337306 -6342 337542 -6106
rect 336986 -6662 337222 -6426
rect 337306 -6662 337542 -6426
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 361826 435218 362062 435454
rect 362146 435218 362382 435454
rect 361826 434898 362062 435134
rect 362146 434898 362382 435134
rect 361826 399218 362062 399454
rect 362146 399218 362382 399454
rect 361826 398898 362062 399134
rect 362146 398898 362382 399134
rect 361826 363218 362062 363454
rect 362146 363218 362382 363454
rect 361826 362898 362062 363134
rect 362146 362898 362382 363134
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 365546 690938 365782 691174
rect 365866 690938 366102 691174
rect 365546 690618 365782 690854
rect 365866 690618 366102 690854
rect 365546 654938 365782 655174
rect 365866 654938 366102 655174
rect 365546 654618 365782 654854
rect 365866 654618 366102 654854
rect 365546 618938 365782 619174
rect 365866 618938 366102 619174
rect 365546 618618 365782 618854
rect 365866 618618 366102 618854
rect 365546 582938 365782 583174
rect 365866 582938 366102 583174
rect 365546 582618 365782 582854
rect 365866 582618 366102 582854
rect 365546 546938 365782 547174
rect 365866 546938 366102 547174
rect 365546 546618 365782 546854
rect 365866 546618 366102 546854
rect 365546 510938 365782 511174
rect 365866 510938 366102 511174
rect 365546 510618 365782 510854
rect 365866 510618 366102 510854
rect 365546 474938 365782 475174
rect 365866 474938 366102 475174
rect 365546 474618 365782 474854
rect 365866 474618 366102 474854
rect 365546 438938 365782 439174
rect 365866 438938 366102 439174
rect 365546 438618 365782 438854
rect 365866 438618 366102 438854
rect 365546 402938 365782 403174
rect 365866 402938 366102 403174
rect 365546 402618 365782 402854
rect 365866 402618 366102 402854
rect 365546 366938 365782 367174
rect 365866 366938 366102 367174
rect 365546 366618 365782 366854
rect 365866 366618 366102 366854
rect 365546 330938 365782 331174
rect 365866 330938 366102 331174
rect 365546 330618 365782 330854
rect 365866 330618 366102 330854
rect 365546 294938 365782 295174
rect 365866 294938 366102 295174
rect 365546 294618 365782 294854
rect 365866 294618 366102 294854
rect 365546 258938 365782 259174
rect 365866 258938 366102 259174
rect 365546 258618 365782 258854
rect 365866 258618 366102 258854
rect 365546 222938 365782 223174
rect 365866 222938 366102 223174
rect 365546 222618 365782 222854
rect 365866 222618 366102 222854
rect 365546 186938 365782 187174
rect 365866 186938 366102 187174
rect 365546 186618 365782 186854
rect 365866 186618 366102 186854
rect 365546 150938 365782 151174
rect 365866 150938 366102 151174
rect 365546 150618 365782 150854
rect 365866 150618 366102 150854
rect 365546 114938 365782 115174
rect 365866 114938 366102 115174
rect 365546 114618 365782 114854
rect 365866 114618 366102 114854
rect 365546 78938 365782 79174
rect 365866 78938 366102 79174
rect 365546 78618 365782 78854
rect 365866 78618 366102 78854
rect 365546 42938 365782 43174
rect 365866 42938 366102 43174
rect 365546 42618 365782 42854
rect 365866 42618 366102 42854
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 365546 -2502 365782 -2266
rect 365866 -2502 366102 -2266
rect 365546 -2822 365782 -2586
rect 365866 -2822 366102 -2586
rect 369266 694658 369502 694894
rect 369586 694658 369822 694894
rect 369266 694338 369502 694574
rect 369586 694338 369822 694574
rect 369266 658658 369502 658894
rect 369586 658658 369822 658894
rect 369266 658338 369502 658574
rect 369586 658338 369822 658574
rect 369266 622658 369502 622894
rect 369586 622658 369822 622894
rect 369266 622338 369502 622574
rect 369586 622338 369822 622574
rect 369266 586658 369502 586894
rect 369586 586658 369822 586894
rect 369266 586338 369502 586574
rect 369586 586338 369822 586574
rect 369266 550658 369502 550894
rect 369586 550658 369822 550894
rect 369266 550338 369502 550574
rect 369586 550338 369822 550574
rect 369266 514658 369502 514894
rect 369586 514658 369822 514894
rect 369266 514338 369502 514574
rect 369586 514338 369822 514574
rect 369266 478658 369502 478894
rect 369586 478658 369822 478894
rect 369266 478338 369502 478574
rect 369586 478338 369822 478574
rect 369266 442658 369502 442894
rect 369586 442658 369822 442894
rect 369266 442338 369502 442574
rect 369586 442338 369822 442574
rect 369266 406658 369502 406894
rect 369586 406658 369822 406894
rect 369266 406338 369502 406574
rect 369586 406338 369822 406574
rect 369266 370658 369502 370894
rect 369586 370658 369822 370894
rect 369266 370338 369502 370574
rect 369586 370338 369822 370574
rect 369266 334658 369502 334894
rect 369586 334658 369822 334894
rect 369266 334338 369502 334574
rect 369586 334338 369822 334574
rect 369266 298658 369502 298894
rect 369586 298658 369822 298894
rect 369266 298338 369502 298574
rect 369586 298338 369822 298574
rect 369266 262658 369502 262894
rect 369586 262658 369822 262894
rect 369266 262338 369502 262574
rect 369586 262338 369822 262574
rect 369266 226658 369502 226894
rect 369586 226658 369822 226894
rect 369266 226338 369502 226574
rect 369586 226338 369822 226574
rect 369266 190658 369502 190894
rect 369586 190658 369822 190894
rect 369266 190338 369502 190574
rect 369586 190338 369822 190574
rect 369266 154658 369502 154894
rect 369586 154658 369822 154894
rect 369266 154338 369502 154574
rect 369586 154338 369822 154574
rect 369266 118658 369502 118894
rect 369586 118658 369822 118894
rect 369266 118338 369502 118574
rect 369586 118338 369822 118574
rect 369266 82658 369502 82894
rect 369586 82658 369822 82894
rect 369266 82338 369502 82574
rect 369586 82338 369822 82574
rect 369266 46658 369502 46894
rect 369586 46658 369822 46894
rect 369266 46338 369502 46574
rect 369586 46338 369822 46574
rect 369266 10658 369502 10894
rect 369586 10658 369822 10894
rect 369266 10338 369502 10574
rect 369586 10338 369822 10574
rect 369266 -4422 369502 -4186
rect 369586 -4422 369822 -4186
rect 369266 -4742 369502 -4506
rect 369586 -4742 369822 -4506
rect 390986 711322 391222 711558
rect 391306 711322 391542 711558
rect 390986 711002 391222 711238
rect 391306 711002 391542 711238
rect 387266 709402 387502 709638
rect 387586 709402 387822 709638
rect 387266 709082 387502 709318
rect 387586 709082 387822 709318
rect 383546 707482 383782 707718
rect 383866 707482 384102 707718
rect 383546 707162 383782 707398
rect 383866 707162 384102 707398
rect 372986 698378 373222 698614
rect 373306 698378 373542 698614
rect 372986 698058 373222 698294
rect 373306 698058 373542 698294
rect 372986 662378 373222 662614
rect 373306 662378 373542 662614
rect 372986 662058 373222 662294
rect 373306 662058 373542 662294
rect 372986 626378 373222 626614
rect 373306 626378 373542 626614
rect 372986 626058 373222 626294
rect 373306 626058 373542 626294
rect 372986 590378 373222 590614
rect 373306 590378 373542 590614
rect 372986 590058 373222 590294
rect 373306 590058 373542 590294
rect 372986 554378 373222 554614
rect 373306 554378 373542 554614
rect 372986 554058 373222 554294
rect 373306 554058 373542 554294
rect 372986 518378 373222 518614
rect 373306 518378 373542 518614
rect 372986 518058 373222 518294
rect 373306 518058 373542 518294
rect 372986 482378 373222 482614
rect 373306 482378 373542 482614
rect 372986 482058 373222 482294
rect 373306 482058 373542 482294
rect 372986 446378 373222 446614
rect 373306 446378 373542 446614
rect 372986 446058 373222 446294
rect 373306 446058 373542 446294
rect 372986 410378 373222 410614
rect 373306 410378 373542 410614
rect 372986 410058 373222 410294
rect 373306 410058 373542 410294
rect 372986 374378 373222 374614
rect 373306 374378 373542 374614
rect 372986 374058 373222 374294
rect 373306 374058 373542 374294
rect 372986 338378 373222 338614
rect 373306 338378 373542 338614
rect 372986 338058 373222 338294
rect 373306 338058 373542 338294
rect 372986 302378 373222 302614
rect 373306 302378 373542 302614
rect 372986 302058 373222 302294
rect 373306 302058 373542 302294
rect 372986 266378 373222 266614
rect 373306 266378 373542 266614
rect 372986 266058 373222 266294
rect 373306 266058 373542 266294
rect 372986 230378 373222 230614
rect 373306 230378 373542 230614
rect 372986 230058 373222 230294
rect 373306 230058 373542 230294
rect 372986 194378 373222 194614
rect 373306 194378 373542 194614
rect 372986 194058 373222 194294
rect 373306 194058 373542 194294
rect 372986 158378 373222 158614
rect 373306 158378 373542 158614
rect 372986 158058 373222 158294
rect 373306 158058 373542 158294
rect 372986 122378 373222 122614
rect 373306 122378 373542 122614
rect 372986 122058 373222 122294
rect 373306 122058 373542 122294
rect 372986 86378 373222 86614
rect 373306 86378 373542 86614
rect 372986 86058 373222 86294
rect 373306 86058 373542 86294
rect 372986 50378 373222 50614
rect 373306 50378 373542 50614
rect 372986 50058 373222 50294
rect 373306 50058 373542 50294
rect 372986 14378 373222 14614
rect 373306 14378 373542 14614
rect 372986 14058 373222 14294
rect 373306 14058 373542 14294
rect 354986 -7302 355222 -7066
rect 355306 -7302 355542 -7066
rect 354986 -7622 355222 -7386
rect 355306 -7622 355542 -7386
rect 379826 705562 380062 705798
rect 380146 705562 380382 705798
rect 379826 705242 380062 705478
rect 380146 705242 380382 705478
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 379826 561218 380062 561454
rect 380146 561218 380382 561454
rect 379826 560898 380062 561134
rect 380146 560898 380382 561134
rect 379826 525218 380062 525454
rect 380146 525218 380382 525454
rect 379826 524898 380062 525134
rect 380146 524898 380382 525134
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 379826 453218 380062 453454
rect 380146 453218 380382 453454
rect 379826 452898 380062 453134
rect 380146 452898 380382 453134
rect 379826 417218 380062 417454
rect 380146 417218 380382 417454
rect 379826 416898 380062 417134
rect 380146 416898 380382 417134
rect 379826 381218 380062 381454
rect 380146 381218 380382 381454
rect 379826 380898 380062 381134
rect 380146 380898 380382 381134
rect 379826 345218 380062 345454
rect 380146 345218 380382 345454
rect 379826 344898 380062 345134
rect 380146 344898 380382 345134
rect 379826 309218 380062 309454
rect 380146 309218 380382 309454
rect 379826 308898 380062 309134
rect 380146 308898 380382 309134
rect 379826 273218 380062 273454
rect 380146 273218 380382 273454
rect 379826 272898 380062 273134
rect 380146 272898 380382 273134
rect 379826 237218 380062 237454
rect 380146 237218 380382 237454
rect 379826 236898 380062 237134
rect 380146 236898 380382 237134
rect 379826 201218 380062 201454
rect 380146 201218 380382 201454
rect 379826 200898 380062 201134
rect 380146 200898 380382 201134
rect 379826 165218 380062 165454
rect 380146 165218 380382 165454
rect 379826 164898 380062 165134
rect 380146 164898 380382 165134
rect 379826 129218 380062 129454
rect 380146 129218 380382 129454
rect 379826 128898 380062 129134
rect 380146 128898 380382 129134
rect 379826 93218 380062 93454
rect 380146 93218 380382 93454
rect 379826 92898 380062 93134
rect 380146 92898 380382 93134
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -1542 380062 -1306
rect 380146 -1542 380382 -1306
rect 379826 -1862 380062 -1626
rect 380146 -1862 380382 -1626
rect 383546 672938 383782 673174
rect 383866 672938 384102 673174
rect 383546 672618 383782 672854
rect 383866 672618 384102 672854
rect 383546 636938 383782 637174
rect 383866 636938 384102 637174
rect 383546 636618 383782 636854
rect 383866 636618 384102 636854
rect 383546 600938 383782 601174
rect 383866 600938 384102 601174
rect 383546 600618 383782 600854
rect 383866 600618 384102 600854
rect 383546 564938 383782 565174
rect 383866 564938 384102 565174
rect 383546 564618 383782 564854
rect 383866 564618 384102 564854
rect 383546 528938 383782 529174
rect 383866 528938 384102 529174
rect 383546 528618 383782 528854
rect 383866 528618 384102 528854
rect 383546 492938 383782 493174
rect 383866 492938 384102 493174
rect 383546 492618 383782 492854
rect 383866 492618 384102 492854
rect 383546 456938 383782 457174
rect 383866 456938 384102 457174
rect 383546 456618 383782 456854
rect 383866 456618 384102 456854
rect 383546 420938 383782 421174
rect 383866 420938 384102 421174
rect 383546 420618 383782 420854
rect 383866 420618 384102 420854
rect 383546 384938 383782 385174
rect 383866 384938 384102 385174
rect 383546 384618 383782 384854
rect 383866 384618 384102 384854
rect 383546 348938 383782 349174
rect 383866 348938 384102 349174
rect 383546 348618 383782 348854
rect 383866 348618 384102 348854
rect 383546 312938 383782 313174
rect 383866 312938 384102 313174
rect 383546 312618 383782 312854
rect 383866 312618 384102 312854
rect 383546 276938 383782 277174
rect 383866 276938 384102 277174
rect 383546 276618 383782 276854
rect 383866 276618 384102 276854
rect 383546 240938 383782 241174
rect 383866 240938 384102 241174
rect 383546 240618 383782 240854
rect 383866 240618 384102 240854
rect 383546 204938 383782 205174
rect 383866 204938 384102 205174
rect 383546 204618 383782 204854
rect 383866 204618 384102 204854
rect 383546 168938 383782 169174
rect 383866 168938 384102 169174
rect 383546 168618 383782 168854
rect 383866 168618 384102 168854
rect 383546 132938 383782 133174
rect 383866 132938 384102 133174
rect 383546 132618 383782 132854
rect 383866 132618 384102 132854
rect 383546 96938 383782 97174
rect 383866 96938 384102 97174
rect 383546 96618 383782 96854
rect 383866 96618 384102 96854
rect 383546 60938 383782 61174
rect 383866 60938 384102 61174
rect 383546 60618 383782 60854
rect 383866 60618 384102 60854
rect 383546 24938 383782 25174
rect 383866 24938 384102 25174
rect 383546 24618 383782 24854
rect 383866 24618 384102 24854
rect 383546 -3462 383782 -3226
rect 383866 -3462 384102 -3226
rect 383546 -3782 383782 -3546
rect 383866 -3782 384102 -3546
rect 387266 676658 387502 676894
rect 387586 676658 387822 676894
rect 387266 676338 387502 676574
rect 387586 676338 387822 676574
rect 387266 640658 387502 640894
rect 387586 640658 387822 640894
rect 387266 640338 387502 640574
rect 387586 640338 387822 640574
rect 387266 604658 387502 604894
rect 387586 604658 387822 604894
rect 387266 604338 387502 604574
rect 387586 604338 387822 604574
rect 387266 568658 387502 568894
rect 387586 568658 387822 568894
rect 387266 568338 387502 568574
rect 387586 568338 387822 568574
rect 387266 532658 387502 532894
rect 387586 532658 387822 532894
rect 387266 532338 387502 532574
rect 387586 532338 387822 532574
rect 387266 496658 387502 496894
rect 387586 496658 387822 496894
rect 387266 496338 387502 496574
rect 387586 496338 387822 496574
rect 387266 460658 387502 460894
rect 387586 460658 387822 460894
rect 387266 460338 387502 460574
rect 387586 460338 387822 460574
rect 387266 424658 387502 424894
rect 387586 424658 387822 424894
rect 387266 424338 387502 424574
rect 387586 424338 387822 424574
rect 387266 388658 387502 388894
rect 387586 388658 387822 388894
rect 387266 388338 387502 388574
rect 387586 388338 387822 388574
rect 387266 352658 387502 352894
rect 387586 352658 387822 352894
rect 387266 352338 387502 352574
rect 387586 352338 387822 352574
rect 387266 316658 387502 316894
rect 387586 316658 387822 316894
rect 387266 316338 387502 316574
rect 387586 316338 387822 316574
rect 387266 280658 387502 280894
rect 387586 280658 387822 280894
rect 387266 280338 387502 280574
rect 387586 280338 387822 280574
rect 387266 244658 387502 244894
rect 387586 244658 387822 244894
rect 387266 244338 387502 244574
rect 387586 244338 387822 244574
rect 387266 208658 387502 208894
rect 387586 208658 387822 208894
rect 387266 208338 387502 208574
rect 387586 208338 387822 208574
rect 387266 172658 387502 172894
rect 387586 172658 387822 172894
rect 387266 172338 387502 172574
rect 387586 172338 387822 172574
rect 387266 136658 387502 136894
rect 387586 136658 387822 136894
rect 387266 136338 387502 136574
rect 387586 136338 387822 136574
rect 387266 100658 387502 100894
rect 387586 100658 387822 100894
rect 387266 100338 387502 100574
rect 387586 100338 387822 100574
rect 387266 64658 387502 64894
rect 387586 64658 387822 64894
rect 387266 64338 387502 64574
rect 387586 64338 387822 64574
rect 387266 28658 387502 28894
rect 387586 28658 387822 28894
rect 387266 28338 387502 28574
rect 387586 28338 387822 28574
rect 387266 -5382 387502 -5146
rect 387586 -5382 387822 -5146
rect 387266 -5702 387502 -5466
rect 387586 -5702 387822 -5466
rect 408986 710362 409222 710598
rect 409306 710362 409542 710598
rect 408986 710042 409222 710278
rect 409306 710042 409542 710278
rect 405266 708442 405502 708678
rect 405586 708442 405822 708678
rect 405266 708122 405502 708358
rect 405586 708122 405822 708358
rect 401546 706522 401782 706758
rect 401866 706522 402102 706758
rect 401546 706202 401782 706438
rect 401866 706202 402102 706438
rect 390986 680378 391222 680614
rect 391306 680378 391542 680614
rect 390986 680058 391222 680294
rect 391306 680058 391542 680294
rect 390986 644378 391222 644614
rect 391306 644378 391542 644614
rect 390986 644058 391222 644294
rect 391306 644058 391542 644294
rect 390986 608378 391222 608614
rect 391306 608378 391542 608614
rect 390986 608058 391222 608294
rect 391306 608058 391542 608294
rect 390986 572378 391222 572614
rect 391306 572378 391542 572614
rect 390986 572058 391222 572294
rect 391306 572058 391542 572294
rect 390986 536378 391222 536614
rect 391306 536378 391542 536614
rect 390986 536058 391222 536294
rect 391306 536058 391542 536294
rect 390986 500378 391222 500614
rect 391306 500378 391542 500614
rect 390986 500058 391222 500294
rect 391306 500058 391542 500294
rect 390986 464378 391222 464614
rect 391306 464378 391542 464614
rect 390986 464058 391222 464294
rect 391306 464058 391542 464294
rect 390986 428378 391222 428614
rect 391306 428378 391542 428614
rect 390986 428058 391222 428294
rect 391306 428058 391542 428294
rect 390986 392378 391222 392614
rect 391306 392378 391542 392614
rect 390986 392058 391222 392294
rect 391306 392058 391542 392294
rect 390986 356378 391222 356614
rect 391306 356378 391542 356614
rect 390986 356058 391222 356294
rect 391306 356058 391542 356294
rect 390986 320378 391222 320614
rect 391306 320378 391542 320614
rect 390986 320058 391222 320294
rect 391306 320058 391542 320294
rect 390986 284378 391222 284614
rect 391306 284378 391542 284614
rect 390986 284058 391222 284294
rect 391306 284058 391542 284294
rect 390986 248378 391222 248614
rect 391306 248378 391542 248614
rect 390986 248058 391222 248294
rect 391306 248058 391542 248294
rect 390986 212378 391222 212614
rect 391306 212378 391542 212614
rect 390986 212058 391222 212294
rect 391306 212058 391542 212294
rect 390986 176378 391222 176614
rect 391306 176378 391542 176614
rect 390986 176058 391222 176294
rect 391306 176058 391542 176294
rect 390986 140378 391222 140614
rect 391306 140378 391542 140614
rect 390986 140058 391222 140294
rect 391306 140058 391542 140294
rect 390986 104378 391222 104614
rect 391306 104378 391542 104614
rect 390986 104058 391222 104294
rect 391306 104058 391542 104294
rect 390986 68378 391222 68614
rect 391306 68378 391542 68614
rect 390986 68058 391222 68294
rect 391306 68058 391542 68294
rect 390986 32378 391222 32614
rect 391306 32378 391542 32614
rect 390986 32058 391222 32294
rect 391306 32058 391542 32294
rect 372986 -6342 373222 -6106
rect 373306 -6342 373542 -6106
rect 372986 -6662 373222 -6426
rect 373306 -6662 373542 -6426
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 690938 401782 691174
rect 401866 690938 402102 691174
rect 401546 690618 401782 690854
rect 401866 690618 402102 690854
rect 401546 654938 401782 655174
rect 401866 654938 402102 655174
rect 401546 654618 401782 654854
rect 401866 654618 402102 654854
rect 401546 618938 401782 619174
rect 401866 618938 402102 619174
rect 401546 618618 401782 618854
rect 401866 618618 402102 618854
rect 401546 582938 401782 583174
rect 401866 582938 402102 583174
rect 401546 582618 401782 582854
rect 401866 582618 402102 582854
rect 401546 546938 401782 547174
rect 401866 546938 402102 547174
rect 401546 546618 401782 546854
rect 401866 546618 402102 546854
rect 401546 510938 401782 511174
rect 401866 510938 402102 511174
rect 401546 510618 401782 510854
rect 401866 510618 402102 510854
rect 401546 474938 401782 475174
rect 401866 474938 402102 475174
rect 401546 474618 401782 474854
rect 401866 474618 402102 474854
rect 401546 438938 401782 439174
rect 401866 438938 402102 439174
rect 401546 438618 401782 438854
rect 401866 438618 402102 438854
rect 401546 402938 401782 403174
rect 401866 402938 402102 403174
rect 401546 402618 401782 402854
rect 401866 402618 402102 402854
rect 401546 366938 401782 367174
rect 401866 366938 402102 367174
rect 401546 366618 401782 366854
rect 401866 366618 402102 366854
rect 401546 330938 401782 331174
rect 401866 330938 402102 331174
rect 401546 330618 401782 330854
rect 401866 330618 402102 330854
rect 401546 294938 401782 295174
rect 401866 294938 402102 295174
rect 401546 294618 401782 294854
rect 401866 294618 402102 294854
rect 401546 258938 401782 259174
rect 401866 258938 402102 259174
rect 401546 258618 401782 258854
rect 401866 258618 402102 258854
rect 401546 222938 401782 223174
rect 401866 222938 402102 223174
rect 401546 222618 401782 222854
rect 401866 222618 402102 222854
rect 401546 186938 401782 187174
rect 401866 186938 402102 187174
rect 401546 186618 401782 186854
rect 401866 186618 402102 186854
rect 401546 150938 401782 151174
rect 401866 150938 402102 151174
rect 401546 150618 401782 150854
rect 401866 150618 402102 150854
rect 401546 114938 401782 115174
rect 401866 114938 402102 115174
rect 401546 114618 401782 114854
rect 401866 114618 402102 114854
rect 401546 78938 401782 79174
rect 401866 78938 402102 79174
rect 401546 78618 401782 78854
rect 401866 78618 402102 78854
rect 401546 42938 401782 43174
rect 401866 42938 402102 43174
rect 401546 42618 401782 42854
rect 401866 42618 402102 42854
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 401546 -2502 401782 -2266
rect 401866 -2502 402102 -2266
rect 401546 -2822 401782 -2586
rect 401866 -2822 402102 -2586
rect 405266 694658 405502 694894
rect 405586 694658 405822 694894
rect 405266 694338 405502 694574
rect 405586 694338 405822 694574
rect 405266 658658 405502 658894
rect 405586 658658 405822 658894
rect 405266 658338 405502 658574
rect 405586 658338 405822 658574
rect 405266 622658 405502 622894
rect 405586 622658 405822 622894
rect 405266 622338 405502 622574
rect 405586 622338 405822 622574
rect 405266 586658 405502 586894
rect 405586 586658 405822 586894
rect 405266 586338 405502 586574
rect 405586 586338 405822 586574
rect 405266 550658 405502 550894
rect 405586 550658 405822 550894
rect 405266 550338 405502 550574
rect 405586 550338 405822 550574
rect 405266 514658 405502 514894
rect 405586 514658 405822 514894
rect 405266 514338 405502 514574
rect 405586 514338 405822 514574
rect 405266 478658 405502 478894
rect 405586 478658 405822 478894
rect 405266 478338 405502 478574
rect 405586 478338 405822 478574
rect 405266 442658 405502 442894
rect 405586 442658 405822 442894
rect 405266 442338 405502 442574
rect 405586 442338 405822 442574
rect 405266 406658 405502 406894
rect 405586 406658 405822 406894
rect 405266 406338 405502 406574
rect 405586 406338 405822 406574
rect 405266 370658 405502 370894
rect 405586 370658 405822 370894
rect 405266 370338 405502 370574
rect 405586 370338 405822 370574
rect 405266 334658 405502 334894
rect 405586 334658 405822 334894
rect 405266 334338 405502 334574
rect 405586 334338 405822 334574
rect 405266 298658 405502 298894
rect 405586 298658 405822 298894
rect 405266 298338 405502 298574
rect 405586 298338 405822 298574
rect 405266 262658 405502 262894
rect 405586 262658 405822 262894
rect 405266 262338 405502 262574
rect 405586 262338 405822 262574
rect 405266 226658 405502 226894
rect 405586 226658 405822 226894
rect 405266 226338 405502 226574
rect 405586 226338 405822 226574
rect 405266 190658 405502 190894
rect 405586 190658 405822 190894
rect 405266 190338 405502 190574
rect 405586 190338 405822 190574
rect 405266 154658 405502 154894
rect 405586 154658 405822 154894
rect 405266 154338 405502 154574
rect 405586 154338 405822 154574
rect 405266 118658 405502 118894
rect 405586 118658 405822 118894
rect 405266 118338 405502 118574
rect 405586 118338 405822 118574
rect 405266 82658 405502 82894
rect 405586 82658 405822 82894
rect 405266 82338 405502 82574
rect 405586 82338 405822 82574
rect 405266 46658 405502 46894
rect 405586 46658 405822 46894
rect 405266 46338 405502 46574
rect 405586 46338 405822 46574
rect 405266 10658 405502 10894
rect 405586 10658 405822 10894
rect 405266 10338 405502 10574
rect 405586 10338 405822 10574
rect 405266 -4422 405502 -4186
rect 405586 -4422 405822 -4186
rect 405266 -4742 405502 -4506
rect 405586 -4742 405822 -4506
rect 426986 711322 427222 711558
rect 427306 711322 427542 711558
rect 426986 711002 427222 711238
rect 427306 711002 427542 711238
rect 423266 709402 423502 709638
rect 423586 709402 423822 709638
rect 423266 709082 423502 709318
rect 423586 709082 423822 709318
rect 419546 707482 419782 707718
rect 419866 707482 420102 707718
rect 419546 707162 419782 707398
rect 419866 707162 420102 707398
rect 408986 698378 409222 698614
rect 409306 698378 409542 698614
rect 408986 698058 409222 698294
rect 409306 698058 409542 698294
rect 408986 662378 409222 662614
rect 409306 662378 409542 662614
rect 408986 662058 409222 662294
rect 409306 662058 409542 662294
rect 408986 626378 409222 626614
rect 409306 626378 409542 626614
rect 408986 626058 409222 626294
rect 409306 626058 409542 626294
rect 408986 590378 409222 590614
rect 409306 590378 409542 590614
rect 408986 590058 409222 590294
rect 409306 590058 409542 590294
rect 408986 554378 409222 554614
rect 409306 554378 409542 554614
rect 408986 554058 409222 554294
rect 409306 554058 409542 554294
rect 408986 518378 409222 518614
rect 409306 518378 409542 518614
rect 408986 518058 409222 518294
rect 409306 518058 409542 518294
rect 408986 482378 409222 482614
rect 409306 482378 409542 482614
rect 408986 482058 409222 482294
rect 409306 482058 409542 482294
rect 408986 446378 409222 446614
rect 409306 446378 409542 446614
rect 408986 446058 409222 446294
rect 409306 446058 409542 446294
rect 408986 410378 409222 410614
rect 409306 410378 409542 410614
rect 408986 410058 409222 410294
rect 409306 410058 409542 410294
rect 408986 374378 409222 374614
rect 409306 374378 409542 374614
rect 408986 374058 409222 374294
rect 409306 374058 409542 374294
rect 408986 338378 409222 338614
rect 409306 338378 409542 338614
rect 408986 338058 409222 338294
rect 409306 338058 409542 338294
rect 408986 302378 409222 302614
rect 409306 302378 409542 302614
rect 408986 302058 409222 302294
rect 409306 302058 409542 302294
rect 408986 266378 409222 266614
rect 409306 266378 409542 266614
rect 408986 266058 409222 266294
rect 409306 266058 409542 266294
rect 408986 230378 409222 230614
rect 409306 230378 409542 230614
rect 408986 230058 409222 230294
rect 409306 230058 409542 230294
rect 408986 194378 409222 194614
rect 409306 194378 409542 194614
rect 408986 194058 409222 194294
rect 409306 194058 409542 194294
rect 408986 158378 409222 158614
rect 409306 158378 409542 158614
rect 408986 158058 409222 158294
rect 409306 158058 409542 158294
rect 408986 122378 409222 122614
rect 409306 122378 409542 122614
rect 408986 122058 409222 122294
rect 409306 122058 409542 122294
rect 408986 86378 409222 86614
rect 409306 86378 409542 86614
rect 408986 86058 409222 86294
rect 409306 86058 409542 86294
rect 408986 50378 409222 50614
rect 409306 50378 409542 50614
rect 408986 50058 409222 50294
rect 409306 50058 409542 50294
rect 408986 14378 409222 14614
rect 409306 14378 409542 14614
rect 408986 14058 409222 14294
rect 409306 14058 409542 14294
rect 390986 -7302 391222 -7066
rect 391306 -7302 391542 -7066
rect 390986 -7622 391222 -7386
rect 391306 -7622 391542 -7386
rect 415826 705562 416062 705798
rect 416146 705562 416382 705798
rect 415826 705242 416062 705478
rect 416146 705242 416382 705478
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 415826 561218 416062 561454
rect 416146 561218 416382 561454
rect 415826 560898 416062 561134
rect 416146 560898 416382 561134
rect 415826 525218 416062 525454
rect 416146 525218 416382 525454
rect 415826 524898 416062 525134
rect 416146 524898 416382 525134
rect 415826 489218 416062 489454
rect 416146 489218 416382 489454
rect 415826 488898 416062 489134
rect 416146 488898 416382 489134
rect 415826 453218 416062 453454
rect 416146 453218 416382 453454
rect 415826 452898 416062 453134
rect 416146 452898 416382 453134
rect 415826 417218 416062 417454
rect 416146 417218 416382 417454
rect 415826 416898 416062 417134
rect 416146 416898 416382 417134
rect 415826 381218 416062 381454
rect 416146 381218 416382 381454
rect 415826 380898 416062 381134
rect 416146 380898 416382 381134
rect 415826 345218 416062 345454
rect 416146 345218 416382 345454
rect 415826 344898 416062 345134
rect 416146 344898 416382 345134
rect 415826 309218 416062 309454
rect 416146 309218 416382 309454
rect 415826 308898 416062 309134
rect 416146 308898 416382 309134
rect 415826 273218 416062 273454
rect 416146 273218 416382 273454
rect 415826 272898 416062 273134
rect 416146 272898 416382 273134
rect 415826 237218 416062 237454
rect 416146 237218 416382 237454
rect 415826 236898 416062 237134
rect 416146 236898 416382 237134
rect 415826 201218 416062 201454
rect 416146 201218 416382 201454
rect 415826 200898 416062 201134
rect 416146 200898 416382 201134
rect 415826 165218 416062 165454
rect 416146 165218 416382 165454
rect 415826 164898 416062 165134
rect 416146 164898 416382 165134
rect 415826 129218 416062 129454
rect 416146 129218 416382 129454
rect 415826 128898 416062 129134
rect 416146 128898 416382 129134
rect 415826 93218 416062 93454
rect 416146 93218 416382 93454
rect 415826 92898 416062 93134
rect 416146 92898 416382 93134
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -1542 416062 -1306
rect 416146 -1542 416382 -1306
rect 415826 -1862 416062 -1626
rect 416146 -1862 416382 -1626
rect 419546 672938 419782 673174
rect 419866 672938 420102 673174
rect 419546 672618 419782 672854
rect 419866 672618 420102 672854
rect 419546 636938 419782 637174
rect 419866 636938 420102 637174
rect 419546 636618 419782 636854
rect 419866 636618 420102 636854
rect 419546 600938 419782 601174
rect 419866 600938 420102 601174
rect 419546 600618 419782 600854
rect 419866 600618 420102 600854
rect 419546 564938 419782 565174
rect 419866 564938 420102 565174
rect 419546 564618 419782 564854
rect 419866 564618 420102 564854
rect 419546 528938 419782 529174
rect 419866 528938 420102 529174
rect 419546 528618 419782 528854
rect 419866 528618 420102 528854
rect 419546 492938 419782 493174
rect 419866 492938 420102 493174
rect 419546 492618 419782 492854
rect 419866 492618 420102 492854
rect 419546 456938 419782 457174
rect 419866 456938 420102 457174
rect 419546 456618 419782 456854
rect 419866 456618 420102 456854
rect 419546 420938 419782 421174
rect 419866 420938 420102 421174
rect 419546 420618 419782 420854
rect 419866 420618 420102 420854
rect 419546 384938 419782 385174
rect 419866 384938 420102 385174
rect 419546 384618 419782 384854
rect 419866 384618 420102 384854
rect 419546 348938 419782 349174
rect 419866 348938 420102 349174
rect 419546 348618 419782 348854
rect 419866 348618 420102 348854
rect 419546 312938 419782 313174
rect 419866 312938 420102 313174
rect 419546 312618 419782 312854
rect 419866 312618 420102 312854
rect 419546 276938 419782 277174
rect 419866 276938 420102 277174
rect 419546 276618 419782 276854
rect 419866 276618 420102 276854
rect 419546 240938 419782 241174
rect 419866 240938 420102 241174
rect 419546 240618 419782 240854
rect 419866 240618 420102 240854
rect 419546 204938 419782 205174
rect 419866 204938 420102 205174
rect 419546 204618 419782 204854
rect 419866 204618 420102 204854
rect 419546 168938 419782 169174
rect 419866 168938 420102 169174
rect 419546 168618 419782 168854
rect 419866 168618 420102 168854
rect 419546 132938 419782 133174
rect 419866 132938 420102 133174
rect 419546 132618 419782 132854
rect 419866 132618 420102 132854
rect 419546 96938 419782 97174
rect 419866 96938 420102 97174
rect 419546 96618 419782 96854
rect 419866 96618 420102 96854
rect 419546 60938 419782 61174
rect 419866 60938 420102 61174
rect 419546 60618 419782 60854
rect 419866 60618 420102 60854
rect 419546 24938 419782 25174
rect 419866 24938 420102 25174
rect 419546 24618 419782 24854
rect 419866 24618 420102 24854
rect 419546 -3462 419782 -3226
rect 419866 -3462 420102 -3226
rect 419546 -3782 419782 -3546
rect 419866 -3782 420102 -3546
rect 423266 676658 423502 676894
rect 423586 676658 423822 676894
rect 423266 676338 423502 676574
rect 423586 676338 423822 676574
rect 423266 640658 423502 640894
rect 423586 640658 423822 640894
rect 423266 640338 423502 640574
rect 423586 640338 423822 640574
rect 423266 604658 423502 604894
rect 423586 604658 423822 604894
rect 423266 604338 423502 604574
rect 423586 604338 423822 604574
rect 423266 568658 423502 568894
rect 423586 568658 423822 568894
rect 423266 568338 423502 568574
rect 423586 568338 423822 568574
rect 423266 532658 423502 532894
rect 423586 532658 423822 532894
rect 423266 532338 423502 532574
rect 423586 532338 423822 532574
rect 423266 496658 423502 496894
rect 423586 496658 423822 496894
rect 423266 496338 423502 496574
rect 423586 496338 423822 496574
rect 423266 460658 423502 460894
rect 423586 460658 423822 460894
rect 423266 460338 423502 460574
rect 423586 460338 423822 460574
rect 423266 424658 423502 424894
rect 423586 424658 423822 424894
rect 423266 424338 423502 424574
rect 423586 424338 423822 424574
rect 423266 388658 423502 388894
rect 423586 388658 423822 388894
rect 423266 388338 423502 388574
rect 423586 388338 423822 388574
rect 423266 352658 423502 352894
rect 423586 352658 423822 352894
rect 423266 352338 423502 352574
rect 423586 352338 423822 352574
rect 423266 316658 423502 316894
rect 423586 316658 423822 316894
rect 423266 316338 423502 316574
rect 423586 316338 423822 316574
rect 423266 280658 423502 280894
rect 423586 280658 423822 280894
rect 423266 280338 423502 280574
rect 423586 280338 423822 280574
rect 423266 244658 423502 244894
rect 423586 244658 423822 244894
rect 423266 244338 423502 244574
rect 423586 244338 423822 244574
rect 423266 208658 423502 208894
rect 423586 208658 423822 208894
rect 423266 208338 423502 208574
rect 423586 208338 423822 208574
rect 423266 172658 423502 172894
rect 423586 172658 423822 172894
rect 423266 172338 423502 172574
rect 423586 172338 423822 172574
rect 423266 136658 423502 136894
rect 423586 136658 423822 136894
rect 423266 136338 423502 136574
rect 423586 136338 423822 136574
rect 423266 100658 423502 100894
rect 423586 100658 423822 100894
rect 423266 100338 423502 100574
rect 423586 100338 423822 100574
rect 423266 64658 423502 64894
rect 423586 64658 423822 64894
rect 423266 64338 423502 64574
rect 423586 64338 423822 64574
rect 423266 28658 423502 28894
rect 423586 28658 423822 28894
rect 423266 28338 423502 28574
rect 423586 28338 423822 28574
rect 423266 -5382 423502 -5146
rect 423586 -5382 423822 -5146
rect 423266 -5702 423502 -5466
rect 423586 -5702 423822 -5466
rect 444986 710362 445222 710598
rect 445306 710362 445542 710598
rect 444986 710042 445222 710278
rect 445306 710042 445542 710278
rect 441266 708442 441502 708678
rect 441586 708442 441822 708678
rect 441266 708122 441502 708358
rect 441586 708122 441822 708358
rect 437546 706522 437782 706758
rect 437866 706522 438102 706758
rect 437546 706202 437782 706438
rect 437866 706202 438102 706438
rect 426986 680378 427222 680614
rect 427306 680378 427542 680614
rect 426986 680058 427222 680294
rect 427306 680058 427542 680294
rect 426986 644378 427222 644614
rect 427306 644378 427542 644614
rect 426986 644058 427222 644294
rect 427306 644058 427542 644294
rect 426986 608378 427222 608614
rect 427306 608378 427542 608614
rect 426986 608058 427222 608294
rect 427306 608058 427542 608294
rect 426986 572378 427222 572614
rect 427306 572378 427542 572614
rect 426986 572058 427222 572294
rect 427306 572058 427542 572294
rect 426986 536378 427222 536614
rect 427306 536378 427542 536614
rect 426986 536058 427222 536294
rect 427306 536058 427542 536294
rect 426986 500378 427222 500614
rect 427306 500378 427542 500614
rect 426986 500058 427222 500294
rect 427306 500058 427542 500294
rect 426986 464378 427222 464614
rect 427306 464378 427542 464614
rect 426986 464058 427222 464294
rect 427306 464058 427542 464294
rect 426986 428378 427222 428614
rect 427306 428378 427542 428614
rect 426986 428058 427222 428294
rect 427306 428058 427542 428294
rect 426986 392378 427222 392614
rect 427306 392378 427542 392614
rect 426986 392058 427222 392294
rect 427306 392058 427542 392294
rect 426986 356378 427222 356614
rect 427306 356378 427542 356614
rect 426986 356058 427222 356294
rect 427306 356058 427542 356294
rect 426986 320378 427222 320614
rect 427306 320378 427542 320614
rect 426986 320058 427222 320294
rect 427306 320058 427542 320294
rect 426986 284378 427222 284614
rect 427306 284378 427542 284614
rect 426986 284058 427222 284294
rect 427306 284058 427542 284294
rect 426986 248378 427222 248614
rect 427306 248378 427542 248614
rect 426986 248058 427222 248294
rect 427306 248058 427542 248294
rect 426986 212378 427222 212614
rect 427306 212378 427542 212614
rect 426986 212058 427222 212294
rect 427306 212058 427542 212294
rect 426986 176378 427222 176614
rect 427306 176378 427542 176614
rect 426986 176058 427222 176294
rect 427306 176058 427542 176294
rect 426986 140378 427222 140614
rect 427306 140378 427542 140614
rect 426986 140058 427222 140294
rect 427306 140058 427542 140294
rect 426986 104378 427222 104614
rect 427306 104378 427542 104614
rect 426986 104058 427222 104294
rect 427306 104058 427542 104294
rect 426986 68378 427222 68614
rect 427306 68378 427542 68614
rect 426986 68058 427222 68294
rect 427306 68058 427542 68294
rect 426986 32378 427222 32614
rect 427306 32378 427542 32614
rect 426986 32058 427222 32294
rect 427306 32058 427542 32294
rect 408986 -6342 409222 -6106
rect 409306 -6342 409542 -6106
rect 408986 -6662 409222 -6426
rect 409306 -6662 409542 -6426
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 433826 435218 434062 435454
rect 434146 435218 434382 435454
rect 433826 434898 434062 435134
rect 434146 434898 434382 435134
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 437546 690938 437782 691174
rect 437866 690938 438102 691174
rect 437546 690618 437782 690854
rect 437866 690618 438102 690854
rect 437546 654938 437782 655174
rect 437866 654938 438102 655174
rect 437546 654618 437782 654854
rect 437866 654618 438102 654854
rect 437546 618938 437782 619174
rect 437866 618938 438102 619174
rect 437546 618618 437782 618854
rect 437866 618618 438102 618854
rect 437546 582938 437782 583174
rect 437866 582938 438102 583174
rect 437546 582618 437782 582854
rect 437866 582618 438102 582854
rect 437546 546938 437782 547174
rect 437866 546938 438102 547174
rect 437546 546618 437782 546854
rect 437866 546618 438102 546854
rect 437546 510938 437782 511174
rect 437866 510938 438102 511174
rect 437546 510618 437782 510854
rect 437866 510618 438102 510854
rect 437546 474938 437782 475174
rect 437866 474938 438102 475174
rect 437546 474618 437782 474854
rect 437866 474618 438102 474854
rect 437546 438938 437782 439174
rect 437866 438938 438102 439174
rect 437546 438618 437782 438854
rect 437866 438618 438102 438854
rect 437546 402938 437782 403174
rect 437866 402938 438102 403174
rect 437546 402618 437782 402854
rect 437866 402618 438102 402854
rect 437546 366938 437782 367174
rect 437866 366938 438102 367174
rect 437546 366618 437782 366854
rect 437866 366618 438102 366854
rect 437546 330938 437782 331174
rect 437866 330938 438102 331174
rect 437546 330618 437782 330854
rect 437866 330618 438102 330854
rect 437546 294938 437782 295174
rect 437866 294938 438102 295174
rect 437546 294618 437782 294854
rect 437866 294618 438102 294854
rect 437546 258938 437782 259174
rect 437866 258938 438102 259174
rect 437546 258618 437782 258854
rect 437866 258618 438102 258854
rect 437546 222938 437782 223174
rect 437866 222938 438102 223174
rect 437546 222618 437782 222854
rect 437866 222618 438102 222854
rect 437546 186938 437782 187174
rect 437866 186938 438102 187174
rect 437546 186618 437782 186854
rect 437866 186618 438102 186854
rect 437546 150938 437782 151174
rect 437866 150938 438102 151174
rect 437546 150618 437782 150854
rect 437866 150618 438102 150854
rect 437546 114938 437782 115174
rect 437866 114938 438102 115174
rect 437546 114618 437782 114854
rect 437866 114618 438102 114854
rect 437546 78938 437782 79174
rect 437866 78938 438102 79174
rect 437546 78618 437782 78854
rect 437866 78618 438102 78854
rect 437546 42938 437782 43174
rect 437866 42938 438102 43174
rect 437546 42618 437782 42854
rect 437866 42618 438102 42854
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 437546 -2502 437782 -2266
rect 437866 -2502 438102 -2266
rect 437546 -2822 437782 -2586
rect 437866 -2822 438102 -2586
rect 441266 694658 441502 694894
rect 441586 694658 441822 694894
rect 441266 694338 441502 694574
rect 441586 694338 441822 694574
rect 441266 658658 441502 658894
rect 441586 658658 441822 658894
rect 441266 658338 441502 658574
rect 441586 658338 441822 658574
rect 441266 622658 441502 622894
rect 441586 622658 441822 622894
rect 441266 622338 441502 622574
rect 441586 622338 441822 622574
rect 441266 586658 441502 586894
rect 441586 586658 441822 586894
rect 441266 586338 441502 586574
rect 441586 586338 441822 586574
rect 441266 550658 441502 550894
rect 441586 550658 441822 550894
rect 441266 550338 441502 550574
rect 441586 550338 441822 550574
rect 441266 514658 441502 514894
rect 441586 514658 441822 514894
rect 441266 514338 441502 514574
rect 441586 514338 441822 514574
rect 441266 478658 441502 478894
rect 441586 478658 441822 478894
rect 441266 478338 441502 478574
rect 441586 478338 441822 478574
rect 441266 442658 441502 442894
rect 441586 442658 441822 442894
rect 441266 442338 441502 442574
rect 441586 442338 441822 442574
rect 441266 406658 441502 406894
rect 441586 406658 441822 406894
rect 441266 406338 441502 406574
rect 441586 406338 441822 406574
rect 441266 370658 441502 370894
rect 441586 370658 441822 370894
rect 441266 370338 441502 370574
rect 441586 370338 441822 370574
rect 441266 334658 441502 334894
rect 441586 334658 441822 334894
rect 441266 334338 441502 334574
rect 441586 334338 441822 334574
rect 441266 298658 441502 298894
rect 441586 298658 441822 298894
rect 441266 298338 441502 298574
rect 441586 298338 441822 298574
rect 441266 262658 441502 262894
rect 441586 262658 441822 262894
rect 441266 262338 441502 262574
rect 441586 262338 441822 262574
rect 441266 226658 441502 226894
rect 441586 226658 441822 226894
rect 441266 226338 441502 226574
rect 441586 226338 441822 226574
rect 441266 190658 441502 190894
rect 441586 190658 441822 190894
rect 441266 190338 441502 190574
rect 441586 190338 441822 190574
rect 441266 154658 441502 154894
rect 441586 154658 441822 154894
rect 441266 154338 441502 154574
rect 441586 154338 441822 154574
rect 441266 118658 441502 118894
rect 441586 118658 441822 118894
rect 441266 118338 441502 118574
rect 441586 118338 441822 118574
rect 441266 82658 441502 82894
rect 441586 82658 441822 82894
rect 441266 82338 441502 82574
rect 441586 82338 441822 82574
rect 441266 46658 441502 46894
rect 441586 46658 441822 46894
rect 441266 46338 441502 46574
rect 441586 46338 441822 46574
rect 441266 10658 441502 10894
rect 441586 10658 441822 10894
rect 441266 10338 441502 10574
rect 441586 10338 441822 10574
rect 441266 -4422 441502 -4186
rect 441586 -4422 441822 -4186
rect 441266 -4742 441502 -4506
rect 441586 -4742 441822 -4506
rect 462986 711322 463222 711558
rect 463306 711322 463542 711558
rect 462986 711002 463222 711238
rect 463306 711002 463542 711238
rect 459266 709402 459502 709638
rect 459586 709402 459822 709638
rect 459266 709082 459502 709318
rect 459586 709082 459822 709318
rect 455546 707482 455782 707718
rect 455866 707482 456102 707718
rect 455546 707162 455782 707398
rect 455866 707162 456102 707398
rect 444986 698378 445222 698614
rect 445306 698378 445542 698614
rect 444986 698058 445222 698294
rect 445306 698058 445542 698294
rect 444986 662378 445222 662614
rect 445306 662378 445542 662614
rect 444986 662058 445222 662294
rect 445306 662058 445542 662294
rect 444986 626378 445222 626614
rect 445306 626378 445542 626614
rect 444986 626058 445222 626294
rect 445306 626058 445542 626294
rect 444986 590378 445222 590614
rect 445306 590378 445542 590614
rect 444986 590058 445222 590294
rect 445306 590058 445542 590294
rect 444986 554378 445222 554614
rect 445306 554378 445542 554614
rect 444986 554058 445222 554294
rect 445306 554058 445542 554294
rect 444986 518378 445222 518614
rect 445306 518378 445542 518614
rect 444986 518058 445222 518294
rect 445306 518058 445542 518294
rect 444986 482378 445222 482614
rect 445306 482378 445542 482614
rect 444986 482058 445222 482294
rect 445306 482058 445542 482294
rect 444986 446378 445222 446614
rect 445306 446378 445542 446614
rect 444986 446058 445222 446294
rect 445306 446058 445542 446294
rect 444986 410378 445222 410614
rect 445306 410378 445542 410614
rect 444986 410058 445222 410294
rect 445306 410058 445542 410294
rect 444986 374378 445222 374614
rect 445306 374378 445542 374614
rect 444986 374058 445222 374294
rect 445306 374058 445542 374294
rect 444986 338378 445222 338614
rect 445306 338378 445542 338614
rect 444986 338058 445222 338294
rect 445306 338058 445542 338294
rect 444986 302378 445222 302614
rect 445306 302378 445542 302614
rect 444986 302058 445222 302294
rect 445306 302058 445542 302294
rect 444986 266378 445222 266614
rect 445306 266378 445542 266614
rect 444986 266058 445222 266294
rect 445306 266058 445542 266294
rect 444986 230378 445222 230614
rect 445306 230378 445542 230614
rect 444986 230058 445222 230294
rect 445306 230058 445542 230294
rect 444986 194378 445222 194614
rect 445306 194378 445542 194614
rect 444986 194058 445222 194294
rect 445306 194058 445542 194294
rect 444986 158378 445222 158614
rect 445306 158378 445542 158614
rect 444986 158058 445222 158294
rect 445306 158058 445542 158294
rect 444986 122378 445222 122614
rect 445306 122378 445542 122614
rect 444986 122058 445222 122294
rect 445306 122058 445542 122294
rect 444986 86378 445222 86614
rect 445306 86378 445542 86614
rect 444986 86058 445222 86294
rect 445306 86058 445542 86294
rect 444986 50378 445222 50614
rect 445306 50378 445542 50614
rect 444986 50058 445222 50294
rect 445306 50058 445542 50294
rect 444986 14378 445222 14614
rect 445306 14378 445542 14614
rect 444986 14058 445222 14294
rect 445306 14058 445542 14294
rect 426986 -7302 427222 -7066
rect 427306 -7302 427542 -7066
rect 426986 -7622 427222 -7386
rect 427306 -7622 427542 -7386
rect 451826 705562 452062 705798
rect 452146 705562 452382 705798
rect 451826 705242 452062 705478
rect 452146 705242 452382 705478
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 451826 453218 452062 453454
rect 452146 453218 452382 453454
rect 451826 452898 452062 453134
rect 452146 452898 452382 453134
rect 451826 417218 452062 417454
rect 452146 417218 452382 417454
rect 451826 416898 452062 417134
rect 452146 416898 452382 417134
rect 451826 381218 452062 381454
rect 452146 381218 452382 381454
rect 451826 380898 452062 381134
rect 452146 380898 452382 381134
rect 451826 345218 452062 345454
rect 452146 345218 452382 345454
rect 451826 344898 452062 345134
rect 452146 344898 452382 345134
rect 451826 309218 452062 309454
rect 452146 309218 452382 309454
rect 451826 308898 452062 309134
rect 452146 308898 452382 309134
rect 451826 273218 452062 273454
rect 452146 273218 452382 273454
rect 451826 272898 452062 273134
rect 452146 272898 452382 273134
rect 451826 237218 452062 237454
rect 452146 237218 452382 237454
rect 451826 236898 452062 237134
rect 452146 236898 452382 237134
rect 451826 201218 452062 201454
rect 452146 201218 452382 201454
rect 451826 200898 452062 201134
rect 452146 200898 452382 201134
rect 451826 165218 452062 165454
rect 452146 165218 452382 165454
rect 451826 164898 452062 165134
rect 452146 164898 452382 165134
rect 451826 129218 452062 129454
rect 452146 129218 452382 129454
rect 451826 128898 452062 129134
rect 452146 128898 452382 129134
rect 451826 93218 452062 93454
rect 452146 93218 452382 93454
rect 451826 92898 452062 93134
rect 452146 92898 452382 93134
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -1542 452062 -1306
rect 452146 -1542 452382 -1306
rect 451826 -1862 452062 -1626
rect 452146 -1862 452382 -1626
rect 455546 672938 455782 673174
rect 455866 672938 456102 673174
rect 455546 672618 455782 672854
rect 455866 672618 456102 672854
rect 455546 636938 455782 637174
rect 455866 636938 456102 637174
rect 455546 636618 455782 636854
rect 455866 636618 456102 636854
rect 455546 600938 455782 601174
rect 455866 600938 456102 601174
rect 455546 600618 455782 600854
rect 455866 600618 456102 600854
rect 455546 564938 455782 565174
rect 455866 564938 456102 565174
rect 455546 564618 455782 564854
rect 455866 564618 456102 564854
rect 455546 528938 455782 529174
rect 455866 528938 456102 529174
rect 455546 528618 455782 528854
rect 455866 528618 456102 528854
rect 455546 492938 455782 493174
rect 455866 492938 456102 493174
rect 455546 492618 455782 492854
rect 455866 492618 456102 492854
rect 455546 456938 455782 457174
rect 455866 456938 456102 457174
rect 455546 456618 455782 456854
rect 455866 456618 456102 456854
rect 455546 420938 455782 421174
rect 455866 420938 456102 421174
rect 455546 420618 455782 420854
rect 455866 420618 456102 420854
rect 455546 384938 455782 385174
rect 455866 384938 456102 385174
rect 455546 384618 455782 384854
rect 455866 384618 456102 384854
rect 455546 348938 455782 349174
rect 455866 348938 456102 349174
rect 455546 348618 455782 348854
rect 455866 348618 456102 348854
rect 455546 312938 455782 313174
rect 455866 312938 456102 313174
rect 455546 312618 455782 312854
rect 455866 312618 456102 312854
rect 455546 276938 455782 277174
rect 455866 276938 456102 277174
rect 455546 276618 455782 276854
rect 455866 276618 456102 276854
rect 455546 240938 455782 241174
rect 455866 240938 456102 241174
rect 455546 240618 455782 240854
rect 455866 240618 456102 240854
rect 455546 204938 455782 205174
rect 455866 204938 456102 205174
rect 455546 204618 455782 204854
rect 455866 204618 456102 204854
rect 455546 168938 455782 169174
rect 455866 168938 456102 169174
rect 455546 168618 455782 168854
rect 455866 168618 456102 168854
rect 455546 132938 455782 133174
rect 455866 132938 456102 133174
rect 455546 132618 455782 132854
rect 455866 132618 456102 132854
rect 455546 96938 455782 97174
rect 455866 96938 456102 97174
rect 455546 96618 455782 96854
rect 455866 96618 456102 96854
rect 455546 60938 455782 61174
rect 455866 60938 456102 61174
rect 455546 60618 455782 60854
rect 455866 60618 456102 60854
rect 455546 24938 455782 25174
rect 455866 24938 456102 25174
rect 455546 24618 455782 24854
rect 455866 24618 456102 24854
rect 455546 -3462 455782 -3226
rect 455866 -3462 456102 -3226
rect 455546 -3782 455782 -3546
rect 455866 -3782 456102 -3546
rect 459266 676658 459502 676894
rect 459586 676658 459822 676894
rect 459266 676338 459502 676574
rect 459586 676338 459822 676574
rect 459266 640658 459502 640894
rect 459586 640658 459822 640894
rect 459266 640338 459502 640574
rect 459586 640338 459822 640574
rect 459266 604658 459502 604894
rect 459586 604658 459822 604894
rect 459266 604338 459502 604574
rect 459586 604338 459822 604574
rect 459266 568658 459502 568894
rect 459586 568658 459822 568894
rect 459266 568338 459502 568574
rect 459586 568338 459822 568574
rect 459266 532658 459502 532894
rect 459586 532658 459822 532894
rect 459266 532338 459502 532574
rect 459586 532338 459822 532574
rect 459266 496658 459502 496894
rect 459586 496658 459822 496894
rect 459266 496338 459502 496574
rect 459586 496338 459822 496574
rect 459266 460658 459502 460894
rect 459586 460658 459822 460894
rect 459266 460338 459502 460574
rect 459586 460338 459822 460574
rect 459266 424658 459502 424894
rect 459586 424658 459822 424894
rect 459266 424338 459502 424574
rect 459586 424338 459822 424574
rect 459266 388658 459502 388894
rect 459586 388658 459822 388894
rect 459266 388338 459502 388574
rect 459586 388338 459822 388574
rect 459266 352658 459502 352894
rect 459586 352658 459822 352894
rect 459266 352338 459502 352574
rect 459586 352338 459822 352574
rect 459266 316658 459502 316894
rect 459586 316658 459822 316894
rect 459266 316338 459502 316574
rect 459586 316338 459822 316574
rect 459266 280658 459502 280894
rect 459586 280658 459822 280894
rect 459266 280338 459502 280574
rect 459586 280338 459822 280574
rect 459266 244658 459502 244894
rect 459586 244658 459822 244894
rect 459266 244338 459502 244574
rect 459586 244338 459822 244574
rect 459266 208658 459502 208894
rect 459586 208658 459822 208894
rect 459266 208338 459502 208574
rect 459586 208338 459822 208574
rect 459266 172658 459502 172894
rect 459586 172658 459822 172894
rect 459266 172338 459502 172574
rect 459586 172338 459822 172574
rect 459266 136658 459502 136894
rect 459586 136658 459822 136894
rect 459266 136338 459502 136574
rect 459586 136338 459822 136574
rect 459266 100658 459502 100894
rect 459586 100658 459822 100894
rect 459266 100338 459502 100574
rect 459586 100338 459822 100574
rect 459266 64658 459502 64894
rect 459586 64658 459822 64894
rect 459266 64338 459502 64574
rect 459586 64338 459822 64574
rect 459266 28658 459502 28894
rect 459586 28658 459822 28894
rect 459266 28338 459502 28574
rect 459586 28338 459822 28574
rect 459266 -5382 459502 -5146
rect 459586 -5382 459822 -5146
rect 459266 -5702 459502 -5466
rect 459586 -5702 459822 -5466
rect 480986 710362 481222 710598
rect 481306 710362 481542 710598
rect 480986 710042 481222 710278
rect 481306 710042 481542 710278
rect 477266 708442 477502 708678
rect 477586 708442 477822 708678
rect 477266 708122 477502 708358
rect 477586 708122 477822 708358
rect 473546 706522 473782 706758
rect 473866 706522 474102 706758
rect 473546 706202 473782 706438
rect 473866 706202 474102 706438
rect 462986 680378 463222 680614
rect 463306 680378 463542 680614
rect 462986 680058 463222 680294
rect 463306 680058 463542 680294
rect 462986 644378 463222 644614
rect 463306 644378 463542 644614
rect 462986 644058 463222 644294
rect 463306 644058 463542 644294
rect 462986 608378 463222 608614
rect 463306 608378 463542 608614
rect 462986 608058 463222 608294
rect 463306 608058 463542 608294
rect 462986 572378 463222 572614
rect 463306 572378 463542 572614
rect 462986 572058 463222 572294
rect 463306 572058 463542 572294
rect 462986 536378 463222 536614
rect 463306 536378 463542 536614
rect 462986 536058 463222 536294
rect 463306 536058 463542 536294
rect 462986 500378 463222 500614
rect 463306 500378 463542 500614
rect 462986 500058 463222 500294
rect 463306 500058 463542 500294
rect 462986 464378 463222 464614
rect 463306 464378 463542 464614
rect 462986 464058 463222 464294
rect 463306 464058 463542 464294
rect 462986 428378 463222 428614
rect 463306 428378 463542 428614
rect 462986 428058 463222 428294
rect 463306 428058 463542 428294
rect 462986 392378 463222 392614
rect 463306 392378 463542 392614
rect 462986 392058 463222 392294
rect 463306 392058 463542 392294
rect 462986 356378 463222 356614
rect 463306 356378 463542 356614
rect 462986 356058 463222 356294
rect 463306 356058 463542 356294
rect 462986 320378 463222 320614
rect 463306 320378 463542 320614
rect 462986 320058 463222 320294
rect 463306 320058 463542 320294
rect 462986 284378 463222 284614
rect 463306 284378 463542 284614
rect 462986 284058 463222 284294
rect 463306 284058 463542 284294
rect 462986 248378 463222 248614
rect 463306 248378 463542 248614
rect 462986 248058 463222 248294
rect 463306 248058 463542 248294
rect 462986 212378 463222 212614
rect 463306 212378 463542 212614
rect 462986 212058 463222 212294
rect 463306 212058 463542 212294
rect 462986 176378 463222 176614
rect 463306 176378 463542 176614
rect 462986 176058 463222 176294
rect 463306 176058 463542 176294
rect 462986 140378 463222 140614
rect 463306 140378 463542 140614
rect 462986 140058 463222 140294
rect 463306 140058 463542 140294
rect 462986 104378 463222 104614
rect 463306 104378 463542 104614
rect 462986 104058 463222 104294
rect 463306 104058 463542 104294
rect 462986 68378 463222 68614
rect 463306 68378 463542 68614
rect 462986 68058 463222 68294
rect 463306 68058 463542 68294
rect 462986 32378 463222 32614
rect 463306 32378 463542 32614
rect 462986 32058 463222 32294
rect 463306 32058 463542 32294
rect 444986 -6342 445222 -6106
rect 445306 -6342 445542 -6106
rect 444986 -6662 445222 -6426
rect 445306 -6662 445542 -6426
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 690938 473782 691174
rect 473866 690938 474102 691174
rect 473546 690618 473782 690854
rect 473866 690618 474102 690854
rect 473546 654938 473782 655174
rect 473866 654938 474102 655174
rect 473546 654618 473782 654854
rect 473866 654618 474102 654854
rect 473546 618938 473782 619174
rect 473866 618938 474102 619174
rect 473546 618618 473782 618854
rect 473866 618618 474102 618854
rect 473546 582938 473782 583174
rect 473866 582938 474102 583174
rect 473546 582618 473782 582854
rect 473866 582618 474102 582854
rect 473546 546938 473782 547174
rect 473866 546938 474102 547174
rect 473546 546618 473782 546854
rect 473866 546618 474102 546854
rect 473546 510938 473782 511174
rect 473866 510938 474102 511174
rect 473546 510618 473782 510854
rect 473866 510618 474102 510854
rect 473546 474938 473782 475174
rect 473866 474938 474102 475174
rect 473546 474618 473782 474854
rect 473866 474618 474102 474854
rect 473546 438938 473782 439174
rect 473866 438938 474102 439174
rect 473546 438618 473782 438854
rect 473866 438618 474102 438854
rect 473546 402938 473782 403174
rect 473866 402938 474102 403174
rect 473546 402618 473782 402854
rect 473866 402618 474102 402854
rect 473546 366938 473782 367174
rect 473866 366938 474102 367174
rect 473546 366618 473782 366854
rect 473866 366618 474102 366854
rect 473546 330938 473782 331174
rect 473866 330938 474102 331174
rect 473546 330618 473782 330854
rect 473866 330618 474102 330854
rect 473546 294938 473782 295174
rect 473866 294938 474102 295174
rect 473546 294618 473782 294854
rect 473866 294618 474102 294854
rect 473546 258938 473782 259174
rect 473866 258938 474102 259174
rect 473546 258618 473782 258854
rect 473866 258618 474102 258854
rect 473546 222938 473782 223174
rect 473866 222938 474102 223174
rect 473546 222618 473782 222854
rect 473866 222618 474102 222854
rect 473546 186938 473782 187174
rect 473866 186938 474102 187174
rect 473546 186618 473782 186854
rect 473866 186618 474102 186854
rect 473546 150938 473782 151174
rect 473866 150938 474102 151174
rect 473546 150618 473782 150854
rect 473866 150618 474102 150854
rect 473546 114938 473782 115174
rect 473866 114938 474102 115174
rect 473546 114618 473782 114854
rect 473866 114618 474102 114854
rect 473546 78938 473782 79174
rect 473866 78938 474102 79174
rect 473546 78618 473782 78854
rect 473866 78618 474102 78854
rect 473546 42938 473782 43174
rect 473866 42938 474102 43174
rect 473546 42618 473782 42854
rect 473866 42618 474102 42854
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -2502 473782 -2266
rect 473866 -2502 474102 -2266
rect 473546 -2822 473782 -2586
rect 473866 -2822 474102 -2586
rect 477266 694658 477502 694894
rect 477586 694658 477822 694894
rect 477266 694338 477502 694574
rect 477586 694338 477822 694574
rect 477266 658658 477502 658894
rect 477586 658658 477822 658894
rect 477266 658338 477502 658574
rect 477586 658338 477822 658574
rect 477266 622658 477502 622894
rect 477586 622658 477822 622894
rect 477266 622338 477502 622574
rect 477586 622338 477822 622574
rect 477266 586658 477502 586894
rect 477586 586658 477822 586894
rect 477266 586338 477502 586574
rect 477586 586338 477822 586574
rect 477266 550658 477502 550894
rect 477586 550658 477822 550894
rect 477266 550338 477502 550574
rect 477586 550338 477822 550574
rect 477266 514658 477502 514894
rect 477586 514658 477822 514894
rect 477266 514338 477502 514574
rect 477586 514338 477822 514574
rect 477266 478658 477502 478894
rect 477586 478658 477822 478894
rect 477266 478338 477502 478574
rect 477586 478338 477822 478574
rect 477266 442658 477502 442894
rect 477586 442658 477822 442894
rect 477266 442338 477502 442574
rect 477586 442338 477822 442574
rect 477266 406658 477502 406894
rect 477586 406658 477822 406894
rect 477266 406338 477502 406574
rect 477586 406338 477822 406574
rect 477266 370658 477502 370894
rect 477586 370658 477822 370894
rect 477266 370338 477502 370574
rect 477586 370338 477822 370574
rect 477266 334658 477502 334894
rect 477586 334658 477822 334894
rect 477266 334338 477502 334574
rect 477586 334338 477822 334574
rect 477266 298658 477502 298894
rect 477586 298658 477822 298894
rect 477266 298338 477502 298574
rect 477586 298338 477822 298574
rect 477266 262658 477502 262894
rect 477586 262658 477822 262894
rect 477266 262338 477502 262574
rect 477586 262338 477822 262574
rect 477266 226658 477502 226894
rect 477586 226658 477822 226894
rect 477266 226338 477502 226574
rect 477586 226338 477822 226574
rect 477266 190658 477502 190894
rect 477586 190658 477822 190894
rect 477266 190338 477502 190574
rect 477586 190338 477822 190574
rect 477266 154658 477502 154894
rect 477586 154658 477822 154894
rect 477266 154338 477502 154574
rect 477586 154338 477822 154574
rect 477266 118658 477502 118894
rect 477586 118658 477822 118894
rect 477266 118338 477502 118574
rect 477586 118338 477822 118574
rect 477266 82658 477502 82894
rect 477586 82658 477822 82894
rect 477266 82338 477502 82574
rect 477586 82338 477822 82574
rect 477266 46658 477502 46894
rect 477586 46658 477822 46894
rect 477266 46338 477502 46574
rect 477586 46338 477822 46574
rect 477266 10658 477502 10894
rect 477586 10658 477822 10894
rect 477266 10338 477502 10574
rect 477586 10338 477822 10574
rect 477266 -4422 477502 -4186
rect 477586 -4422 477822 -4186
rect 477266 -4742 477502 -4506
rect 477586 -4742 477822 -4506
rect 498986 711322 499222 711558
rect 499306 711322 499542 711558
rect 498986 711002 499222 711238
rect 499306 711002 499542 711238
rect 495266 709402 495502 709638
rect 495586 709402 495822 709638
rect 495266 709082 495502 709318
rect 495586 709082 495822 709318
rect 491546 707482 491782 707718
rect 491866 707482 492102 707718
rect 491546 707162 491782 707398
rect 491866 707162 492102 707398
rect 480986 698378 481222 698614
rect 481306 698378 481542 698614
rect 480986 698058 481222 698294
rect 481306 698058 481542 698294
rect 480986 662378 481222 662614
rect 481306 662378 481542 662614
rect 480986 662058 481222 662294
rect 481306 662058 481542 662294
rect 480986 626378 481222 626614
rect 481306 626378 481542 626614
rect 480986 626058 481222 626294
rect 481306 626058 481542 626294
rect 480986 590378 481222 590614
rect 481306 590378 481542 590614
rect 480986 590058 481222 590294
rect 481306 590058 481542 590294
rect 480986 554378 481222 554614
rect 481306 554378 481542 554614
rect 480986 554058 481222 554294
rect 481306 554058 481542 554294
rect 480986 518378 481222 518614
rect 481306 518378 481542 518614
rect 480986 518058 481222 518294
rect 481306 518058 481542 518294
rect 480986 482378 481222 482614
rect 481306 482378 481542 482614
rect 480986 482058 481222 482294
rect 481306 482058 481542 482294
rect 480986 446378 481222 446614
rect 481306 446378 481542 446614
rect 480986 446058 481222 446294
rect 481306 446058 481542 446294
rect 480986 410378 481222 410614
rect 481306 410378 481542 410614
rect 480986 410058 481222 410294
rect 481306 410058 481542 410294
rect 480986 374378 481222 374614
rect 481306 374378 481542 374614
rect 480986 374058 481222 374294
rect 481306 374058 481542 374294
rect 480986 338378 481222 338614
rect 481306 338378 481542 338614
rect 480986 338058 481222 338294
rect 481306 338058 481542 338294
rect 480986 302378 481222 302614
rect 481306 302378 481542 302614
rect 480986 302058 481222 302294
rect 481306 302058 481542 302294
rect 480986 266378 481222 266614
rect 481306 266378 481542 266614
rect 480986 266058 481222 266294
rect 481306 266058 481542 266294
rect 480986 230378 481222 230614
rect 481306 230378 481542 230614
rect 480986 230058 481222 230294
rect 481306 230058 481542 230294
rect 480986 194378 481222 194614
rect 481306 194378 481542 194614
rect 480986 194058 481222 194294
rect 481306 194058 481542 194294
rect 480986 158378 481222 158614
rect 481306 158378 481542 158614
rect 480986 158058 481222 158294
rect 481306 158058 481542 158294
rect 480986 122378 481222 122614
rect 481306 122378 481542 122614
rect 480986 122058 481222 122294
rect 481306 122058 481542 122294
rect 480986 86378 481222 86614
rect 481306 86378 481542 86614
rect 480986 86058 481222 86294
rect 481306 86058 481542 86294
rect 480986 50378 481222 50614
rect 481306 50378 481542 50614
rect 480986 50058 481222 50294
rect 481306 50058 481542 50294
rect 480986 14378 481222 14614
rect 481306 14378 481542 14614
rect 480986 14058 481222 14294
rect 481306 14058 481542 14294
rect 462986 -7302 463222 -7066
rect 463306 -7302 463542 -7066
rect 462986 -7622 463222 -7386
rect 463306 -7622 463542 -7386
rect 487826 705562 488062 705798
rect 488146 705562 488382 705798
rect 487826 705242 488062 705478
rect 488146 705242 488382 705478
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 487826 453218 488062 453454
rect 488146 453218 488382 453454
rect 487826 452898 488062 453134
rect 488146 452898 488382 453134
rect 487826 417218 488062 417454
rect 488146 417218 488382 417454
rect 487826 416898 488062 417134
rect 488146 416898 488382 417134
rect 487826 381218 488062 381454
rect 488146 381218 488382 381454
rect 487826 380898 488062 381134
rect 488146 380898 488382 381134
rect 487826 345218 488062 345454
rect 488146 345218 488382 345454
rect 487826 344898 488062 345134
rect 488146 344898 488382 345134
rect 487826 309218 488062 309454
rect 488146 309218 488382 309454
rect 487826 308898 488062 309134
rect 488146 308898 488382 309134
rect 487826 273218 488062 273454
rect 488146 273218 488382 273454
rect 487826 272898 488062 273134
rect 488146 272898 488382 273134
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 487826 129218 488062 129454
rect 488146 129218 488382 129454
rect 487826 128898 488062 129134
rect 488146 128898 488382 129134
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -1542 488062 -1306
rect 488146 -1542 488382 -1306
rect 487826 -1862 488062 -1626
rect 488146 -1862 488382 -1626
rect 491546 672938 491782 673174
rect 491866 672938 492102 673174
rect 491546 672618 491782 672854
rect 491866 672618 492102 672854
rect 491546 636938 491782 637174
rect 491866 636938 492102 637174
rect 491546 636618 491782 636854
rect 491866 636618 492102 636854
rect 491546 600938 491782 601174
rect 491866 600938 492102 601174
rect 491546 600618 491782 600854
rect 491866 600618 492102 600854
rect 491546 564938 491782 565174
rect 491866 564938 492102 565174
rect 491546 564618 491782 564854
rect 491866 564618 492102 564854
rect 491546 528938 491782 529174
rect 491866 528938 492102 529174
rect 491546 528618 491782 528854
rect 491866 528618 492102 528854
rect 491546 492938 491782 493174
rect 491866 492938 492102 493174
rect 491546 492618 491782 492854
rect 491866 492618 492102 492854
rect 491546 456938 491782 457174
rect 491866 456938 492102 457174
rect 491546 456618 491782 456854
rect 491866 456618 492102 456854
rect 491546 420938 491782 421174
rect 491866 420938 492102 421174
rect 491546 420618 491782 420854
rect 491866 420618 492102 420854
rect 491546 384938 491782 385174
rect 491866 384938 492102 385174
rect 491546 384618 491782 384854
rect 491866 384618 492102 384854
rect 491546 348938 491782 349174
rect 491866 348938 492102 349174
rect 491546 348618 491782 348854
rect 491866 348618 492102 348854
rect 491546 312938 491782 313174
rect 491866 312938 492102 313174
rect 491546 312618 491782 312854
rect 491866 312618 492102 312854
rect 491546 276938 491782 277174
rect 491866 276938 492102 277174
rect 491546 276618 491782 276854
rect 491866 276618 492102 276854
rect 491546 240938 491782 241174
rect 491866 240938 492102 241174
rect 491546 240618 491782 240854
rect 491866 240618 492102 240854
rect 491546 204938 491782 205174
rect 491866 204938 492102 205174
rect 491546 204618 491782 204854
rect 491866 204618 492102 204854
rect 491546 168938 491782 169174
rect 491866 168938 492102 169174
rect 491546 168618 491782 168854
rect 491866 168618 492102 168854
rect 491546 132938 491782 133174
rect 491866 132938 492102 133174
rect 491546 132618 491782 132854
rect 491866 132618 492102 132854
rect 491546 96938 491782 97174
rect 491866 96938 492102 97174
rect 491546 96618 491782 96854
rect 491866 96618 492102 96854
rect 491546 60938 491782 61174
rect 491866 60938 492102 61174
rect 491546 60618 491782 60854
rect 491866 60618 492102 60854
rect 491546 24938 491782 25174
rect 491866 24938 492102 25174
rect 491546 24618 491782 24854
rect 491866 24618 492102 24854
rect 491546 -3462 491782 -3226
rect 491866 -3462 492102 -3226
rect 491546 -3782 491782 -3546
rect 491866 -3782 492102 -3546
rect 495266 676658 495502 676894
rect 495586 676658 495822 676894
rect 495266 676338 495502 676574
rect 495586 676338 495822 676574
rect 495266 640658 495502 640894
rect 495586 640658 495822 640894
rect 495266 640338 495502 640574
rect 495586 640338 495822 640574
rect 495266 604658 495502 604894
rect 495586 604658 495822 604894
rect 495266 604338 495502 604574
rect 495586 604338 495822 604574
rect 495266 568658 495502 568894
rect 495586 568658 495822 568894
rect 495266 568338 495502 568574
rect 495586 568338 495822 568574
rect 495266 532658 495502 532894
rect 495586 532658 495822 532894
rect 495266 532338 495502 532574
rect 495586 532338 495822 532574
rect 495266 496658 495502 496894
rect 495586 496658 495822 496894
rect 495266 496338 495502 496574
rect 495586 496338 495822 496574
rect 495266 460658 495502 460894
rect 495586 460658 495822 460894
rect 495266 460338 495502 460574
rect 495586 460338 495822 460574
rect 495266 424658 495502 424894
rect 495586 424658 495822 424894
rect 495266 424338 495502 424574
rect 495586 424338 495822 424574
rect 495266 388658 495502 388894
rect 495586 388658 495822 388894
rect 495266 388338 495502 388574
rect 495586 388338 495822 388574
rect 495266 352658 495502 352894
rect 495586 352658 495822 352894
rect 495266 352338 495502 352574
rect 495586 352338 495822 352574
rect 495266 316658 495502 316894
rect 495586 316658 495822 316894
rect 495266 316338 495502 316574
rect 495586 316338 495822 316574
rect 495266 280658 495502 280894
rect 495586 280658 495822 280894
rect 495266 280338 495502 280574
rect 495586 280338 495822 280574
rect 495266 244658 495502 244894
rect 495586 244658 495822 244894
rect 495266 244338 495502 244574
rect 495586 244338 495822 244574
rect 495266 208658 495502 208894
rect 495586 208658 495822 208894
rect 495266 208338 495502 208574
rect 495586 208338 495822 208574
rect 495266 172658 495502 172894
rect 495586 172658 495822 172894
rect 495266 172338 495502 172574
rect 495586 172338 495822 172574
rect 495266 136658 495502 136894
rect 495586 136658 495822 136894
rect 495266 136338 495502 136574
rect 495586 136338 495822 136574
rect 495266 100658 495502 100894
rect 495586 100658 495822 100894
rect 495266 100338 495502 100574
rect 495586 100338 495822 100574
rect 495266 64658 495502 64894
rect 495586 64658 495822 64894
rect 495266 64338 495502 64574
rect 495586 64338 495822 64574
rect 495266 28658 495502 28894
rect 495586 28658 495822 28894
rect 495266 28338 495502 28574
rect 495586 28338 495822 28574
rect 495266 -5382 495502 -5146
rect 495586 -5382 495822 -5146
rect 495266 -5702 495502 -5466
rect 495586 -5702 495822 -5466
rect 516986 710362 517222 710598
rect 517306 710362 517542 710598
rect 516986 710042 517222 710278
rect 517306 710042 517542 710278
rect 513266 708442 513502 708678
rect 513586 708442 513822 708678
rect 513266 708122 513502 708358
rect 513586 708122 513822 708358
rect 509546 706522 509782 706758
rect 509866 706522 510102 706758
rect 509546 706202 509782 706438
rect 509866 706202 510102 706438
rect 498986 680378 499222 680614
rect 499306 680378 499542 680614
rect 498986 680058 499222 680294
rect 499306 680058 499542 680294
rect 498986 644378 499222 644614
rect 499306 644378 499542 644614
rect 498986 644058 499222 644294
rect 499306 644058 499542 644294
rect 498986 608378 499222 608614
rect 499306 608378 499542 608614
rect 498986 608058 499222 608294
rect 499306 608058 499542 608294
rect 498986 572378 499222 572614
rect 499306 572378 499542 572614
rect 498986 572058 499222 572294
rect 499306 572058 499542 572294
rect 498986 536378 499222 536614
rect 499306 536378 499542 536614
rect 498986 536058 499222 536294
rect 499306 536058 499542 536294
rect 498986 500378 499222 500614
rect 499306 500378 499542 500614
rect 498986 500058 499222 500294
rect 499306 500058 499542 500294
rect 498986 464378 499222 464614
rect 499306 464378 499542 464614
rect 498986 464058 499222 464294
rect 499306 464058 499542 464294
rect 498986 428378 499222 428614
rect 499306 428378 499542 428614
rect 498986 428058 499222 428294
rect 499306 428058 499542 428294
rect 498986 392378 499222 392614
rect 499306 392378 499542 392614
rect 498986 392058 499222 392294
rect 499306 392058 499542 392294
rect 498986 356378 499222 356614
rect 499306 356378 499542 356614
rect 498986 356058 499222 356294
rect 499306 356058 499542 356294
rect 498986 320378 499222 320614
rect 499306 320378 499542 320614
rect 498986 320058 499222 320294
rect 499306 320058 499542 320294
rect 498986 284378 499222 284614
rect 499306 284378 499542 284614
rect 498986 284058 499222 284294
rect 499306 284058 499542 284294
rect 498986 248378 499222 248614
rect 499306 248378 499542 248614
rect 498986 248058 499222 248294
rect 499306 248058 499542 248294
rect 498986 212378 499222 212614
rect 499306 212378 499542 212614
rect 498986 212058 499222 212294
rect 499306 212058 499542 212294
rect 498986 176378 499222 176614
rect 499306 176378 499542 176614
rect 498986 176058 499222 176294
rect 499306 176058 499542 176294
rect 498986 140378 499222 140614
rect 499306 140378 499542 140614
rect 498986 140058 499222 140294
rect 499306 140058 499542 140294
rect 498986 104378 499222 104614
rect 499306 104378 499542 104614
rect 498986 104058 499222 104294
rect 499306 104058 499542 104294
rect 498986 68378 499222 68614
rect 499306 68378 499542 68614
rect 498986 68058 499222 68294
rect 499306 68058 499542 68294
rect 498986 32378 499222 32614
rect 499306 32378 499542 32614
rect 498986 32058 499222 32294
rect 499306 32058 499542 32294
rect 480986 -6342 481222 -6106
rect 481306 -6342 481542 -6106
rect 480986 -6662 481222 -6426
rect 481306 -6662 481542 -6426
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 690938 509782 691174
rect 509866 690938 510102 691174
rect 509546 690618 509782 690854
rect 509866 690618 510102 690854
rect 509546 654938 509782 655174
rect 509866 654938 510102 655174
rect 509546 654618 509782 654854
rect 509866 654618 510102 654854
rect 509546 618938 509782 619174
rect 509866 618938 510102 619174
rect 509546 618618 509782 618854
rect 509866 618618 510102 618854
rect 509546 582938 509782 583174
rect 509866 582938 510102 583174
rect 509546 582618 509782 582854
rect 509866 582618 510102 582854
rect 509546 546938 509782 547174
rect 509866 546938 510102 547174
rect 509546 546618 509782 546854
rect 509866 546618 510102 546854
rect 509546 510938 509782 511174
rect 509866 510938 510102 511174
rect 509546 510618 509782 510854
rect 509866 510618 510102 510854
rect 509546 474938 509782 475174
rect 509866 474938 510102 475174
rect 509546 474618 509782 474854
rect 509866 474618 510102 474854
rect 509546 438938 509782 439174
rect 509866 438938 510102 439174
rect 509546 438618 509782 438854
rect 509866 438618 510102 438854
rect 509546 402938 509782 403174
rect 509866 402938 510102 403174
rect 509546 402618 509782 402854
rect 509866 402618 510102 402854
rect 509546 366938 509782 367174
rect 509866 366938 510102 367174
rect 509546 366618 509782 366854
rect 509866 366618 510102 366854
rect 509546 330938 509782 331174
rect 509866 330938 510102 331174
rect 509546 330618 509782 330854
rect 509866 330618 510102 330854
rect 509546 294938 509782 295174
rect 509866 294938 510102 295174
rect 509546 294618 509782 294854
rect 509866 294618 510102 294854
rect 509546 258938 509782 259174
rect 509866 258938 510102 259174
rect 509546 258618 509782 258854
rect 509866 258618 510102 258854
rect 509546 222938 509782 223174
rect 509866 222938 510102 223174
rect 509546 222618 509782 222854
rect 509866 222618 510102 222854
rect 509546 186938 509782 187174
rect 509866 186938 510102 187174
rect 509546 186618 509782 186854
rect 509866 186618 510102 186854
rect 509546 150938 509782 151174
rect 509866 150938 510102 151174
rect 509546 150618 509782 150854
rect 509866 150618 510102 150854
rect 509546 114938 509782 115174
rect 509866 114938 510102 115174
rect 509546 114618 509782 114854
rect 509866 114618 510102 114854
rect 509546 78938 509782 79174
rect 509866 78938 510102 79174
rect 509546 78618 509782 78854
rect 509866 78618 510102 78854
rect 509546 42938 509782 43174
rect 509866 42938 510102 43174
rect 509546 42618 509782 42854
rect 509866 42618 510102 42854
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -2502 509782 -2266
rect 509866 -2502 510102 -2266
rect 509546 -2822 509782 -2586
rect 509866 -2822 510102 -2586
rect 513266 694658 513502 694894
rect 513586 694658 513822 694894
rect 513266 694338 513502 694574
rect 513586 694338 513822 694574
rect 513266 658658 513502 658894
rect 513586 658658 513822 658894
rect 513266 658338 513502 658574
rect 513586 658338 513822 658574
rect 513266 622658 513502 622894
rect 513586 622658 513822 622894
rect 513266 622338 513502 622574
rect 513586 622338 513822 622574
rect 513266 586658 513502 586894
rect 513586 586658 513822 586894
rect 513266 586338 513502 586574
rect 513586 586338 513822 586574
rect 513266 550658 513502 550894
rect 513586 550658 513822 550894
rect 513266 550338 513502 550574
rect 513586 550338 513822 550574
rect 513266 514658 513502 514894
rect 513586 514658 513822 514894
rect 513266 514338 513502 514574
rect 513586 514338 513822 514574
rect 513266 478658 513502 478894
rect 513586 478658 513822 478894
rect 513266 478338 513502 478574
rect 513586 478338 513822 478574
rect 513266 442658 513502 442894
rect 513586 442658 513822 442894
rect 513266 442338 513502 442574
rect 513586 442338 513822 442574
rect 513266 406658 513502 406894
rect 513586 406658 513822 406894
rect 513266 406338 513502 406574
rect 513586 406338 513822 406574
rect 513266 370658 513502 370894
rect 513586 370658 513822 370894
rect 513266 370338 513502 370574
rect 513586 370338 513822 370574
rect 513266 334658 513502 334894
rect 513586 334658 513822 334894
rect 513266 334338 513502 334574
rect 513586 334338 513822 334574
rect 513266 298658 513502 298894
rect 513586 298658 513822 298894
rect 513266 298338 513502 298574
rect 513586 298338 513822 298574
rect 513266 262658 513502 262894
rect 513586 262658 513822 262894
rect 513266 262338 513502 262574
rect 513586 262338 513822 262574
rect 513266 226658 513502 226894
rect 513586 226658 513822 226894
rect 513266 226338 513502 226574
rect 513586 226338 513822 226574
rect 513266 190658 513502 190894
rect 513586 190658 513822 190894
rect 513266 190338 513502 190574
rect 513586 190338 513822 190574
rect 513266 154658 513502 154894
rect 513586 154658 513822 154894
rect 513266 154338 513502 154574
rect 513586 154338 513822 154574
rect 513266 118658 513502 118894
rect 513586 118658 513822 118894
rect 513266 118338 513502 118574
rect 513586 118338 513822 118574
rect 513266 82658 513502 82894
rect 513586 82658 513822 82894
rect 513266 82338 513502 82574
rect 513586 82338 513822 82574
rect 513266 46658 513502 46894
rect 513586 46658 513822 46894
rect 513266 46338 513502 46574
rect 513586 46338 513822 46574
rect 513266 10658 513502 10894
rect 513586 10658 513822 10894
rect 513266 10338 513502 10574
rect 513586 10338 513822 10574
rect 513266 -4422 513502 -4186
rect 513586 -4422 513822 -4186
rect 513266 -4742 513502 -4506
rect 513586 -4742 513822 -4506
rect 534986 711322 535222 711558
rect 535306 711322 535542 711558
rect 534986 711002 535222 711238
rect 535306 711002 535542 711238
rect 531266 709402 531502 709638
rect 531586 709402 531822 709638
rect 531266 709082 531502 709318
rect 531586 709082 531822 709318
rect 527546 707482 527782 707718
rect 527866 707482 528102 707718
rect 527546 707162 527782 707398
rect 527866 707162 528102 707398
rect 516986 698378 517222 698614
rect 517306 698378 517542 698614
rect 516986 698058 517222 698294
rect 517306 698058 517542 698294
rect 516986 662378 517222 662614
rect 517306 662378 517542 662614
rect 516986 662058 517222 662294
rect 517306 662058 517542 662294
rect 516986 626378 517222 626614
rect 517306 626378 517542 626614
rect 516986 626058 517222 626294
rect 517306 626058 517542 626294
rect 516986 590378 517222 590614
rect 517306 590378 517542 590614
rect 516986 590058 517222 590294
rect 517306 590058 517542 590294
rect 516986 554378 517222 554614
rect 517306 554378 517542 554614
rect 516986 554058 517222 554294
rect 517306 554058 517542 554294
rect 516986 518378 517222 518614
rect 517306 518378 517542 518614
rect 516986 518058 517222 518294
rect 517306 518058 517542 518294
rect 516986 482378 517222 482614
rect 517306 482378 517542 482614
rect 516986 482058 517222 482294
rect 517306 482058 517542 482294
rect 516986 446378 517222 446614
rect 517306 446378 517542 446614
rect 516986 446058 517222 446294
rect 517306 446058 517542 446294
rect 516986 410378 517222 410614
rect 517306 410378 517542 410614
rect 516986 410058 517222 410294
rect 517306 410058 517542 410294
rect 516986 374378 517222 374614
rect 517306 374378 517542 374614
rect 516986 374058 517222 374294
rect 517306 374058 517542 374294
rect 516986 338378 517222 338614
rect 517306 338378 517542 338614
rect 516986 338058 517222 338294
rect 517306 338058 517542 338294
rect 516986 302378 517222 302614
rect 517306 302378 517542 302614
rect 516986 302058 517222 302294
rect 517306 302058 517542 302294
rect 516986 266378 517222 266614
rect 517306 266378 517542 266614
rect 516986 266058 517222 266294
rect 517306 266058 517542 266294
rect 516986 230378 517222 230614
rect 517306 230378 517542 230614
rect 516986 230058 517222 230294
rect 517306 230058 517542 230294
rect 516986 194378 517222 194614
rect 517306 194378 517542 194614
rect 516986 194058 517222 194294
rect 517306 194058 517542 194294
rect 516986 158378 517222 158614
rect 517306 158378 517542 158614
rect 516986 158058 517222 158294
rect 517306 158058 517542 158294
rect 516986 122378 517222 122614
rect 517306 122378 517542 122614
rect 516986 122058 517222 122294
rect 517306 122058 517542 122294
rect 516986 86378 517222 86614
rect 517306 86378 517542 86614
rect 516986 86058 517222 86294
rect 517306 86058 517542 86294
rect 516986 50378 517222 50614
rect 517306 50378 517542 50614
rect 516986 50058 517222 50294
rect 517306 50058 517542 50294
rect 516986 14378 517222 14614
rect 517306 14378 517542 14614
rect 516986 14058 517222 14294
rect 517306 14058 517542 14294
rect 498986 -7302 499222 -7066
rect 499306 -7302 499542 -7066
rect 498986 -7622 499222 -7386
rect 499306 -7622 499542 -7386
rect 523826 705562 524062 705798
rect 524146 705562 524382 705798
rect 523826 705242 524062 705478
rect 524146 705242 524382 705478
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -1542 524062 -1306
rect 524146 -1542 524382 -1306
rect 523826 -1862 524062 -1626
rect 524146 -1862 524382 -1626
rect 527546 672938 527782 673174
rect 527866 672938 528102 673174
rect 527546 672618 527782 672854
rect 527866 672618 528102 672854
rect 527546 636938 527782 637174
rect 527866 636938 528102 637174
rect 527546 636618 527782 636854
rect 527866 636618 528102 636854
rect 527546 600938 527782 601174
rect 527866 600938 528102 601174
rect 527546 600618 527782 600854
rect 527866 600618 528102 600854
rect 527546 564938 527782 565174
rect 527866 564938 528102 565174
rect 527546 564618 527782 564854
rect 527866 564618 528102 564854
rect 527546 528938 527782 529174
rect 527866 528938 528102 529174
rect 527546 528618 527782 528854
rect 527866 528618 528102 528854
rect 527546 492938 527782 493174
rect 527866 492938 528102 493174
rect 527546 492618 527782 492854
rect 527866 492618 528102 492854
rect 527546 456938 527782 457174
rect 527866 456938 528102 457174
rect 527546 456618 527782 456854
rect 527866 456618 528102 456854
rect 527546 420938 527782 421174
rect 527866 420938 528102 421174
rect 527546 420618 527782 420854
rect 527866 420618 528102 420854
rect 527546 384938 527782 385174
rect 527866 384938 528102 385174
rect 527546 384618 527782 384854
rect 527866 384618 528102 384854
rect 527546 348938 527782 349174
rect 527866 348938 528102 349174
rect 527546 348618 527782 348854
rect 527866 348618 528102 348854
rect 527546 312938 527782 313174
rect 527866 312938 528102 313174
rect 527546 312618 527782 312854
rect 527866 312618 528102 312854
rect 527546 276938 527782 277174
rect 527866 276938 528102 277174
rect 527546 276618 527782 276854
rect 527866 276618 528102 276854
rect 527546 240938 527782 241174
rect 527866 240938 528102 241174
rect 527546 240618 527782 240854
rect 527866 240618 528102 240854
rect 527546 204938 527782 205174
rect 527866 204938 528102 205174
rect 527546 204618 527782 204854
rect 527866 204618 528102 204854
rect 527546 168938 527782 169174
rect 527866 168938 528102 169174
rect 527546 168618 527782 168854
rect 527866 168618 528102 168854
rect 527546 132938 527782 133174
rect 527866 132938 528102 133174
rect 527546 132618 527782 132854
rect 527866 132618 528102 132854
rect 527546 96938 527782 97174
rect 527866 96938 528102 97174
rect 527546 96618 527782 96854
rect 527866 96618 528102 96854
rect 527546 60938 527782 61174
rect 527866 60938 528102 61174
rect 527546 60618 527782 60854
rect 527866 60618 528102 60854
rect 527546 24938 527782 25174
rect 527866 24938 528102 25174
rect 527546 24618 527782 24854
rect 527866 24618 528102 24854
rect 527546 -3462 527782 -3226
rect 527866 -3462 528102 -3226
rect 527546 -3782 527782 -3546
rect 527866 -3782 528102 -3546
rect 531266 676658 531502 676894
rect 531586 676658 531822 676894
rect 531266 676338 531502 676574
rect 531586 676338 531822 676574
rect 531266 640658 531502 640894
rect 531586 640658 531822 640894
rect 531266 640338 531502 640574
rect 531586 640338 531822 640574
rect 531266 604658 531502 604894
rect 531586 604658 531822 604894
rect 531266 604338 531502 604574
rect 531586 604338 531822 604574
rect 531266 568658 531502 568894
rect 531586 568658 531822 568894
rect 531266 568338 531502 568574
rect 531586 568338 531822 568574
rect 531266 532658 531502 532894
rect 531586 532658 531822 532894
rect 531266 532338 531502 532574
rect 531586 532338 531822 532574
rect 531266 496658 531502 496894
rect 531586 496658 531822 496894
rect 531266 496338 531502 496574
rect 531586 496338 531822 496574
rect 531266 460658 531502 460894
rect 531586 460658 531822 460894
rect 531266 460338 531502 460574
rect 531586 460338 531822 460574
rect 531266 424658 531502 424894
rect 531586 424658 531822 424894
rect 531266 424338 531502 424574
rect 531586 424338 531822 424574
rect 531266 388658 531502 388894
rect 531586 388658 531822 388894
rect 531266 388338 531502 388574
rect 531586 388338 531822 388574
rect 531266 352658 531502 352894
rect 531586 352658 531822 352894
rect 531266 352338 531502 352574
rect 531586 352338 531822 352574
rect 531266 316658 531502 316894
rect 531586 316658 531822 316894
rect 531266 316338 531502 316574
rect 531586 316338 531822 316574
rect 531266 280658 531502 280894
rect 531586 280658 531822 280894
rect 531266 280338 531502 280574
rect 531586 280338 531822 280574
rect 531266 244658 531502 244894
rect 531586 244658 531822 244894
rect 531266 244338 531502 244574
rect 531586 244338 531822 244574
rect 531266 208658 531502 208894
rect 531586 208658 531822 208894
rect 531266 208338 531502 208574
rect 531586 208338 531822 208574
rect 531266 172658 531502 172894
rect 531586 172658 531822 172894
rect 531266 172338 531502 172574
rect 531586 172338 531822 172574
rect 531266 136658 531502 136894
rect 531586 136658 531822 136894
rect 531266 136338 531502 136574
rect 531586 136338 531822 136574
rect 531266 100658 531502 100894
rect 531586 100658 531822 100894
rect 531266 100338 531502 100574
rect 531586 100338 531822 100574
rect 531266 64658 531502 64894
rect 531586 64658 531822 64894
rect 531266 64338 531502 64574
rect 531586 64338 531822 64574
rect 531266 28658 531502 28894
rect 531586 28658 531822 28894
rect 531266 28338 531502 28574
rect 531586 28338 531822 28574
rect 531266 -5382 531502 -5146
rect 531586 -5382 531822 -5146
rect 531266 -5702 531502 -5466
rect 531586 -5702 531822 -5466
rect 552986 710362 553222 710598
rect 553306 710362 553542 710598
rect 552986 710042 553222 710278
rect 553306 710042 553542 710278
rect 549266 708442 549502 708678
rect 549586 708442 549822 708678
rect 549266 708122 549502 708358
rect 549586 708122 549822 708358
rect 545546 706522 545782 706758
rect 545866 706522 546102 706758
rect 545546 706202 545782 706438
rect 545866 706202 546102 706438
rect 534986 680378 535222 680614
rect 535306 680378 535542 680614
rect 534986 680058 535222 680294
rect 535306 680058 535542 680294
rect 534986 644378 535222 644614
rect 535306 644378 535542 644614
rect 534986 644058 535222 644294
rect 535306 644058 535542 644294
rect 534986 608378 535222 608614
rect 535306 608378 535542 608614
rect 534986 608058 535222 608294
rect 535306 608058 535542 608294
rect 534986 572378 535222 572614
rect 535306 572378 535542 572614
rect 534986 572058 535222 572294
rect 535306 572058 535542 572294
rect 534986 536378 535222 536614
rect 535306 536378 535542 536614
rect 534986 536058 535222 536294
rect 535306 536058 535542 536294
rect 534986 500378 535222 500614
rect 535306 500378 535542 500614
rect 534986 500058 535222 500294
rect 535306 500058 535542 500294
rect 534986 464378 535222 464614
rect 535306 464378 535542 464614
rect 534986 464058 535222 464294
rect 535306 464058 535542 464294
rect 534986 428378 535222 428614
rect 535306 428378 535542 428614
rect 534986 428058 535222 428294
rect 535306 428058 535542 428294
rect 534986 392378 535222 392614
rect 535306 392378 535542 392614
rect 534986 392058 535222 392294
rect 535306 392058 535542 392294
rect 534986 356378 535222 356614
rect 535306 356378 535542 356614
rect 534986 356058 535222 356294
rect 535306 356058 535542 356294
rect 534986 320378 535222 320614
rect 535306 320378 535542 320614
rect 534986 320058 535222 320294
rect 535306 320058 535542 320294
rect 534986 284378 535222 284614
rect 535306 284378 535542 284614
rect 534986 284058 535222 284294
rect 535306 284058 535542 284294
rect 534986 248378 535222 248614
rect 535306 248378 535542 248614
rect 534986 248058 535222 248294
rect 535306 248058 535542 248294
rect 534986 212378 535222 212614
rect 535306 212378 535542 212614
rect 534986 212058 535222 212294
rect 535306 212058 535542 212294
rect 534986 176378 535222 176614
rect 535306 176378 535542 176614
rect 534986 176058 535222 176294
rect 535306 176058 535542 176294
rect 534986 140378 535222 140614
rect 535306 140378 535542 140614
rect 534986 140058 535222 140294
rect 535306 140058 535542 140294
rect 534986 104378 535222 104614
rect 535306 104378 535542 104614
rect 534986 104058 535222 104294
rect 535306 104058 535542 104294
rect 534986 68378 535222 68614
rect 535306 68378 535542 68614
rect 534986 68058 535222 68294
rect 535306 68058 535542 68294
rect 534986 32378 535222 32614
rect 535306 32378 535542 32614
rect 534986 32058 535222 32294
rect 535306 32058 535542 32294
rect 516986 -6342 517222 -6106
rect 517306 -6342 517542 -6106
rect 516986 -6662 517222 -6426
rect 517306 -6662 517542 -6426
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 690938 545782 691174
rect 545866 690938 546102 691174
rect 545546 690618 545782 690854
rect 545866 690618 546102 690854
rect 545546 654938 545782 655174
rect 545866 654938 546102 655174
rect 545546 654618 545782 654854
rect 545866 654618 546102 654854
rect 545546 618938 545782 619174
rect 545866 618938 546102 619174
rect 545546 618618 545782 618854
rect 545866 618618 546102 618854
rect 545546 582938 545782 583174
rect 545866 582938 546102 583174
rect 545546 582618 545782 582854
rect 545866 582618 546102 582854
rect 545546 546938 545782 547174
rect 545866 546938 546102 547174
rect 545546 546618 545782 546854
rect 545866 546618 546102 546854
rect 545546 510938 545782 511174
rect 545866 510938 546102 511174
rect 545546 510618 545782 510854
rect 545866 510618 546102 510854
rect 545546 474938 545782 475174
rect 545866 474938 546102 475174
rect 545546 474618 545782 474854
rect 545866 474618 546102 474854
rect 545546 438938 545782 439174
rect 545866 438938 546102 439174
rect 545546 438618 545782 438854
rect 545866 438618 546102 438854
rect 545546 402938 545782 403174
rect 545866 402938 546102 403174
rect 545546 402618 545782 402854
rect 545866 402618 546102 402854
rect 545546 366938 545782 367174
rect 545866 366938 546102 367174
rect 545546 366618 545782 366854
rect 545866 366618 546102 366854
rect 545546 330938 545782 331174
rect 545866 330938 546102 331174
rect 545546 330618 545782 330854
rect 545866 330618 546102 330854
rect 545546 294938 545782 295174
rect 545866 294938 546102 295174
rect 545546 294618 545782 294854
rect 545866 294618 546102 294854
rect 545546 258938 545782 259174
rect 545866 258938 546102 259174
rect 545546 258618 545782 258854
rect 545866 258618 546102 258854
rect 545546 222938 545782 223174
rect 545866 222938 546102 223174
rect 545546 222618 545782 222854
rect 545866 222618 546102 222854
rect 545546 186938 545782 187174
rect 545866 186938 546102 187174
rect 545546 186618 545782 186854
rect 545866 186618 546102 186854
rect 545546 150938 545782 151174
rect 545866 150938 546102 151174
rect 545546 150618 545782 150854
rect 545866 150618 546102 150854
rect 545546 114938 545782 115174
rect 545866 114938 546102 115174
rect 545546 114618 545782 114854
rect 545866 114618 546102 114854
rect 545546 78938 545782 79174
rect 545866 78938 546102 79174
rect 545546 78618 545782 78854
rect 545866 78618 546102 78854
rect 545546 42938 545782 43174
rect 545866 42938 546102 43174
rect 545546 42618 545782 42854
rect 545866 42618 546102 42854
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -2502 545782 -2266
rect 545866 -2502 546102 -2266
rect 545546 -2822 545782 -2586
rect 545866 -2822 546102 -2586
rect 549266 694658 549502 694894
rect 549586 694658 549822 694894
rect 549266 694338 549502 694574
rect 549586 694338 549822 694574
rect 549266 658658 549502 658894
rect 549586 658658 549822 658894
rect 549266 658338 549502 658574
rect 549586 658338 549822 658574
rect 549266 622658 549502 622894
rect 549586 622658 549822 622894
rect 549266 622338 549502 622574
rect 549586 622338 549822 622574
rect 549266 586658 549502 586894
rect 549586 586658 549822 586894
rect 549266 586338 549502 586574
rect 549586 586338 549822 586574
rect 549266 550658 549502 550894
rect 549586 550658 549822 550894
rect 549266 550338 549502 550574
rect 549586 550338 549822 550574
rect 549266 514658 549502 514894
rect 549586 514658 549822 514894
rect 549266 514338 549502 514574
rect 549586 514338 549822 514574
rect 549266 478658 549502 478894
rect 549586 478658 549822 478894
rect 549266 478338 549502 478574
rect 549586 478338 549822 478574
rect 549266 442658 549502 442894
rect 549586 442658 549822 442894
rect 549266 442338 549502 442574
rect 549586 442338 549822 442574
rect 549266 406658 549502 406894
rect 549586 406658 549822 406894
rect 549266 406338 549502 406574
rect 549586 406338 549822 406574
rect 549266 370658 549502 370894
rect 549586 370658 549822 370894
rect 549266 370338 549502 370574
rect 549586 370338 549822 370574
rect 549266 334658 549502 334894
rect 549586 334658 549822 334894
rect 549266 334338 549502 334574
rect 549586 334338 549822 334574
rect 549266 298658 549502 298894
rect 549586 298658 549822 298894
rect 549266 298338 549502 298574
rect 549586 298338 549822 298574
rect 549266 262658 549502 262894
rect 549586 262658 549822 262894
rect 549266 262338 549502 262574
rect 549586 262338 549822 262574
rect 549266 226658 549502 226894
rect 549586 226658 549822 226894
rect 549266 226338 549502 226574
rect 549586 226338 549822 226574
rect 549266 190658 549502 190894
rect 549586 190658 549822 190894
rect 549266 190338 549502 190574
rect 549586 190338 549822 190574
rect 549266 154658 549502 154894
rect 549586 154658 549822 154894
rect 549266 154338 549502 154574
rect 549586 154338 549822 154574
rect 549266 118658 549502 118894
rect 549586 118658 549822 118894
rect 549266 118338 549502 118574
rect 549586 118338 549822 118574
rect 549266 82658 549502 82894
rect 549586 82658 549822 82894
rect 549266 82338 549502 82574
rect 549586 82338 549822 82574
rect 549266 46658 549502 46894
rect 549586 46658 549822 46894
rect 549266 46338 549502 46574
rect 549586 46338 549822 46574
rect 549266 10658 549502 10894
rect 549586 10658 549822 10894
rect 549266 10338 549502 10574
rect 549586 10338 549822 10574
rect 549266 -4422 549502 -4186
rect 549586 -4422 549822 -4186
rect 549266 -4742 549502 -4506
rect 549586 -4742 549822 -4506
rect 570986 711322 571222 711558
rect 571306 711322 571542 711558
rect 570986 711002 571222 711238
rect 571306 711002 571542 711238
rect 567266 709402 567502 709638
rect 567586 709402 567822 709638
rect 567266 709082 567502 709318
rect 567586 709082 567822 709318
rect 563546 707482 563782 707718
rect 563866 707482 564102 707718
rect 563546 707162 563782 707398
rect 563866 707162 564102 707398
rect 552986 698378 553222 698614
rect 553306 698378 553542 698614
rect 552986 698058 553222 698294
rect 553306 698058 553542 698294
rect 552986 662378 553222 662614
rect 553306 662378 553542 662614
rect 552986 662058 553222 662294
rect 553306 662058 553542 662294
rect 552986 626378 553222 626614
rect 553306 626378 553542 626614
rect 552986 626058 553222 626294
rect 553306 626058 553542 626294
rect 552986 590378 553222 590614
rect 553306 590378 553542 590614
rect 552986 590058 553222 590294
rect 553306 590058 553542 590294
rect 552986 554378 553222 554614
rect 553306 554378 553542 554614
rect 552986 554058 553222 554294
rect 553306 554058 553542 554294
rect 552986 518378 553222 518614
rect 553306 518378 553542 518614
rect 552986 518058 553222 518294
rect 553306 518058 553542 518294
rect 552986 482378 553222 482614
rect 553306 482378 553542 482614
rect 552986 482058 553222 482294
rect 553306 482058 553542 482294
rect 552986 446378 553222 446614
rect 553306 446378 553542 446614
rect 552986 446058 553222 446294
rect 553306 446058 553542 446294
rect 552986 410378 553222 410614
rect 553306 410378 553542 410614
rect 552986 410058 553222 410294
rect 553306 410058 553542 410294
rect 552986 374378 553222 374614
rect 553306 374378 553542 374614
rect 552986 374058 553222 374294
rect 553306 374058 553542 374294
rect 552986 338378 553222 338614
rect 553306 338378 553542 338614
rect 552986 338058 553222 338294
rect 553306 338058 553542 338294
rect 552986 302378 553222 302614
rect 553306 302378 553542 302614
rect 552986 302058 553222 302294
rect 553306 302058 553542 302294
rect 552986 266378 553222 266614
rect 553306 266378 553542 266614
rect 552986 266058 553222 266294
rect 553306 266058 553542 266294
rect 552986 230378 553222 230614
rect 553306 230378 553542 230614
rect 552986 230058 553222 230294
rect 553306 230058 553542 230294
rect 552986 194378 553222 194614
rect 553306 194378 553542 194614
rect 552986 194058 553222 194294
rect 553306 194058 553542 194294
rect 552986 158378 553222 158614
rect 553306 158378 553542 158614
rect 552986 158058 553222 158294
rect 553306 158058 553542 158294
rect 552986 122378 553222 122614
rect 553306 122378 553542 122614
rect 552986 122058 553222 122294
rect 553306 122058 553542 122294
rect 552986 86378 553222 86614
rect 553306 86378 553542 86614
rect 552986 86058 553222 86294
rect 553306 86058 553542 86294
rect 552986 50378 553222 50614
rect 553306 50378 553542 50614
rect 552986 50058 553222 50294
rect 553306 50058 553542 50294
rect 552986 14378 553222 14614
rect 553306 14378 553542 14614
rect 552986 14058 553222 14294
rect 553306 14058 553542 14294
rect 534986 -7302 535222 -7066
rect 535306 -7302 535542 -7066
rect 534986 -7622 535222 -7386
rect 535306 -7622 535542 -7386
rect 559826 705562 560062 705798
rect 560146 705562 560382 705798
rect 559826 705242 560062 705478
rect 560146 705242 560382 705478
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -1542 560062 -1306
rect 560146 -1542 560382 -1306
rect 559826 -1862 560062 -1626
rect 560146 -1862 560382 -1626
rect 563546 672938 563782 673174
rect 563866 672938 564102 673174
rect 563546 672618 563782 672854
rect 563866 672618 564102 672854
rect 563546 636938 563782 637174
rect 563866 636938 564102 637174
rect 563546 636618 563782 636854
rect 563866 636618 564102 636854
rect 563546 600938 563782 601174
rect 563866 600938 564102 601174
rect 563546 600618 563782 600854
rect 563866 600618 564102 600854
rect 563546 564938 563782 565174
rect 563866 564938 564102 565174
rect 563546 564618 563782 564854
rect 563866 564618 564102 564854
rect 563546 528938 563782 529174
rect 563866 528938 564102 529174
rect 563546 528618 563782 528854
rect 563866 528618 564102 528854
rect 563546 492938 563782 493174
rect 563866 492938 564102 493174
rect 563546 492618 563782 492854
rect 563866 492618 564102 492854
rect 563546 456938 563782 457174
rect 563866 456938 564102 457174
rect 563546 456618 563782 456854
rect 563866 456618 564102 456854
rect 563546 420938 563782 421174
rect 563866 420938 564102 421174
rect 563546 420618 563782 420854
rect 563866 420618 564102 420854
rect 563546 384938 563782 385174
rect 563866 384938 564102 385174
rect 563546 384618 563782 384854
rect 563866 384618 564102 384854
rect 563546 348938 563782 349174
rect 563866 348938 564102 349174
rect 563546 348618 563782 348854
rect 563866 348618 564102 348854
rect 563546 312938 563782 313174
rect 563866 312938 564102 313174
rect 563546 312618 563782 312854
rect 563866 312618 564102 312854
rect 563546 276938 563782 277174
rect 563866 276938 564102 277174
rect 563546 276618 563782 276854
rect 563866 276618 564102 276854
rect 563546 240938 563782 241174
rect 563866 240938 564102 241174
rect 563546 240618 563782 240854
rect 563866 240618 564102 240854
rect 563546 204938 563782 205174
rect 563866 204938 564102 205174
rect 563546 204618 563782 204854
rect 563866 204618 564102 204854
rect 563546 168938 563782 169174
rect 563866 168938 564102 169174
rect 563546 168618 563782 168854
rect 563866 168618 564102 168854
rect 563546 132938 563782 133174
rect 563866 132938 564102 133174
rect 563546 132618 563782 132854
rect 563866 132618 564102 132854
rect 563546 96938 563782 97174
rect 563866 96938 564102 97174
rect 563546 96618 563782 96854
rect 563866 96618 564102 96854
rect 563546 60938 563782 61174
rect 563866 60938 564102 61174
rect 563546 60618 563782 60854
rect 563866 60618 564102 60854
rect 563546 24938 563782 25174
rect 563866 24938 564102 25174
rect 563546 24618 563782 24854
rect 563866 24618 564102 24854
rect 563546 -3462 563782 -3226
rect 563866 -3462 564102 -3226
rect 563546 -3782 563782 -3546
rect 563866 -3782 564102 -3546
rect 567266 676658 567502 676894
rect 567586 676658 567822 676894
rect 567266 676338 567502 676574
rect 567586 676338 567822 676574
rect 567266 640658 567502 640894
rect 567586 640658 567822 640894
rect 567266 640338 567502 640574
rect 567586 640338 567822 640574
rect 567266 604658 567502 604894
rect 567586 604658 567822 604894
rect 567266 604338 567502 604574
rect 567586 604338 567822 604574
rect 567266 568658 567502 568894
rect 567586 568658 567822 568894
rect 567266 568338 567502 568574
rect 567586 568338 567822 568574
rect 567266 532658 567502 532894
rect 567586 532658 567822 532894
rect 567266 532338 567502 532574
rect 567586 532338 567822 532574
rect 567266 496658 567502 496894
rect 567586 496658 567822 496894
rect 567266 496338 567502 496574
rect 567586 496338 567822 496574
rect 567266 460658 567502 460894
rect 567586 460658 567822 460894
rect 567266 460338 567502 460574
rect 567586 460338 567822 460574
rect 567266 424658 567502 424894
rect 567586 424658 567822 424894
rect 567266 424338 567502 424574
rect 567586 424338 567822 424574
rect 567266 388658 567502 388894
rect 567586 388658 567822 388894
rect 567266 388338 567502 388574
rect 567586 388338 567822 388574
rect 567266 352658 567502 352894
rect 567586 352658 567822 352894
rect 567266 352338 567502 352574
rect 567586 352338 567822 352574
rect 567266 316658 567502 316894
rect 567586 316658 567822 316894
rect 567266 316338 567502 316574
rect 567586 316338 567822 316574
rect 567266 280658 567502 280894
rect 567586 280658 567822 280894
rect 567266 280338 567502 280574
rect 567586 280338 567822 280574
rect 567266 244658 567502 244894
rect 567586 244658 567822 244894
rect 567266 244338 567502 244574
rect 567586 244338 567822 244574
rect 567266 208658 567502 208894
rect 567586 208658 567822 208894
rect 567266 208338 567502 208574
rect 567586 208338 567822 208574
rect 567266 172658 567502 172894
rect 567586 172658 567822 172894
rect 567266 172338 567502 172574
rect 567586 172338 567822 172574
rect 567266 136658 567502 136894
rect 567586 136658 567822 136894
rect 567266 136338 567502 136574
rect 567586 136338 567822 136574
rect 567266 100658 567502 100894
rect 567586 100658 567822 100894
rect 567266 100338 567502 100574
rect 567586 100338 567822 100574
rect 567266 64658 567502 64894
rect 567586 64658 567822 64894
rect 567266 64338 567502 64574
rect 567586 64338 567822 64574
rect 567266 28658 567502 28894
rect 567586 28658 567822 28894
rect 567266 28338 567502 28574
rect 567586 28338 567822 28574
rect 567266 -5382 567502 -5146
rect 567586 -5382 567822 -5146
rect 567266 -5702 567502 -5466
rect 567586 -5702 567822 -5466
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 581546 706522 581782 706758
rect 581866 706522 582102 706758
rect 581546 706202 581782 706438
rect 581866 706202 582102 706438
rect 570986 680378 571222 680614
rect 571306 680378 571542 680614
rect 570986 680058 571222 680294
rect 571306 680058 571542 680294
rect 570986 644378 571222 644614
rect 571306 644378 571542 644614
rect 570986 644058 571222 644294
rect 571306 644058 571542 644294
rect 570986 608378 571222 608614
rect 571306 608378 571542 608614
rect 570986 608058 571222 608294
rect 571306 608058 571542 608294
rect 570986 572378 571222 572614
rect 571306 572378 571542 572614
rect 570986 572058 571222 572294
rect 571306 572058 571542 572294
rect 570986 536378 571222 536614
rect 571306 536378 571542 536614
rect 570986 536058 571222 536294
rect 571306 536058 571542 536294
rect 570986 500378 571222 500614
rect 571306 500378 571542 500614
rect 570986 500058 571222 500294
rect 571306 500058 571542 500294
rect 570986 464378 571222 464614
rect 571306 464378 571542 464614
rect 570986 464058 571222 464294
rect 571306 464058 571542 464294
rect 570986 428378 571222 428614
rect 571306 428378 571542 428614
rect 570986 428058 571222 428294
rect 571306 428058 571542 428294
rect 570986 392378 571222 392614
rect 571306 392378 571542 392614
rect 570986 392058 571222 392294
rect 571306 392058 571542 392294
rect 570986 356378 571222 356614
rect 571306 356378 571542 356614
rect 570986 356058 571222 356294
rect 571306 356058 571542 356294
rect 570986 320378 571222 320614
rect 571306 320378 571542 320614
rect 570986 320058 571222 320294
rect 571306 320058 571542 320294
rect 570986 284378 571222 284614
rect 571306 284378 571542 284614
rect 570986 284058 571222 284294
rect 571306 284058 571542 284294
rect 570986 248378 571222 248614
rect 571306 248378 571542 248614
rect 570986 248058 571222 248294
rect 571306 248058 571542 248294
rect 570986 212378 571222 212614
rect 571306 212378 571542 212614
rect 570986 212058 571222 212294
rect 571306 212058 571542 212294
rect 570986 176378 571222 176614
rect 571306 176378 571542 176614
rect 570986 176058 571222 176294
rect 571306 176058 571542 176294
rect 570986 140378 571222 140614
rect 571306 140378 571542 140614
rect 570986 140058 571222 140294
rect 571306 140058 571542 140294
rect 570986 104378 571222 104614
rect 571306 104378 571542 104614
rect 570986 104058 571222 104294
rect 571306 104058 571542 104294
rect 570986 68378 571222 68614
rect 571306 68378 571542 68614
rect 570986 68058 571222 68294
rect 571306 68058 571542 68294
rect 570986 32378 571222 32614
rect 571306 32378 571542 32614
rect 570986 32058 571222 32294
rect 571306 32058 571542 32294
rect 552986 -6342 553222 -6106
rect 553306 -6342 553542 -6106
rect 552986 -6662 553222 -6426
rect 553306 -6662 553542 -6426
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 669218 586538 669454
rect 586622 669218 586858 669454
rect 586302 668898 586538 669134
rect 586622 668898 586858 669134
rect 586302 633218 586538 633454
rect 586622 633218 586858 633454
rect 586302 632898 586538 633134
rect 586622 632898 586858 633134
rect 586302 597218 586538 597454
rect 586622 597218 586858 597454
rect 586302 596898 586538 597134
rect 586622 596898 586858 597134
rect 586302 561218 586538 561454
rect 586622 561218 586858 561454
rect 586302 560898 586538 561134
rect 586622 560898 586858 561134
rect 586302 525218 586538 525454
rect 586622 525218 586858 525454
rect 586302 524898 586538 525134
rect 586622 524898 586858 525134
rect 586302 489218 586538 489454
rect 586622 489218 586858 489454
rect 586302 488898 586538 489134
rect 586622 488898 586858 489134
rect 586302 453218 586538 453454
rect 586622 453218 586858 453454
rect 586302 452898 586538 453134
rect 586622 452898 586858 453134
rect 586302 417218 586538 417454
rect 586622 417218 586858 417454
rect 586302 416898 586538 417134
rect 586622 416898 586858 417134
rect 586302 381218 586538 381454
rect 586622 381218 586858 381454
rect 586302 380898 586538 381134
rect 586622 380898 586858 381134
rect 586302 345218 586538 345454
rect 586622 345218 586858 345454
rect 586302 344898 586538 345134
rect 586622 344898 586858 345134
rect 586302 309218 586538 309454
rect 586622 309218 586858 309454
rect 586302 308898 586538 309134
rect 586622 308898 586858 309134
rect 586302 273218 586538 273454
rect 586622 273218 586858 273454
rect 586302 272898 586538 273134
rect 586622 272898 586858 273134
rect 586302 237218 586538 237454
rect 586622 237218 586858 237454
rect 586302 236898 586538 237134
rect 586622 236898 586858 237134
rect 586302 201218 586538 201454
rect 586622 201218 586858 201454
rect 586302 200898 586538 201134
rect 586622 200898 586858 201134
rect 586302 165218 586538 165454
rect 586622 165218 586858 165454
rect 586302 164898 586538 165134
rect 586622 164898 586858 165134
rect 586302 129218 586538 129454
rect 586622 129218 586858 129454
rect 586302 128898 586538 129134
rect 586622 128898 586858 129134
rect 586302 93218 586538 93454
rect 586622 93218 586858 93454
rect 586302 92898 586538 93134
rect 586622 92898 586858 93134
rect 586302 57218 586538 57454
rect 586622 57218 586858 57454
rect 586302 56898 586538 57134
rect 586622 56898 586858 57134
rect 586302 21218 586538 21454
rect 586622 21218 586858 21454
rect 586302 20898 586538 21134
rect 586622 20898 586858 21134
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 690938 587498 691174
rect 587582 690938 587818 691174
rect 587262 690618 587498 690854
rect 587582 690618 587818 690854
rect 587262 654938 587498 655174
rect 587582 654938 587818 655174
rect 587262 654618 587498 654854
rect 587582 654618 587818 654854
rect 587262 618938 587498 619174
rect 587582 618938 587818 619174
rect 587262 618618 587498 618854
rect 587582 618618 587818 618854
rect 587262 582938 587498 583174
rect 587582 582938 587818 583174
rect 587262 582618 587498 582854
rect 587582 582618 587818 582854
rect 587262 546938 587498 547174
rect 587582 546938 587818 547174
rect 587262 546618 587498 546854
rect 587582 546618 587818 546854
rect 587262 510938 587498 511174
rect 587582 510938 587818 511174
rect 587262 510618 587498 510854
rect 587582 510618 587818 510854
rect 587262 474938 587498 475174
rect 587582 474938 587818 475174
rect 587262 474618 587498 474854
rect 587582 474618 587818 474854
rect 587262 438938 587498 439174
rect 587582 438938 587818 439174
rect 587262 438618 587498 438854
rect 587582 438618 587818 438854
rect 587262 402938 587498 403174
rect 587582 402938 587818 403174
rect 587262 402618 587498 402854
rect 587582 402618 587818 402854
rect 587262 366938 587498 367174
rect 587582 366938 587818 367174
rect 587262 366618 587498 366854
rect 587582 366618 587818 366854
rect 587262 330938 587498 331174
rect 587582 330938 587818 331174
rect 587262 330618 587498 330854
rect 587582 330618 587818 330854
rect 587262 294938 587498 295174
rect 587582 294938 587818 295174
rect 587262 294618 587498 294854
rect 587582 294618 587818 294854
rect 587262 258938 587498 259174
rect 587582 258938 587818 259174
rect 587262 258618 587498 258854
rect 587582 258618 587818 258854
rect 587262 222938 587498 223174
rect 587582 222938 587818 223174
rect 587262 222618 587498 222854
rect 587582 222618 587818 222854
rect 587262 186938 587498 187174
rect 587582 186938 587818 187174
rect 587262 186618 587498 186854
rect 587582 186618 587818 186854
rect 587262 150938 587498 151174
rect 587582 150938 587818 151174
rect 587262 150618 587498 150854
rect 587582 150618 587818 150854
rect 587262 114938 587498 115174
rect 587582 114938 587818 115174
rect 587262 114618 587498 114854
rect 587582 114618 587818 114854
rect 587262 78938 587498 79174
rect 587582 78938 587818 79174
rect 587262 78618 587498 78854
rect 587582 78618 587818 78854
rect 587262 42938 587498 43174
rect 587582 42938 587818 43174
rect 587262 42618 587498 42854
rect 587582 42618 587818 42854
rect 587262 6938 587498 7174
rect 587582 6938 587818 7174
rect 587262 6618 587498 6854
rect 587582 6618 587818 6854
rect 581546 -2502 581782 -2266
rect 581866 -2502 582102 -2266
rect 581546 -2822 581782 -2586
rect 581866 -2822 582102 -2586
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 672938 588458 673174
rect 588542 672938 588778 673174
rect 588222 672618 588458 672854
rect 588542 672618 588778 672854
rect 588222 636938 588458 637174
rect 588542 636938 588778 637174
rect 588222 636618 588458 636854
rect 588542 636618 588778 636854
rect 588222 600938 588458 601174
rect 588542 600938 588778 601174
rect 588222 600618 588458 600854
rect 588542 600618 588778 600854
rect 588222 564938 588458 565174
rect 588542 564938 588778 565174
rect 588222 564618 588458 564854
rect 588542 564618 588778 564854
rect 588222 528938 588458 529174
rect 588542 528938 588778 529174
rect 588222 528618 588458 528854
rect 588542 528618 588778 528854
rect 588222 492938 588458 493174
rect 588542 492938 588778 493174
rect 588222 492618 588458 492854
rect 588542 492618 588778 492854
rect 588222 456938 588458 457174
rect 588542 456938 588778 457174
rect 588222 456618 588458 456854
rect 588542 456618 588778 456854
rect 588222 420938 588458 421174
rect 588542 420938 588778 421174
rect 588222 420618 588458 420854
rect 588542 420618 588778 420854
rect 588222 384938 588458 385174
rect 588542 384938 588778 385174
rect 588222 384618 588458 384854
rect 588542 384618 588778 384854
rect 588222 348938 588458 349174
rect 588542 348938 588778 349174
rect 588222 348618 588458 348854
rect 588542 348618 588778 348854
rect 588222 312938 588458 313174
rect 588542 312938 588778 313174
rect 588222 312618 588458 312854
rect 588542 312618 588778 312854
rect 588222 276938 588458 277174
rect 588542 276938 588778 277174
rect 588222 276618 588458 276854
rect 588542 276618 588778 276854
rect 588222 240938 588458 241174
rect 588542 240938 588778 241174
rect 588222 240618 588458 240854
rect 588542 240618 588778 240854
rect 588222 204938 588458 205174
rect 588542 204938 588778 205174
rect 588222 204618 588458 204854
rect 588542 204618 588778 204854
rect 588222 168938 588458 169174
rect 588542 168938 588778 169174
rect 588222 168618 588458 168854
rect 588542 168618 588778 168854
rect 588222 132938 588458 133174
rect 588542 132938 588778 133174
rect 588222 132618 588458 132854
rect 588542 132618 588778 132854
rect 588222 96938 588458 97174
rect 588542 96938 588778 97174
rect 588222 96618 588458 96854
rect 588542 96618 588778 96854
rect 588222 60938 588458 61174
rect 588542 60938 588778 61174
rect 588222 60618 588458 60854
rect 588542 60618 588778 60854
rect 588222 24938 588458 25174
rect 588542 24938 588778 25174
rect 588222 24618 588458 24854
rect 588542 24618 588778 24854
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 694658 589418 694894
rect 589502 694658 589738 694894
rect 589182 694338 589418 694574
rect 589502 694338 589738 694574
rect 589182 658658 589418 658894
rect 589502 658658 589738 658894
rect 589182 658338 589418 658574
rect 589502 658338 589738 658574
rect 589182 622658 589418 622894
rect 589502 622658 589738 622894
rect 589182 622338 589418 622574
rect 589502 622338 589738 622574
rect 589182 586658 589418 586894
rect 589502 586658 589738 586894
rect 589182 586338 589418 586574
rect 589502 586338 589738 586574
rect 589182 550658 589418 550894
rect 589502 550658 589738 550894
rect 589182 550338 589418 550574
rect 589502 550338 589738 550574
rect 589182 514658 589418 514894
rect 589502 514658 589738 514894
rect 589182 514338 589418 514574
rect 589502 514338 589738 514574
rect 589182 478658 589418 478894
rect 589502 478658 589738 478894
rect 589182 478338 589418 478574
rect 589502 478338 589738 478574
rect 589182 442658 589418 442894
rect 589502 442658 589738 442894
rect 589182 442338 589418 442574
rect 589502 442338 589738 442574
rect 589182 406658 589418 406894
rect 589502 406658 589738 406894
rect 589182 406338 589418 406574
rect 589502 406338 589738 406574
rect 589182 370658 589418 370894
rect 589502 370658 589738 370894
rect 589182 370338 589418 370574
rect 589502 370338 589738 370574
rect 589182 334658 589418 334894
rect 589502 334658 589738 334894
rect 589182 334338 589418 334574
rect 589502 334338 589738 334574
rect 589182 298658 589418 298894
rect 589502 298658 589738 298894
rect 589182 298338 589418 298574
rect 589502 298338 589738 298574
rect 589182 262658 589418 262894
rect 589502 262658 589738 262894
rect 589182 262338 589418 262574
rect 589502 262338 589738 262574
rect 589182 226658 589418 226894
rect 589502 226658 589738 226894
rect 589182 226338 589418 226574
rect 589502 226338 589738 226574
rect 589182 190658 589418 190894
rect 589502 190658 589738 190894
rect 589182 190338 589418 190574
rect 589502 190338 589738 190574
rect 589182 154658 589418 154894
rect 589502 154658 589738 154894
rect 589182 154338 589418 154574
rect 589502 154338 589738 154574
rect 589182 118658 589418 118894
rect 589502 118658 589738 118894
rect 589182 118338 589418 118574
rect 589502 118338 589738 118574
rect 589182 82658 589418 82894
rect 589502 82658 589738 82894
rect 589182 82338 589418 82574
rect 589502 82338 589738 82574
rect 589182 46658 589418 46894
rect 589502 46658 589738 46894
rect 589182 46338 589418 46574
rect 589502 46338 589738 46574
rect 589182 10658 589418 10894
rect 589502 10658 589738 10894
rect 589182 10338 589418 10574
rect 589502 10338 589738 10574
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 676658 590378 676894
rect 590462 676658 590698 676894
rect 590142 676338 590378 676574
rect 590462 676338 590698 676574
rect 590142 640658 590378 640894
rect 590462 640658 590698 640894
rect 590142 640338 590378 640574
rect 590462 640338 590698 640574
rect 590142 604658 590378 604894
rect 590462 604658 590698 604894
rect 590142 604338 590378 604574
rect 590462 604338 590698 604574
rect 590142 568658 590378 568894
rect 590462 568658 590698 568894
rect 590142 568338 590378 568574
rect 590462 568338 590698 568574
rect 590142 532658 590378 532894
rect 590462 532658 590698 532894
rect 590142 532338 590378 532574
rect 590462 532338 590698 532574
rect 590142 496658 590378 496894
rect 590462 496658 590698 496894
rect 590142 496338 590378 496574
rect 590462 496338 590698 496574
rect 590142 460658 590378 460894
rect 590462 460658 590698 460894
rect 590142 460338 590378 460574
rect 590462 460338 590698 460574
rect 590142 424658 590378 424894
rect 590462 424658 590698 424894
rect 590142 424338 590378 424574
rect 590462 424338 590698 424574
rect 590142 388658 590378 388894
rect 590462 388658 590698 388894
rect 590142 388338 590378 388574
rect 590462 388338 590698 388574
rect 590142 352658 590378 352894
rect 590462 352658 590698 352894
rect 590142 352338 590378 352574
rect 590462 352338 590698 352574
rect 590142 316658 590378 316894
rect 590462 316658 590698 316894
rect 590142 316338 590378 316574
rect 590462 316338 590698 316574
rect 590142 280658 590378 280894
rect 590462 280658 590698 280894
rect 590142 280338 590378 280574
rect 590462 280338 590698 280574
rect 590142 244658 590378 244894
rect 590462 244658 590698 244894
rect 590142 244338 590378 244574
rect 590462 244338 590698 244574
rect 590142 208658 590378 208894
rect 590462 208658 590698 208894
rect 590142 208338 590378 208574
rect 590462 208338 590698 208574
rect 590142 172658 590378 172894
rect 590462 172658 590698 172894
rect 590142 172338 590378 172574
rect 590462 172338 590698 172574
rect 590142 136658 590378 136894
rect 590462 136658 590698 136894
rect 590142 136338 590378 136574
rect 590462 136338 590698 136574
rect 590142 100658 590378 100894
rect 590462 100658 590698 100894
rect 590142 100338 590378 100574
rect 590462 100338 590698 100574
rect 590142 64658 590378 64894
rect 590462 64658 590698 64894
rect 590142 64338 590378 64574
rect 590462 64338 590698 64574
rect 590142 28658 590378 28894
rect 590462 28658 590698 28894
rect 590142 28338 590378 28574
rect 590462 28338 590698 28574
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 698378 591338 698614
rect 591422 698378 591658 698614
rect 591102 698058 591338 698294
rect 591422 698058 591658 698294
rect 591102 662378 591338 662614
rect 591422 662378 591658 662614
rect 591102 662058 591338 662294
rect 591422 662058 591658 662294
rect 591102 626378 591338 626614
rect 591422 626378 591658 626614
rect 591102 626058 591338 626294
rect 591422 626058 591658 626294
rect 591102 590378 591338 590614
rect 591422 590378 591658 590614
rect 591102 590058 591338 590294
rect 591422 590058 591658 590294
rect 591102 554378 591338 554614
rect 591422 554378 591658 554614
rect 591102 554058 591338 554294
rect 591422 554058 591658 554294
rect 591102 518378 591338 518614
rect 591422 518378 591658 518614
rect 591102 518058 591338 518294
rect 591422 518058 591658 518294
rect 591102 482378 591338 482614
rect 591422 482378 591658 482614
rect 591102 482058 591338 482294
rect 591422 482058 591658 482294
rect 591102 446378 591338 446614
rect 591422 446378 591658 446614
rect 591102 446058 591338 446294
rect 591422 446058 591658 446294
rect 591102 410378 591338 410614
rect 591422 410378 591658 410614
rect 591102 410058 591338 410294
rect 591422 410058 591658 410294
rect 591102 374378 591338 374614
rect 591422 374378 591658 374614
rect 591102 374058 591338 374294
rect 591422 374058 591658 374294
rect 591102 338378 591338 338614
rect 591422 338378 591658 338614
rect 591102 338058 591338 338294
rect 591422 338058 591658 338294
rect 591102 302378 591338 302614
rect 591422 302378 591658 302614
rect 591102 302058 591338 302294
rect 591422 302058 591658 302294
rect 591102 266378 591338 266614
rect 591422 266378 591658 266614
rect 591102 266058 591338 266294
rect 591422 266058 591658 266294
rect 591102 230378 591338 230614
rect 591422 230378 591658 230614
rect 591102 230058 591338 230294
rect 591422 230058 591658 230294
rect 591102 194378 591338 194614
rect 591422 194378 591658 194614
rect 591102 194058 591338 194294
rect 591422 194058 591658 194294
rect 591102 158378 591338 158614
rect 591422 158378 591658 158614
rect 591102 158058 591338 158294
rect 591422 158058 591658 158294
rect 591102 122378 591338 122614
rect 591422 122378 591658 122614
rect 591102 122058 591338 122294
rect 591422 122058 591658 122294
rect 591102 86378 591338 86614
rect 591422 86378 591658 86614
rect 591102 86058 591338 86294
rect 591422 86058 591658 86294
rect 591102 50378 591338 50614
rect 591422 50378 591658 50614
rect 591102 50058 591338 50294
rect 591422 50058 591658 50294
rect 591102 14378 591338 14614
rect 591422 14378 591658 14614
rect 591102 14058 591338 14294
rect 591422 14058 591658 14294
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 680378 592298 680614
rect 592382 680378 592618 680614
rect 592062 680058 592298 680294
rect 592382 680058 592618 680294
rect 592062 644378 592298 644614
rect 592382 644378 592618 644614
rect 592062 644058 592298 644294
rect 592382 644058 592618 644294
rect 592062 608378 592298 608614
rect 592382 608378 592618 608614
rect 592062 608058 592298 608294
rect 592382 608058 592618 608294
rect 592062 572378 592298 572614
rect 592382 572378 592618 572614
rect 592062 572058 592298 572294
rect 592382 572058 592618 572294
rect 592062 536378 592298 536614
rect 592382 536378 592618 536614
rect 592062 536058 592298 536294
rect 592382 536058 592618 536294
rect 592062 500378 592298 500614
rect 592382 500378 592618 500614
rect 592062 500058 592298 500294
rect 592382 500058 592618 500294
rect 592062 464378 592298 464614
rect 592382 464378 592618 464614
rect 592062 464058 592298 464294
rect 592382 464058 592618 464294
rect 592062 428378 592298 428614
rect 592382 428378 592618 428614
rect 592062 428058 592298 428294
rect 592382 428058 592618 428294
rect 592062 392378 592298 392614
rect 592382 392378 592618 392614
rect 592062 392058 592298 392294
rect 592382 392058 592618 392294
rect 592062 356378 592298 356614
rect 592382 356378 592618 356614
rect 592062 356058 592298 356294
rect 592382 356058 592618 356294
rect 592062 320378 592298 320614
rect 592382 320378 592618 320614
rect 592062 320058 592298 320294
rect 592382 320058 592618 320294
rect 592062 284378 592298 284614
rect 592382 284378 592618 284614
rect 592062 284058 592298 284294
rect 592382 284058 592618 284294
rect 592062 248378 592298 248614
rect 592382 248378 592618 248614
rect 592062 248058 592298 248294
rect 592382 248058 592618 248294
rect 592062 212378 592298 212614
rect 592382 212378 592618 212614
rect 592062 212058 592298 212294
rect 592382 212058 592618 212294
rect 592062 176378 592298 176614
rect 592382 176378 592618 176614
rect 592062 176058 592298 176294
rect 592382 176058 592618 176294
rect 592062 140378 592298 140614
rect 592382 140378 592618 140614
rect 592062 140058 592298 140294
rect 592382 140058 592618 140294
rect 592062 104378 592298 104614
rect 592382 104378 592618 104614
rect 592062 104058 592298 104294
rect 592382 104058 592618 104294
rect 592062 68378 592298 68614
rect 592382 68378 592618 68614
rect 592062 68058 592298 68294
rect 592382 68058 592618 68294
rect 592062 32378 592298 32614
rect 592382 32378 592618 32614
rect 592062 32058 592298 32294
rect 592382 32058 592618 32294
rect 570986 -7302 571222 -7066
rect 571306 -7302 571542 -7066
rect 570986 -7622 571222 -7386
rect 571306 -7622 571542 -7386
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 592650 698294
rect -8726 698026 592650 698058
rect -6806 694894 590730 694926
rect -6806 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 590730 694894
rect -6806 694574 590730 694658
rect -6806 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 590730 694574
rect -6806 694306 590730 694338
rect -4886 691174 588810 691206
rect -4886 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 588810 691174
rect -4886 690854 588810 690938
rect -4886 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 588810 690854
rect -4886 690586 588810 690618
rect -2966 687454 586890 687486
rect -2966 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 586890 687454
rect -2966 687134 586890 687218
rect -2966 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 586890 687134
rect -2966 686866 586890 686898
rect -8726 680614 592650 680646
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect -8726 680294 592650 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect -8726 680026 592650 680058
rect -6806 676894 590730 676926
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect -6806 676574 590730 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect -6806 676306 590730 676338
rect -4886 673174 588810 673206
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect -4886 672854 588810 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect -4886 672586 588810 672618
rect -2966 669454 586890 669486
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect -2966 669134 586890 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect -2966 668866 586890 668898
rect -8726 662614 592650 662646
rect -8726 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 592650 662294
rect -8726 662026 592650 662058
rect -6806 658894 590730 658926
rect -6806 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 590730 658894
rect -6806 658574 590730 658658
rect -6806 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 590730 658574
rect -6806 658306 590730 658338
rect -4886 655174 588810 655206
rect -4886 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 588810 655174
rect -4886 654854 588810 654938
rect -4886 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 588810 654854
rect -4886 654586 588810 654618
rect -2966 651454 586890 651486
rect -2966 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 586890 651454
rect -2966 651134 586890 651218
rect -2966 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 586890 651134
rect -2966 650866 586890 650898
rect -8726 644614 592650 644646
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect -8726 644294 592650 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect -8726 644026 592650 644058
rect -6806 640894 590730 640926
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect -6806 640574 590730 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect -6806 640306 590730 640338
rect -4886 637174 588810 637206
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect -4886 636854 588810 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect -4886 636586 588810 636618
rect -2966 633454 586890 633486
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect -2966 633134 586890 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect -2966 632866 586890 632898
rect -8726 626614 592650 626646
rect -8726 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 592650 626294
rect -8726 626026 592650 626058
rect -6806 622894 590730 622926
rect -6806 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 590730 622894
rect -6806 622574 590730 622658
rect -6806 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 590730 622574
rect -6806 622306 590730 622338
rect -4886 619174 588810 619206
rect -4886 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 588810 619174
rect -4886 618854 588810 618938
rect -4886 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 588810 618854
rect -4886 618586 588810 618618
rect -2966 615454 586890 615486
rect -2966 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 586890 615454
rect -2966 615134 586890 615218
rect -2966 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 586890 615134
rect -2966 614866 586890 614898
rect -8726 608614 592650 608646
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect -8726 608294 592650 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect -8726 608026 592650 608058
rect -6806 604894 590730 604926
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect -6806 604574 590730 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect -6806 604306 590730 604338
rect -4886 601174 588810 601206
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect -4886 600854 588810 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect -4886 600586 588810 600618
rect -2966 597454 586890 597486
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect -2966 597134 586890 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect -2966 596866 586890 596898
rect -8726 590614 592650 590646
rect -8726 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 592650 590294
rect -8726 590026 592650 590058
rect -6806 586894 590730 586926
rect -6806 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 590730 586894
rect -6806 586574 590730 586658
rect -6806 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 590730 586574
rect -6806 586306 590730 586338
rect -4886 583174 588810 583206
rect -4886 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 77546 583174
rect 77782 582938 77866 583174
rect 78102 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 588810 583174
rect -4886 582854 588810 582938
rect -4886 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 77546 582854
rect 77782 582618 77866 582854
rect 78102 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 588810 582854
rect -4886 582586 588810 582618
rect -2966 579454 586890 579486
rect -2966 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 586890 579454
rect -2966 579134 586890 579218
rect -2966 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 586890 579134
rect -2966 578866 586890 578898
rect -8726 572614 592650 572646
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect -8726 572294 592650 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect -8726 572026 592650 572058
rect -6806 568894 590730 568926
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect -6806 568574 590730 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect -6806 568306 590730 568338
rect -4886 565174 588810 565206
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 95546 565174
rect 95782 564938 95866 565174
rect 96102 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect -4886 564854 588810 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 95546 564854
rect 95782 564618 95866 564854
rect 96102 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect -4886 564586 588810 564618
rect -2966 561454 586890 561486
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect -2966 561134 586890 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect -2966 560866 586890 560898
rect -8726 554614 592650 554646
rect -8726 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 84986 554614
rect 85222 554378 85306 554614
rect 85542 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 84986 554294
rect 85222 554058 85306 554294
rect 85542 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 592650 554294
rect -8726 554026 592650 554058
rect -6806 550894 590730 550926
rect -6806 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 81266 550894
rect 81502 550658 81586 550894
rect 81822 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 590730 550894
rect -6806 550574 590730 550658
rect -6806 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 81266 550574
rect 81502 550338 81586 550574
rect 81822 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 590730 550574
rect -6806 550306 590730 550338
rect -4886 547174 588810 547206
rect -4886 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 77546 547174
rect 77782 546938 77866 547174
rect 78102 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 588810 547174
rect -4886 546854 588810 546938
rect -4886 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 77546 546854
rect 77782 546618 77866 546854
rect 78102 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 588810 546854
rect -4886 546586 588810 546618
rect -2966 543454 586890 543486
rect -2966 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 586890 543454
rect -2966 543134 586890 543218
rect -2966 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 586890 543134
rect -2966 542866 586890 542898
rect -8726 536614 592650 536646
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 174986 536614
rect 175222 536378 175306 536614
rect 175542 536378 210986 536614
rect 211222 536378 211306 536614
rect 211542 536378 246986 536614
rect 247222 536378 247306 536614
rect 247542 536378 282986 536614
rect 283222 536378 283306 536614
rect 283542 536378 318986 536614
rect 319222 536378 319306 536614
rect 319542 536378 354986 536614
rect 355222 536378 355306 536614
rect 355542 536378 390986 536614
rect 391222 536378 391306 536614
rect 391542 536378 426986 536614
rect 427222 536378 427306 536614
rect 427542 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect -8726 536294 592650 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 174986 536294
rect 175222 536058 175306 536294
rect 175542 536058 210986 536294
rect 211222 536058 211306 536294
rect 211542 536058 246986 536294
rect 247222 536058 247306 536294
rect 247542 536058 282986 536294
rect 283222 536058 283306 536294
rect 283542 536058 318986 536294
rect 319222 536058 319306 536294
rect 319542 536058 354986 536294
rect 355222 536058 355306 536294
rect 355542 536058 390986 536294
rect 391222 536058 391306 536294
rect 391542 536058 426986 536294
rect 427222 536058 427306 536294
rect 427542 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect -8726 536026 592650 536058
rect -6806 532894 590730 532926
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 171266 532894
rect 171502 532658 171586 532894
rect 171822 532658 207266 532894
rect 207502 532658 207586 532894
rect 207822 532658 243266 532894
rect 243502 532658 243586 532894
rect 243822 532658 279266 532894
rect 279502 532658 279586 532894
rect 279822 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 351266 532894
rect 351502 532658 351586 532894
rect 351822 532658 387266 532894
rect 387502 532658 387586 532894
rect 387822 532658 423266 532894
rect 423502 532658 423586 532894
rect 423822 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect -6806 532574 590730 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 171266 532574
rect 171502 532338 171586 532574
rect 171822 532338 207266 532574
rect 207502 532338 207586 532574
rect 207822 532338 243266 532574
rect 243502 532338 243586 532574
rect 243822 532338 279266 532574
rect 279502 532338 279586 532574
rect 279822 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 351266 532574
rect 351502 532338 351586 532574
rect 351822 532338 387266 532574
rect 387502 532338 387586 532574
rect 387822 532338 423266 532574
rect 423502 532338 423586 532574
rect 423822 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect -6806 532306 590730 532338
rect -4886 529174 588810 529206
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 167546 529174
rect 167782 528938 167866 529174
rect 168102 528938 203546 529174
rect 203782 528938 203866 529174
rect 204102 528938 239546 529174
rect 239782 528938 239866 529174
rect 240102 528938 275546 529174
rect 275782 528938 275866 529174
rect 276102 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 347546 529174
rect 347782 528938 347866 529174
rect 348102 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 419546 529174
rect 419782 528938 419866 529174
rect 420102 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect -4886 528854 588810 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 167546 528854
rect 167782 528618 167866 528854
rect 168102 528618 203546 528854
rect 203782 528618 203866 528854
rect 204102 528618 239546 528854
rect 239782 528618 239866 528854
rect 240102 528618 275546 528854
rect 275782 528618 275866 528854
rect 276102 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 347546 528854
rect 347782 528618 347866 528854
rect 348102 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 419546 528854
rect 419782 528618 419866 528854
rect 420102 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect -4886 528586 588810 528618
rect -2966 525454 586890 525486
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect -2966 525134 586890 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect -2966 524866 586890 524898
rect -8726 518614 592650 518646
rect -8726 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 592650 518294
rect -8726 518026 592650 518058
rect -6806 514894 590730 514926
rect -6806 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 590730 514894
rect -6806 514574 590730 514658
rect -6806 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 590730 514574
rect -6806 514306 590730 514338
rect -4886 511174 588810 511206
rect -4886 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 588810 511174
rect -4886 510854 588810 510938
rect -4886 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 588810 510854
rect -4886 510586 588810 510618
rect -2966 507454 586890 507486
rect -2966 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 586890 507454
rect -2966 507134 586890 507218
rect -2966 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 586890 507134
rect -2966 506866 586890 506898
rect -8726 500614 592650 500646
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 138986 500614
rect 139222 500378 139306 500614
rect 139542 500378 174986 500614
rect 175222 500378 175306 500614
rect 175542 500378 210986 500614
rect 211222 500378 211306 500614
rect 211542 500378 246986 500614
rect 247222 500378 247306 500614
rect 247542 500378 282986 500614
rect 283222 500378 283306 500614
rect 283542 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect -8726 500294 592650 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 138986 500294
rect 139222 500058 139306 500294
rect 139542 500058 174986 500294
rect 175222 500058 175306 500294
rect 175542 500058 210986 500294
rect 211222 500058 211306 500294
rect 211542 500058 246986 500294
rect 247222 500058 247306 500294
rect 247542 500058 282986 500294
rect 283222 500058 283306 500294
rect 283542 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect -8726 500026 592650 500058
rect -6806 496894 590730 496926
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 171266 496894
rect 171502 496658 171586 496894
rect 171822 496658 207266 496894
rect 207502 496658 207586 496894
rect 207822 496658 243266 496894
rect 243502 496658 243586 496894
rect 243822 496658 279266 496894
rect 279502 496658 279586 496894
rect 279822 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect -6806 496574 590730 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 171266 496574
rect 171502 496338 171586 496574
rect 171822 496338 207266 496574
rect 207502 496338 207586 496574
rect 207822 496338 243266 496574
rect 243502 496338 243586 496574
rect 243822 496338 279266 496574
rect 279502 496338 279586 496574
rect 279822 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect -6806 496306 590730 496338
rect -4886 493174 588810 493206
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 167546 493174
rect 167782 492938 167866 493174
rect 168102 492938 203546 493174
rect 203782 492938 203866 493174
rect 204102 492938 239546 493174
rect 239782 492938 239866 493174
rect 240102 492938 275546 493174
rect 275782 492938 275866 493174
rect 276102 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect -4886 492854 588810 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 167546 492854
rect 167782 492618 167866 492854
rect 168102 492618 203546 492854
rect 203782 492618 203866 492854
rect 204102 492618 239546 492854
rect 239782 492618 239866 492854
rect 240102 492618 275546 492854
rect 275782 492618 275866 492854
rect 276102 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect -4886 492586 588810 492618
rect -2966 489454 586890 489486
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect -2966 489134 586890 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect -2966 488866 586890 488898
rect -8726 482614 592650 482646
rect -8726 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 592650 482294
rect -8726 482026 592650 482058
rect -6806 478894 590730 478926
rect -6806 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 590730 478894
rect -6806 478574 590730 478658
rect -6806 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 590730 478574
rect -6806 478306 590730 478338
rect -4886 475174 588810 475206
rect -4886 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 588810 475174
rect -4886 474854 588810 474938
rect -4886 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 588810 474854
rect -4886 474586 588810 474618
rect -2966 471454 586890 471486
rect -2966 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 586890 471454
rect -2966 471134 586890 471218
rect -2966 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 586890 471134
rect -2966 470866 586890 470898
rect -8726 464614 592650 464646
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 102986 464614
rect 103222 464378 103306 464614
rect 103542 464378 138986 464614
rect 139222 464378 139306 464614
rect 139542 464378 174986 464614
rect 175222 464378 175306 464614
rect 175542 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 246986 464614
rect 247222 464378 247306 464614
rect 247542 464378 282986 464614
rect 283222 464378 283306 464614
rect 283542 464378 318986 464614
rect 319222 464378 319306 464614
rect 319542 464378 354986 464614
rect 355222 464378 355306 464614
rect 355542 464378 390986 464614
rect 391222 464378 391306 464614
rect 391542 464378 426986 464614
rect 427222 464378 427306 464614
rect 427542 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect -8726 464294 592650 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 102986 464294
rect 103222 464058 103306 464294
rect 103542 464058 138986 464294
rect 139222 464058 139306 464294
rect 139542 464058 174986 464294
rect 175222 464058 175306 464294
rect 175542 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 246986 464294
rect 247222 464058 247306 464294
rect 247542 464058 282986 464294
rect 283222 464058 283306 464294
rect 283542 464058 318986 464294
rect 319222 464058 319306 464294
rect 319542 464058 354986 464294
rect 355222 464058 355306 464294
rect 355542 464058 390986 464294
rect 391222 464058 391306 464294
rect 391542 464058 426986 464294
rect 427222 464058 427306 464294
rect 427542 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect -8726 464026 592650 464058
rect -6806 460894 590730 460926
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 99266 460894
rect 99502 460658 99586 460894
rect 99822 460658 135266 460894
rect 135502 460658 135586 460894
rect 135822 460658 171266 460894
rect 171502 460658 171586 460894
rect 171822 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 243266 460894
rect 243502 460658 243586 460894
rect 243822 460658 279266 460894
rect 279502 460658 279586 460894
rect 279822 460658 315266 460894
rect 315502 460658 315586 460894
rect 315822 460658 351266 460894
rect 351502 460658 351586 460894
rect 351822 460658 387266 460894
rect 387502 460658 387586 460894
rect 387822 460658 423266 460894
rect 423502 460658 423586 460894
rect 423822 460658 459266 460894
rect 459502 460658 459586 460894
rect 459822 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect -6806 460574 590730 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 99266 460574
rect 99502 460338 99586 460574
rect 99822 460338 135266 460574
rect 135502 460338 135586 460574
rect 135822 460338 171266 460574
rect 171502 460338 171586 460574
rect 171822 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 243266 460574
rect 243502 460338 243586 460574
rect 243822 460338 279266 460574
rect 279502 460338 279586 460574
rect 279822 460338 315266 460574
rect 315502 460338 315586 460574
rect 315822 460338 351266 460574
rect 351502 460338 351586 460574
rect 351822 460338 387266 460574
rect 387502 460338 387586 460574
rect 387822 460338 423266 460574
rect 423502 460338 423586 460574
rect 423822 460338 459266 460574
rect 459502 460338 459586 460574
rect 459822 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect -6806 460306 590730 460338
rect -4886 457174 588810 457206
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 95546 457174
rect 95782 456938 95866 457174
rect 96102 456938 131546 457174
rect 131782 456938 131866 457174
rect 132102 456938 167546 457174
rect 167782 456938 167866 457174
rect 168102 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 239546 457174
rect 239782 456938 239866 457174
rect 240102 456938 275546 457174
rect 275782 456938 275866 457174
rect 276102 456938 311546 457174
rect 311782 456938 311866 457174
rect 312102 456938 347546 457174
rect 347782 456938 347866 457174
rect 348102 456938 383546 457174
rect 383782 456938 383866 457174
rect 384102 456938 419546 457174
rect 419782 456938 419866 457174
rect 420102 456938 455546 457174
rect 455782 456938 455866 457174
rect 456102 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect -4886 456854 588810 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 95546 456854
rect 95782 456618 95866 456854
rect 96102 456618 131546 456854
rect 131782 456618 131866 456854
rect 132102 456618 167546 456854
rect 167782 456618 167866 456854
rect 168102 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 239546 456854
rect 239782 456618 239866 456854
rect 240102 456618 275546 456854
rect 275782 456618 275866 456854
rect 276102 456618 311546 456854
rect 311782 456618 311866 456854
rect 312102 456618 347546 456854
rect 347782 456618 347866 456854
rect 348102 456618 383546 456854
rect 383782 456618 383866 456854
rect 384102 456618 419546 456854
rect 419782 456618 419866 456854
rect 420102 456618 455546 456854
rect 455782 456618 455866 456854
rect 456102 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect -4886 456586 588810 456618
rect -2966 453454 586890 453486
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect -2966 453134 586890 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect -2966 452866 586890 452898
rect -8726 446614 592650 446646
rect -8726 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 84986 446614
rect 85222 446378 85306 446614
rect 85542 446378 120986 446614
rect 121222 446378 121306 446614
rect 121542 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 192986 446614
rect 193222 446378 193306 446614
rect 193542 446378 228986 446614
rect 229222 446378 229306 446614
rect 229542 446378 264986 446614
rect 265222 446378 265306 446614
rect 265542 446378 300986 446614
rect 301222 446378 301306 446614
rect 301542 446378 336986 446614
rect 337222 446378 337306 446614
rect 337542 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 84986 446294
rect 85222 446058 85306 446294
rect 85542 446058 120986 446294
rect 121222 446058 121306 446294
rect 121542 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 192986 446294
rect 193222 446058 193306 446294
rect 193542 446058 228986 446294
rect 229222 446058 229306 446294
rect 229542 446058 264986 446294
rect 265222 446058 265306 446294
rect 265542 446058 300986 446294
rect 301222 446058 301306 446294
rect 301542 446058 336986 446294
rect 337222 446058 337306 446294
rect 337542 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 592650 446294
rect -8726 446026 592650 446058
rect -6806 442894 590730 442926
rect -6806 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 81266 442894
rect 81502 442658 81586 442894
rect 81822 442658 117266 442894
rect 117502 442658 117586 442894
rect 117822 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 225266 442894
rect 225502 442658 225586 442894
rect 225822 442658 261266 442894
rect 261502 442658 261586 442894
rect 261822 442658 297266 442894
rect 297502 442658 297586 442894
rect 297822 442658 333266 442894
rect 333502 442658 333586 442894
rect 333822 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 441266 442894
rect 441502 442658 441586 442894
rect 441822 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 590730 442894
rect -6806 442574 590730 442658
rect -6806 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 81266 442574
rect 81502 442338 81586 442574
rect 81822 442338 117266 442574
rect 117502 442338 117586 442574
rect 117822 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 225266 442574
rect 225502 442338 225586 442574
rect 225822 442338 261266 442574
rect 261502 442338 261586 442574
rect 261822 442338 297266 442574
rect 297502 442338 297586 442574
rect 297822 442338 333266 442574
rect 333502 442338 333586 442574
rect 333822 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 441266 442574
rect 441502 442338 441586 442574
rect 441822 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 590730 442574
rect -6806 442306 590730 442338
rect -4886 439174 588810 439206
rect -4886 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 77546 439174
rect 77782 438938 77866 439174
rect 78102 438938 113546 439174
rect 113782 438938 113866 439174
rect 114102 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 221546 439174
rect 221782 438938 221866 439174
rect 222102 438938 257546 439174
rect 257782 438938 257866 439174
rect 258102 438938 293546 439174
rect 293782 438938 293866 439174
rect 294102 438938 329546 439174
rect 329782 438938 329866 439174
rect 330102 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 588810 439174
rect -4886 438854 588810 438938
rect -4886 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 77546 438854
rect 77782 438618 77866 438854
rect 78102 438618 113546 438854
rect 113782 438618 113866 438854
rect 114102 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 221546 438854
rect 221782 438618 221866 438854
rect 222102 438618 257546 438854
rect 257782 438618 257866 438854
rect 258102 438618 293546 438854
rect 293782 438618 293866 438854
rect 294102 438618 329546 438854
rect 329782 438618 329866 438854
rect 330102 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 588810 438854
rect -4886 438586 588810 438618
rect -2966 435454 586890 435486
rect -2966 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 586890 435454
rect -2966 435134 586890 435218
rect -2966 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 586890 435134
rect -2966 434866 586890 434898
rect -8726 428614 592650 428646
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 66986 428614
rect 67222 428378 67306 428614
rect 67542 428378 102986 428614
rect 103222 428378 103306 428614
rect 103542 428378 138986 428614
rect 139222 428378 139306 428614
rect 139542 428378 174986 428614
rect 175222 428378 175306 428614
rect 175542 428378 210986 428614
rect 211222 428378 211306 428614
rect 211542 428378 246986 428614
rect 247222 428378 247306 428614
rect 247542 428378 282986 428614
rect 283222 428378 283306 428614
rect 283542 428378 318986 428614
rect 319222 428378 319306 428614
rect 319542 428378 354986 428614
rect 355222 428378 355306 428614
rect 355542 428378 390986 428614
rect 391222 428378 391306 428614
rect 391542 428378 426986 428614
rect 427222 428378 427306 428614
rect 427542 428378 462986 428614
rect 463222 428378 463306 428614
rect 463542 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect -8726 428294 592650 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 66986 428294
rect 67222 428058 67306 428294
rect 67542 428058 102986 428294
rect 103222 428058 103306 428294
rect 103542 428058 138986 428294
rect 139222 428058 139306 428294
rect 139542 428058 174986 428294
rect 175222 428058 175306 428294
rect 175542 428058 210986 428294
rect 211222 428058 211306 428294
rect 211542 428058 246986 428294
rect 247222 428058 247306 428294
rect 247542 428058 282986 428294
rect 283222 428058 283306 428294
rect 283542 428058 318986 428294
rect 319222 428058 319306 428294
rect 319542 428058 354986 428294
rect 355222 428058 355306 428294
rect 355542 428058 390986 428294
rect 391222 428058 391306 428294
rect 391542 428058 426986 428294
rect 427222 428058 427306 428294
rect 427542 428058 462986 428294
rect 463222 428058 463306 428294
rect 463542 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect -8726 428026 592650 428058
rect -6806 424894 590730 424926
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 99266 424894
rect 99502 424658 99586 424894
rect 99822 424658 135266 424894
rect 135502 424658 135586 424894
rect 135822 424658 171266 424894
rect 171502 424658 171586 424894
rect 171822 424658 207266 424894
rect 207502 424658 207586 424894
rect 207822 424658 243266 424894
rect 243502 424658 243586 424894
rect 243822 424658 279266 424894
rect 279502 424658 279586 424894
rect 279822 424658 315266 424894
rect 315502 424658 315586 424894
rect 315822 424658 351266 424894
rect 351502 424658 351586 424894
rect 351822 424658 387266 424894
rect 387502 424658 387586 424894
rect 387822 424658 423266 424894
rect 423502 424658 423586 424894
rect 423822 424658 459266 424894
rect 459502 424658 459586 424894
rect 459822 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect -6806 424574 590730 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 99266 424574
rect 99502 424338 99586 424574
rect 99822 424338 135266 424574
rect 135502 424338 135586 424574
rect 135822 424338 171266 424574
rect 171502 424338 171586 424574
rect 171822 424338 207266 424574
rect 207502 424338 207586 424574
rect 207822 424338 243266 424574
rect 243502 424338 243586 424574
rect 243822 424338 279266 424574
rect 279502 424338 279586 424574
rect 279822 424338 315266 424574
rect 315502 424338 315586 424574
rect 315822 424338 351266 424574
rect 351502 424338 351586 424574
rect 351822 424338 387266 424574
rect 387502 424338 387586 424574
rect 387822 424338 423266 424574
rect 423502 424338 423586 424574
rect 423822 424338 459266 424574
rect 459502 424338 459586 424574
rect 459822 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect -6806 424306 590730 424338
rect -4886 421174 588810 421206
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 95546 421174
rect 95782 420938 95866 421174
rect 96102 420938 131546 421174
rect 131782 420938 131866 421174
rect 132102 420938 167546 421174
rect 167782 420938 167866 421174
rect 168102 420938 203546 421174
rect 203782 420938 203866 421174
rect 204102 420938 239546 421174
rect 239782 420938 239866 421174
rect 240102 420938 275546 421174
rect 275782 420938 275866 421174
rect 276102 420938 311546 421174
rect 311782 420938 311866 421174
rect 312102 420938 347546 421174
rect 347782 420938 347866 421174
rect 348102 420938 383546 421174
rect 383782 420938 383866 421174
rect 384102 420938 419546 421174
rect 419782 420938 419866 421174
rect 420102 420938 455546 421174
rect 455782 420938 455866 421174
rect 456102 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect -4886 420854 588810 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 95546 420854
rect 95782 420618 95866 420854
rect 96102 420618 131546 420854
rect 131782 420618 131866 420854
rect 132102 420618 167546 420854
rect 167782 420618 167866 420854
rect 168102 420618 203546 420854
rect 203782 420618 203866 420854
rect 204102 420618 239546 420854
rect 239782 420618 239866 420854
rect 240102 420618 275546 420854
rect 275782 420618 275866 420854
rect 276102 420618 311546 420854
rect 311782 420618 311866 420854
rect 312102 420618 347546 420854
rect 347782 420618 347866 420854
rect 348102 420618 383546 420854
rect 383782 420618 383866 420854
rect 384102 420618 419546 420854
rect 419782 420618 419866 420854
rect 420102 420618 455546 420854
rect 455782 420618 455866 420854
rect 456102 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect -4886 420586 588810 420618
rect -2966 417454 586890 417486
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect -2966 417134 586890 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect -2966 416866 586890 416898
rect -8726 410614 592650 410646
rect -8726 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 84986 410614
rect 85222 410378 85306 410614
rect 85542 410378 120986 410614
rect 121222 410378 121306 410614
rect 121542 410378 156986 410614
rect 157222 410378 157306 410614
rect 157542 410378 192986 410614
rect 193222 410378 193306 410614
rect 193542 410378 228986 410614
rect 229222 410378 229306 410614
rect 229542 410378 264986 410614
rect 265222 410378 265306 410614
rect 265542 410378 300986 410614
rect 301222 410378 301306 410614
rect 301542 410378 336986 410614
rect 337222 410378 337306 410614
rect 337542 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 84986 410294
rect 85222 410058 85306 410294
rect 85542 410058 120986 410294
rect 121222 410058 121306 410294
rect 121542 410058 156986 410294
rect 157222 410058 157306 410294
rect 157542 410058 192986 410294
rect 193222 410058 193306 410294
rect 193542 410058 228986 410294
rect 229222 410058 229306 410294
rect 229542 410058 264986 410294
rect 265222 410058 265306 410294
rect 265542 410058 300986 410294
rect 301222 410058 301306 410294
rect 301542 410058 336986 410294
rect 337222 410058 337306 410294
rect 337542 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 592650 410294
rect -8726 410026 592650 410058
rect -6806 406894 590730 406926
rect -6806 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 81266 406894
rect 81502 406658 81586 406894
rect 81822 406658 117266 406894
rect 117502 406658 117586 406894
rect 117822 406658 153266 406894
rect 153502 406658 153586 406894
rect 153822 406658 189266 406894
rect 189502 406658 189586 406894
rect 189822 406658 225266 406894
rect 225502 406658 225586 406894
rect 225822 406658 261266 406894
rect 261502 406658 261586 406894
rect 261822 406658 297266 406894
rect 297502 406658 297586 406894
rect 297822 406658 333266 406894
rect 333502 406658 333586 406894
rect 333822 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 590730 406894
rect -6806 406574 590730 406658
rect -6806 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 81266 406574
rect 81502 406338 81586 406574
rect 81822 406338 117266 406574
rect 117502 406338 117586 406574
rect 117822 406338 153266 406574
rect 153502 406338 153586 406574
rect 153822 406338 189266 406574
rect 189502 406338 189586 406574
rect 189822 406338 225266 406574
rect 225502 406338 225586 406574
rect 225822 406338 261266 406574
rect 261502 406338 261586 406574
rect 261822 406338 297266 406574
rect 297502 406338 297586 406574
rect 297822 406338 333266 406574
rect 333502 406338 333586 406574
rect 333822 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 590730 406574
rect -6806 406306 590730 406338
rect -4886 403174 588810 403206
rect -4886 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 77546 403174
rect 77782 402938 77866 403174
rect 78102 402938 113546 403174
rect 113782 402938 113866 403174
rect 114102 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 185546 403174
rect 185782 402938 185866 403174
rect 186102 402938 221546 403174
rect 221782 402938 221866 403174
rect 222102 402938 257546 403174
rect 257782 402938 257866 403174
rect 258102 402938 293546 403174
rect 293782 402938 293866 403174
rect 294102 402938 329546 403174
rect 329782 402938 329866 403174
rect 330102 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 588810 403174
rect -4886 402854 588810 402938
rect -4886 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 77546 402854
rect 77782 402618 77866 402854
rect 78102 402618 113546 402854
rect 113782 402618 113866 402854
rect 114102 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 185546 402854
rect 185782 402618 185866 402854
rect 186102 402618 221546 402854
rect 221782 402618 221866 402854
rect 222102 402618 257546 402854
rect 257782 402618 257866 402854
rect 258102 402618 293546 402854
rect 293782 402618 293866 402854
rect 294102 402618 329546 402854
rect 329782 402618 329866 402854
rect 330102 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 588810 402854
rect -4886 402586 588810 402618
rect -2966 399454 586890 399486
rect -2966 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 586890 399454
rect -2966 399134 586890 399218
rect -2966 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 586890 399134
rect -2966 398866 586890 398898
rect -8726 392614 592650 392646
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 66986 392614
rect 67222 392378 67306 392614
rect 67542 392378 102986 392614
rect 103222 392378 103306 392614
rect 103542 392378 138986 392614
rect 139222 392378 139306 392614
rect 139542 392378 174986 392614
rect 175222 392378 175306 392614
rect 175542 392378 210986 392614
rect 211222 392378 211306 392614
rect 211542 392378 246986 392614
rect 247222 392378 247306 392614
rect 247542 392378 282986 392614
rect 283222 392378 283306 392614
rect 283542 392378 318986 392614
rect 319222 392378 319306 392614
rect 319542 392378 354986 392614
rect 355222 392378 355306 392614
rect 355542 392378 390986 392614
rect 391222 392378 391306 392614
rect 391542 392378 426986 392614
rect 427222 392378 427306 392614
rect 427542 392378 462986 392614
rect 463222 392378 463306 392614
rect 463542 392378 498986 392614
rect 499222 392378 499306 392614
rect 499542 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect -8726 392294 592650 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 66986 392294
rect 67222 392058 67306 392294
rect 67542 392058 102986 392294
rect 103222 392058 103306 392294
rect 103542 392058 138986 392294
rect 139222 392058 139306 392294
rect 139542 392058 174986 392294
rect 175222 392058 175306 392294
rect 175542 392058 210986 392294
rect 211222 392058 211306 392294
rect 211542 392058 246986 392294
rect 247222 392058 247306 392294
rect 247542 392058 282986 392294
rect 283222 392058 283306 392294
rect 283542 392058 318986 392294
rect 319222 392058 319306 392294
rect 319542 392058 354986 392294
rect 355222 392058 355306 392294
rect 355542 392058 390986 392294
rect 391222 392058 391306 392294
rect 391542 392058 426986 392294
rect 427222 392058 427306 392294
rect 427542 392058 462986 392294
rect 463222 392058 463306 392294
rect 463542 392058 498986 392294
rect 499222 392058 499306 392294
rect 499542 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect -8726 392026 592650 392058
rect -6806 388894 590730 388926
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 99266 388894
rect 99502 388658 99586 388894
rect 99822 388658 135266 388894
rect 135502 388658 135586 388894
rect 135822 388658 171266 388894
rect 171502 388658 171586 388894
rect 171822 388658 207266 388894
rect 207502 388658 207586 388894
rect 207822 388658 243266 388894
rect 243502 388658 243586 388894
rect 243822 388658 279266 388894
rect 279502 388658 279586 388894
rect 279822 388658 315266 388894
rect 315502 388658 315586 388894
rect 315822 388658 351266 388894
rect 351502 388658 351586 388894
rect 351822 388658 387266 388894
rect 387502 388658 387586 388894
rect 387822 388658 423266 388894
rect 423502 388658 423586 388894
rect 423822 388658 459266 388894
rect 459502 388658 459586 388894
rect 459822 388658 495266 388894
rect 495502 388658 495586 388894
rect 495822 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect -6806 388574 590730 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 99266 388574
rect 99502 388338 99586 388574
rect 99822 388338 135266 388574
rect 135502 388338 135586 388574
rect 135822 388338 171266 388574
rect 171502 388338 171586 388574
rect 171822 388338 207266 388574
rect 207502 388338 207586 388574
rect 207822 388338 243266 388574
rect 243502 388338 243586 388574
rect 243822 388338 279266 388574
rect 279502 388338 279586 388574
rect 279822 388338 315266 388574
rect 315502 388338 315586 388574
rect 315822 388338 351266 388574
rect 351502 388338 351586 388574
rect 351822 388338 387266 388574
rect 387502 388338 387586 388574
rect 387822 388338 423266 388574
rect 423502 388338 423586 388574
rect 423822 388338 459266 388574
rect 459502 388338 459586 388574
rect 459822 388338 495266 388574
rect 495502 388338 495586 388574
rect 495822 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect -6806 388306 590730 388338
rect -4886 385174 588810 385206
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 59546 385174
rect 59782 384938 59866 385174
rect 60102 384938 95546 385174
rect 95782 384938 95866 385174
rect 96102 384938 131546 385174
rect 131782 384938 131866 385174
rect 132102 384938 167546 385174
rect 167782 384938 167866 385174
rect 168102 384938 203546 385174
rect 203782 384938 203866 385174
rect 204102 384938 239546 385174
rect 239782 384938 239866 385174
rect 240102 384938 275546 385174
rect 275782 384938 275866 385174
rect 276102 384938 311546 385174
rect 311782 384938 311866 385174
rect 312102 384938 347546 385174
rect 347782 384938 347866 385174
rect 348102 384938 383546 385174
rect 383782 384938 383866 385174
rect 384102 384938 419546 385174
rect 419782 384938 419866 385174
rect 420102 384938 455546 385174
rect 455782 384938 455866 385174
rect 456102 384938 491546 385174
rect 491782 384938 491866 385174
rect 492102 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect -4886 384854 588810 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 59546 384854
rect 59782 384618 59866 384854
rect 60102 384618 95546 384854
rect 95782 384618 95866 384854
rect 96102 384618 131546 384854
rect 131782 384618 131866 384854
rect 132102 384618 167546 384854
rect 167782 384618 167866 384854
rect 168102 384618 203546 384854
rect 203782 384618 203866 384854
rect 204102 384618 239546 384854
rect 239782 384618 239866 384854
rect 240102 384618 275546 384854
rect 275782 384618 275866 384854
rect 276102 384618 311546 384854
rect 311782 384618 311866 384854
rect 312102 384618 347546 384854
rect 347782 384618 347866 384854
rect 348102 384618 383546 384854
rect 383782 384618 383866 384854
rect 384102 384618 419546 384854
rect 419782 384618 419866 384854
rect 420102 384618 455546 384854
rect 455782 384618 455866 384854
rect 456102 384618 491546 384854
rect 491782 384618 491866 384854
rect 492102 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect -4886 384586 588810 384618
rect -2966 381454 586890 381486
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect -2966 381134 586890 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect -2966 380866 586890 380898
rect -8726 374614 592650 374646
rect -8726 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 264986 374614
rect 265222 374378 265306 374614
rect 265542 374378 300986 374614
rect 301222 374378 301306 374614
rect 301542 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 264986 374294
rect 265222 374058 265306 374294
rect 265542 374058 300986 374294
rect 301222 374058 301306 374294
rect 301542 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 592650 374294
rect -8726 374026 592650 374058
rect -6806 370894 590730 370926
rect -6806 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 261266 370894
rect 261502 370658 261586 370894
rect 261822 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 590730 370894
rect -6806 370574 590730 370658
rect -6806 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 261266 370574
rect 261502 370338 261586 370574
rect 261822 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 590730 370574
rect -6806 370306 590730 370338
rect -4886 367174 588810 367206
rect -4886 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 257546 367174
rect 257782 366938 257866 367174
rect 258102 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 588810 367174
rect -4886 366854 588810 366938
rect -4886 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 257546 366854
rect 257782 366618 257866 366854
rect 258102 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 588810 366854
rect -4886 366586 588810 366618
rect -2966 363454 586890 363486
rect -2966 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 586890 363454
rect -2966 363134 586890 363218
rect -2966 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 586890 363134
rect -2966 362866 586890 362898
rect -8726 356614 592650 356646
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 102986 356614
rect 103222 356378 103306 356614
rect 103542 356378 138986 356614
rect 139222 356378 139306 356614
rect 139542 356378 174986 356614
rect 175222 356378 175306 356614
rect 175542 356378 210986 356614
rect 211222 356378 211306 356614
rect 211542 356378 246986 356614
rect 247222 356378 247306 356614
rect 247542 356378 282986 356614
rect 283222 356378 283306 356614
rect 283542 356378 318986 356614
rect 319222 356378 319306 356614
rect 319542 356378 354986 356614
rect 355222 356378 355306 356614
rect 355542 356378 390986 356614
rect 391222 356378 391306 356614
rect 391542 356378 426986 356614
rect 427222 356378 427306 356614
rect 427542 356378 462986 356614
rect 463222 356378 463306 356614
rect 463542 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect -8726 356294 592650 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 102986 356294
rect 103222 356058 103306 356294
rect 103542 356058 138986 356294
rect 139222 356058 139306 356294
rect 139542 356058 174986 356294
rect 175222 356058 175306 356294
rect 175542 356058 210986 356294
rect 211222 356058 211306 356294
rect 211542 356058 246986 356294
rect 247222 356058 247306 356294
rect 247542 356058 282986 356294
rect 283222 356058 283306 356294
rect 283542 356058 318986 356294
rect 319222 356058 319306 356294
rect 319542 356058 354986 356294
rect 355222 356058 355306 356294
rect 355542 356058 390986 356294
rect 391222 356058 391306 356294
rect 391542 356058 426986 356294
rect 427222 356058 427306 356294
rect 427542 356058 462986 356294
rect 463222 356058 463306 356294
rect 463542 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect -8726 356026 592650 356058
rect -6806 352894 590730 352926
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 63266 352894
rect 63502 352658 63586 352894
rect 63822 352658 99266 352894
rect 99502 352658 99586 352894
rect 99822 352658 135266 352894
rect 135502 352658 135586 352894
rect 135822 352658 171266 352894
rect 171502 352658 171586 352894
rect 171822 352658 207266 352894
rect 207502 352658 207586 352894
rect 207822 352658 243266 352894
rect 243502 352658 243586 352894
rect 243822 352658 279266 352894
rect 279502 352658 279586 352894
rect 279822 352658 315266 352894
rect 315502 352658 315586 352894
rect 315822 352658 351266 352894
rect 351502 352658 351586 352894
rect 351822 352658 387266 352894
rect 387502 352658 387586 352894
rect 387822 352658 423266 352894
rect 423502 352658 423586 352894
rect 423822 352658 459266 352894
rect 459502 352658 459586 352894
rect 459822 352658 495266 352894
rect 495502 352658 495586 352894
rect 495822 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect -6806 352574 590730 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 63266 352574
rect 63502 352338 63586 352574
rect 63822 352338 99266 352574
rect 99502 352338 99586 352574
rect 99822 352338 135266 352574
rect 135502 352338 135586 352574
rect 135822 352338 171266 352574
rect 171502 352338 171586 352574
rect 171822 352338 207266 352574
rect 207502 352338 207586 352574
rect 207822 352338 243266 352574
rect 243502 352338 243586 352574
rect 243822 352338 279266 352574
rect 279502 352338 279586 352574
rect 279822 352338 315266 352574
rect 315502 352338 315586 352574
rect 315822 352338 351266 352574
rect 351502 352338 351586 352574
rect 351822 352338 387266 352574
rect 387502 352338 387586 352574
rect 387822 352338 423266 352574
rect 423502 352338 423586 352574
rect 423822 352338 459266 352574
rect 459502 352338 459586 352574
rect 459822 352338 495266 352574
rect 495502 352338 495586 352574
rect 495822 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect -6806 352306 590730 352338
rect -4886 349174 588810 349206
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 59546 349174
rect 59782 348938 59866 349174
rect 60102 348938 95546 349174
rect 95782 348938 95866 349174
rect 96102 348938 131546 349174
rect 131782 348938 131866 349174
rect 132102 348938 167546 349174
rect 167782 348938 167866 349174
rect 168102 348938 203546 349174
rect 203782 348938 203866 349174
rect 204102 348938 239546 349174
rect 239782 348938 239866 349174
rect 240102 348938 275546 349174
rect 275782 348938 275866 349174
rect 276102 348938 311546 349174
rect 311782 348938 311866 349174
rect 312102 348938 347546 349174
rect 347782 348938 347866 349174
rect 348102 348938 383546 349174
rect 383782 348938 383866 349174
rect 384102 348938 419546 349174
rect 419782 348938 419866 349174
rect 420102 348938 455546 349174
rect 455782 348938 455866 349174
rect 456102 348938 491546 349174
rect 491782 348938 491866 349174
rect 492102 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect -4886 348854 588810 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 59546 348854
rect 59782 348618 59866 348854
rect 60102 348618 95546 348854
rect 95782 348618 95866 348854
rect 96102 348618 131546 348854
rect 131782 348618 131866 348854
rect 132102 348618 167546 348854
rect 167782 348618 167866 348854
rect 168102 348618 203546 348854
rect 203782 348618 203866 348854
rect 204102 348618 239546 348854
rect 239782 348618 239866 348854
rect 240102 348618 275546 348854
rect 275782 348618 275866 348854
rect 276102 348618 311546 348854
rect 311782 348618 311866 348854
rect 312102 348618 347546 348854
rect 347782 348618 347866 348854
rect 348102 348618 383546 348854
rect 383782 348618 383866 348854
rect 384102 348618 419546 348854
rect 419782 348618 419866 348854
rect 420102 348618 455546 348854
rect 455782 348618 455866 348854
rect 456102 348618 491546 348854
rect 491782 348618 491866 348854
rect 492102 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect -4886 348586 588810 348618
rect -2966 345454 586890 345486
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect -2966 345134 586890 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect -2966 344866 586890 344898
rect -8726 338614 592650 338646
rect -8726 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 84986 338614
rect 85222 338378 85306 338614
rect 85542 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 192986 338614
rect 193222 338378 193306 338614
rect 193542 338378 228986 338614
rect 229222 338378 229306 338614
rect 229542 338378 264986 338614
rect 265222 338378 265306 338614
rect 265542 338378 300986 338614
rect 301222 338378 301306 338614
rect 301542 338378 336986 338614
rect 337222 338378 337306 338614
rect 337542 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 84986 338294
rect 85222 338058 85306 338294
rect 85542 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 192986 338294
rect 193222 338058 193306 338294
rect 193542 338058 228986 338294
rect 229222 338058 229306 338294
rect 229542 338058 264986 338294
rect 265222 338058 265306 338294
rect 265542 338058 300986 338294
rect 301222 338058 301306 338294
rect 301542 338058 336986 338294
rect 337222 338058 337306 338294
rect 337542 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 592650 338294
rect -8726 338026 592650 338058
rect -6806 334894 590730 334926
rect -6806 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 189266 334894
rect 189502 334658 189586 334894
rect 189822 334658 225266 334894
rect 225502 334658 225586 334894
rect 225822 334658 261266 334894
rect 261502 334658 261586 334894
rect 261822 334658 297266 334894
rect 297502 334658 297586 334894
rect 297822 334658 333266 334894
rect 333502 334658 333586 334894
rect 333822 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 590730 334894
rect -6806 334574 590730 334658
rect -6806 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 189266 334574
rect 189502 334338 189586 334574
rect 189822 334338 225266 334574
rect 225502 334338 225586 334574
rect 225822 334338 261266 334574
rect 261502 334338 261586 334574
rect 261822 334338 297266 334574
rect 297502 334338 297586 334574
rect 297822 334338 333266 334574
rect 333502 334338 333586 334574
rect 333822 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 590730 334574
rect -6806 334306 590730 334338
rect -4886 331174 588810 331206
rect -4886 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 113546 331174
rect 113782 330938 113866 331174
rect 114102 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 221546 331174
rect 221782 330938 221866 331174
rect 222102 330938 257546 331174
rect 257782 330938 257866 331174
rect 258102 330938 293546 331174
rect 293782 330938 293866 331174
rect 294102 330938 329546 331174
rect 329782 330938 329866 331174
rect 330102 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 588810 331174
rect -4886 330854 588810 330938
rect -4886 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 113546 330854
rect 113782 330618 113866 330854
rect 114102 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 221546 330854
rect 221782 330618 221866 330854
rect 222102 330618 257546 330854
rect 257782 330618 257866 330854
rect 258102 330618 293546 330854
rect 293782 330618 293866 330854
rect 294102 330618 329546 330854
rect 329782 330618 329866 330854
rect 330102 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 588810 330854
rect -4886 330586 588810 330618
rect -2966 327454 586890 327486
rect -2966 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 586890 327454
rect -2966 327134 586890 327218
rect -2966 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 586890 327134
rect -2966 326866 586890 326898
rect -8726 320614 592650 320646
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 66986 320614
rect 67222 320378 67306 320614
rect 67542 320378 102986 320614
rect 103222 320378 103306 320614
rect 103542 320378 138986 320614
rect 139222 320378 139306 320614
rect 139542 320378 174986 320614
rect 175222 320378 175306 320614
rect 175542 320378 210986 320614
rect 211222 320378 211306 320614
rect 211542 320378 246986 320614
rect 247222 320378 247306 320614
rect 247542 320378 282986 320614
rect 283222 320378 283306 320614
rect 283542 320378 318986 320614
rect 319222 320378 319306 320614
rect 319542 320378 354986 320614
rect 355222 320378 355306 320614
rect 355542 320378 390986 320614
rect 391222 320378 391306 320614
rect 391542 320378 426986 320614
rect 427222 320378 427306 320614
rect 427542 320378 462986 320614
rect 463222 320378 463306 320614
rect 463542 320378 498986 320614
rect 499222 320378 499306 320614
rect 499542 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect -8726 320294 592650 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 66986 320294
rect 67222 320058 67306 320294
rect 67542 320058 102986 320294
rect 103222 320058 103306 320294
rect 103542 320058 138986 320294
rect 139222 320058 139306 320294
rect 139542 320058 174986 320294
rect 175222 320058 175306 320294
rect 175542 320058 210986 320294
rect 211222 320058 211306 320294
rect 211542 320058 246986 320294
rect 247222 320058 247306 320294
rect 247542 320058 282986 320294
rect 283222 320058 283306 320294
rect 283542 320058 318986 320294
rect 319222 320058 319306 320294
rect 319542 320058 354986 320294
rect 355222 320058 355306 320294
rect 355542 320058 390986 320294
rect 391222 320058 391306 320294
rect 391542 320058 426986 320294
rect 427222 320058 427306 320294
rect 427542 320058 462986 320294
rect 463222 320058 463306 320294
rect 463542 320058 498986 320294
rect 499222 320058 499306 320294
rect 499542 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect -8726 320026 592650 320058
rect -6806 316894 590730 316926
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 63266 316894
rect 63502 316658 63586 316894
rect 63822 316658 99266 316894
rect 99502 316658 99586 316894
rect 99822 316658 135266 316894
rect 135502 316658 135586 316894
rect 135822 316658 171266 316894
rect 171502 316658 171586 316894
rect 171822 316658 207266 316894
rect 207502 316658 207586 316894
rect 207822 316658 243266 316894
rect 243502 316658 243586 316894
rect 243822 316658 279266 316894
rect 279502 316658 279586 316894
rect 279822 316658 315266 316894
rect 315502 316658 315586 316894
rect 315822 316658 351266 316894
rect 351502 316658 351586 316894
rect 351822 316658 387266 316894
rect 387502 316658 387586 316894
rect 387822 316658 423266 316894
rect 423502 316658 423586 316894
rect 423822 316658 459266 316894
rect 459502 316658 459586 316894
rect 459822 316658 495266 316894
rect 495502 316658 495586 316894
rect 495822 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect -6806 316574 590730 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 63266 316574
rect 63502 316338 63586 316574
rect 63822 316338 99266 316574
rect 99502 316338 99586 316574
rect 99822 316338 135266 316574
rect 135502 316338 135586 316574
rect 135822 316338 171266 316574
rect 171502 316338 171586 316574
rect 171822 316338 207266 316574
rect 207502 316338 207586 316574
rect 207822 316338 243266 316574
rect 243502 316338 243586 316574
rect 243822 316338 279266 316574
rect 279502 316338 279586 316574
rect 279822 316338 315266 316574
rect 315502 316338 315586 316574
rect 315822 316338 351266 316574
rect 351502 316338 351586 316574
rect 351822 316338 387266 316574
rect 387502 316338 387586 316574
rect 387822 316338 423266 316574
rect 423502 316338 423586 316574
rect 423822 316338 459266 316574
rect 459502 316338 459586 316574
rect 459822 316338 495266 316574
rect 495502 316338 495586 316574
rect 495822 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect -6806 316306 590730 316338
rect -4886 313174 588810 313206
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 59546 313174
rect 59782 312938 59866 313174
rect 60102 312938 95546 313174
rect 95782 312938 95866 313174
rect 96102 312938 131546 313174
rect 131782 312938 131866 313174
rect 132102 312938 167546 313174
rect 167782 312938 167866 313174
rect 168102 312938 203546 313174
rect 203782 312938 203866 313174
rect 204102 312938 239546 313174
rect 239782 312938 239866 313174
rect 240102 312938 275546 313174
rect 275782 312938 275866 313174
rect 276102 312938 311546 313174
rect 311782 312938 311866 313174
rect 312102 312938 347546 313174
rect 347782 312938 347866 313174
rect 348102 312938 383546 313174
rect 383782 312938 383866 313174
rect 384102 312938 419546 313174
rect 419782 312938 419866 313174
rect 420102 312938 455546 313174
rect 455782 312938 455866 313174
rect 456102 312938 491546 313174
rect 491782 312938 491866 313174
rect 492102 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect -4886 312854 588810 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 59546 312854
rect 59782 312618 59866 312854
rect 60102 312618 95546 312854
rect 95782 312618 95866 312854
rect 96102 312618 131546 312854
rect 131782 312618 131866 312854
rect 132102 312618 167546 312854
rect 167782 312618 167866 312854
rect 168102 312618 203546 312854
rect 203782 312618 203866 312854
rect 204102 312618 239546 312854
rect 239782 312618 239866 312854
rect 240102 312618 275546 312854
rect 275782 312618 275866 312854
rect 276102 312618 311546 312854
rect 311782 312618 311866 312854
rect 312102 312618 347546 312854
rect 347782 312618 347866 312854
rect 348102 312618 383546 312854
rect 383782 312618 383866 312854
rect 384102 312618 419546 312854
rect 419782 312618 419866 312854
rect 420102 312618 455546 312854
rect 455782 312618 455866 312854
rect 456102 312618 491546 312854
rect 491782 312618 491866 312854
rect 492102 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect -4886 312586 588810 312618
rect -2966 309454 586890 309486
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect -2966 309134 586890 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect -2966 308866 586890 308898
rect -8726 302614 592650 302646
rect -8726 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 84986 302614
rect 85222 302378 85306 302614
rect 85542 302378 120986 302614
rect 121222 302378 121306 302614
rect 121542 302378 156986 302614
rect 157222 302378 157306 302614
rect 157542 302378 192986 302614
rect 193222 302378 193306 302614
rect 193542 302378 228986 302614
rect 229222 302378 229306 302614
rect 229542 302378 264986 302614
rect 265222 302378 265306 302614
rect 265542 302378 300986 302614
rect 301222 302378 301306 302614
rect 301542 302378 336986 302614
rect 337222 302378 337306 302614
rect 337542 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 84986 302294
rect 85222 302058 85306 302294
rect 85542 302058 120986 302294
rect 121222 302058 121306 302294
rect 121542 302058 156986 302294
rect 157222 302058 157306 302294
rect 157542 302058 192986 302294
rect 193222 302058 193306 302294
rect 193542 302058 228986 302294
rect 229222 302058 229306 302294
rect 229542 302058 264986 302294
rect 265222 302058 265306 302294
rect 265542 302058 300986 302294
rect 301222 302058 301306 302294
rect 301542 302058 336986 302294
rect 337222 302058 337306 302294
rect 337542 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 592650 302294
rect -8726 302026 592650 302058
rect -6806 298894 590730 298926
rect -6806 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 81266 298894
rect 81502 298658 81586 298894
rect 81822 298658 117266 298894
rect 117502 298658 117586 298894
rect 117822 298658 153266 298894
rect 153502 298658 153586 298894
rect 153822 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 225266 298894
rect 225502 298658 225586 298894
rect 225822 298658 261266 298894
rect 261502 298658 261586 298894
rect 261822 298658 297266 298894
rect 297502 298658 297586 298894
rect 297822 298658 333266 298894
rect 333502 298658 333586 298894
rect 333822 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 590730 298894
rect -6806 298574 590730 298658
rect -6806 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 81266 298574
rect 81502 298338 81586 298574
rect 81822 298338 117266 298574
rect 117502 298338 117586 298574
rect 117822 298338 153266 298574
rect 153502 298338 153586 298574
rect 153822 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 225266 298574
rect 225502 298338 225586 298574
rect 225822 298338 261266 298574
rect 261502 298338 261586 298574
rect 261822 298338 297266 298574
rect 297502 298338 297586 298574
rect 297822 298338 333266 298574
rect 333502 298338 333586 298574
rect 333822 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 590730 298574
rect -6806 298306 590730 298338
rect -4886 295174 588810 295206
rect -4886 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 77546 295174
rect 77782 294938 77866 295174
rect 78102 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 149546 295174
rect 149782 294938 149866 295174
rect 150102 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 221546 295174
rect 221782 294938 221866 295174
rect 222102 294938 257546 295174
rect 257782 294938 257866 295174
rect 258102 294938 293546 295174
rect 293782 294938 293866 295174
rect 294102 294938 329546 295174
rect 329782 294938 329866 295174
rect 330102 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 588810 295174
rect -4886 294854 588810 294938
rect -4886 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 77546 294854
rect 77782 294618 77866 294854
rect 78102 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 149546 294854
rect 149782 294618 149866 294854
rect 150102 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 221546 294854
rect 221782 294618 221866 294854
rect 222102 294618 257546 294854
rect 257782 294618 257866 294854
rect 258102 294618 293546 294854
rect 293782 294618 293866 294854
rect 294102 294618 329546 294854
rect 329782 294618 329866 294854
rect 330102 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 588810 294854
rect -4886 294586 588810 294618
rect -2966 291454 586890 291486
rect -2966 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 586890 291454
rect -2966 291134 586890 291218
rect -2966 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 586890 291134
rect -2966 290866 586890 290898
rect -8726 284614 592650 284646
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 66986 284614
rect 67222 284378 67306 284614
rect 67542 284378 102986 284614
rect 103222 284378 103306 284614
rect 103542 284378 138986 284614
rect 139222 284378 139306 284614
rect 139542 284378 174986 284614
rect 175222 284378 175306 284614
rect 175542 284378 210986 284614
rect 211222 284378 211306 284614
rect 211542 284378 246986 284614
rect 247222 284378 247306 284614
rect 247542 284378 282986 284614
rect 283222 284378 283306 284614
rect 283542 284378 318986 284614
rect 319222 284378 319306 284614
rect 319542 284378 354986 284614
rect 355222 284378 355306 284614
rect 355542 284378 390986 284614
rect 391222 284378 391306 284614
rect 391542 284378 426986 284614
rect 427222 284378 427306 284614
rect 427542 284378 462986 284614
rect 463222 284378 463306 284614
rect 463542 284378 498986 284614
rect 499222 284378 499306 284614
rect 499542 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect -8726 284294 592650 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 66986 284294
rect 67222 284058 67306 284294
rect 67542 284058 102986 284294
rect 103222 284058 103306 284294
rect 103542 284058 138986 284294
rect 139222 284058 139306 284294
rect 139542 284058 174986 284294
rect 175222 284058 175306 284294
rect 175542 284058 210986 284294
rect 211222 284058 211306 284294
rect 211542 284058 246986 284294
rect 247222 284058 247306 284294
rect 247542 284058 282986 284294
rect 283222 284058 283306 284294
rect 283542 284058 318986 284294
rect 319222 284058 319306 284294
rect 319542 284058 354986 284294
rect 355222 284058 355306 284294
rect 355542 284058 390986 284294
rect 391222 284058 391306 284294
rect 391542 284058 426986 284294
rect 427222 284058 427306 284294
rect 427542 284058 462986 284294
rect 463222 284058 463306 284294
rect 463542 284058 498986 284294
rect 499222 284058 499306 284294
rect 499542 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect -8726 284026 592650 284058
rect -6806 280894 590730 280926
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 63266 280894
rect 63502 280658 63586 280894
rect 63822 280658 99266 280894
rect 99502 280658 99586 280894
rect 99822 280658 135266 280894
rect 135502 280658 135586 280894
rect 135822 280658 171266 280894
rect 171502 280658 171586 280894
rect 171822 280658 207266 280894
rect 207502 280658 207586 280894
rect 207822 280658 243266 280894
rect 243502 280658 243586 280894
rect 243822 280658 279266 280894
rect 279502 280658 279586 280894
rect 279822 280658 315266 280894
rect 315502 280658 315586 280894
rect 315822 280658 351266 280894
rect 351502 280658 351586 280894
rect 351822 280658 387266 280894
rect 387502 280658 387586 280894
rect 387822 280658 423266 280894
rect 423502 280658 423586 280894
rect 423822 280658 459266 280894
rect 459502 280658 459586 280894
rect 459822 280658 495266 280894
rect 495502 280658 495586 280894
rect 495822 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect -6806 280574 590730 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 63266 280574
rect 63502 280338 63586 280574
rect 63822 280338 99266 280574
rect 99502 280338 99586 280574
rect 99822 280338 135266 280574
rect 135502 280338 135586 280574
rect 135822 280338 171266 280574
rect 171502 280338 171586 280574
rect 171822 280338 207266 280574
rect 207502 280338 207586 280574
rect 207822 280338 243266 280574
rect 243502 280338 243586 280574
rect 243822 280338 279266 280574
rect 279502 280338 279586 280574
rect 279822 280338 315266 280574
rect 315502 280338 315586 280574
rect 315822 280338 351266 280574
rect 351502 280338 351586 280574
rect 351822 280338 387266 280574
rect 387502 280338 387586 280574
rect 387822 280338 423266 280574
rect 423502 280338 423586 280574
rect 423822 280338 459266 280574
rect 459502 280338 459586 280574
rect 459822 280338 495266 280574
rect 495502 280338 495586 280574
rect 495822 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect -6806 280306 590730 280338
rect -4886 277174 588810 277206
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 59546 277174
rect 59782 276938 59866 277174
rect 60102 276938 95546 277174
rect 95782 276938 95866 277174
rect 96102 276938 131546 277174
rect 131782 276938 131866 277174
rect 132102 276938 167546 277174
rect 167782 276938 167866 277174
rect 168102 276938 203546 277174
rect 203782 276938 203866 277174
rect 204102 276938 239546 277174
rect 239782 276938 239866 277174
rect 240102 276938 275546 277174
rect 275782 276938 275866 277174
rect 276102 276938 311546 277174
rect 311782 276938 311866 277174
rect 312102 276938 347546 277174
rect 347782 276938 347866 277174
rect 348102 276938 383546 277174
rect 383782 276938 383866 277174
rect 384102 276938 419546 277174
rect 419782 276938 419866 277174
rect 420102 276938 455546 277174
rect 455782 276938 455866 277174
rect 456102 276938 491546 277174
rect 491782 276938 491866 277174
rect 492102 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect -4886 276854 588810 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 59546 276854
rect 59782 276618 59866 276854
rect 60102 276618 95546 276854
rect 95782 276618 95866 276854
rect 96102 276618 131546 276854
rect 131782 276618 131866 276854
rect 132102 276618 167546 276854
rect 167782 276618 167866 276854
rect 168102 276618 203546 276854
rect 203782 276618 203866 276854
rect 204102 276618 239546 276854
rect 239782 276618 239866 276854
rect 240102 276618 275546 276854
rect 275782 276618 275866 276854
rect 276102 276618 311546 276854
rect 311782 276618 311866 276854
rect 312102 276618 347546 276854
rect 347782 276618 347866 276854
rect 348102 276618 383546 276854
rect 383782 276618 383866 276854
rect 384102 276618 419546 276854
rect 419782 276618 419866 276854
rect 420102 276618 455546 276854
rect 455782 276618 455866 276854
rect 456102 276618 491546 276854
rect 491782 276618 491866 276854
rect 492102 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect -4886 276586 588810 276618
rect -2966 273454 586890 273486
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect -2966 273134 586890 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect -2966 272866 586890 272898
rect -8726 266614 592650 266646
rect -8726 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 84986 266614
rect 85222 266378 85306 266614
rect 85542 266378 120986 266614
rect 121222 266378 121306 266614
rect 121542 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 192986 266614
rect 193222 266378 193306 266614
rect 193542 266378 228986 266614
rect 229222 266378 229306 266614
rect 229542 266378 264986 266614
rect 265222 266378 265306 266614
rect 265542 266378 300986 266614
rect 301222 266378 301306 266614
rect 301542 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 84986 266294
rect 85222 266058 85306 266294
rect 85542 266058 120986 266294
rect 121222 266058 121306 266294
rect 121542 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 192986 266294
rect 193222 266058 193306 266294
rect 193542 266058 228986 266294
rect 229222 266058 229306 266294
rect 229542 266058 264986 266294
rect 265222 266058 265306 266294
rect 265542 266058 300986 266294
rect 301222 266058 301306 266294
rect 301542 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 592650 266294
rect -8726 266026 592650 266058
rect -6806 262894 590730 262926
rect -6806 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 81266 262894
rect 81502 262658 81586 262894
rect 81822 262658 117266 262894
rect 117502 262658 117586 262894
rect 117822 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 225266 262894
rect 225502 262658 225586 262894
rect 225822 262658 261266 262894
rect 261502 262658 261586 262894
rect 261822 262658 297266 262894
rect 297502 262658 297586 262894
rect 297822 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 590730 262894
rect -6806 262574 590730 262658
rect -6806 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 81266 262574
rect 81502 262338 81586 262574
rect 81822 262338 117266 262574
rect 117502 262338 117586 262574
rect 117822 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 225266 262574
rect 225502 262338 225586 262574
rect 225822 262338 261266 262574
rect 261502 262338 261586 262574
rect 261822 262338 297266 262574
rect 297502 262338 297586 262574
rect 297822 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 590730 262574
rect -6806 262306 590730 262338
rect -4886 259174 588810 259206
rect -4886 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 77546 259174
rect 77782 258938 77866 259174
rect 78102 258938 113546 259174
rect 113782 258938 113866 259174
rect 114102 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 221546 259174
rect 221782 258938 221866 259174
rect 222102 258938 257546 259174
rect 257782 258938 257866 259174
rect 258102 258938 293546 259174
rect 293782 258938 293866 259174
rect 294102 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 588810 259174
rect -4886 258854 588810 258938
rect -4886 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 77546 258854
rect 77782 258618 77866 258854
rect 78102 258618 113546 258854
rect 113782 258618 113866 258854
rect 114102 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 221546 258854
rect 221782 258618 221866 258854
rect 222102 258618 257546 258854
rect 257782 258618 257866 258854
rect 258102 258618 293546 258854
rect 293782 258618 293866 258854
rect 294102 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 588810 258854
rect -4886 258586 588810 258618
rect -2966 255454 586890 255486
rect -2966 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 586890 255454
rect -2966 255134 586890 255218
rect -2966 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 586890 255134
rect -2966 254866 586890 254898
rect -8726 248614 592650 248646
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 66986 248614
rect 67222 248378 67306 248614
rect 67542 248378 102986 248614
rect 103222 248378 103306 248614
rect 103542 248378 138986 248614
rect 139222 248378 139306 248614
rect 139542 248378 174986 248614
rect 175222 248378 175306 248614
rect 175542 248378 210986 248614
rect 211222 248378 211306 248614
rect 211542 248378 246986 248614
rect 247222 248378 247306 248614
rect 247542 248378 282986 248614
rect 283222 248378 283306 248614
rect 283542 248378 318986 248614
rect 319222 248378 319306 248614
rect 319542 248378 354986 248614
rect 355222 248378 355306 248614
rect 355542 248378 390986 248614
rect 391222 248378 391306 248614
rect 391542 248378 426986 248614
rect 427222 248378 427306 248614
rect 427542 248378 462986 248614
rect 463222 248378 463306 248614
rect 463542 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect -8726 248294 592650 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 66986 248294
rect 67222 248058 67306 248294
rect 67542 248058 102986 248294
rect 103222 248058 103306 248294
rect 103542 248058 138986 248294
rect 139222 248058 139306 248294
rect 139542 248058 174986 248294
rect 175222 248058 175306 248294
rect 175542 248058 210986 248294
rect 211222 248058 211306 248294
rect 211542 248058 246986 248294
rect 247222 248058 247306 248294
rect 247542 248058 282986 248294
rect 283222 248058 283306 248294
rect 283542 248058 318986 248294
rect 319222 248058 319306 248294
rect 319542 248058 354986 248294
rect 355222 248058 355306 248294
rect 355542 248058 390986 248294
rect 391222 248058 391306 248294
rect 391542 248058 426986 248294
rect 427222 248058 427306 248294
rect 427542 248058 462986 248294
rect 463222 248058 463306 248294
rect 463542 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect -8726 248026 592650 248058
rect -6806 244894 590730 244926
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 99266 244894
rect 99502 244658 99586 244894
rect 99822 244658 135266 244894
rect 135502 244658 135586 244894
rect 135822 244658 171266 244894
rect 171502 244658 171586 244894
rect 171822 244658 207266 244894
rect 207502 244658 207586 244894
rect 207822 244658 243266 244894
rect 243502 244658 243586 244894
rect 243822 244658 279266 244894
rect 279502 244658 279586 244894
rect 279822 244658 315266 244894
rect 315502 244658 315586 244894
rect 315822 244658 351266 244894
rect 351502 244658 351586 244894
rect 351822 244658 387266 244894
rect 387502 244658 387586 244894
rect 387822 244658 423266 244894
rect 423502 244658 423586 244894
rect 423822 244658 459266 244894
rect 459502 244658 459586 244894
rect 459822 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect -6806 244574 590730 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 99266 244574
rect 99502 244338 99586 244574
rect 99822 244338 135266 244574
rect 135502 244338 135586 244574
rect 135822 244338 171266 244574
rect 171502 244338 171586 244574
rect 171822 244338 207266 244574
rect 207502 244338 207586 244574
rect 207822 244338 243266 244574
rect 243502 244338 243586 244574
rect 243822 244338 279266 244574
rect 279502 244338 279586 244574
rect 279822 244338 315266 244574
rect 315502 244338 315586 244574
rect 315822 244338 351266 244574
rect 351502 244338 351586 244574
rect 351822 244338 387266 244574
rect 387502 244338 387586 244574
rect 387822 244338 423266 244574
rect 423502 244338 423586 244574
rect 423822 244338 459266 244574
rect 459502 244338 459586 244574
rect 459822 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect -6806 244306 590730 244338
rect -4886 241174 588810 241206
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 95546 241174
rect 95782 240938 95866 241174
rect 96102 240938 131546 241174
rect 131782 240938 131866 241174
rect 132102 240938 167546 241174
rect 167782 240938 167866 241174
rect 168102 240938 203546 241174
rect 203782 240938 203866 241174
rect 204102 240938 239546 241174
rect 239782 240938 239866 241174
rect 240102 240938 275546 241174
rect 275782 240938 275866 241174
rect 276102 240938 311546 241174
rect 311782 240938 311866 241174
rect 312102 240938 347546 241174
rect 347782 240938 347866 241174
rect 348102 240938 383546 241174
rect 383782 240938 383866 241174
rect 384102 240938 419546 241174
rect 419782 240938 419866 241174
rect 420102 240938 455546 241174
rect 455782 240938 455866 241174
rect 456102 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect -4886 240854 588810 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 95546 240854
rect 95782 240618 95866 240854
rect 96102 240618 131546 240854
rect 131782 240618 131866 240854
rect 132102 240618 167546 240854
rect 167782 240618 167866 240854
rect 168102 240618 203546 240854
rect 203782 240618 203866 240854
rect 204102 240618 239546 240854
rect 239782 240618 239866 240854
rect 240102 240618 275546 240854
rect 275782 240618 275866 240854
rect 276102 240618 311546 240854
rect 311782 240618 311866 240854
rect 312102 240618 347546 240854
rect 347782 240618 347866 240854
rect 348102 240618 383546 240854
rect 383782 240618 383866 240854
rect 384102 240618 419546 240854
rect 419782 240618 419866 240854
rect 420102 240618 455546 240854
rect 455782 240618 455866 240854
rect 456102 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect -4886 240586 588810 240618
rect -2966 237454 586890 237486
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect -2966 237134 586890 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect -2966 236866 586890 236898
rect -8726 230614 592650 230646
rect -8726 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 156986 230614
rect 157222 230378 157306 230614
rect 157542 230378 192986 230614
rect 193222 230378 193306 230614
rect 193542 230378 228986 230614
rect 229222 230378 229306 230614
rect 229542 230378 264986 230614
rect 265222 230378 265306 230614
rect 265542 230378 300986 230614
rect 301222 230378 301306 230614
rect 301542 230378 336986 230614
rect 337222 230378 337306 230614
rect 337542 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 156986 230294
rect 157222 230058 157306 230294
rect 157542 230058 192986 230294
rect 193222 230058 193306 230294
rect 193542 230058 228986 230294
rect 229222 230058 229306 230294
rect 229542 230058 264986 230294
rect 265222 230058 265306 230294
rect 265542 230058 300986 230294
rect 301222 230058 301306 230294
rect 301542 230058 336986 230294
rect 337222 230058 337306 230294
rect 337542 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 592650 230294
rect -8726 230026 592650 230058
rect -6806 226894 590730 226926
rect -6806 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 81266 226894
rect 81502 226658 81586 226894
rect 81822 226658 117266 226894
rect 117502 226658 117586 226894
rect 117822 226658 153266 226894
rect 153502 226658 153586 226894
rect 153822 226658 189266 226894
rect 189502 226658 189586 226894
rect 189822 226658 225266 226894
rect 225502 226658 225586 226894
rect 225822 226658 261266 226894
rect 261502 226658 261586 226894
rect 261822 226658 297266 226894
rect 297502 226658 297586 226894
rect 297822 226658 333266 226894
rect 333502 226658 333586 226894
rect 333822 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 590730 226894
rect -6806 226574 590730 226658
rect -6806 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 81266 226574
rect 81502 226338 81586 226574
rect 81822 226338 117266 226574
rect 117502 226338 117586 226574
rect 117822 226338 153266 226574
rect 153502 226338 153586 226574
rect 153822 226338 189266 226574
rect 189502 226338 189586 226574
rect 189822 226338 225266 226574
rect 225502 226338 225586 226574
rect 225822 226338 261266 226574
rect 261502 226338 261586 226574
rect 261822 226338 297266 226574
rect 297502 226338 297586 226574
rect 297822 226338 333266 226574
rect 333502 226338 333586 226574
rect 333822 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 590730 226574
rect -6806 226306 590730 226338
rect -4886 223174 588810 223206
rect -4886 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 113546 223174
rect 113782 222938 113866 223174
rect 114102 222938 149546 223174
rect 149782 222938 149866 223174
rect 150102 222938 185546 223174
rect 185782 222938 185866 223174
rect 186102 222938 221546 223174
rect 221782 222938 221866 223174
rect 222102 222938 257546 223174
rect 257782 222938 257866 223174
rect 258102 222938 293546 223174
rect 293782 222938 293866 223174
rect 294102 222938 329546 223174
rect 329782 222938 329866 223174
rect 330102 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 588810 223174
rect -4886 222854 588810 222938
rect -4886 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 113546 222854
rect 113782 222618 113866 222854
rect 114102 222618 149546 222854
rect 149782 222618 149866 222854
rect 150102 222618 185546 222854
rect 185782 222618 185866 222854
rect 186102 222618 221546 222854
rect 221782 222618 221866 222854
rect 222102 222618 257546 222854
rect 257782 222618 257866 222854
rect 258102 222618 293546 222854
rect 293782 222618 293866 222854
rect 294102 222618 329546 222854
rect 329782 222618 329866 222854
rect 330102 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 588810 222854
rect -4886 222586 588810 222618
rect -2966 219454 586890 219486
rect -2966 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 586890 219454
rect -2966 219134 586890 219218
rect -2966 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 586890 219134
rect -2966 218866 586890 218898
rect -8726 212614 592650 212646
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 66986 212614
rect 67222 212378 67306 212614
rect 67542 212378 102986 212614
rect 103222 212378 103306 212614
rect 103542 212378 138986 212614
rect 139222 212378 139306 212614
rect 139542 212378 174986 212614
rect 175222 212378 175306 212614
rect 175542 212378 210986 212614
rect 211222 212378 211306 212614
rect 211542 212378 246986 212614
rect 247222 212378 247306 212614
rect 247542 212378 282986 212614
rect 283222 212378 283306 212614
rect 283542 212378 318986 212614
rect 319222 212378 319306 212614
rect 319542 212378 354986 212614
rect 355222 212378 355306 212614
rect 355542 212378 390986 212614
rect 391222 212378 391306 212614
rect 391542 212378 426986 212614
rect 427222 212378 427306 212614
rect 427542 212378 462986 212614
rect 463222 212378 463306 212614
rect 463542 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect -8726 212294 592650 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 66986 212294
rect 67222 212058 67306 212294
rect 67542 212058 102986 212294
rect 103222 212058 103306 212294
rect 103542 212058 138986 212294
rect 139222 212058 139306 212294
rect 139542 212058 174986 212294
rect 175222 212058 175306 212294
rect 175542 212058 210986 212294
rect 211222 212058 211306 212294
rect 211542 212058 246986 212294
rect 247222 212058 247306 212294
rect 247542 212058 282986 212294
rect 283222 212058 283306 212294
rect 283542 212058 318986 212294
rect 319222 212058 319306 212294
rect 319542 212058 354986 212294
rect 355222 212058 355306 212294
rect 355542 212058 390986 212294
rect 391222 212058 391306 212294
rect 391542 212058 426986 212294
rect 427222 212058 427306 212294
rect 427542 212058 462986 212294
rect 463222 212058 463306 212294
rect 463542 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect -8726 212026 592650 212058
rect -6806 208894 590730 208926
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 63266 208894
rect 63502 208658 63586 208894
rect 63822 208658 99266 208894
rect 99502 208658 99586 208894
rect 99822 208658 135266 208894
rect 135502 208658 135586 208894
rect 135822 208658 171266 208894
rect 171502 208658 171586 208894
rect 171822 208658 207266 208894
rect 207502 208658 207586 208894
rect 207822 208658 243266 208894
rect 243502 208658 243586 208894
rect 243822 208658 279266 208894
rect 279502 208658 279586 208894
rect 279822 208658 315266 208894
rect 315502 208658 315586 208894
rect 315822 208658 351266 208894
rect 351502 208658 351586 208894
rect 351822 208658 387266 208894
rect 387502 208658 387586 208894
rect 387822 208658 423266 208894
rect 423502 208658 423586 208894
rect 423822 208658 459266 208894
rect 459502 208658 459586 208894
rect 459822 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect -6806 208574 590730 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 63266 208574
rect 63502 208338 63586 208574
rect 63822 208338 99266 208574
rect 99502 208338 99586 208574
rect 99822 208338 135266 208574
rect 135502 208338 135586 208574
rect 135822 208338 171266 208574
rect 171502 208338 171586 208574
rect 171822 208338 207266 208574
rect 207502 208338 207586 208574
rect 207822 208338 243266 208574
rect 243502 208338 243586 208574
rect 243822 208338 279266 208574
rect 279502 208338 279586 208574
rect 279822 208338 315266 208574
rect 315502 208338 315586 208574
rect 315822 208338 351266 208574
rect 351502 208338 351586 208574
rect 351822 208338 387266 208574
rect 387502 208338 387586 208574
rect 387822 208338 423266 208574
rect 423502 208338 423586 208574
rect 423822 208338 459266 208574
rect 459502 208338 459586 208574
rect 459822 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect -6806 208306 590730 208338
rect -4886 205174 588810 205206
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 59546 205174
rect 59782 204938 59866 205174
rect 60102 204938 95546 205174
rect 95782 204938 95866 205174
rect 96102 204938 131546 205174
rect 131782 204938 131866 205174
rect 132102 204938 167546 205174
rect 167782 204938 167866 205174
rect 168102 204938 203546 205174
rect 203782 204938 203866 205174
rect 204102 204938 239546 205174
rect 239782 204938 239866 205174
rect 240102 204938 275546 205174
rect 275782 204938 275866 205174
rect 276102 204938 311546 205174
rect 311782 204938 311866 205174
rect 312102 204938 347546 205174
rect 347782 204938 347866 205174
rect 348102 204938 383546 205174
rect 383782 204938 383866 205174
rect 384102 204938 419546 205174
rect 419782 204938 419866 205174
rect 420102 204938 455546 205174
rect 455782 204938 455866 205174
rect 456102 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect -4886 204854 588810 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 59546 204854
rect 59782 204618 59866 204854
rect 60102 204618 95546 204854
rect 95782 204618 95866 204854
rect 96102 204618 131546 204854
rect 131782 204618 131866 204854
rect 132102 204618 167546 204854
rect 167782 204618 167866 204854
rect 168102 204618 203546 204854
rect 203782 204618 203866 204854
rect 204102 204618 239546 204854
rect 239782 204618 239866 204854
rect 240102 204618 275546 204854
rect 275782 204618 275866 204854
rect 276102 204618 311546 204854
rect 311782 204618 311866 204854
rect 312102 204618 347546 204854
rect 347782 204618 347866 204854
rect 348102 204618 383546 204854
rect 383782 204618 383866 204854
rect 384102 204618 419546 204854
rect 419782 204618 419866 204854
rect 420102 204618 455546 204854
rect 455782 204618 455866 204854
rect 456102 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect -4886 204586 588810 204618
rect -2966 201454 586890 201486
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect -2966 201134 586890 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect -2966 200866 586890 200898
rect -8726 194614 592650 194646
rect -8726 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 120986 194614
rect 121222 194378 121306 194614
rect 121542 194378 156986 194614
rect 157222 194378 157306 194614
rect 157542 194378 192986 194614
rect 193222 194378 193306 194614
rect 193542 194378 336986 194614
rect 337222 194378 337306 194614
rect 337542 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 120986 194294
rect 121222 194058 121306 194294
rect 121542 194058 156986 194294
rect 157222 194058 157306 194294
rect 157542 194058 192986 194294
rect 193222 194058 193306 194294
rect 193542 194058 336986 194294
rect 337222 194058 337306 194294
rect 337542 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 592650 194294
rect -8726 194026 592650 194058
rect -6806 190894 590730 190926
rect -6806 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 117266 190894
rect 117502 190658 117586 190894
rect 117822 190658 153266 190894
rect 153502 190658 153586 190894
rect 153822 190658 189266 190894
rect 189502 190658 189586 190894
rect 189822 190658 333266 190894
rect 333502 190658 333586 190894
rect 333822 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 590730 190894
rect -6806 190574 590730 190658
rect -6806 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 117266 190574
rect 117502 190338 117586 190574
rect 117822 190338 153266 190574
rect 153502 190338 153586 190574
rect 153822 190338 189266 190574
rect 189502 190338 189586 190574
rect 189822 190338 333266 190574
rect 333502 190338 333586 190574
rect 333822 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 590730 190574
rect -6806 190306 590730 190338
rect -4886 187174 588810 187206
rect -4886 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 149546 187174
rect 149782 186938 149866 187174
rect 150102 186938 185546 187174
rect 185782 186938 185866 187174
rect 186102 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 588810 187174
rect -4886 186854 588810 186938
rect -4886 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 149546 186854
rect 149782 186618 149866 186854
rect 150102 186618 185546 186854
rect 185782 186618 185866 186854
rect 186102 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 588810 186854
rect -4886 186586 588810 186618
rect -2966 183454 586890 183486
rect -2966 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 162285 183454
rect 162521 183218 164882 183454
rect 165118 183218 167479 183454
rect 167715 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 204250 183454
rect 204486 183218 234970 183454
rect 235206 183218 265690 183454
rect 265926 183218 296410 183454
rect 296646 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 586890 183454
rect -2966 183134 586890 183218
rect -2966 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 162285 183134
rect 162521 182898 164882 183134
rect 165118 182898 167479 183134
rect 167715 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 204250 183134
rect 204486 182898 234970 183134
rect 235206 182898 265690 183134
rect 265926 182898 296410 183134
rect 296646 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 586890 183134
rect -2966 182866 586890 182898
rect -8726 176614 592650 176646
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 66986 176614
rect 67222 176378 67306 176614
rect 67542 176378 102986 176614
rect 103222 176378 103306 176614
rect 103542 176378 138986 176614
rect 139222 176378 139306 176614
rect 139542 176378 174986 176614
rect 175222 176378 175306 176614
rect 175542 176378 318986 176614
rect 319222 176378 319306 176614
rect 319542 176378 354986 176614
rect 355222 176378 355306 176614
rect 355542 176378 390986 176614
rect 391222 176378 391306 176614
rect 391542 176378 426986 176614
rect 427222 176378 427306 176614
rect 427542 176378 462986 176614
rect 463222 176378 463306 176614
rect 463542 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect -8726 176294 592650 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 66986 176294
rect 67222 176058 67306 176294
rect 67542 176058 102986 176294
rect 103222 176058 103306 176294
rect 103542 176058 138986 176294
rect 139222 176058 139306 176294
rect 139542 176058 174986 176294
rect 175222 176058 175306 176294
rect 175542 176058 318986 176294
rect 319222 176058 319306 176294
rect 319542 176058 354986 176294
rect 355222 176058 355306 176294
rect 355542 176058 390986 176294
rect 391222 176058 391306 176294
rect 391542 176058 426986 176294
rect 427222 176058 427306 176294
rect 427542 176058 462986 176294
rect 463222 176058 463306 176294
rect 463542 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect -8726 176026 592650 176058
rect -6806 172894 590730 172926
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 63266 172894
rect 63502 172658 63586 172894
rect 63822 172658 99266 172894
rect 99502 172658 99586 172894
rect 99822 172658 135266 172894
rect 135502 172658 135586 172894
rect 135822 172658 315266 172894
rect 315502 172658 315586 172894
rect 315822 172658 351266 172894
rect 351502 172658 351586 172894
rect 351822 172658 387266 172894
rect 387502 172658 387586 172894
rect 387822 172658 423266 172894
rect 423502 172658 423586 172894
rect 423822 172658 459266 172894
rect 459502 172658 459586 172894
rect 459822 172658 495266 172894
rect 495502 172658 495586 172894
rect 495822 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect -6806 172574 590730 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 63266 172574
rect 63502 172338 63586 172574
rect 63822 172338 99266 172574
rect 99502 172338 99586 172574
rect 99822 172338 135266 172574
rect 135502 172338 135586 172574
rect 135822 172338 315266 172574
rect 315502 172338 315586 172574
rect 315822 172338 351266 172574
rect 351502 172338 351586 172574
rect 351822 172338 387266 172574
rect 387502 172338 387586 172574
rect 387822 172338 423266 172574
rect 423502 172338 423586 172574
rect 423822 172338 459266 172574
rect 459502 172338 459586 172574
rect 459822 172338 495266 172574
rect 495502 172338 495586 172574
rect 495822 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect -6806 172306 590730 172338
rect -4886 169174 588810 169206
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 59546 169174
rect 59782 168938 59866 169174
rect 60102 168938 95546 169174
rect 95782 168938 95866 169174
rect 96102 168938 131546 169174
rect 131782 168938 131866 169174
rect 132102 168938 311546 169174
rect 311782 168938 311866 169174
rect 312102 168938 347546 169174
rect 347782 168938 347866 169174
rect 348102 168938 383546 169174
rect 383782 168938 383866 169174
rect 384102 168938 419546 169174
rect 419782 168938 419866 169174
rect 420102 168938 455546 169174
rect 455782 168938 455866 169174
rect 456102 168938 491546 169174
rect 491782 168938 491866 169174
rect 492102 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect -4886 168854 588810 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 59546 168854
rect 59782 168618 59866 168854
rect 60102 168618 95546 168854
rect 95782 168618 95866 168854
rect 96102 168618 131546 168854
rect 131782 168618 131866 168854
rect 132102 168618 311546 168854
rect 311782 168618 311866 168854
rect 312102 168618 347546 168854
rect 347782 168618 347866 168854
rect 348102 168618 383546 168854
rect 383782 168618 383866 168854
rect 384102 168618 419546 168854
rect 419782 168618 419866 168854
rect 420102 168618 455546 168854
rect 455782 168618 455866 168854
rect 456102 168618 491546 168854
rect 491782 168618 491866 168854
rect 492102 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect -4886 168586 588810 168618
rect -2966 165454 586890 165486
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 163583 165454
rect 163819 165218 166180 165454
rect 166416 165218 219610 165454
rect 219846 165218 250330 165454
rect 250566 165218 281050 165454
rect 281286 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect -2966 165134 586890 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 163583 165134
rect 163819 164898 166180 165134
rect 166416 164898 219610 165134
rect 219846 164898 250330 165134
rect 250566 164898 281050 165134
rect 281286 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect -2966 164866 586890 164898
rect -8726 158614 592650 158646
rect -8726 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 84986 158614
rect 85222 158378 85306 158614
rect 85542 158378 120986 158614
rect 121222 158378 121306 158614
rect 121542 158378 156986 158614
rect 157222 158378 157306 158614
rect 157542 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 84986 158294
rect 85222 158058 85306 158294
rect 85542 158058 120986 158294
rect 121222 158058 121306 158294
rect 121542 158058 156986 158294
rect 157222 158058 157306 158294
rect 157542 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 592650 158294
rect -8726 158026 592650 158058
rect -6806 154894 590730 154926
rect -6806 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 81266 154894
rect 81502 154658 81586 154894
rect 81822 154658 117266 154894
rect 117502 154658 117586 154894
rect 117822 154658 153266 154894
rect 153502 154658 153586 154894
rect 153822 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 590730 154894
rect -6806 154574 590730 154658
rect -6806 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 81266 154574
rect 81502 154338 81586 154574
rect 81822 154338 117266 154574
rect 117502 154338 117586 154574
rect 117822 154338 153266 154574
rect 153502 154338 153586 154574
rect 153822 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 590730 154574
rect -6806 154306 590730 154338
rect -4886 151174 588810 151206
rect -4886 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 77546 151174
rect 77782 150938 77866 151174
rect 78102 150938 113546 151174
rect 113782 150938 113866 151174
rect 114102 150938 149546 151174
rect 149782 150938 149866 151174
rect 150102 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 588810 151174
rect -4886 150854 588810 150938
rect -4886 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 77546 150854
rect 77782 150618 77866 150854
rect 78102 150618 113546 150854
rect 113782 150618 113866 150854
rect 114102 150618 149546 150854
rect 149782 150618 149866 150854
rect 150102 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 588810 150854
rect -4886 150586 588810 150618
rect -2966 147454 586890 147486
rect -2966 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 162285 147454
rect 162521 147218 164882 147454
rect 165118 147218 167479 147454
rect 167715 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 204250 147454
rect 204486 147218 234970 147454
rect 235206 147218 265690 147454
rect 265926 147218 296410 147454
rect 296646 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 586890 147454
rect -2966 147134 586890 147218
rect -2966 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 162285 147134
rect 162521 146898 164882 147134
rect 165118 146898 167479 147134
rect 167715 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 204250 147134
rect 204486 146898 234970 147134
rect 235206 146898 265690 147134
rect 265926 146898 296410 147134
rect 296646 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 586890 147134
rect -2966 146866 586890 146898
rect -8726 140614 592650 140646
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 66986 140614
rect 67222 140378 67306 140614
rect 67542 140378 102986 140614
rect 103222 140378 103306 140614
rect 103542 140378 138986 140614
rect 139222 140378 139306 140614
rect 139542 140378 174986 140614
rect 175222 140378 175306 140614
rect 175542 140378 318986 140614
rect 319222 140378 319306 140614
rect 319542 140378 354986 140614
rect 355222 140378 355306 140614
rect 355542 140378 390986 140614
rect 391222 140378 391306 140614
rect 391542 140378 426986 140614
rect 427222 140378 427306 140614
rect 427542 140378 462986 140614
rect 463222 140378 463306 140614
rect 463542 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect -8726 140294 592650 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 66986 140294
rect 67222 140058 67306 140294
rect 67542 140058 102986 140294
rect 103222 140058 103306 140294
rect 103542 140058 138986 140294
rect 139222 140058 139306 140294
rect 139542 140058 174986 140294
rect 175222 140058 175306 140294
rect 175542 140058 318986 140294
rect 319222 140058 319306 140294
rect 319542 140058 354986 140294
rect 355222 140058 355306 140294
rect 355542 140058 390986 140294
rect 391222 140058 391306 140294
rect 391542 140058 426986 140294
rect 427222 140058 427306 140294
rect 427542 140058 462986 140294
rect 463222 140058 463306 140294
rect 463542 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect -8726 140026 592650 140058
rect -6806 136894 590730 136926
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 63266 136894
rect 63502 136658 63586 136894
rect 63822 136658 99266 136894
rect 99502 136658 99586 136894
rect 99822 136658 135266 136894
rect 135502 136658 135586 136894
rect 135822 136658 315266 136894
rect 315502 136658 315586 136894
rect 315822 136658 351266 136894
rect 351502 136658 351586 136894
rect 351822 136658 387266 136894
rect 387502 136658 387586 136894
rect 387822 136658 423266 136894
rect 423502 136658 423586 136894
rect 423822 136658 459266 136894
rect 459502 136658 459586 136894
rect 459822 136658 495266 136894
rect 495502 136658 495586 136894
rect 495822 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect -6806 136574 590730 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 63266 136574
rect 63502 136338 63586 136574
rect 63822 136338 99266 136574
rect 99502 136338 99586 136574
rect 99822 136338 135266 136574
rect 135502 136338 135586 136574
rect 135822 136338 315266 136574
rect 315502 136338 315586 136574
rect 315822 136338 351266 136574
rect 351502 136338 351586 136574
rect 351822 136338 387266 136574
rect 387502 136338 387586 136574
rect 387822 136338 423266 136574
rect 423502 136338 423586 136574
rect 423822 136338 459266 136574
rect 459502 136338 459586 136574
rect 459822 136338 495266 136574
rect 495502 136338 495586 136574
rect 495822 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect -6806 136306 590730 136338
rect -4886 133174 588810 133206
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 59546 133174
rect 59782 132938 59866 133174
rect 60102 132938 95546 133174
rect 95782 132938 95866 133174
rect 96102 132938 131546 133174
rect 131782 132938 131866 133174
rect 132102 132938 311546 133174
rect 311782 132938 311866 133174
rect 312102 132938 347546 133174
rect 347782 132938 347866 133174
rect 348102 132938 383546 133174
rect 383782 132938 383866 133174
rect 384102 132938 419546 133174
rect 419782 132938 419866 133174
rect 420102 132938 455546 133174
rect 455782 132938 455866 133174
rect 456102 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect -4886 132854 588810 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 59546 132854
rect 59782 132618 59866 132854
rect 60102 132618 95546 132854
rect 95782 132618 95866 132854
rect 96102 132618 131546 132854
rect 131782 132618 131866 132854
rect 132102 132618 311546 132854
rect 311782 132618 311866 132854
rect 312102 132618 347546 132854
rect 347782 132618 347866 132854
rect 348102 132618 383546 132854
rect 383782 132618 383866 132854
rect 384102 132618 419546 132854
rect 419782 132618 419866 132854
rect 420102 132618 455546 132854
rect 455782 132618 455866 132854
rect 456102 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect -4886 132586 588810 132618
rect -2966 129454 586890 129486
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 127826 129454
rect 128062 129218 128146 129454
rect 128382 129218 163583 129454
rect 163819 129218 166180 129454
rect 166416 129218 219610 129454
rect 219846 129218 250330 129454
rect 250566 129218 281050 129454
rect 281286 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect -2966 129134 586890 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 127826 129134
rect 128062 128898 128146 129134
rect 128382 128898 163583 129134
rect 163819 128898 166180 129134
rect 166416 128898 219610 129134
rect 219846 128898 250330 129134
rect 250566 128898 281050 129134
rect 281286 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect -2966 128866 586890 128898
rect -8726 122614 592650 122646
rect -8726 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 84986 122614
rect 85222 122378 85306 122614
rect 85542 122378 120986 122614
rect 121222 122378 121306 122614
rect 121542 122378 156986 122614
rect 157222 122378 157306 122614
rect 157542 122378 192986 122614
rect 193222 122378 193306 122614
rect 193542 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 84986 122294
rect 85222 122058 85306 122294
rect 85542 122058 120986 122294
rect 121222 122058 121306 122294
rect 121542 122058 156986 122294
rect 157222 122058 157306 122294
rect 157542 122058 192986 122294
rect 193222 122058 193306 122294
rect 193542 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 592650 122294
rect -8726 122026 592650 122058
rect -6806 118894 590730 118926
rect -6806 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 81266 118894
rect 81502 118658 81586 118894
rect 81822 118658 117266 118894
rect 117502 118658 117586 118894
rect 117822 118658 153266 118894
rect 153502 118658 153586 118894
rect 153822 118658 189266 118894
rect 189502 118658 189586 118894
rect 189822 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 590730 118894
rect -6806 118574 590730 118658
rect -6806 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 81266 118574
rect 81502 118338 81586 118574
rect 81822 118338 117266 118574
rect 117502 118338 117586 118574
rect 117822 118338 153266 118574
rect 153502 118338 153586 118574
rect 153822 118338 189266 118574
rect 189502 118338 189586 118574
rect 189822 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 590730 118574
rect -6806 118306 590730 118338
rect -4886 115174 588810 115206
rect -4886 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 77546 115174
rect 77782 114938 77866 115174
rect 78102 114938 113546 115174
rect 113782 114938 113866 115174
rect 114102 114938 149546 115174
rect 149782 114938 149866 115174
rect 150102 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 588810 115174
rect -4886 114854 588810 114938
rect -4886 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 77546 114854
rect 77782 114618 77866 114854
rect 78102 114618 113546 114854
rect 113782 114618 113866 114854
rect 114102 114618 149546 114854
rect 149782 114618 149866 114854
rect 150102 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 588810 114854
rect -4886 114586 588810 114618
rect -2966 111454 586890 111486
rect -2966 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 204250 111454
rect 204486 111218 234970 111454
rect 235206 111218 265690 111454
rect 265926 111218 296410 111454
rect 296646 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 586890 111454
rect -2966 111134 586890 111218
rect -2966 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 204250 111134
rect 204486 110898 234970 111134
rect 235206 110898 265690 111134
rect 265926 110898 296410 111134
rect 296646 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 586890 111134
rect -2966 110866 586890 110898
rect -8726 104614 592650 104646
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 66986 104614
rect 67222 104378 67306 104614
rect 67542 104378 102986 104614
rect 103222 104378 103306 104614
rect 103542 104378 138986 104614
rect 139222 104378 139306 104614
rect 139542 104378 174986 104614
rect 175222 104378 175306 104614
rect 175542 104378 318986 104614
rect 319222 104378 319306 104614
rect 319542 104378 354986 104614
rect 355222 104378 355306 104614
rect 355542 104378 390986 104614
rect 391222 104378 391306 104614
rect 391542 104378 426986 104614
rect 427222 104378 427306 104614
rect 427542 104378 462986 104614
rect 463222 104378 463306 104614
rect 463542 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect -8726 104294 592650 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 66986 104294
rect 67222 104058 67306 104294
rect 67542 104058 102986 104294
rect 103222 104058 103306 104294
rect 103542 104058 138986 104294
rect 139222 104058 139306 104294
rect 139542 104058 174986 104294
rect 175222 104058 175306 104294
rect 175542 104058 318986 104294
rect 319222 104058 319306 104294
rect 319542 104058 354986 104294
rect 355222 104058 355306 104294
rect 355542 104058 390986 104294
rect 391222 104058 391306 104294
rect 391542 104058 426986 104294
rect 427222 104058 427306 104294
rect 427542 104058 462986 104294
rect 463222 104058 463306 104294
rect 463542 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect -8726 104026 592650 104058
rect -6806 100894 590730 100926
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 63266 100894
rect 63502 100658 63586 100894
rect 63822 100658 99266 100894
rect 99502 100658 99586 100894
rect 99822 100658 135266 100894
rect 135502 100658 135586 100894
rect 135822 100658 171266 100894
rect 171502 100658 171586 100894
rect 171822 100658 315266 100894
rect 315502 100658 315586 100894
rect 315822 100658 351266 100894
rect 351502 100658 351586 100894
rect 351822 100658 387266 100894
rect 387502 100658 387586 100894
rect 387822 100658 423266 100894
rect 423502 100658 423586 100894
rect 423822 100658 459266 100894
rect 459502 100658 459586 100894
rect 459822 100658 495266 100894
rect 495502 100658 495586 100894
rect 495822 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect -6806 100574 590730 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 63266 100574
rect 63502 100338 63586 100574
rect 63822 100338 99266 100574
rect 99502 100338 99586 100574
rect 99822 100338 135266 100574
rect 135502 100338 135586 100574
rect 135822 100338 171266 100574
rect 171502 100338 171586 100574
rect 171822 100338 315266 100574
rect 315502 100338 315586 100574
rect 315822 100338 351266 100574
rect 351502 100338 351586 100574
rect 351822 100338 387266 100574
rect 387502 100338 387586 100574
rect 387822 100338 423266 100574
rect 423502 100338 423586 100574
rect 423822 100338 459266 100574
rect 459502 100338 459586 100574
rect 459822 100338 495266 100574
rect 495502 100338 495586 100574
rect 495822 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect -6806 100306 590730 100338
rect -4886 97174 588810 97206
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 59546 97174
rect 59782 96938 59866 97174
rect 60102 96938 95546 97174
rect 95782 96938 95866 97174
rect 96102 96938 131546 97174
rect 131782 96938 131866 97174
rect 132102 96938 167546 97174
rect 167782 96938 167866 97174
rect 168102 96938 203546 97174
rect 203782 96938 203866 97174
rect 204102 96938 239546 97174
rect 239782 96938 239866 97174
rect 240102 96938 275546 97174
rect 275782 96938 275866 97174
rect 276102 96938 311546 97174
rect 311782 96938 311866 97174
rect 312102 96938 347546 97174
rect 347782 96938 347866 97174
rect 348102 96938 383546 97174
rect 383782 96938 383866 97174
rect 384102 96938 419546 97174
rect 419782 96938 419866 97174
rect 420102 96938 455546 97174
rect 455782 96938 455866 97174
rect 456102 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect -4886 96854 588810 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 59546 96854
rect 59782 96618 59866 96854
rect 60102 96618 95546 96854
rect 95782 96618 95866 96854
rect 96102 96618 131546 96854
rect 131782 96618 131866 96854
rect 132102 96618 167546 96854
rect 167782 96618 167866 96854
rect 168102 96618 203546 96854
rect 203782 96618 203866 96854
rect 204102 96618 239546 96854
rect 239782 96618 239866 96854
rect 240102 96618 275546 96854
rect 275782 96618 275866 96854
rect 276102 96618 311546 96854
rect 311782 96618 311866 96854
rect 312102 96618 347546 96854
rect 347782 96618 347866 96854
rect 348102 96618 383546 96854
rect 383782 96618 383866 96854
rect 384102 96618 419546 96854
rect 419782 96618 419866 96854
rect 420102 96618 455546 96854
rect 455782 96618 455866 96854
rect 456102 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect -4886 96586 588810 96618
rect -2966 93454 586890 93486
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 127826 93454
rect 128062 93218 128146 93454
rect 128382 93218 163826 93454
rect 164062 93218 164146 93454
rect 164382 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect -2966 93134 586890 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 127826 93134
rect 128062 92898 128146 93134
rect 128382 92898 163826 93134
rect 164062 92898 164146 93134
rect 164382 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect -2966 92866 586890 92898
rect -8726 86614 592650 86646
rect -8726 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 120986 86614
rect 121222 86378 121306 86614
rect 121542 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 192986 86614
rect 193222 86378 193306 86614
rect 193542 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 120986 86294
rect 121222 86058 121306 86294
rect 121542 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 192986 86294
rect 193222 86058 193306 86294
rect 193542 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 592650 86294
rect -8726 86026 592650 86058
rect -6806 82894 590730 82926
rect -6806 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 117266 82894
rect 117502 82658 117586 82894
rect 117822 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 189266 82894
rect 189502 82658 189586 82894
rect 189822 82658 225266 82894
rect 225502 82658 225586 82894
rect 225822 82658 261266 82894
rect 261502 82658 261586 82894
rect 261822 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 590730 82894
rect -6806 82574 590730 82658
rect -6806 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 117266 82574
rect 117502 82338 117586 82574
rect 117822 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 189266 82574
rect 189502 82338 189586 82574
rect 189822 82338 225266 82574
rect 225502 82338 225586 82574
rect 225822 82338 261266 82574
rect 261502 82338 261586 82574
rect 261822 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 590730 82574
rect -6806 82306 590730 82338
rect -4886 79174 588810 79206
rect -4886 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 588810 79174
rect -4886 78854 588810 78938
rect -4886 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 588810 78854
rect -4886 78586 588810 78618
rect -2966 75454 586890 75486
rect -2966 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 586890 75454
rect -2966 75134 586890 75218
rect -2966 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 586890 75134
rect -2966 74866 586890 74898
rect -8726 68614 592650 68646
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 66986 68614
rect 67222 68378 67306 68614
rect 67542 68378 102986 68614
rect 103222 68378 103306 68614
rect 103542 68378 138986 68614
rect 139222 68378 139306 68614
rect 139542 68378 174986 68614
rect 175222 68378 175306 68614
rect 175542 68378 210986 68614
rect 211222 68378 211306 68614
rect 211542 68378 246986 68614
rect 247222 68378 247306 68614
rect 247542 68378 282986 68614
rect 283222 68378 283306 68614
rect 283542 68378 318986 68614
rect 319222 68378 319306 68614
rect 319542 68378 354986 68614
rect 355222 68378 355306 68614
rect 355542 68378 390986 68614
rect 391222 68378 391306 68614
rect 391542 68378 426986 68614
rect 427222 68378 427306 68614
rect 427542 68378 462986 68614
rect 463222 68378 463306 68614
rect 463542 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect -8726 68294 592650 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 66986 68294
rect 67222 68058 67306 68294
rect 67542 68058 102986 68294
rect 103222 68058 103306 68294
rect 103542 68058 138986 68294
rect 139222 68058 139306 68294
rect 139542 68058 174986 68294
rect 175222 68058 175306 68294
rect 175542 68058 210986 68294
rect 211222 68058 211306 68294
rect 211542 68058 246986 68294
rect 247222 68058 247306 68294
rect 247542 68058 282986 68294
rect 283222 68058 283306 68294
rect 283542 68058 318986 68294
rect 319222 68058 319306 68294
rect 319542 68058 354986 68294
rect 355222 68058 355306 68294
rect 355542 68058 390986 68294
rect 391222 68058 391306 68294
rect 391542 68058 426986 68294
rect 427222 68058 427306 68294
rect 427542 68058 462986 68294
rect 463222 68058 463306 68294
rect 463542 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect -8726 68026 592650 68058
rect -6806 64894 590730 64926
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 63266 64894
rect 63502 64658 63586 64894
rect 63822 64658 99266 64894
rect 99502 64658 99586 64894
rect 99822 64658 135266 64894
rect 135502 64658 135586 64894
rect 135822 64658 171266 64894
rect 171502 64658 171586 64894
rect 171822 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 243266 64894
rect 243502 64658 243586 64894
rect 243822 64658 279266 64894
rect 279502 64658 279586 64894
rect 279822 64658 315266 64894
rect 315502 64658 315586 64894
rect 315822 64658 351266 64894
rect 351502 64658 351586 64894
rect 351822 64658 387266 64894
rect 387502 64658 387586 64894
rect 387822 64658 423266 64894
rect 423502 64658 423586 64894
rect 423822 64658 459266 64894
rect 459502 64658 459586 64894
rect 459822 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect -6806 64574 590730 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 63266 64574
rect 63502 64338 63586 64574
rect 63822 64338 99266 64574
rect 99502 64338 99586 64574
rect 99822 64338 135266 64574
rect 135502 64338 135586 64574
rect 135822 64338 171266 64574
rect 171502 64338 171586 64574
rect 171822 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 243266 64574
rect 243502 64338 243586 64574
rect 243822 64338 279266 64574
rect 279502 64338 279586 64574
rect 279822 64338 315266 64574
rect 315502 64338 315586 64574
rect 315822 64338 351266 64574
rect 351502 64338 351586 64574
rect 351822 64338 387266 64574
rect 387502 64338 387586 64574
rect 387822 64338 423266 64574
rect 423502 64338 423586 64574
rect 423822 64338 459266 64574
rect 459502 64338 459586 64574
rect 459822 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect -6806 64306 590730 64338
rect -4886 61174 588810 61206
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 59546 61174
rect 59782 60938 59866 61174
rect 60102 60938 95546 61174
rect 95782 60938 95866 61174
rect 96102 60938 131546 61174
rect 131782 60938 131866 61174
rect 132102 60938 167546 61174
rect 167782 60938 167866 61174
rect 168102 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 239546 61174
rect 239782 60938 239866 61174
rect 240102 60938 275546 61174
rect 275782 60938 275866 61174
rect 276102 60938 311546 61174
rect 311782 60938 311866 61174
rect 312102 60938 347546 61174
rect 347782 60938 347866 61174
rect 348102 60938 383546 61174
rect 383782 60938 383866 61174
rect 384102 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect -4886 60854 588810 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 59546 60854
rect 59782 60618 59866 60854
rect 60102 60618 95546 60854
rect 95782 60618 95866 60854
rect 96102 60618 131546 60854
rect 131782 60618 131866 60854
rect 132102 60618 167546 60854
rect 167782 60618 167866 60854
rect 168102 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 239546 60854
rect 239782 60618 239866 60854
rect 240102 60618 275546 60854
rect 275782 60618 275866 60854
rect 276102 60618 311546 60854
rect 311782 60618 311866 60854
rect 312102 60618 347546 60854
rect 347782 60618 347866 60854
rect 348102 60618 383546 60854
rect 383782 60618 383866 60854
rect 384102 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect -4886 60586 588810 60618
rect -2966 57454 586890 57486
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect -2966 57134 586890 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect -2966 56866 586890 56898
rect -8726 50614 592650 50646
rect -8726 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 592650 50294
rect -8726 50026 592650 50058
rect -6806 46894 590730 46926
rect -6806 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 590730 46894
rect -6806 46574 590730 46658
rect -6806 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 590730 46574
rect -6806 46306 590730 46338
rect -4886 43174 588810 43206
rect -4886 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 588810 43174
rect -4886 42854 588810 42938
rect -4886 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 588810 42854
rect -4886 42586 588810 42618
rect -2966 39454 586890 39486
rect -2966 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 586890 39454
rect -2966 39134 586890 39218
rect -2966 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 586890 39134
rect -2966 38866 586890 38898
rect -8726 32614 592650 32646
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect -8726 32294 592650 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect -8726 32026 592650 32058
rect -6806 28894 590730 28926
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect -6806 28574 590730 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect -6806 28306 590730 28338
rect -4886 25174 588810 25206
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect -4886 24854 588810 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect -4886 24586 588810 24618
rect -2966 21454 586890 21486
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect -2966 21134 586890 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect -2966 20866 586890 20898
rect -8726 14614 592650 14646
rect -8726 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 592650 14294
rect -8726 14026 592650 14058
rect -6806 10894 590730 10926
rect -6806 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 590730 10894
rect -6806 10574 590730 10658
rect -6806 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 590730 10574
rect -6806 10306 590730 10338
rect -4886 7174 588810 7206
rect -4886 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 588810 7174
rect -4886 6854 588810 6938
rect -4886 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 588810 6854
rect -4886 6586 588810 6618
rect -2966 3454 586890 3486
rect -2966 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 586890 3454
rect -2966 3134 586890 3218
rect -2966 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 586890 3134
rect -2966 2866 586890 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use ringosc_macro  ring1
timestamp 1635131530
transform 1 0 160000 0 1 160000
box 934 0 10000 29504
use collapsering_macro  ring0
timestamp 1635131530
transform 1 0 160000 0 1 124000
box 934 0 10000 29776
use digitalcore_macro  digitalcore
timestamp 1635131530
transform 1 0 200000 0 1 100000
box 0 0 99898 100000
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 38866 586890 39486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 74866 586890 75486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 110866 586890 111486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 146866 586890 147486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 182866 586890 183486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 218866 586890 219486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 254866 586890 255486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 290866 586890 291486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 326866 586890 327486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 362866 586890 363486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 398866 586890 399486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 434866 586890 435486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 470866 586890 471486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 506866 586890 507486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 542866 586890 543486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 578866 586890 579486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 614866 586890 615486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 650866 586890 651486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 686866 586890 687486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 -1894 218414 98000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 -1894 254414 98000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 -1894 290414 98000 6 vccd1
port 531 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 1794 -1894 2414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 -1894 38414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 -1894 74414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 -1894 110414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 -1894 146414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 -1894 182414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 202000 218414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 202000 254414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 202000 290414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 -1894 326414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 -1894 362414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 -1894 398414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 -1894 434414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 -1894 470414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 -1894 506414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 -1894 542414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 577794 -1894 578414 705830 6 vccd1
port 531 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 532 nsew power input
rlabel metal5 s -4886 6586 588810 7206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 42586 588810 43206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 78586 588810 79206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 114586 588810 115206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 150586 588810 151206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 186586 588810 187206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 222586 588810 223206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 258586 588810 259206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 294586 588810 295206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 330586 588810 331206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 366586 588810 367206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 402586 588810 403206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 438586 588810 439206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 474586 588810 475206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 510586 588810 511206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 546586 588810 547206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 582586 588810 583206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 618586 588810 619206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 654586 588810 655206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 690586 588810 691206 6 vccd2
port 532 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 -3814 222134 98000 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 -3814 258134 98000 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 -3814 294134 98000 6 vccd2
port 532 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 532 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 5514 -3814 6134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 41514 -3814 42134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 -3814 78134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 -3814 114134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 -3814 150134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 -3814 186134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 202000 222134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 202000 258134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 202000 294134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 -3814 330134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 -3814 366134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 -3814 402134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 -3814 438134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 -3814 474134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 -3814 510134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 545514 -3814 546134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 581514 -3814 582134 707750 6 vccd2
port 532 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 533 nsew power input
rlabel metal5 s -6806 10306 590730 10926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 46306 590730 46926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 82306 590730 82926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 118306 590730 118926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 154306 590730 154926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 190306 590730 190926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 226306 590730 226926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 262306 590730 262926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 298306 590730 298926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 334306 590730 334926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 370306 590730 370926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 406306 590730 406926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 442306 590730 442926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 478306 590730 478926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 514306 590730 514926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 550306 590730 550926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 586306 590730 586926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 622306 590730 622926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 658306 590730 658926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 694306 590730 694926 6 vdda1
port 533 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 -5734 225854 98000 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 -5734 261854 98000 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 -5734 297854 98000 6 vdda1
port 533 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 533 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 9234 -5734 9854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 45234 -5734 45854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 -5734 81854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 -5734 117854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 -5734 153854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 -5734 189854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 202000 225854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 202000 261854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 202000 297854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 -5734 333854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 -5734 369854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 -5734 405854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 -5734 441854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 -5734 477854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 -5734 513854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 549234 -5734 549854 709670 6 vdda1
port 533 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 534 nsew power input
rlabel metal5 s -8726 14026 592650 14646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 50026 592650 50646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 86026 592650 86646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 122026 592650 122646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 158026 592650 158646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 194026 592650 194646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 230026 592650 230646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 266026 592650 266646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 302026 592650 302646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 338026 592650 338646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 374026 592650 374646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 410026 592650 410646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 446026 592650 446646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 482026 592650 482646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 518026 592650 518646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 554026 592650 554646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 590026 592650 590646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 626026 592650 626646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 662026 592650 662646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 698026 592650 698646 6 vdda2
port 534 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 -7654 229574 98000 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 -7654 265574 98000 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 -7654 301574 98000 6 vdda2
port 534 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 534 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 12954 -7654 13574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 -7654 49574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 -7654 85574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 -7654 121574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 -7654 157574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 -7654 193574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 202000 229574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 202000 265574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 202000 301574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 -7654 337574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 -7654 373574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 -7654 409574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 -7654 445574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 -7654 481574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 -7654 517574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 552954 -7654 553574 711590 6 vdda2
port 534 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 28306 590730 28926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 64306 590730 64926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 100306 590730 100926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 136306 590730 136926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 172306 590730 172926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 208306 590730 208926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 244306 590730 244926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 280306 590730 280926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 316306 590730 316926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 352306 590730 352926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 388306 590730 388926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 424306 590730 424926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 460306 590730 460926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 496306 590730 496926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 532306 590730 532926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 568306 590730 568926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 604306 590730 604926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 640306 590730 640926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 676306 590730 676926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 -5734 207854 98000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 -5734 243854 98000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 -5734 279854 98000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 -5734 171854 122000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 156000 171854 158000 6 vssa1
port 535 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 535 nsew ground input
rlabel metal4 s 27234 -5734 27854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 -5734 63854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 -5734 99854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 -5734 135854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 192000 171854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 202000 207854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 202000 243854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 202000 279854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 -5734 315854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 -5734 351854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 -5734 387854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 -5734 423854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 -5734 459854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 -5734 495854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 -5734 531854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 567234 -5734 567854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 32026 592650 32646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 68026 592650 68646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 104026 592650 104646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 140026 592650 140646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 176026 592650 176646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 212026 592650 212646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 248026 592650 248646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 284026 592650 284646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 320026 592650 320646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 356026 592650 356646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 392026 592650 392646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 428026 592650 428646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 464026 592650 464646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 500026 592650 500646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 536026 592650 536646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 572026 592650 572646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 608026 592650 608646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 644026 592650 644646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 680026 592650 680646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 -7654 211574 98000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 -7654 247574 98000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 -7654 283574 98000 6 vssa2
port 536 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 536 nsew ground input
rlabel metal4 s 30954 -7654 31574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 -7654 67574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 -7654 103574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 -7654 139574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 -7654 175574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 202000 211574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 202000 247574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 202000 283574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 -7654 319574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 -7654 355574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 -7654 391574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 -7654 427574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 -7654 463574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 -7654 499574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 -7654 535574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 570954 -7654 571574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 20866 586890 21486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 56866 586890 57486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 92866 586890 93486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 128866 586890 129486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 164866 586890 165486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 200866 586890 201486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 236866 586890 237486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 272866 586890 273486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 308866 586890 309486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 344866 586890 345486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 380866 586890 381486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 416866 586890 417486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 452866 586890 453486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 488866 586890 489486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 524866 586890 525486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 560866 586890 561486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 596866 586890 597486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 632866 586890 633486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 668866 586890 669486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 -1894 200414 98000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 -1894 236414 98000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 -1894 272414 98000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 -1894 164414 122000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 156000 164414 158000 6 vssd1
port 537 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 537 nsew ground input
rlabel metal4 s 19794 -1894 20414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 -1894 56414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 -1894 92414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 -1894 128414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 192000 164414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 202000 200414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 202000 236414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 202000 272414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 -1894 308414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 -1894 344414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 -1894 380414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 -1894 416414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 -1894 452414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 -1894 488414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 -1894 524414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 559794 -1894 560414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 24586 588810 25206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 60586 588810 61206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 96586 588810 97206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 132586 588810 133206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 168586 588810 169206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 204586 588810 205206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 240586 588810 241206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 276586 588810 277206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 312586 588810 313206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 348586 588810 349206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 384586 588810 385206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 420586 588810 421206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 456586 588810 457206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 492586 588810 493206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 528586 588810 529206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 564586 588810 565206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 600586 588810 601206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 636586 588810 637206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 672586 588810 673206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 -3814 204134 98000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 -3814 240134 98000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 -3814 276134 98000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 -3814 168134 122000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 156000 168134 158000 6 vssd2
port 538 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 538 nsew ground input
rlabel metal4 s 23514 -3814 24134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 -3814 60134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 -3814 96134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 -3814 132134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 192000 168134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 202000 204134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 202000 240134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 202000 276134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 -3814 312134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 -3814 348134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 -3814 384134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 -3814 420134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 -3814 456134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 -3814 492134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 -3814 528134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 563514 -3814 564134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 539 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 540 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 541 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 542 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 543 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 544 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 545 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 546 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 547 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 548 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 549 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 550 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 551 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 552 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 553 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 554 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 555 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 556 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 557 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 558 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 559 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 560 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 561 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 562 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 563 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 564 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 565 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 566 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 567 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 568 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 569 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 570 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 571 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 572 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 573 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 574 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 575 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 576 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 577 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 578 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 579 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 580 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 581 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 582 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 583 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 584 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 585 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 586 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 587 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 588 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 589 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 590 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 591 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 592 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 593 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 594 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 595 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 596 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 597 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 598 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 599 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 600 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 601 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 602 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 603 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 604 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 605 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 606 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 607 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 608 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 609 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 610 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 611 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 612 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 613 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 614 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 615 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 616 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 617 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 618 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 619 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 620 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 621 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 622 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 623 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 624 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 625 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 626 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 627 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 628 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 629 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 630 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 631 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 632 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 633 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 634 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 635 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 636 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 637 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 638 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 639 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 640 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 641 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 642 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 643 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
