magic
tech sky130A
magscale 1 2
timestamp 1636514986
<< viali >>
rect 7113 27489 7147 27523
rect 7573 27421 7607 27455
rect 7021 27353 7055 27387
rect 6469 27285 6503 27319
rect 8033 27285 8067 27319
rect 6561 27081 6595 27115
rect 6377 26945 6411 26979
rect 7573 26945 7607 26979
rect 8033 26945 8067 26979
rect 7021 26877 7055 26911
rect 7113 26809 7147 26843
rect 5273 26537 5307 26571
rect 6837 26469 6871 26503
rect 5365 26333 5399 26367
rect 5917 26333 5951 26367
rect 6101 26333 6135 26367
rect 6837 26333 6871 26367
rect 8125 26333 8159 26367
rect 6837 25925 6871 25959
rect 7113 25925 7147 25959
rect 5825 25857 5859 25891
rect 7757 25857 7791 25891
rect 6837 25381 6871 25415
rect 7205 25245 7239 25279
rect 8125 25245 8159 25279
rect 6101 25109 6135 25143
rect 7665 24837 7699 24871
rect 7113 24769 7147 24803
rect 7021 24701 7055 24735
rect 7573 24701 7607 24735
rect 8125 24701 8159 24735
rect 6469 24565 6503 24599
rect 6101 24225 6135 24259
rect 6561 24157 6595 24191
rect 7389 24157 7423 24191
rect 8125 24157 8159 24191
rect 7205 24089 7239 24123
rect 6745 24021 6779 24055
rect 5825 23817 5859 23851
rect 6929 23817 6963 23851
rect 7573 23749 7607 23783
rect 7021 23681 7055 23715
rect 7665 23681 7699 23715
rect 8125 23681 8159 23715
rect 5641 23205 5675 23239
rect 6101 23069 6135 23103
rect 6745 23069 6779 23103
rect 7665 23069 7699 23103
rect 6929 23001 6963 23035
rect 6285 22933 6319 22967
rect 6837 22661 6871 22695
rect 6929 22661 6963 22695
rect 7849 22661 7883 22695
rect 8033 22661 8067 22695
rect 5825 22593 5859 22627
rect 5181 22525 5215 22559
rect 7389 22525 7423 22559
rect 5733 22389 5767 22423
rect 6377 21981 6411 22015
rect 7849 21981 7883 22015
rect 7941 21913 7975 21947
rect 5365 21845 5399 21879
rect 5917 21845 5951 21879
rect 6837 21573 6871 21607
rect 6929 21573 6963 21607
rect 7941 21573 7975 21607
rect 5641 21505 5675 21539
rect 7389 21437 7423 21471
rect 8125 21369 8159 21403
rect 5181 21301 5215 21335
rect 5733 21301 5767 21335
rect 6285 21029 6319 21063
rect 6193 20961 6227 20995
rect 5181 20893 5215 20927
rect 6745 20893 6779 20927
rect 8125 20893 8159 20927
rect 5641 20825 5675 20859
rect 5733 20825 5767 20859
rect 7205 20825 7239 20859
rect 7389 20825 7423 20859
rect 4721 20757 4755 20791
rect 5181 20553 5215 20587
rect 5641 20553 5675 20587
rect 6561 20485 6595 20519
rect 5825 20417 5859 20451
rect 7205 20417 7239 20451
rect 8125 20417 8159 20451
rect 6009 20009 6043 20043
rect 6561 19805 6595 19839
rect 7481 19805 7515 19839
rect 8125 19805 8159 19839
rect 7205 19737 7239 19771
rect 5549 19669 5583 19703
rect 7941 19669 7975 19703
rect 8033 19465 8067 19499
rect 7205 19397 7239 19431
rect 7297 19397 7331 19431
rect 7941 19329 7975 19363
rect 6745 19261 6779 19295
rect 6745 18921 6779 18955
rect 7205 18717 7239 18751
rect 7849 18649 7883 18683
rect 7297 18581 7331 18615
rect 6377 18241 6411 18275
rect 7849 18241 7883 18275
rect 7849 18105 7883 18139
rect 5733 18037 5767 18071
rect 5365 17697 5399 17731
rect 5825 17697 5859 17731
rect 6285 17697 6319 17731
rect 7389 17697 7423 17731
rect 6837 17629 6871 17663
rect 8125 17629 8159 17663
rect 6377 17561 6411 17595
rect 7297 17561 7331 17595
rect 7941 17493 7975 17527
rect 6561 17221 6595 17255
rect 7205 17153 7239 17187
rect 8125 17153 8159 17187
rect 5825 16949 5859 16983
rect 5181 16745 5215 16779
rect 6653 16677 6687 16711
rect 5733 16609 5767 16643
rect 6193 16609 6227 16643
rect 7389 16541 7423 16575
rect 8125 16541 8159 16575
rect 6745 16473 6779 16507
rect 7205 16473 7239 16507
rect 8033 16201 8067 16235
rect 6561 16133 6595 16167
rect 7941 16133 7975 16167
rect 5641 16065 5675 16099
rect 6745 16065 6779 16099
rect 7481 16065 7515 16099
rect 5181 15997 5215 16031
rect 5825 15861 5859 15895
rect 4813 15657 4847 15691
rect 6561 15589 6595 15623
rect 5365 15521 5399 15555
rect 6469 15521 6503 15555
rect 7021 15521 7055 15555
rect 8033 15521 8067 15555
rect 6009 15453 6043 15487
rect 7573 15453 7607 15487
rect 5825 15385 5859 15419
rect 7481 15385 7515 15419
rect 5089 15113 5123 15147
rect 5733 15113 5767 15147
rect 5641 15045 5675 15079
rect 6561 14977 6595 15011
rect 6745 14977 6779 15011
rect 7205 14977 7239 15011
rect 7389 14977 7423 15011
rect 8125 14977 8159 15011
rect 4537 14841 4571 14875
rect 6469 14773 6503 14807
rect 5549 14501 5583 14535
rect 7389 14501 7423 14535
rect 5641 14433 5675 14467
rect 5089 14365 5123 14399
rect 6101 14365 6135 14399
rect 7021 14365 7055 14399
rect 6561 13889 6595 13923
rect 7481 13889 7515 13923
rect 7849 13753 7883 13787
rect 5825 13685 5859 13719
rect 5733 13481 5767 13515
rect 7113 13481 7147 13515
rect 7665 13413 7699 13447
rect 6929 13277 6963 13311
rect 8125 13277 8159 13311
rect 7573 13209 7607 13243
rect 6377 13141 6411 13175
rect 7297 12937 7331 12971
rect 7389 12937 7423 12971
rect 8033 12801 8067 12835
rect 6745 12733 6779 12767
rect 7849 12597 7883 12631
rect 6745 12325 6779 12359
rect 7757 12257 7791 12291
rect 6377 12189 6411 12223
rect 7205 12189 7239 12223
rect 7665 12121 7699 12155
rect 5825 12053 5859 12087
rect 6745 12053 6779 12087
rect 7021 11781 7055 11815
rect 6837 11713 6871 11747
rect 7573 11713 7607 11747
rect 7481 11645 7515 11679
rect 8033 11645 8067 11679
rect 5825 11577 5859 11611
rect 5457 11305 5491 11339
rect 6009 11305 6043 11339
rect 6837 11237 6871 11271
rect 7205 11101 7239 11135
rect 8125 11101 8159 11135
rect 6101 11033 6135 11067
rect 7297 10693 7331 10727
rect 6469 10625 6503 10659
rect 6653 10625 6687 10659
rect 7113 10625 7147 10659
rect 8033 10625 8067 10659
rect 5825 10557 5859 10591
rect 7573 10081 7607 10115
rect 7113 10013 7147 10047
rect 7665 10013 7699 10047
rect 8125 10013 8159 10047
rect 6929 9945 6963 9979
rect 6469 9877 6503 9911
rect 5825 9537 5859 9571
rect 6469 9537 6503 9571
rect 7113 9537 7147 9571
rect 7389 9537 7423 9571
rect 8033 9537 8067 9571
rect 7849 9333 7883 9367
rect 5549 9129 5583 9163
rect 7113 9061 7147 9095
rect 6653 8993 6687 9027
rect 7205 8993 7239 9027
rect 6193 8925 6227 8959
rect 7757 8857 7791 8891
rect 4997 8789 5031 8823
rect 6101 8789 6135 8823
rect 7849 8789 7883 8823
rect 4813 8585 4847 8619
rect 5825 8517 5859 8551
rect 4629 8449 4663 8483
rect 7205 8449 7239 8483
rect 8125 8449 8159 8483
rect 5273 8381 5307 8415
rect 5733 8381 5767 8415
rect 6561 8381 6595 8415
rect 4169 8313 4203 8347
rect 4905 8041 4939 8075
rect 5549 7973 5583 8007
rect 3249 7905 3283 7939
rect 4813 7837 4847 7871
rect 5733 7837 5767 7871
rect 7389 7837 7423 7871
rect 8125 7837 8159 7871
rect 4353 7769 4387 7803
rect 7205 7769 7239 7803
rect 5733 7497 5767 7531
rect 5733 7361 5767 7395
rect 6377 7361 6411 7395
rect 7849 7361 7883 7395
rect 3985 7293 4019 7327
rect 4537 7293 4571 7327
rect 7849 7225 7883 7259
rect 5089 7157 5123 7191
rect 5089 6817 5123 6851
rect 7389 6817 7423 6851
rect 4445 6749 4479 6783
rect 7941 6749 7975 6783
rect 4537 6681 4571 6715
rect 5365 6681 5399 6715
rect 7481 6681 7515 6715
rect 6837 6613 6871 6647
rect 5641 6341 5675 6375
rect 5089 6273 5123 6307
rect 8125 6273 8159 6307
rect 5825 6205 5859 6239
rect 6929 6205 6963 6239
rect 7481 6205 7515 6239
rect 3893 6137 3927 6171
rect 4445 6137 4479 6171
rect 7389 6137 7423 6171
rect 7941 6137 7975 6171
rect 4997 6069 5031 6103
rect 6377 6069 6411 6103
rect 5273 5729 5307 5763
rect 4537 5661 4571 5695
rect 6377 5661 6411 5695
rect 6837 5661 6871 5695
rect 7757 5661 7791 5695
rect 3249 5593 3283 5627
rect 5825 5593 5859 5627
rect 5917 5593 5951 5627
rect 7021 5593 7055 5627
rect 4077 5525 4111 5559
rect 4721 5525 4755 5559
rect 5365 5525 5399 5559
rect 2605 5321 2639 5355
rect 5089 5321 5123 5355
rect 6561 5321 6595 5355
rect 7389 5253 7423 5287
rect 4353 5185 4387 5219
rect 5181 5185 5215 5219
rect 6653 5185 6687 5219
rect 7205 5185 7239 5219
rect 8125 5185 8159 5219
rect 4905 5117 4939 5151
rect 3617 5049 3651 5083
rect 5549 5049 5583 5083
rect 3157 4981 3191 5015
rect 4261 4981 4295 5015
rect 4353 4641 4387 4675
rect 7573 4641 7607 4675
rect 4445 4573 4479 4607
rect 4721 4573 4755 4607
rect 7113 4573 7147 4607
rect 8125 4573 8159 4607
rect 4169 4505 4203 4539
rect 6837 4505 6871 4539
rect 7665 4505 7699 4539
rect 2697 4437 2731 4471
rect 3157 4437 3191 4471
rect 5365 4437 5399 4471
rect 3341 4233 3375 4267
rect 4629 4233 4663 4267
rect 5457 4233 5491 4267
rect 6561 4165 6595 4199
rect 2789 4097 2823 4131
rect 3157 4097 3191 4131
rect 4261 4097 4295 4131
rect 7205 4097 7239 4131
rect 8125 4097 8159 4131
rect 3249 4029 3283 4063
rect 4077 4029 4111 4063
rect 4169 4029 4203 4063
rect 5549 4029 5583 4063
rect 5641 4029 5675 4063
rect 2237 3961 2271 3995
rect 1777 3893 1811 3927
rect 5089 3893 5123 3927
rect 7205 3689 7239 3723
rect 2697 3621 2731 3655
rect 4997 3553 5031 3587
rect 5457 3553 5491 3587
rect 7849 3553 7883 3587
rect 4353 3485 4387 3519
rect 4629 3485 4663 3519
rect 4813 3485 4847 3519
rect 5733 3417 5767 3451
rect 8033 3417 8067 3451
rect 3157 3349 3191 3383
rect 3893 3349 3927 3383
rect 4997 3145 5031 3179
rect 5365 3145 5399 3179
rect 5457 3145 5491 3179
rect 4353 3077 4387 3111
rect 4261 3009 4295 3043
rect 6561 3009 6595 3043
rect 7481 3009 7515 3043
rect 3709 2941 3743 2975
rect 5549 2941 5583 2975
rect 7849 2873 7883 2907
rect 2697 2805 2731 2839
rect 3249 2805 3283 2839
rect 3157 2601 3191 2635
rect 6469 2601 6503 2635
rect 5181 2465 5215 2499
rect 5733 2465 5767 2499
rect 7205 2465 7239 2499
rect 4537 2397 4571 2431
rect 4813 2397 4847 2431
rect 4997 2397 5031 2431
rect 5641 2397 5675 2431
rect 6561 2397 6595 2431
rect 7113 2397 7147 2431
rect 7665 2397 7699 2431
rect 4077 2329 4111 2363
<< metal1 >>
rect 1104 27770 8832 27792
rect 1104 27718 2248 27770
rect 2300 27718 2312 27770
rect 2364 27718 2376 27770
rect 2428 27718 2440 27770
rect 2492 27718 2504 27770
rect 2556 27718 4846 27770
rect 4898 27718 4910 27770
rect 4962 27718 4974 27770
rect 5026 27718 5038 27770
rect 5090 27718 5102 27770
rect 5154 27718 7443 27770
rect 7495 27718 7507 27770
rect 7559 27718 7571 27770
rect 7623 27718 7635 27770
rect 7687 27718 7699 27770
rect 7751 27718 8832 27770
rect 1104 27696 8832 27718
rect 7006 27480 7012 27532
rect 7064 27520 7070 27532
rect 7101 27523 7159 27529
rect 7101 27520 7113 27523
rect 7064 27492 7113 27520
rect 7064 27480 7070 27492
rect 7101 27489 7113 27492
rect 7147 27489 7159 27523
rect 7101 27483 7159 27489
rect 7561 27455 7619 27461
rect 7561 27421 7573 27455
rect 7607 27452 7619 27455
rect 7607 27424 7880 27452
rect 7607 27421 7619 27424
rect 7561 27415 7619 27421
rect 6546 27344 6552 27396
rect 6604 27384 6610 27396
rect 7009 27387 7067 27393
rect 7009 27384 7021 27387
rect 6604 27356 7021 27384
rect 6604 27344 6610 27356
rect 7009 27353 7021 27356
rect 7055 27353 7067 27387
rect 7009 27347 7067 27353
rect 7852 27328 7880 27424
rect 5902 27276 5908 27328
rect 5960 27316 5966 27328
rect 6457 27319 6515 27325
rect 6457 27316 6469 27319
rect 5960 27288 6469 27316
rect 5960 27276 5966 27288
rect 6457 27285 6469 27288
rect 6503 27285 6515 27319
rect 6457 27279 6515 27285
rect 7834 27276 7840 27328
rect 7892 27316 7898 27328
rect 8021 27319 8079 27325
rect 8021 27316 8033 27319
rect 7892 27288 8033 27316
rect 7892 27276 7898 27288
rect 8021 27285 8033 27288
rect 8067 27285 8079 27319
rect 8021 27279 8079 27285
rect 1104 27226 8832 27248
rect 1104 27174 3547 27226
rect 3599 27174 3611 27226
rect 3663 27174 3675 27226
rect 3727 27174 3739 27226
rect 3791 27174 3803 27226
rect 3855 27174 6144 27226
rect 6196 27174 6208 27226
rect 6260 27174 6272 27226
rect 6324 27174 6336 27226
rect 6388 27174 6400 27226
rect 6452 27174 8832 27226
rect 1104 27152 8832 27174
rect 6546 27112 6552 27124
rect 6507 27084 6552 27112
rect 6546 27072 6552 27084
rect 6604 27072 6610 27124
rect 5902 27004 5908 27056
rect 5960 27044 5966 27056
rect 5960 27016 7604 27044
rect 5960 27004 5966 27016
rect 6362 26976 6368 26988
rect 6323 26948 6368 26976
rect 6362 26936 6368 26948
rect 6420 26936 6426 26988
rect 7576 26985 7604 27016
rect 7561 26979 7619 26985
rect 7561 26945 7573 26979
rect 7607 26976 7619 26979
rect 8021 26979 8079 26985
rect 8021 26976 8033 26979
rect 7607 26948 8033 26976
rect 7607 26945 7619 26948
rect 7561 26939 7619 26945
rect 8021 26945 8033 26948
rect 8067 26976 8079 26979
rect 8110 26976 8116 26988
rect 8067 26948 8116 26976
rect 8067 26945 8079 26948
rect 8021 26939 8079 26945
rect 8110 26936 8116 26948
rect 8168 26936 8174 26988
rect 5258 26868 5264 26920
rect 5316 26908 5322 26920
rect 7009 26911 7067 26917
rect 7009 26908 7021 26911
rect 5316 26880 7021 26908
rect 5316 26868 5322 26880
rect 7009 26877 7021 26880
rect 7055 26877 7067 26911
rect 7009 26871 7067 26877
rect 7098 26840 7104 26852
rect 7059 26812 7104 26840
rect 7098 26800 7104 26812
rect 7156 26800 7162 26852
rect 1104 26682 8832 26704
rect 1104 26630 2248 26682
rect 2300 26630 2312 26682
rect 2364 26630 2376 26682
rect 2428 26630 2440 26682
rect 2492 26630 2504 26682
rect 2556 26630 4846 26682
rect 4898 26630 4910 26682
rect 4962 26630 4974 26682
rect 5026 26630 5038 26682
rect 5090 26630 5102 26682
rect 5154 26630 7443 26682
rect 7495 26630 7507 26682
rect 7559 26630 7571 26682
rect 7623 26630 7635 26682
rect 7687 26630 7699 26682
rect 7751 26630 8832 26682
rect 1104 26608 8832 26630
rect 5258 26568 5264 26580
rect 5219 26540 5264 26568
rect 5258 26528 5264 26540
rect 5316 26528 5322 26580
rect 6825 26503 6883 26509
rect 6825 26469 6837 26503
rect 6871 26500 6883 26503
rect 7098 26500 7104 26512
rect 6871 26472 7104 26500
rect 6871 26469 6883 26472
rect 6825 26463 6883 26469
rect 7098 26460 7104 26472
rect 7156 26500 7162 26512
rect 8018 26500 8024 26512
rect 7156 26472 8024 26500
rect 7156 26460 7162 26472
rect 8018 26460 8024 26472
rect 8076 26460 8082 26512
rect 7006 26432 7012 26444
rect 5368 26404 7012 26432
rect 5368 26373 5396 26404
rect 7006 26392 7012 26404
rect 7064 26392 7070 26444
rect 5353 26367 5411 26373
rect 5353 26333 5365 26367
rect 5399 26333 5411 26367
rect 5905 26367 5963 26373
rect 5905 26364 5917 26367
rect 5353 26327 5411 26333
rect 5828 26336 5917 26364
rect 5828 26234 5856 26336
rect 5905 26333 5917 26336
rect 5951 26333 5963 26367
rect 5905 26327 5963 26333
rect 6089 26367 6147 26373
rect 6089 26333 6101 26367
rect 6135 26364 6147 26367
rect 6362 26364 6368 26376
rect 6135 26336 6368 26364
rect 6135 26333 6147 26336
rect 6089 26327 6147 26333
rect 6362 26324 6368 26336
rect 6420 26364 6426 26376
rect 6822 26364 6828 26376
rect 6420 26336 6828 26364
rect 6420 26324 6426 26336
rect 6822 26324 6828 26336
rect 6880 26324 6886 26376
rect 8110 26364 8116 26376
rect 8071 26336 8116 26364
rect 8110 26324 8116 26336
rect 8168 26324 8174 26376
rect 5828 26228 5948 26234
rect 6914 26228 6920 26240
rect 5828 26206 6920 26228
rect 5920 26200 6920 26206
rect 6914 26188 6920 26200
rect 6972 26188 6978 26240
rect 1104 26138 8832 26160
rect 1104 26086 3547 26138
rect 3599 26086 3611 26138
rect 3663 26086 3675 26138
rect 3727 26086 3739 26138
rect 3791 26086 3803 26138
rect 3855 26086 6144 26138
rect 6196 26086 6208 26138
rect 6260 26086 6272 26138
rect 6324 26086 6336 26138
rect 6388 26086 6400 26138
rect 6452 26086 8832 26138
rect 1104 26064 8832 26086
rect 6822 25956 6828 25968
rect 6783 25928 6828 25956
rect 6822 25916 6828 25928
rect 6880 25916 6886 25968
rect 7098 25956 7104 25968
rect 7059 25928 7104 25956
rect 7098 25916 7104 25928
rect 7156 25916 7162 25968
rect 5813 25891 5871 25897
rect 5813 25857 5825 25891
rect 5859 25888 5871 25891
rect 7745 25891 7803 25897
rect 7745 25888 7757 25891
rect 5859 25860 7757 25888
rect 5859 25857 5871 25860
rect 5813 25851 5871 25857
rect 7745 25857 7757 25860
rect 7791 25888 7803 25891
rect 7834 25888 7840 25900
rect 7791 25860 7840 25888
rect 7791 25857 7803 25860
rect 7745 25851 7803 25857
rect 7834 25848 7840 25860
rect 7892 25848 7898 25900
rect 1104 25594 8832 25616
rect 1104 25542 2248 25594
rect 2300 25542 2312 25594
rect 2364 25542 2376 25594
rect 2428 25542 2440 25594
rect 2492 25542 2504 25594
rect 2556 25542 4846 25594
rect 4898 25542 4910 25594
rect 4962 25542 4974 25594
rect 5026 25542 5038 25594
rect 5090 25542 5102 25594
rect 5154 25542 7443 25594
rect 7495 25542 7507 25594
rect 7559 25542 7571 25594
rect 7623 25542 7635 25594
rect 7687 25542 7699 25594
rect 7751 25542 8832 25594
rect 1104 25520 8832 25542
rect 6825 25415 6883 25421
rect 6825 25381 6837 25415
rect 6871 25412 6883 25415
rect 6914 25412 6920 25424
rect 6871 25384 6920 25412
rect 6871 25381 6883 25384
rect 6825 25375 6883 25381
rect 6914 25372 6920 25384
rect 6972 25412 6978 25424
rect 7650 25412 7656 25424
rect 6972 25384 7656 25412
rect 6972 25372 6978 25384
rect 7650 25372 7656 25384
rect 7708 25372 7714 25424
rect 7190 25276 7196 25288
rect 7151 25248 7196 25276
rect 7190 25236 7196 25248
rect 7248 25236 7254 25288
rect 8113 25279 8171 25285
rect 8113 25245 8125 25279
rect 8159 25245 8171 25279
rect 8113 25239 8171 25245
rect 6089 25143 6147 25149
rect 6089 25109 6101 25143
rect 6135 25140 6147 25143
rect 6638 25140 6644 25152
rect 6135 25112 6644 25140
rect 6135 25109 6147 25112
rect 6089 25103 6147 25109
rect 6638 25100 6644 25112
rect 6696 25140 6702 25152
rect 8128 25140 8156 25239
rect 6696 25112 8156 25140
rect 6696 25100 6702 25112
rect 1104 25050 8832 25072
rect 1104 24998 3547 25050
rect 3599 24998 3611 25050
rect 3663 24998 3675 25050
rect 3727 24998 3739 25050
rect 3791 24998 3803 25050
rect 3855 24998 6144 25050
rect 6196 24998 6208 25050
rect 6260 24998 6272 25050
rect 6324 24998 6336 25050
rect 6388 24998 6400 25050
rect 6452 24998 8832 25050
rect 1104 24976 8832 24998
rect 7650 24868 7656 24880
rect 7611 24840 7656 24868
rect 7650 24828 7656 24840
rect 7708 24828 7714 24880
rect 7098 24800 7104 24812
rect 7059 24772 7104 24800
rect 7098 24760 7104 24772
rect 7156 24760 7162 24812
rect 7009 24735 7067 24741
rect 7009 24701 7021 24735
rect 7055 24732 7067 24735
rect 7561 24735 7619 24741
rect 7561 24732 7573 24735
rect 7055 24704 7573 24732
rect 7055 24701 7067 24704
rect 7009 24695 7067 24701
rect 7561 24701 7573 24704
rect 7607 24701 7619 24735
rect 7561 24695 7619 24701
rect 8113 24735 8171 24741
rect 8113 24701 8125 24735
rect 8159 24701 8171 24735
rect 8113 24695 8171 24701
rect 6457 24599 6515 24605
rect 6457 24565 6469 24599
rect 6503 24596 6515 24599
rect 6638 24596 6644 24608
rect 6503 24568 6644 24596
rect 6503 24565 6515 24568
rect 6457 24559 6515 24565
rect 6638 24556 6644 24568
rect 6696 24596 6702 24608
rect 8128 24596 8156 24695
rect 6696 24568 8156 24596
rect 6696 24556 6702 24568
rect 1104 24506 8832 24528
rect 1104 24454 2248 24506
rect 2300 24454 2312 24506
rect 2364 24454 2376 24506
rect 2428 24454 2440 24506
rect 2492 24454 2504 24506
rect 2556 24454 4846 24506
rect 4898 24454 4910 24506
rect 4962 24454 4974 24506
rect 5026 24454 5038 24506
rect 5090 24454 5102 24506
rect 5154 24454 7443 24506
rect 7495 24454 7507 24506
rect 7559 24454 7571 24506
rect 7623 24454 7635 24506
rect 7687 24454 7699 24506
rect 7751 24454 8832 24506
rect 1104 24432 8832 24454
rect 5810 24216 5816 24268
rect 5868 24256 5874 24268
rect 6089 24259 6147 24265
rect 6089 24256 6101 24259
rect 5868 24228 6101 24256
rect 5868 24216 5874 24228
rect 6089 24225 6101 24228
rect 6135 24256 6147 24259
rect 6135 24228 8156 24256
rect 6135 24225 6147 24228
rect 6089 24219 6147 24225
rect 8128 24200 8156 24228
rect 6549 24191 6607 24197
rect 6549 24157 6561 24191
rect 6595 24188 6607 24191
rect 6595 24160 6914 24188
rect 6595 24157 6607 24160
rect 6549 24151 6607 24157
rect 6886 24120 6914 24160
rect 7098 24148 7104 24200
rect 7156 24188 7162 24200
rect 7377 24191 7435 24197
rect 7377 24188 7389 24191
rect 7156 24160 7389 24188
rect 7156 24148 7162 24160
rect 7377 24157 7389 24160
rect 7423 24157 7435 24191
rect 8110 24188 8116 24200
rect 8071 24160 8116 24188
rect 7377 24151 7435 24157
rect 8110 24148 8116 24160
rect 8168 24148 8174 24200
rect 7190 24120 7196 24132
rect 6886 24092 7196 24120
rect 7190 24080 7196 24092
rect 7248 24080 7254 24132
rect 6733 24055 6791 24061
rect 6733 24021 6745 24055
rect 6779 24052 6791 24055
rect 7558 24052 7564 24064
rect 6779 24024 7564 24052
rect 6779 24021 6791 24024
rect 6733 24015 6791 24021
rect 7558 24012 7564 24024
rect 7616 24012 7622 24064
rect 1104 23962 8832 23984
rect 1104 23910 3547 23962
rect 3599 23910 3611 23962
rect 3663 23910 3675 23962
rect 3727 23910 3739 23962
rect 3791 23910 3803 23962
rect 3855 23910 6144 23962
rect 6196 23910 6208 23962
rect 6260 23910 6272 23962
rect 6324 23910 6336 23962
rect 6388 23910 6400 23962
rect 6452 23910 8832 23962
rect 1104 23888 8832 23910
rect 5810 23848 5816 23860
rect 5771 23820 5816 23848
rect 5810 23808 5816 23820
rect 5868 23808 5874 23860
rect 6917 23851 6975 23857
rect 6917 23817 6929 23851
rect 6963 23848 6975 23851
rect 7190 23848 7196 23860
rect 6963 23820 7196 23848
rect 6963 23817 6975 23820
rect 6917 23811 6975 23817
rect 7190 23808 7196 23820
rect 7248 23808 7254 23860
rect 7558 23780 7564 23792
rect 7519 23752 7564 23780
rect 7558 23740 7564 23752
rect 7616 23740 7622 23792
rect 6546 23672 6552 23724
rect 6604 23712 6610 23724
rect 7009 23715 7067 23721
rect 7009 23712 7021 23715
rect 6604 23684 7021 23712
rect 6604 23672 6610 23684
rect 7009 23681 7021 23684
rect 7055 23681 7067 23715
rect 7009 23675 7067 23681
rect 7098 23672 7104 23724
rect 7156 23712 7162 23724
rect 7653 23715 7711 23721
rect 7653 23712 7665 23715
rect 7156 23684 7665 23712
rect 7156 23672 7162 23684
rect 7653 23681 7665 23684
rect 7699 23681 7711 23715
rect 8110 23712 8116 23724
rect 8071 23684 8116 23712
rect 7653 23675 7711 23681
rect 8110 23672 8116 23684
rect 8168 23672 8174 23724
rect 1104 23418 8832 23440
rect 1104 23366 2248 23418
rect 2300 23366 2312 23418
rect 2364 23366 2376 23418
rect 2428 23366 2440 23418
rect 2492 23366 2504 23418
rect 2556 23366 4846 23418
rect 4898 23366 4910 23418
rect 4962 23366 4974 23418
rect 5026 23366 5038 23418
rect 5090 23366 5102 23418
rect 5154 23366 7443 23418
rect 7495 23366 7507 23418
rect 7559 23366 7571 23418
rect 7623 23366 7635 23418
rect 7687 23366 7699 23418
rect 7751 23366 8832 23418
rect 1104 23344 8832 23366
rect 5629 23239 5687 23245
rect 5629 23205 5641 23239
rect 5675 23236 5687 23239
rect 6730 23236 6736 23248
rect 5675 23208 6736 23236
rect 5675 23205 5687 23208
rect 5629 23199 5687 23205
rect 6730 23196 6736 23208
rect 6788 23236 6794 23248
rect 6788 23208 7696 23236
rect 6788 23196 6794 23208
rect 6089 23103 6147 23109
rect 6089 23069 6101 23103
rect 6135 23100 6147 23103
rect 6733 23103 6791 23109
rect 6733 23100 6745 23103
rect 6135 23072 6745 23100
rect 6135 23069 6147 23072
rect 6089 23063 6147 23069
rect 6733 23069 6745 23072
rect 6779 23100 6791 23103
rect 7558 23100 7564 23112
rect 6779 23072 7564 23100
rect 6779 23069 6791 23072
rect 6733 23063 6791 23069
rect 7558 23060 7564 23072
rect 7616 23060 7622 23112
rect 7668 23109 7696 23208
rect 7653 23103 7711 23109
rect 7653 23069 7665 23103
rect 7699 23069 7711 23103
rect 7653 23063 7711 23069
rect 6914 22992 6920 23044
rect 6972 23032 6978 23044
rect 6972 23004 7017 23032
rect 6972 22992 6978 23004
rect 6273 22967 6331 22973
rect 6273 22933 6285 22967
rect 6319 22964 6331 22967
rect 6822 22964 6828 22976
rect 6319 22936 6828 22964
rect 6319 22933 6331 22936
rect 6273 22927 6331 22933
rect 6822 22924 6828 22936
rect 6880 22924 6886 22976
rect 1104 22874 8832 22896
rect 1104 22822 3547 22874
rect 3599 22822 3611 22874
rect 3663 22822 3675 22874
rect 3727 22822 3739 22874
rect 3791 22822 3803 22874
rect 3855 22822 6144 22874
rect 6196 22822 6208 22874
rect 6260 22822 6272 22874
rect 6324 22822 6336 22874
rect 6388 22822 6400 22874
rect 6452 22822 8832 22874
rect 1104 22800 8832 22822
rect 6822 22692 6828 22704
rect 6783 22664 6828 22692
rect 6822 22652 6828 22664
rect 6880 22652 6886 22704
rect 6914 22652 6920 22704
rect 6972 22692 6978 22704
rect 6972 22664 7017 22692
rect 6972 22652 6978 22664
rect 7558 22652 7564 22704
rect 7616 22692 7622 22704
rect 7834 22692 7840 22704
rect 7616 22664 7840 22692
rect 7616 22652 7622 22664
rect 7834 22652 7840 22664
rect 7892 22652 7898 22704
rect 8018 22692 8024 22704
rect 7979 22664 8024 22692
rect 8018 22652 8024 22664
rect 8076 22652 8082 22704
rect 5813 22627 5871 22633
rect 5813 22593 5825 22627
rect 5859 22624 5871 22627
rect 6932 22624 6960 22652
rect 5859 22596 6960 22624
rect 5859 22593 5871 22596
rect 5813 22587 5871 22593
rect 5169 22559 5227 22565
rect 5169 22525 5181 22559
rect 5215 22556 5227 22559
rect 6730 22556 6736 22568
rect 5215 22528 6736 22556
rect 5215 22525 5227 22528
rect 5169 22519 5227 22525
rect 6730 22516 6736 22528
rect 6788 22556 6794 22568
rect 7377 22559 7435 22565
rect 7377 22556 7389 22559
rect 6788 22528 7389 22556
rect 6788 22516 6794 22528
rect 7377 22525 7389 22528
rect 7423 22525 7435 22559
rect 7377 22519 7435 22525
rect 5718 22420 5724 22432
rect 5679 22392 5724 22420
rect 5718 22380 5724 22392
rect 5776 22380 5782 22432
rect 1104 22330 8832 22352
rect 1104 22278 2248 22330
rect 2300 22278 2312 22330
rect 2364 22278 2376 22330
rect 2428 22278 2440 22330
rect 2492 22278 2504 22330
rect 2556 22278 4846 22330
rect 4898 22278 4910 22330
rect 4962 22278 4974 22330
rect 5026 22278 5038 22330
rect 5090 22278 5102 22330
rect 5154 22278 7443 22330
rect 7495 22278 7507 22330
rect 7559 22278 7571 22330
rect 7623 22278 7635 22330
rect 7687 22278 7699 22330
rect 7751 22278 8832 22330
rect 1104 22256 8832 22278
rect 6365 22015 6423 22021
rect 6365 22012 6377 22015
rect 6012 21984 6377 22012
rect 6012 21888 6040 21984
rect 6365 21981 6377 21984
rect 6411 21981 6423 22015
rect 7834 22012 7840 22024
rect 7795 21984 7840 22012
rect 6365 21975 6423 21981
rect 7834 21972 7840 21984
rect 7892 21972 7898 22024
rect 7926 21944 7932 21956
rect 7887 21916 7932 21944
rect 7926 21904 7932 21916
rect 7984 21904 7990 21956
rect 5353 21879 5411 21885
rect 5353 21845 5365 21879
rect 5399 21876 5411 21879
rect 5905 21879 5963 21885
rect 5905 21876 5917 21879
rect 5399 21848 5917 21876
rect 5399 21845 5411 21848
rect 5353 21839 5411 21845
rect 5905 21845 5917 21848
rect 5951 21876 5963 21879
rect 5994 21876 6000 21888
rect 5951 21848 6000 21876
rect 5951 21845 5963 21848
rect 5905 21839 5963 21845
rect 5994 21836 6000 21848
rect 6052 21836 6058 21888
rect 1104 21786 8832 21808
rect 1104 21734 3547 21786
rect 3599 21734 3611 21786
rect 3663 21734 3675 21786
rect 3727 21734 3739 21786
rect 3791 21734 3803 21786
rect 3855 21734 6144 21786
rect 6196 21734 6208 21786
rect 6260 21734 6272 21786
rect 6324 21734 6336 21786
rect 6388 21734 6400 21786
rect 6452 21734 8832 21786
rect 1104 21712 8832 21734
rect 5718 21564 5724 21616
rect 5776 21604 5782 21616
rect 6825 21607 6883 21613
rect 6825 21604 6837 21607
rect 5776 21576 6837 21604
rect 5776 21564 5782 21576
rect 6825 21573 6837 21576
rect 6871 21573 6883 21607
rect 6825 21567 6883 21573
rect 6917 21607 6975 21613
rect 6917 21573 6929 21607
rect 6963 21604 6975 21607
rect 7926 21604 7932 21616
rect 6963 21576 7932 21604
rect 6963 21573 6975 21576
rect 6917 21567 6975 21573
rect 7926 21564 7932 21576
rect 7984 21564 7990 21616
rect 5626 21536 5632 21548
rect 5587 21508 5632 21536
rect 5626 21496 5632 21508
rect 5684 21496 5690 21548
rect 5994 21428 6000 21480
rect 6052 21468 6058 21480
rect 7377 21471 7435 21477
rect 7377 21468 7389 21471
rect 6052 21440 7389 21468
rect 6052 21428 6058 21440
rect 7377 21437 7389 21440
rect 7423 21437 7435 21471
rect 7377 21431 7435 21437
rect 8110 21400 8116 21412
rect 8071 21372 8116 21400
rect 8110 21360 8116 21372
rect 8168 21360 8174 21412
rect 5166 21332 5172 21344
rect 5127 21304 5172 21332
rect 5166 21292 5172 21304
rect 5224 21292 5230 21344
rect 5721 21335 5779 21341
rect 5721 21301 5733 21335
rect 5767 21332 5779 21335
rect 6178 21332 6184 21344
rect 5767 21304 6184 21332
rect 5767 21301 5779 21304
rect 5721 21295 5779 21301
rect 6178 21292 6184 21304
rect 6236 21292 6242 21344
rect 1104 21242 8832 21264
rect 1104 21190 2248 21242
rect 2300 21190 2312 21242
rect 2364 21190 2376 21242
rect 2428 21190 2440 21242
rect 2492 21190 2504 21242
rect 2556 21190 4846 21242
rect 4898 21190 4910 21242
rect 4962 21190 4974 21242
rect 5026 21190 5038 21242
rect 5090 21190 5102 21242
rect 5154 21190 7443 21242
rect 7495 21190 7507 21242
rect 7559 21190 7571 21242
rect 7623 21190 7635 21242
rect 7687 21190 7699 21242
rect 7751 21190 8832 21242
rect 1104 21168 8832 21190
rect 6273 21063 6331 21069
rect 6273 21029 6285 21063
rect 6319 21060 6331 21063
rect 6546 21060 6552 21072
rect 6319 21032 6552 21060
rect 6319 21029 6331 21032
rect 6273 21023 6331 21029
rect 6546 21020 6552 21032
rect 6604 21020 6610 21072
rect 6178 20992 6184 21004
rect 6139 20964 6184 20992
rect 6178 20952 6184 20964
rect 6236 20952 6242 21004
rect 6380 20964 8156 20992
rect 5166 20924 5172 20936
rect 5079 20896 5172 20924
rect 5166 20884 5172 20896
rect 5224 20924 5230 20936
rect 6380 20924 6408 20964
rect 5224 20896 6408 20924
rect 5224 20884 5230 20896
rect 6638 20884 6644 20936
rect 6696 20924 6702 20936
rect 8128 20933 8156 20964
rect 6733 20927 6791 20933
rect 6733 20924 6745 20927
rect 6696 20896 6745 20924
rect 6696 20884 6702 20896
rect 6733 20893 6745 20896
rect 6779 20893 6791 20927
rect 6733 20887 6791 20893
rect 8113 20927 8171 20933
rect 8113 20893 8125 20927
rect 8159 20924 8171 20927
rect 8202 20924 8208 20936
rect 8159 20896 8208 20924
rect 8159 20893 8171 20896
rect 8113 20887 8171 20893
rect 8202 20884 8208 20896
rect 8260 20884 8266 20936
rect 5626 20856 5632 20868
rect 5539 20828 5632 20856
rect 5626 20816 5632 20828
rect 5684 20816 5690 20868
rect 5718 20816 5724 20868
rect 5776 20856 5782 20868
rect 7190 20856 7196 20868
rect 5776 20828 5821 20856
rect 7151 20828 7196 20856
rect 5776 20816 5782 20828
rect 7190 20816 7196 20828
rect 7248 20816 7254 20868
rect 7377 20859 7435 20865
rect 7377 20825 7389 20859
rect 7423 20825 7435 20859
rect 7377 20819 7435 20825
rect 4709 20791 4767 20797
rect 4709 20757 4721 20791
rect 4755 20788 4767 20791
rect 5258 20788 5264 20800
rect 4755 20760 5264 20788
rect 4755 20757 4767 20760
rect 4709 20751 4767 20757
rect 5258 20748 5264 20760
rect 5316 20748 5322 20800
rect 5644 20788 5672 20816
rect 7392 20788 7420 20819
rect 5644 20760 7420 20788
rect 1104 20698 8832 20720
rect 1104 20646 3547 20698
rect 3599 20646 3611 20698
rect 3663 20646 3675 20698
rect 3727 20646 3739 20698
rect 3791 20646 3803 20698
rect 3855 20646 6144 20698
rect 6196 20646 6208 20698
rect 6260 20646 6272 20698
rect 6324 20646 6336 20698
rect 6388 20646 6400 20698
rect 6452 20646 8832 20698
rect 1104 20624 8832 20646
rect 5166 20584 5172 20596
rect 5127 20556 5172 20584
rect 5166 20544 5172 20556
rect 5224 20544 5230 20596
rect 5629 20587 5687 20593
rect 5629 20553 5641 20587
rect 5675 20584 5687 20587
rect 5718 20584 5724 20596
rect 5675 20556 5724 20584
rect 5675 20553 5687 20556
rect 5629 20547 5687 20553
rect 5718 20544 5724 20556
rect 5776 20544 5782 20596
rect 6546 20516 6552 20528
rect 6507 20488 6552 20516
rect 6546 20476 6552 20488
rect 6604 20476 6610 20528
rect 6638 20476 6644 20528
rect 6696 20516 6702 20528
rect 6696 20488 8156 20516
rect 6696 20476 6702 20488
rect 5813 20451 5871 20457
rect 5813 20417 5825 20451
rect 5859 20448 5871 20451
rect 7190 20448 7196 20460
rect 5859 20420 7196 20448
rect 5859 20417 5871 20420
rect 5813 20411 5871 20417
rect 7190 20408 7196 20420
rect 7248 20448 7254 20460
rect 8018 20448 8024 20460
rect 7248 20420 8024 20448
rect 7248 20408 7254 20420
rect 8018 20408 8024 20420
rect 8076 20408 8082 20460
rect 8128 20457 8156 20488
rect 8113 20451 8171 20457
rect 8113 20417 8125 20451
rect 8159 20417 8171 20451
rect 8113 20411 8171 20417
rect 1104 20154 8832 20176
rect 1104 20102 2248 20154
rect 2300 20102 2312 20154
rect 2364 20102 2376 20154
rect 2428 20102 2440 20154
rect 2492 20102 2504 20154
rect 2556 20102 4846 20154
rect 4898 20102 4910 20154
rect 4962 20102 4974 20154
rect 5026 20102 5038 20154
rect 5090 20102 5102 20154
rect 5154 20102 7443 20154
rect 7495 20102 7507 20154
rect 7559 20102 7571 20154
rect 7623 20102 7635 20154
rect 7687 20102 7699 20154
rect 7751 20102 8832 20154
rect 1104 20080 8832 20102
rect 5534 20000 5540 20052
rect 5592 20040 5598 20052
rect 5997 20043 6055 20049
rect 5997 20040 6009 20043
rect 5592 20012 6009 20040
rect 5592 20000 5598 20012
rect 5997 20009 6009 20012
rect 6043 20009 6055 20043
rect 5997 20003 6055 20009
rect 6012 19836 6040 20003
rect 6549 19839 6607 19845
rect 6549 19836 6561 19839
rect 6012 19808 6561 19836
rect 6549 19805 6561 19808
rect 6595 19836 6607 19839
rect 6730 19836 6736 19848
rect 6595 19808 6736 19836
rect 6595 19805 6607 19808
rect 6549 19799 6607 19805
rect 6730 19796 6736 19808
rect 6788 19796 6794 19848
rect 7469 19839 7527 19845
rect 7469 19805 7481 19839
rect 7515 19836 7527 19839
rect 8110 19836 8116 19848
rect 7515 19808 8116 19836
rect 7515 19805 7527 19808
rect 7469 19799 7527 19805
rect 8110 19796 8116 19808
rect 8168 19796 8174 19848
rect 7190 19768 7196 19780
rect 7151 19740 7196 19768
rect 7190 19728 7196 19740
rect 7248 19728 7254 19780
rect 5258 19660 5264 19712
rect 5316 19700 5322 19712
rect 5537 19703 5595 19709
rect 5537 19700 5549 19703
rect 5316 19672 5549 19700
rect 5316 19660 5322 19672
rect 5537 19669 5549 19672
rect 5583 19700 5595 19703
rect 6638 19700 6644 19712
rect 5583 19672 6644 19700
rect 5583 19669 5595 19672
rect 5537 19663 5595 19669
rect 6638 19660 6644 19672
rect 6696 19660 6702 19712
rect 7282 19660 7288 19712
rect 7340 19700 7346 19712
rect 7929 19703 7987 19709
rect 7929 19700 7941 19703
rect 7340 19672 7941 19700
rect 7340 19660 7346 19672
rect 7929 19669 7941 19672
rect 7975 19669 7987 19703
rect 7929 19663 7987 19669
rect 1104 19610 8832 19632
rect 1104 19558 3547 19610
rect 3599 19558 3611 19610
rect 3663 19558 3675 19610
rect 3727 19558 3739 19610
rect 3791 19558 3803 19610
rect 3855 19558 6144 19610
rect 6196 19558 6208 19610
rect 6260 19558 6272 19610
rect 6324 19558 6336 19610
rect 6388 19558 6400 19610
rect 6452 19558 8832 19610
rect 1104 19536 8832 19558
rect 8018 19496 8024 19508
rect 7979 19468 8024 19496
rect 8018 19456 8024 19468
rect 8076 19456 8082 19508
rect 7190 19428 7196 19440
rect 7151 19400 7196 19428
rect 7190 19388 7196 19400
rect 7248 19388 7254 19440
rect 7282 19388 7288 19440
rect 7340 19428 7346 19440
rect 7340 19400 7385 19428
rect 7340 19388 7346 19400
rect 6546 19320 6552 19372
rect 6604 19360 6610 19372
rect 7929 19363 7987 19369
rect 7929 19360 7941 19363
rect 6604 19332 7941 19360
rect 6604 19320 6610 19332
rect 7929 19329 7941 19332
rect 7975 19329 7987 19363
rect 7929 19323 7987 19329
rect 6730 19292 6736 19304
rect 6691 19264 6736 19292
rect 6730 19252 6736 19264
rect 6788 19252 6794 19304
rect 5626 19116 5632 19168
rect 5684 19156 5690 19168
rect 6822 19156 6828 19168
rect 5684 19128 6828 19156
rect 5684 19116 5690 19128
rect 6822 19116 6828 19128
rect 6880 19116 6886 19168
rect 1104 19066 8832 19088
rect 1104 19014 2248 19066
rect 2300 19014 2312 19066
rect 2364 19014 2376 19066
rect 2428 19014 2440 19066
rect 2492 19014 2504 19066
rect 2556 19014 4846 19066
rect 4898 19014 4910 19066
rect 4962 19014 4974 19066
rect 5026 19014 5038 19066
rect 5090 19014 5102 19066
rect 5154 19014 7443 19066
rect 7495 19014 7507 19066
rect 7559 19014 7571 19066
rect 7623 19014 7635 19066
rect 7687 19014 7699 19066
rect 7751 19014 8832 19066
rect 1104 18992 8832 19014
rect 6730 18952 6736 18964
rect 6691 18924 6736 18952
rect 6730 18912 6736 18924
rect 6788 18912 6794 18964
rect 7190 18748 7196 18760
rect 7151 18720 7196 18748
rect 7190 18708 7196 18720
rect 7248 18708 7254 18760
rect 6730 18640 6736 18692
rect 6788 18680 6794 18692
rect 7837 18683 7895 18689
rect 7837 18680 7849 18683
rect 6788 18652 7849 18680
rect 6788 18640 6794 18652
rect 7837 18649 7849 18652
rect 7883 18649 7895 18683
rect 7837 18643 7895 18649
rect 7282 18612 7288 18624
rect 7243 18584 7288 18612
rect 7282 18572 7288 18584
rect 7340 18572 7346 18624
rect 1104 18522 8832 18544
rect 1104 18470 3547 18522
rect 3599 18470 3611 18522
rect 3663 18470 3675 18522
rect 3727 18470 3739 18522
rect 3791 18470 3803 18522
rect 3855 18470 6144 18522
rect 6196 18470 6208 18522
rect 6260 18470 6272 18522
rect 6324 18470 6336 18522
rect 6388 18470 6400 18522
rect 6452 18470 8832 18522
rect 1104 18448 8832 18470
rect 5718 18232 5724 18284
rect 5776 18272 5782 18284
rect 6365 18275 6423 18281
rect 6365 18272 6377 18275
rect 5776 18244 6377 18272
rect 5776 18232 5782 18244
rect 6365 18241 6377 18244
rect 6411 18272 6423 18275
rect 6730 18272 6736 18284
rect 6411 18244 6736 18272
rect 6411 18241 6423 18244
rect 6365 18235 6423 18241
rect 6730 18232 6736 18244
rect 6788 18232 6794 18284
rect 7837 18275 7895 18281
rect 7837 18241 7849 18275
rect 7883 18272 7895 18275
rect 8110 18272 8116 18284
rect 7883 18244 8116 18272
rect 7883 18241 7895 18244
rect 7837 18235 7895 18241
rect 8110 18232 8116 18244
rect 8168 18232 8174 18284
rect 7834 18136 7840 18148
rect 7795 18108 7840 18136
rect 7834 18096 7840 18108
rect 7892 18096 7898 18148
rect 5718 18068 5724 18080
rect 5679 18040 5724 18068
rect 5718 18028 5724 18040
rect 5776 18028 5782 18080
rect 1104 17978 8832 18000
rect 1104 17926 2248 17978
rect 2300 17926 2312 17978
rect 2364 17926 2376 17978
rect 2428 17926 2440 17978
rect 2492 17926 2504 17978
rect 2556 17926 4846 17978
rect 4898 17926 4910 17978
rect 4962 17926 4974 17978
rect 5026 17926 5038 17978
rect 5090 17926 5102 17978
rect 5154 17926 7443 17978
rect 7495 17926 7507 17978
rect 7559 17926 7571 17978
rect 7623 17926 7635 17978
rect 7687 17926 7699 17978
rect 7751 17926 8832 17978
rect 1104 17904 8832 17926
rect 5353 17731 5411 17737
rect 5353 17697 5365 17731
rect 5399 17728 5411 17731
rect 5534 17728 5540 17740
rect 5399 17700 5540 17728
rect 5399 17697 5411 17700
rect 5353 17691 5411 17697
rect 5534 17688 5540 17700
rect 5592 17728 5598 17740
rect 5810 17728 5816 17740
rect 5592 17700 5816 17728
rect 5592 17688 5598 17700
rect 5810 17688 5816 17700
rect 5868 17688 5874 17740
rect 6273 17731 6331 17737
rect 6273 17697 6285 17731
rect 6319 17728 6331 17731
rect 7098 17728 7104 17740
rect 6319 17700 7104 17728
rect 6319 17697 6331 17700
rect 6273 17691 6331 17697
rect 7098 17688 7104 17700
rect 7156 17688 7162 17740
rect 7282 17688 7288 17740
rect 7340 17728 7346 17740
rect 7377 17731 7435 17737
rect 7377 17728 7389 17731
rect 7340 17700 7389 17728
rect 7340 17688 7346 17700
rect 7377 17697 7389 17700
rect 7423 17697 7435 17731
rect 7377 17691 7435 17697
rect 6825 17663 6883 17669
rect 6825 17660 6837 17663
rect 6288 17632 6837 17660
rect 5718 17552 5724 17604
rect 5776 17592 5782 17604
rect 6288 17592 6316 17632
rect 6825 17629 6837 17632
rect 6871 17629 6883 17663
rect 6825 17623 6883 17629
rect 7190 17620 7196 17672
rect 7248 17660 7254 17672
rect 8113 17663 8171 17669
rect 8113 17660 8125 17663
rect 7248 17632 8125 17660
rect 7248 17620 7254 17632
rect 8113 17629 8125 17632
rect 8159 17629 8171 17663
rect 8113 17623 8171 17629
rect 5776 17564 6316 17592
rect 6365 17595 6423 17601
rect 5776 17552 5782 17564
rect 6365 17561 6377 17595
rect 6411 17561 6423 17595
rect 6365 17555 6423 17561
rect 6380 17524 6408 17555
rect 6914 17552 6920 17604
rect 6972 17592 6978 17604
rect 7285 17595 7343 17601
rect 7285 17592 7297 17595
rect 6972 17564 7297 17592
rect 6972 17552 6978 17564
rect 7285 17561 7297 17564
rect 7331 17592 7343 17595
rect 7834 17592 7840 17604
rect 7331 17564 7840 17592
rect 7331 17561 7343 17564
rect 7285 17555 7343 17561
rect 7834 17552 7840 17564
rect 7892 17552 7898 17604
rect 7929 17527 7987 17533
rect 7929 17524 7941 17527
rect 6380 17496 7941 17524
rect 7929 17493 7941 17496
rect 7975 17493 7987 17527
rect 7929 17487 7987 17493
rect 1104 17434 8832 17456
rect 1104 17382 3547 17434
rect 3599 17382 3611 17434
rect 3663 17382 3675 17434
rect 3727 17382 3739 17434
rect 3791 17382 3803 17434
rect 3855 17382 6144 17434
rect 6196 17382 6208 17434
rect 6260 17382 6272 17434
rect 6324 17382 6336 17434
rect 6388 17382 6400 17434
rect 6452 17382 8832 17434
rect 1104 17360 8832 17382
rect 5902 17280 5908 17332
rect 5960 17320 5966 17332
rect 6638 17320 6644 17332
rect 5960 17292 6644 17320
rect 5960 17280 5966 17292
rect 6638 17280 6644 17292
rect 6696 17280 6702 17332
rect 6546 17252 6552 17264
rect 6507 17224 6552 17252
rect 6546 17212 6552 17224
rect 6604 17212 6610 17264
rect 7190 17184 7196 17196
rect 7151 17156 7196 17184
rect 7190 17144 7196 17156
rect 7248 17144 7254 17196
rect 8113 17187 8171 17193
rect 8113 17153 8125 17187
rect 8159 17153 8171 17187
rect 8113 17147 8171 17153
rect 8128 17116 8156 17147
rect 5828 17088 8156 17116
rect 5828 16992 5856 17088
rect 5810 16980 5816 16992
rect 5771 16952 5816 16980
rect 5810 16940 5816 16952
rect 5868 16940 5874 16992
rect 1104 16890 8832 16912
rect 1104 16838 2248 16890
rect 2300 16838 2312 16890
rect 2364 16838 2376 16890
rect 2428 16838 2440 16890
rect 2492 16838 2504 16890
rect 2556 16838 4846 16890
rect 4898 16838 4910 16890
rect 4962 16838 4974 16890
rect 5026 16838 5038 16890
rect 5090 16838 5102 16890
rect 5154 16838 7443 16890
rect 7495 16838 7507 16890
rect 7559 16838 7571 16890
rect 7623 16838 7635 16890
rect 7687 16838 7699 16890
rect 7751 16838 8832 16890
rect 1104 16816 8832 16838
rect 5169 16779 5227 16785
rect 5169 16745 5181 16779
rect 5215 16776 5227 16779
rect 5534 16776 5540 16788
rect 5215 16748 5540 16776
rect 5215 16745 5227 16748
rect 5169 16739 5227 16745
rect 5534 16736 5540 16748
rect 5592 16776 5598 16788
rect 5592 16748 6914 16776
rect 5592 16736 5598 16748
rect 6546 16668 6552 16720
rect 6604 16708 6610 16720
rect 6641 16711 6699 16717
rect 6641 16708 6653 16711
rect 6604 16680 6653 16708
rect 6604 16668 6610 16680
rect 6641 16677 6653 16680
rect 6687 16677 6699 16711
rect 6641 16671 6699 16677
rect 5721 16643 5779 16649
rect 5721 16609 5733 16643
rect 5767 16640 5779 16643
rect 5810 16640 5816 16652
rect 5767 16612 5816 16640
rect 5767 16609 5779 16612
rect 5721 16603 5779 16609
rect 5810 16600 5816 16612
rect 5868 16640 5874 16652
rect 6181 16643 6239 16649
rect 6181 16640 6193 16643
rect 5868 16612 6193 16640
rect 5868 16600 5874 16612
rect 6181 16609 6193 16612
rect 6227 16640 6239 16643
rect 6886 16640 6914 16748
rect 6227 16612 6592 16640
rect 6886 16612 7512 16640
rect 6227 16609 6239 16612
rect 6181 16603 6239 16609
rect 6564 16448 6592 16612
rect 7098 16532 7104 16584
rect 7156 16572 7162 16584
rect 7377 16575 7435 16581
rect 7377 16572 7389 16575
rect 7156 16544 7389 16572
rect 7156 16532 7162 16544
rect 7377 16541 7389 16544
rect 7423 16541 7435 16575
rect 7484 16572 7512 16612
rect 8113 16575 8171 16581
rect 8113 16572 8125 16575
rect 7484 16544 8125 16572
rect 7377 16535 7435 16541
rect 8113 16541 8125 16544
rect 8159 16541 8171 16575
rect 8113 16535 8171 16541
rect 6730 16464 6736 16516
rect 6788 16504 6794 16516
rect 7190 16504 7196 16516
rect 6788 16476 6833 16504
rect 7151 16476 7196 16504
rect 6788 16464 6794 16476
rect 7190 16464 7196 16476
rect 7248 16464 7254 16516
rect 6546 16396 6552 16448
rect 6604 16396 6610 16448
rect 1104 16346 8832 16368
rect 1104 16294 3547 16346
rect 3599 16294 3611 16346
rect 3663 16294 3675 16346
rect 3727 16294 3739 16346
rect 3791 16294 3803 16346
rect 3855 16294 6144 16346
rect 6196 16294 6208 16346
rect 6260 16294 6272 16346
rect 6324 16294 6336 16346
rect 6388 16294 6400 16346
rect 6452 16294 8832 16346
rect 1104 16272 8832 16294
rect 6730 16192 6736 16244
rect 6788 16232 6794 16244
rect 8021 16235 8079 16241
rect 8021 16232 8033 16235
rect 6788 16204 8033 16232
rect 6788 16192 6794 16204
rect 8021 16201 8033 16204
rect 8067 16201 8079 16235
rect 8021 16195 8079 16201
rect 6549 16167 6607 16173
rect 6549 16133 6561 16167
rect 6595 16164 6607 16167
rect 6914 16164 6920 16176
rect 6595 16136 6920 16164
rect 6595 16133 6607 16136
rect 6549 16127 6607 16133
rect 5629 16099 5687 16105
rect 5629 16065 5641 16099
rect 5675 16096 5687 16099
rect 6564 16096 6592 16127
rect 6914 16124 6920 16136
rect 6972 16124 6978 16176
rect 7098 16124 7104 16176
rect 7156 16164 7162 16176
rect 7929 16167 7987 16173
rect 7929 16164 7941 16167
rect 7156 16136 7941 16164
rect 7156 16124 7162 16136
rect 7929 16133 7941 16136
rect 7975 16133 7987 16167
rect 7929 16127 7987 16133
rect 6730 16096 6736 16108
rect 5675 16068 6592 16096
rect 6691 16068 6736 16096
rect 5675 16065 5687 16068
rect 5629 16059 5687 16065
rect 6730 16056 6736 16068
rect 6788 16056 6794 16108
rect 7006 16056 7012 16108
rect 7064 16096 7070 16108
rect 7469 16099 7527 16105
rect 7469 16096 7481 16099
rect 7064 16068 7481 16096
rect 7064 16056 7070 16068
rect 7469 16065 7481 16068
rect 7515 16096 7527 16099
rect 7834 16096 7840 16108
rect 7515 16068 7840 16096
rect 7515 16065 7527 16068
rect 7469 16059 7527 16065
rect 7834 16056 7840 16068
rect 7892 16056 7898 16108
rect 5166 16028 5172 16040
rect 5079 16000 5172 16028
rect 5166 15988 5172 16000
rect 5224 16028 5230 16040
rect 7024 16028 7052 16056
rect 5224 16000 7052 16028
rect 5224 15988 5230 16000
rect 5813 15895 5871 15901
rect 5813 15861 5825 15895
rect 5859 15892 5871 15895
rect 6454 15892 6460 15904
rect 5859 15864 6460 15892
rect 5859 15861 5871 15864
rect 5813 15855 5871 15861
rect 6454 15852 6460 15864
rect 6512 15852 6518 15904
rect 1104 15802 8832 15824
rect 1104 15750 2248 15802
rect 2300 15750 2312 15802
rect 2364 15750 2376 15802
rect 2428 15750 2440 15802
rect 2492 15750 2504 15802
rect 2556 15750 4846 15802
rect 4898 15750 4910 15802
rect 4962 15750 4974 15802
rect 5026 15750 5038 15802
rect 5090 15750 5102 15802
rect 5154 15750 7443 15802
rect 7495 15750 7507 15802
rect 7559 15750 7571 15802
rect 7623 15750 7635 15802
rect 7687 15750 7699 15802
rect 7751 15750 8832 15802
rect 1104 15728 8832 15750
rect 4801 15691 4859 15697
rect 4801 15657 4813 15691
rect 4847 15688 4859 15691
rect 5166 15688 5172 15700
rect 4847 15660 5172 15688
rect 4847 15657 4859 15660
rect 4801 15651 4859 15657
rect 5166 15648 5172 15660
rect 5224 15648 5230 15700
rect 5350 15648 5356 15700
rect 5408 15688 5414 15700
rect 5408 15660 8064 15688
rect 5408 15648 5414 15660
rect 6549 15623 6607 15629
rect 6549 15589 6561 15623
rect 6595 15620 6607 15623
rect 6730 15620 6736 15632
rect 6595 15592 6736 15620
rect 6595 15589 6607 15592
rect 6549 15583 6607 15589
rect 5350 15552 5356 15564
rect 5311 15524 5356 15552
rect 5350 15512 5356 15524
rect 5408 15512 5414 15564
rect 6454 15552 6460 15564
rect 6415 15524 6460 15552
rect 6454 15512 6460 15524
rect 6512 15512 6518 15564
rect 5997 15487 6055 15493
rect 5997 15453 6009 15487
rect 6043 15484 6055 15487
rect 6564 15484 6592 15583
rect 6730 15580 6736 15592
rect 6788 15580 6794 15632
rect 7006 15552 7012 15564
rect 6967 15524 7012 15552
rect 7006 15512 7012 15524
rect 7064 15512 7070 15564
rect 8036 15561 8064 15660
rect 8021 15555 8079 15561
rect 8021 15521 8033 15555
rect 8067 15552 8079 15555
rect 8110 15552 8116 15564
rect 8067 15524 8116 15552
rect 8067 15521 8079 15524
rect 8021 15515 8079 15521
rect 8110 15512 8116 15524
rect 8168 15512 8174 15564
rect 6043 15456 6592 15484
rect 6043 15453 6055 15456
rect 5997 15447 6055 15453
rect 7282 15444 7288 15496
rect 7340 15484 7346 15496
rect 7561 15487 7619 15493
rect 7561 15484 7573 15487
rect 7340 15456 7573 15484
rect 7340 15444 7346 15456
rect 7561 15453 7573 15456
rect 7607 15453 7619 15487
rect 7561 15447 7619 15453
rect 5810 15416 5816 15428
rect 5771 15388 5816 15416
rect 5810 15376 5816 15388
rect 5868 15376 5874 15428
rect 7098 15376 7104 15428
rect 7156 15416 7162 15428
rect 7469 15419 7527 15425
rect 7469 15416 7481 15419
rect 7156 15388 7481 15416
rect 7156 15376 7162 15388
rect 7469 15385 7481 15388
rect 7515 15385 7527 15419
rect 7469 15379 7527 15385
rect 1104 15258 8832 15280
rect 1104 15206 3547 15258
rect 3599 15206 3611 15258
rect 3663 15206 3675 15258
rect 3727 15206 3739 15258
rect 3791 15206 3803 15258
rect 3855 15206 6144 15258
rect 6196 15206 6208 15258
rect 6260 15206 6272 15258
rect 6324 15206 6336 15258
rect 6388 15206 6400 15258
rect 6452 15206 8832 15258
rect 1104 15184 8832 15206
rect 5077 15147 5135 15153
rect 5077 15113 5089 15147
rect 5123 15144 5135 15147
rect 5350 15144 5356 15156
rect 5123 15116 5356 15144
rect 5123 15113 5135 15116
rect 5077 15107 5135 15113
rect 5350 15104 5356 15116
rect 5408 15104 5414 15156
rect 5721 15147 5779 15153
rect 5721 15113 5733 15147
rect 5767 15144 5779 15147
rect 7190 15144 7196 15156
rect 5767 15116 7196 15144
rect 5767 15113 5779 15116
rect 5721 15107 5779 15113
rect 7190 15104 7196 15116
rect 7248 15104 7254 15156
rect 5629 15079 5687 15085
rect 5629 15045 5641 15079
rect 5675 15076 5687 15079
rect 7834 15076 7840 15088
rect 5675 15048 7840 15076
rect 5675 15045 5687 15048
rect 5629 15039 5687 15045
rect 7834 15036 7840 15048
rect 7892 15036 7898 15088
rect 6549 15011 6607 15017
rect 6549 14977 6561 15011
rect 6595 14977 6607 15011
rect 6730 15008 6736 15020
rect 6691 14980 6736 15008
rect 6549 14971 6607 14977
rect 6564 14884 6592 14971
rect 6730 14968 6736 14980
rect 6788 14968 6794 15020
rect 7006 14968 7012 15020
rect 7064 15008 7070 15020
rect 7193 15011 7251 15017
rect 7193 15008 7205 15011
rect 7064 14980 7205 15008
rect 7064 14968 7070 14980
rect 7193 14977 7205 14980
rect 7239 14977 7251 15011
rect 7193 14971 7251 14977
rect 7282 14968 7288 15020
rect 7340 15008 7346 15020
rect 7377 15011 7435 15017
rect 7377 15008 7389 15011
rect 7340 14980 7389 15008
rect 7340 14968 7346 14980
rect 7377 14977 7389 14980
rect 7423 14977 7435 15011
rect 8110 15008 8116 15020
rect 8071 14980 8116 15008
rect 7377 14971 7435 14977
rect 8110 14968 8116 14980
rect 8168 14968 8174 15020
rect 4525 14875 4583 14881
rect 4525 14841 4537 14875
rect 4571 14872 4583 14875
rect 5534 14872 5540 14884
rect 4571 14844 5540 14872
rect 4571 14841 4583 14844
rect 4525 14835 4583 14841
rect 5534 14832 5540 14844
rect 5592 14832 5598 14884
rect 6546 14832 6552 14884
rect 6604 14832 6610 14884
rect 6086 14764 6092 14816
rect 6144 14804 6150 14816
rect 6457 14807 6515 14813
rect 6457 14804 6469 14807
rect 6144 14776 6469 14804
rect 6144 14764 6150 14776
rect 6457 14773 6469 14776
rect 6503 14773 6515 14807
rect 6457 14767 6515 14773
rect 1104 14714 8832 14736
rect 1104 14662 2248 14714
rect 2300 14662 2312 14714
rect 2364 14662 2376 14714
rect 2428 14662 2440 14714
rect 2492 14662 2504 14714
rect 2556 14662 4846 14714
rect 4898 14662 4910 14714
rect 4962 14662 4974 14714
rect 5026 14662 5038 14714
rect 5090 14662 5102 14714
rect 5154 14662 7443 14714
rect 7495 14662 7507 14714
rect 7559 14662 7571 14714
rect 7623 14662 7635 14714
rect 7687 14662 7699 14714
rect 7751 14662 8832 14714
rect 1104 14640 8832 14662
rect 5537 14535 5595 14541
rect 5537 14501 5549 14535
rect 5583 14532 5595 14535
rect 7190 14532 7196 14544
rect 5583 14504 7196 14532
rect 5583 14501 5595 14504
rect 5537 14495 5595 14501
rect 7190 14492 7196 14504
rect 7248 14532 7254 14544
rect 7377 14535 7435 14541
rect 7377 14532 7389 14535
rect 7248 14504 7389 14532
rect 7248 14492 7254 14504
rect 7377 14501 7389 14504
rect 7423 14501 7435 14535
rect 7377 14495 7435 14501
rect 5629 14467 5687 14473
rect 5629 14433 5641 14467
rect 5675 14464 5687 14467
rect 5810 14464 5816 14476
rect 5675 14436 5816 14464
rect 5675 14433 5687 14436
rect 5629 14427 5687 14433
rect 5810 14424 5816 14436
rect 5868 14424 5874 14476
rect 6730 14464 6736 14476
rect 5920 14436 6736 14464
rect 5077 14399 5135 14405
rect 5077 14365 5089 14399
rect 5123 14396 5135 14399
rect 5534 14396 5540 14408
rect 5123 14368 5540 14396
rect 5123 14365 5135 14368
rect 5077 14359 5135 14365
rect 5534 14356 5540 14368
rect 5592 14396 5598 14408
rect 5920 14396 5948 14436
rect 6730 14424 6736 14436
rect 6788 14424 6794 14476
rect 6086 14396 6092 14408
rect 5592 14368 5948 14396
rect 6047 14368 6092 14396
rect 5592 14356 5598 14368
rect 6086 14356 6092 14368
rect 6144 14356 6150 14408
rect 6914 14356 6920 14408
rect 6972 14396 6978 14408
rect 7009 14399 7067 14405
rect 7009 14396 7021 14399
rect 6972 14368 7021 14396
rect 6972 14356 6978 14368
rect 7009 14365 7021 14368
rect 7055 14365 7067 14399
rect 7009 14359 7067 14365
rect 6454 14288 6460 14340
rect 6512 14328 6518 14340
rect 6730 14328 6736 14340
rect 6512 14300 6736 14328
rect 6512 14288 6518 14300
rect 6730 14288 6736 14300
rect 6788 14288 6794 14340
rect 1104 14170 8832 14192
rect 1104 14118 3547 14170
rect 3599 14118 3611 14170
rect 3663 14118 3675 14170
rect 3727 14118 3739 14170
rect 3791 14118 3803 14170
rect 3855 14118 6144 14170
rect 6196 14118 6208 14170
rect 6260 14118 6272 14170
rect 6324 14118 6336 14170
rect 6388 14118 6400 14170
rect 6452 14118 8832 14170
rect 1104 14096 8832 14118
rect 5994 13880 6000 13932
rect 6052 13920 6058 13932
rect 6549 13923 6607 13929
rect 6549 13920 6561 13923
rect 6052 13892 6561 13920
rect 6052 13880 6058 13892
rect 6549 13889 6561 13892
rect 6595 13889 6607 13923
rect 6549 13883 6607 13889
rect 7006 13880 7012 13932
rect 7064 13920 7070 13932
rect 7469 13923 7527 13929
rect 7469 13920 7481 13923
rect 7064 13892 7481 13920
rect 7064 13880 7070 13892
rect 7469 13889 7481 13892
rect 7515 13889 7527 13923
rect 7469 13883 7527 13889
rect 7834 13784 7840 13796
rect 7795 13756 7840 13784
rect 7834 13744 7840 13756
rect 7892 13744 7898 13796
rect 5813 13719 5871 13725
rect 5813 13685 5825 13719
rect 5859 13716 5871 13719
rect 5994 13716 6000 13728
rect 5859 13688 6000 13716
rect 5859 13685 5871 13688
rect 5813 13679 5871 13685
rect 5994 13676 6000 13688
rect 6052 13676 6058 13728
rect 1104 13626 8832 13648
rect 1104 13574 2248 13626
rect 2300 13574 2312 13626
rect 2364 13574 2376 13626
rect 2428 13574 2440 13626
rect 2492 13574 2504 13626
rect 2556 13574 4846 13626
rect 4898 13574 4910 13626
rect 4962 13574 4974 13626
rect 5026 13574 5038 13626
rect 5090 13574 5102 13626
rect 5154 13574 7443 13626
rect 7495 13574 7507 13626
rect 7559 13574 7571 13626
rect 7623 13574 7635 13626
rect 7687 13574 7699 13626
rect 7751 13574 8832 13626
rect 1104 13552 8832 13574
rect 5534 13472 5540 13524
rect 5592 13512 5598 13524
rect 5721 13515 5779 13521
rect 5721 13512 5733 13515
rect 5592 13484 5733 13512
rect 5592 13472 5598 13484
rect 5721 13481 5733 13484
rect 5767 13481 5779 13515
rect 7098 13512 7104 13524
rect 7059 13484 7104 13512
rect 5721 13475 5779 13481
rect 7098 13472 7104 13484
rect 7156 13472 7162 13524
rect 7653 13447 7711 13453
rect 7653 13413 7665 13447
rect 7699 13444 7711 13447
rect 7834 13444 7840 13456
rect 7699 13416 7840 13444
rect 7699 13413 7711 13416
rect 7653 13407 7711 13413
rect 7834 13404 7840 13416
rect 7892 13404 7898 13456
rect 6917 13311 6975 13317
rect 6917 13277 6929 13311
rect 6963 13308 6975 13311
rect 7006 13308 7012 13320
rect 6963 13280 7012 13308
rect 6963 13277 6975 13280
rect 6917 13271 6975 13277
rect 7006 13268 7012 13280
rect 7064 13268 7070 13320
rect 8113 13311 8171 13317
rect 8113 13277 8125 13311
rect 8159 13277 8171 13311
rect 8113 13271 8171 13277
rect 7282 13200 7288 13252
rect 7340 13240 7346 13252
rect 7561 13243 7619 13249
rect 7561 13240 7573 13243
rect 7340 13212 7573 13240
rect 7340 13200 7346 13212
rect 7561 13209 7573 13212
rect 7607 13209 7619 13243
rect 7561 13203 7619 13209
rect 5994 13132 6000 13184
rect 6052 13172 6058 13184
rect 6365 13175 6423 13181
rect 6365 13172 6377 13175
rect 6052 13144 6377 13172
rect 6052 13132 6058 13144
rect 6365 13141 6377 13144
rect 6411 13172 6423 13175
rect 8128 13172 8156 13271
rect 6411 13144 8156 13172
rect 6411 13141 6423 13144
rect 6365 13135 6423 13141
rect 1104 13082 8832 13104
rect 1104 13030 3547 13082
rect 3599 13030 3611 13082
rect 3663 13030 3675 13082
rect 3727 13030 3739 13082
rect 3791 13030 3803 13082
rect 3855 13030 6144 13082
rect 6196 13030 6208 13082
rect 6260 13030 6272 13082
rect 6324 13030 6336 13082
rect 6388 13030 6400 13082
rect 6452 13030 8832 13082
rect 1104 13008 8832 13030
rect 6822 12928 6828 12980
rect 6880 12928 6886 12980
rect 7282 12968 7288 12980
rect 7243 12940 7288 12968
rect 7282 12928 7288 12940
rect 7340 12928 7346 12980
rect 7374 12928 7380 12980
rect 7432 12968 7438 12980
rect 7432 12940 7477 12968
rect 7432 12928 7438 12940
rect 6840 12900 6868 12928
rect 8202 12900 8208 12912
rect 6840 12872 8208 12900
rect 8202 12860 8208 12872
rect 8260 12860 8266 12912
rect 5534 12792 5540 12844
rect 5592 12832 5598 12844
rect 6178 12832 6184 12844
rect 5592 12804 6184 12832
rect 5592 12792 5598 12804
rect 6178 12792 6184 12804
rect 6236 12792 6242 12844
rect 7190 12792 7196 12844
rect 7248 12832 7254 12844
rect 8021 12835 8079 12841
rect 8021 12832 8033 12835
rect 7248 12804 8033 12832
rect 7248 12792 7254 12804
rect 8021 12801 8033 12804
rect 8067 12801 8079 12835
rect 8021 12795 8079 12801
rect 6730 12764 6736 12776
rect 6691 12736 6736 12764
rect 6730 12724 6736 12736
rect 6788 12724 6794 12776
rect 7834 12628 7840 12640
rect 7795 12600 7840 12628
rect 7834 12588 7840 12600
rect 7892 12588 7898 12640
rect 1104 12538 8832 12560
rect 1104 12486 2248 12538
rect 2300 12486 2312 12538
rect 2364 12486 2376 12538
rect 2428 12486 2440 12538
rect 2492 12486 2504 12538
rect 2556 12486 4846 12538
rect 4898 12486 4910 12538
rect 4962 12486 4974 12538
rect 5026 12486 5038 12538
rect 5090 12486 5102 12538
rect 5154 12486 7443 12538
rect 7495 12486 7507 12538
rect 7559 12486 7571 12538
rect 7623 12486 7635 12538
rect 7687 12486 7699 12538
rect 7751 12486 8832 12538
rect 1104 12464 8832 12486
rect 5258 12384 5264 12436
rect 5316 12424 5322 12436
rect 5718 12424 5724 12436
rect 5316 12396 5724 12424
rect 5316 12384 5322 12396
rect 5718 12384 5724 12396
rect 5776 12384 5782 12436
rect 6730 12356 6736 12368
rect 6691 12328 6736 12356
rect 6730 12316 6736 12328
rect 6788 12316 6794 12368
rect 6546 12248 6552 12300
rect 6604 12248 6610 12300
rect 7745 12291 7803 12297
rect 7745 12257 7757 12291
rect 7791 12288 7803 12291
rect 7834 12288 7840 12300
rect 7791 12260 7840 12288
rect 7791 12257 7803 12260
rect 7745 12251 7803 12257
rect 7834 12248 7840 12260
rect 7892 12248 7898 12300
rect 5534 12180 5540 12232
rect 5592 12220 5598 12232
rect 5810 12220 5816 12232
rect 5592 12192 5816 12220
rect 5592 12180 5598 12192
rect 5810 12180 5816 12192
rect 5868 12180 5874 12232
rect 5902 12180 5908 12232
rect 5960 12220 5966 12232
rect 6365 12223 6423 12229
rect 6365 12220 6377 12223
rect 5960 12192 6377 12220
rect 5960 12180 5966 12192
rect 6365 12189 6377 12192
rect 6411 12220 6423 12223
rect 6564 12220 6592 12248
rect 6411 12192 6592 12220
rect 7193 12223 7251 12229
rect 6411 12189 6423 12192
rect 6365 12183 6423 12189
rect 7193 12189 7205 12223
rect 7239 12189 7251 12223
rect 7193 12183 7251 12189
rect 6178 12152 6184 12164
rect 5828 12124 6184 12152
rect 5828 12096 5856 12124
rect 6178 12112 6184 12124
rect 6236 12152 6242 12164
rect 7208 12152 7236 12183
rect 6236 12124 7236 12152
rect 6236 12112 6242 12124
rect 7282 12112 7288 12164
rect 7340 12152 7346 12164
rect 7653 12155 7711 12161
rect 7653 12152 7665 12155
rect 7340 12124 7665 12152
rect 7340 12112 7346 12124
rect 7653 12121 7665 12124
rect 7699 12121 7711 12155
rect 7653 12115 7711 12121
rect 5810 12084 5816 12096
rect 5771 12056 5816 12084
rect 5810 12044 5816 12056
rect 5868 12044 5874 12096
rect 6733 12087 6791 12093
rect 6733 12053 6745 12087
rect 6779 12084 6791 12087
rect 6914 12084 6920 12096
rect 6779 12056 6920 12084
rect 6779 12053 6791 12056
rect 6733 12047 6791 12053
rect 6914 12044 6920 12056
rect 6972 12084 6978 12096
rect 7098 12084 7104 12096
rect 6972 12056 7104 12084
rect 6972 12044 6978 12056
rect 7098 12044 7104 12056
rect 7156 12044 7162 12096
rect 1104 11994 8832 12016
rect 1104 11942 3547 11994
rect 3599 11942 3611 11994
rect 3663 11942 3675 11994
rect 3727 11942 3739 11994
rect 3791 11942 3803 11994
rect 3855 11942 6144 11994
rect 6196 11942 6208 11994
rect 6260 11942 6272 11994
rect 6324 11942 6336 11994
rect 6388 11942 6400 11994
rect 6452 11942 8832 11994
rect 1104 11920 8832 11942
rect 7006 11812 7012 11824
rect 6967 11784 7012 11812
rect 7006 11772 7012 11784
rect 7064 11772 7070 11824
rect 6822 11744 6828 11756
rect 6735 11716 6828 11744
rect 6822 11704 6828 11716
rect 6880 11744 6886 11756
rect 7561 11747 7619 11753
rect 7561 11744 7573 11747
rect 6880 11716 7573 11744
rect 6880 11704 6886 11716
rect 7561 11713 7573 11716
rect 7607 11713 7619 11747
rect 7561 11707 7619 11713
rect 5994 11636 6000 11688
rect 6052 11676 6058 11688
rect 7469 11679 7527 11685
rect 7469 11676 7481 11679
rect 6052 11648 7481 11676
rect 6052 11636 6058 11648
rect 7469 11645 7481 11648
rect 7515 11645 7527 11679
rect 7469 11639 7527 11645
rect 8021 11679 8079 11685
rect 8021 11645 8033 11679
rect 8067 11676 8079 11679
rect 8294 11676 8300 11688
rect 8067 11648 8300 11676
rect 8067 11645 8079 11648
rect 8021 11639 8079 11645
rect 5813 11611 5871 11617
rect 5813 11577 5825 11611
rect 5859 11608 5871 11611
rect 8036 11608 8064 11639
rect 8294 11636 8300 11648
rect 8352 11636 8358 11688
rect 5859 11580 8064 11608
rect 5859 11577 5871 11580
rect 5813 11571 5871 11577
rect 5534 11500 5540 11552
rect 5592 11540 5598 11552
rect 5828 11540 5856 11571
rect 5592 11512 5856 11540
rect 5592 11500 5598 11512
rect 1104 11450 8832 11472
rect 1104 11398 2248 11450
rect 2300 11398 2312 11450
rect 2364 11398 2376 11450
rect 2428 11398 2440 11450
rect 2492 11398 2504 11450
rect 2556 11398 4846 11450
rect 4898 11398 4910 11450
rect 4962 11398 4974 11450
rect 5026 11398 5038 11450
rect 5090 11398 5102 11450
rect 5154 11398 7443 11450
rect 7495 11398 7507 11450
rect 7559 11398 7571 11450
rect 7623 11398 7635 11450
rect 7687 11398 7699 11450
rect 7751 11398 8832 11450
rect 1104 11376 8832 11398
rect 5445 11339 5503 11345
rect 5445 11305 5457 11339
rect 5491 11336 5503 11339
rect 5534 11336 5540 11348
rect 5491 11308 5540 11336
rect 5491 11305 5503 11308
rect 5445 11299 5503 11305
rect 5534 11296 5540 11308
rect 5592 11296 5598 11348
rect 5994 11336 6000 11348
rect 5955 11308 6000 11336
rect 5994 11296 6000 11308
rect 6052 11296 6058 11348
rect 6822 11268 6828 11280
rect 6783 11240 6828 11268
rect 6822 11228 6828 11240
rect 6880 11228 6886 11280
rect 7190 11132 7196 11144
rect 7151 11104 7196 11132
rect 7190 11092 7196 11104
rect 7248 11092 7254 11144
rect 8113 11135 8171 11141
rect 8113 11101 8125 11135
rect 8159 11132 8171 11135
rect 8294 11132 8300 11144
rect 8159 11104 8300 11132
rect 8159 11101 8171 11104
rect 8113 11095 8171 11101
rect 8294 11092 8300 11104
rect 8352 11092 8358 11144
rect 6089 11067 6147 11073
rect 6089 11033 6101 11067
rect 6135 11064 6147 11067
rect 7282 11064 7288 11076
rect 6135 11036 7288 11064
rect 6135 11033 6147 11036
rect 6089 11027 6147 11033
rect 7282 11024 7288 11036
rect 7340 11024 7346 11076
rect 1104 10906 8832 10928
rect 1104 10854 3547 10906
rect 3599 10854 3611 10906
rect 3663 10854 3675 10906
rect 3727 10854 3739 10906
rect 3791 10854 3803 10906
rect 3855 10854 6144 10906
rect 6196 10854 6208 10906
rect 6260 10854 6272 10906
rect 6324 10854 6336 10906
rect 6388 10854 6400 10906
rect 6452 10854 8832 10906
rect 1104 10832 8832 10854
rect 6638 10752 6644 10804
rect 6696 10792 6702 10804
rect 7926 10792 7932 10804
rect 6696 10764 7932 10792
rect 6696 10752 6702 10764
rect 7926 10752 7932 10764
rect 7984 10752 7990 10804
rect 7282 10724 7288 10736
rect 7243 10696 7288 10724
rect 7282 10684 7288 10696
rect 7340 10684 7346 10736
rect 6457 10659 6515 10665
rect 6457 10625 6469 10659
rect 6503 10656 6515 10659
rect 6546 10656 6552 10668
rect 6503 10628 6552 10656
rect 6503 10625 6515 10628
rect 6457 10619 6515 10625
rect 6546 10616 6552 10628
rect 6604 10616 6610 10668
rect 6641 10659 6699 10665
rect 6641 10625 6653 10659
rect 6687 10656 6699 10659
rect 7101 10659 7159 10665
rect 7101 10656 7113 10659
rect 6687 10628 7113 10656
rect 6687 10625 6699 10628
rect 6641 10619 6699 10625
rect 7101 10625 7113 10628
rect 7147 10656 7159 10659
rect 7190 10656 7196 10668
rect 7147 10628 7196 10656
rect 7147 10625 7159 10628
rect 7101 10619 7159 10625
rect 7190 10616 7196 10628
rect 7248 10616 7254 10668
rect 8021 10659 8079 10665
rect 8021 10625 8033 10659
rect 8067 10625 8079 10659
rect 8021 10619 8079 10625
rect 5810 10588 5816 10600
rect 5723 10560 5816 10588
rect 5810 10548 5816 10560
rect 5868 10588 5874 10600
rect 8036 10588 8064 10619
rect 5868 10560 8064 10588
rect 5868 10548 5874 10560
rect 1104 10362 8832 10384
rect 1104 10310 2248 10362
rect 2300 10310 2312 10362
rect 2364 10310 2376 10362
rect 2428 10310 2440 10362
rect 2492 10310 2504 10362
rect 2556 10310 4846 10362
rect 4898 10310 4910 10362
rect 4962 10310 4974 10362
rect 5026 10310 5038 10362
rect 5090 10310 5102 10362
rect 5154 10310 7443 10362
rect 7495 10310 7507 10362
rect 7559 10310 7571 10362
rect 7623 10310 7635 10362
rect 7687 10310 7699 10362
rect 7751 10310 8832 10362
rect 1104 10288 8832 10310
rect 5534 10072 5540 10124
rect 5592 10112 5598 10124
rect 7561 10115 7619 10121
rect 7561 10112 7573 10115
rect 5592 10084 7573 10112
rect 5592 10072 5598 10084
rect 7561 10081 7573 10084
rect 7607 10081 7619 10115
rect 7561 10075 7619 10081
rect 7101 10047 7159 10053
rect 7101 10013 7113 10047
rect 7147 10044 7159 10047
rect 7282 10044 7288 10056
rect 7147 10016 7288 10044
rect 7147 10013 7159 10016
rect 7101 10007 7159 10013
rect 7282 10004 7288 10016
rect 7340 10044 7346 10056
rect 7653 10047 7711 10053
rect 7653 10044 7665 10047
rect 7340 10016 7665 10044
rect 7340 10004 7346 10016
rect 7653 10013 7665 10016
rect 7699 10013 7711 10047
rect 8113 10047 8171 10053
rect 8113 10044 8125 10047
rect 7653 10007 7711 10013
rect 7944 10016 8125 10044
rect 6914 9976 6920 9988
rect 6875 9948 6920 9976
rect 6914 9936 6920 9948
rect 6972 9936 6978 9988
rect 7944 9920 7972 10016
rect 8113 10013 8125 10016
rect 8159 10044 8171 10047
rect 8202 10044 8208 10056
rect 8159 10016 8208 10044
rect 8159 10013 8171 10016
rect 8113 10007 8171 10013
rect 8202 10004 8208 10016
rect 8260 10004 8266 10056
rect 5442 9868 5448 9920
rect 5500 9908 5506 9920
rect 5626 9908 5632 9920
rect 5500 9880 5632 9908
rect 5500 9868 5506 9880
rect 5626 9868 5632 9880
rect 5684 9868 5690 9920
rect 6457 9911 6515 9917
rect 6457 9877 6469 9911
rect 6503 9908 6515 9911
rect 7926 9908 7932 9920
rect 6503 9880 7932 9908
rect 6503 9877 6515 9880
rect 6457 9871 6515 9877
rect 7926 9868 7932 9880
rect 7984 9868 7990 9920
rect 1104 9818 8832 9840
rect 1104 9766 3547 9818
rect 3599 9766 3611 9818
rect 3663 9766 3675 9818
rect 3727 9766 3739 9818
rect 3791 9766 3803 9818
rect 3855 9766 6144 9818
rect 6196 9766 6208 9818
rect 6260 9766 6272 9818
rect 6324 9766 6336 9818
rect 6388 9766 6400 9818
rect 6452 9766 8832 9818
rect 1104 9744 8832 9766
rect 5810 9568 5816 9580
rect 5723 9540 5816 9568
rect 5810 9528 5816 9540
rect 5868 9568 5874 9580
rect 6457 9571 6515 9577
rect 6457 9568 6469 9571
rect 5868 9540 6469 9568
rect 5868 9528 5874 9540
rect 6457 9537 6469 9540
rect 6503 9568 6515 9571
rect 6638 9568 6644 9580
rect 6503 9540 6644 9568
rect 6503 9537 6515 9540
rect 6457 9531 6515 9537
rect 6638 9528 6644 9540
rect 6696 9528 6702 9580
rect 7098 9568 7104 9580
rect 7059 9540 7104 9568
rect 7098 9528 7104 9540
rect 7156 9528 7162 9580
rect 7377 9571 7435 9577
rect 7377 9537 7389 9571
rect 7423 9568 7435 9571
rect 7834 9568 7840 9580
rect 7423 9540 7840 9568
rect 7423 9537 7435 9540
rect 7377 9531 7435 9537
rect 7834 9528 7840 9540
rect 7892 9568 7898 9580
rect 8021 9571 8079 9577
rect 8021 9568 8033 9571
rect 7892 9540 8033 9568
rect 7892 9528 7898 9540
rect 8021 9537 8033 9540
rect 8067 9537 8079 9571
rect 8021 9531 8079 9537
rect 7190 9324 7196 9376
rect 7248 9364 7254 9376
rect 7837 9367 7895 9373
rect 7837 9364 7849 9367
rect 7248 9336 7849 9364
rect 7248 9324 7254 9336
rect 7837 9333 7849 9336
rect 7883 9333 7895 9367
rect 7837 9327 7895 9333
rect 1104 9274 8832 9296
rect 1104 9222 2248 9274
rect 2300 9222 2312 9274
rect 2364 9222 2376 9274
rect 2428 9222 2440 9274
rect 2492 9222 2504 9274
rect 2556 9222 4846 9274
rect 4898 9222 4910 9274
rect 4962 9222 4974 9274
rect 5026 9222 5038 9274
rect 5090 9222 5102 9274
rect 5154 9222 7443 9274
rect 7495 9222 7507 9274
rect 7559 9222 7571 9274
rect 7623 9222 7635 9274
rect 7687 9222 7699 9274
rect 7751 9222 8832 9274
rect 1104 9200 8832 9222
rect 5537 9163 5595 9169
rect 5537 9129 5549 9163
rect 5583 9160 5595 9163
rect 5810 9160 5816 9172
rect 5583 9132 5816 9160
rect 5583 9129 5595 9132
rect 5537 9123 5595 9129
rect 5810 9120 5816 9132
rect 5868 9120 5874 9172
rect 7098 9092 7104 9104
rect 6196 9064 7104 9092
rect 6196 8965 6224 9064
rect 7098 9052 7104 9064
rect 7156 9052 7162 9104
rect 6638 9024 6644 9036
rect 6599 8996 6644 9024
rect 6638 8984 6644 8996
rect 6696 8984 6702 9036
rect 7190 9024 7196 9036
rect 7151 8996 7196 9024
rect 7190 8984 7196 8996
rect 7248 8984 7254 9036
rect 6181 8959 6239 8965
rect 6181 8925 6193 8959
rect 6227 8925 6239 8959
rect 6181 8919 6239 8925
rect 7098 8848 7104 8900
rect 7156 8888 7162 8900
rect 7745 8891 7803 8897
rect 7745 8888 7757 8891
rect 7156 8860 7757 8888
rect 7156 8848 7162 8860
rect 7745 8857 7757 8860
rect 7791 8857 7803 8891
rect 7745 8851 7803 8857
rect 4985 8823 5043 8829
rect 4985 8789 4997 8823
rect 5031 8820 5043 8823
rect 5810 8820 5816 8832
rect 5031 8792 5816 8820
rect 5031 8789 5043 8792
rect 4985 8783 5043 8789
rect 5810 8780 5816 8792
rect 5868 8780 5874 8832
rect 6089 8823 6147 8829
rect 6089 8789 6101 8823
rect 6135 8820 6147 8823
rect 6822 8820 6828 8832
rect 6135 8792 6828 8820
rect 6135 8789 6147 8792
rect 6089 8783 6147 8789
rect 6822 8780 6828 8792
rect 6880 8780 6886 8832
rect 7834 8820 7840 8832
rect 7795 8792 7840 8820
rect 7834 8780 7840 8792
rect 7892 8780 7898 8832
rect 1104 8730 8832 8752
rect 1104 8678 3547 8730
rect 3599 8678 3611 8730
rect 3663 8678 3675 8730
rect 3727 8678 3739 8730
rect 3791 8678 3803 8730
rect 3855 8678 6144 8730
rect 6196 8678 6208 8730
rect 6260 8678 6272 8730
rect 6324 8678 6336 8730
rect 6388 8678 6400 8730
rect 6452 8678 8832 8730
rect 1104 8656 8832 8678
rect 4801 8619 4859 8625
rect 4801 8585 4813 8619
rect 4847 8616 4859 8619
rect 5534 8616 5540 8628
rect 4847 8588 5540 8616
rect 4847 8585 4859 8588
rect 4801 8579 4859 8585
rect 5534 8576 5540 8588
rect 5592 8576 5598 8628
rect 5813 8551 5871 8557
rect 5813 8517 5825 8551
rect 5859 8548 5871 8551
rect 6914 8548 6920 8560
rect 5859 8520 6920 8548
rect 5859 8517 5871 8520
rect 5813 8511 5871 8517
rect 6914 8508 6920 8520
rect 6972 8508 6978 8560
rect 4617 8483 4675 8489
rect 4617 8449 4629 8483
rect 4663 8480 4675 8483
rect 7190 8480 7196 8492
rect 4663 8452 7196 8480
rect 4663 8449 4675 8452
rect 4617 8443 4675 8449
rect 7190 8440 7196 8452
rect 7248 8440 7254 8492
rect 8113 8483 8171 8489
rect 8113 8449 8125 8483
rect 8159 8449 8171 8483
rect 8113 8443 8171 8449
rect 5261 8415 5319 8421
rect 5261 8381 5273 8415
rect 5307 8381 5319 8415
rect 5261 8375 5319 8381
rect 5721 8415 5779 8421
rect 5721 8381 5733 8415
rect 5767 8412 5779 8415
rect 6546 8412 6552 8424
rect 5767 8384 6552 8412
rect 5767 8381 5779 8384
rect 5721 8375 5779 8381
rect 4157 8347 4215 8353
rect 4157 8313 4169 8347
rect 4203 8344 4215 8347
rect 5276 8344 5304 8375
rect 6546 8372 6552 8384
rect 6604 8372 6610 8424
rect 5810 8344 5816 8356
rect 4203 8316 5816 8344
rect 4203 8313 4215 8316
rect 4157 8307 4215 8313
rect 5810 8304 5816 8316
rect 5868 8344 5874 8356
rect 6454 8344 6460 8356
rect 5868 8316 6460 8344
rect 5868 8304 5874 8316
rect 6454 8304 6460 8316
rect 6512 8344 6518 8356
rect 8128 8344 8156 8443
rect 6512 8316 8156 8344
rect 6512 8304 6518 8316
rect 1104 8186 8832 8208
rect 1104 8134 2248 8186
rect 2300 8134 2312 8186
rect 2364 8134 2376 8186
rect 2428 8134 2440 8186
rect 2492 8134 2504 8186
rect 2556 8134 4846 8186
rect 4898 8134 4910 8186
rect 4962 8134 4974 8186
rect 5026 8134 5038 8186
rect 5090 8134 5102 8186
rect 5154 8134 7443 8186
rect 7495 8134 7507 8186
rect 7559 8134 7571 8186
rect 7623 8134 7635 8186
rect 7687 8134 7699 8186
rect 7751 8134 8832 8186
rect 1104 8112 8832 8134
rect 4893 8075 4951 8081
rect 4893 8041 4905 8075
rect 4939 8072 4951 8075
rect 5902 8072 5908 8084
rect 4939 8044 5908 8072
rect 4939 8041 4951 8044
rect 4893 8035 4951 8041
rect 5902 8032 5908 8044
rect 5960 8032 5966 8084
rect 5534 8004 5540 8016
rect 5495 7976 5540 8004
rect 5534 7964 5540 7976
rect 5592 7964 5598 8016
rect 3237 7939 3295 7945
rect 3237 7905 3249 7939
rect 3283 7936 3295 7939
rect 7926 7936 7932 7948
rect 3283 7908 7932 7936
rect 3283 7905 3295 7908
rect 3237 7899 3295 7905
rect 7926 7896 7932 7908
rect 7984 7936 7990 7948
rect 7984 7908 8156 7936
rect 7984 7896 7990 7908
rect 4801 7871 4859 7877
rect 4801 7837 4813 7871
rect 4847 7837 4859 7871
rect 5718 7868 5724 7880
rect 5679 7840 5724 7868
rect 4801 7831 4859 7837
rect 4341 7803 4399 7809
rect 4341 7769 4353 7803
rect 4387 7800 4399 7803
rect 4816 7800 4844 7831
rect 5718 7828 5724 7840
rect 5776 7828 5782 7880
rect 7282 7828 7288 7880
rect 7340 7868 7346 7880
rect 8128 7877 8156 7908
rect 7377 7871 7435 7877
rect 7377 7868 7389 7871
rect 7340 7840 7389 7868
rect 7340 7828 7346 7840
rect 7377 7837 7389 7840
rect 7423 7837 7435 7871
rect 7377 7831 7435 7837
rect 8113 7871 8171 7877
rect 8113 7837 8125 7871
rect 8159 7837 8171 7871
rect 8113 7831 8171 7837
rect 5626 7800 5632 7812
rect 4387 7772 5632 7800
rect 4387 7769 4399 7772
rect 4341 7763 4399 7769
rect 5626 7760 5632 7772
rect 5684 7760 5690 7812
rect 7190 7800 7196 7812
rect 7103 7772 7196 7800
rect 7190 7760 7196 7772
rect 7248 7800 7254 7812
rect 7248 7772 7328 7800
rect 7248 7760 7254 7772
rect 7300 7744 7328 7772
rect 7282 7692 7288 7744
rect 7340 7692 7346 7744
rect 1104 7642 8832 7664
rect 1104 7590 3547 7642
rect 3599 7590 3611 7642
rect 3663 7590 3675 7642
rect 3727 7590 3739 7642
rect 3791 7590 3803 7642
rect 3855 7590 6144 7642
rect 6196 7590 6208 7642
rect 6260 7590 6272 7642
rect 6324 7590 6336 7642
rect 6388 7590 6400 7642
rect 6452 7590 8832 7642
rect 1104 7568 8832 7590
rect 5718 7528 5724 7540
rect 5679 7500 5724 7528
rect 5718 7488 5724 7500
rect 5776 7488 5782 7540
rect 7098 7460 7104 7472
rect 5736 7432 7104 7460
rect 5736 7401 5764 7432
rect 7098 7420 7104 7432
rect 7156 7420 7162 7472
rect 5721 7395 5779 7401
rect 5721 7361 5733 7395
rect 5767 7361 5779 7395
rect 5721 7355 5779 7361
rect 6365 7395 6423 7401
rect 6365 7361 6377 7395
rect 6411 7361 6423 7395
rect 7834 7392 7840 7404
rect 7795 7364 7840 7392
rect 6365 7355 6423 7361
rect 3973 7327 4031 7333
rect 3973 7293 3985 7327
rect 4019 7324 4031 7327
rect 4525 7327 4583 7333
rect 4525 7324 4537 7327
rect 4019 7296 4537 7324
rect 4019 7293 4031 7296
rect 3973 7287 4031 7293
rect 4525 7293 4537 7296
rect 4571 7324 4583 7327
rect 6380 7324 6408 7355
rect 7834 7352 7840 7364
rect 7892 7352 7898 7404
rect 7926 7324 7932 7336
rect 4571 7296 7932 7324
rect 4571 7293 4583 7296
rect 4525 7287 4583 7293
rect 7926 7284 7932 7296
rect 7984 7284 7990 7336
rect 7834 7256 7840 7268
rect 7795 7228 7840 7256
rect 7834 7216 7840 7228
rect 7892 7216 7898 7268
rect 5077 7191 5135 7197
rect 5077 7157 5089 7191
rect 5123 7188 5135 7191
rect 5626 7188 5632 7200
rect 5123 7160 5632 7188
rect 5123 7157 5135 7160
rect 5077 7151 5135 7157
rect 5626 7148 5632 7160
rect 5684 7188 5690 7200
rect 6454 7188 6460 7200
rect 5684 7160 6460 7188
rect 5684 7148 5690 7160
rect 6454 7148 6460 7160
rect 6512 7148 6518 7200
rect 1104 7098 8832 7120
rect 1104 7046 2248 7098
rect 2300 7046 2312 7098
rect 2364 7046 2376 7098
rect 2428 7046 2440 7098
rect 2492 7046 2504 7098
rect 2556 7046 4846 7098
rect 4898 7046 4910 7098
rect 4962 7046 4974 7098
rect 5026 7046 5038 7098
rect 5090 7046 5102 7098
rect 5154 7046 7443 7098
rect 7495 7046 7507 7098
rect 7559 7046 7571 7098
rect 7623 7046 7635 7098
rect 7687 7046 7699 7098
rect 7751 7046 8832 7098
rect 1104 7024 8832 7046
rect 5077 6851 5135 6857
rect 5077 6817 5089 6851
rect 5123 6848 5135 6851
rect 5442 6848 5448 6860
rect 5123 6820 5448 6848
rect 5123 6817 5135 6820
rect 5077 6811 5135 6817
rect 5442 6808 5448 6820
rect 5500 6808 5506 6860
rect 6822 6808 6828 6860
rect 6880 6848 6886 6860
rect 7377 6851 7435 6857
rect 7377 6848 7389 6851
rect 6880 6820 7389 6848
rect 6880 6808 6886 6820
rect 7377 6817 7389 6820
rect 7423 6817 7435 6851
rect 7377 6811 7435 6817
rect 4430 6780 4436 6792
rect 4391 6752 4436 6780
rect 4430 6740 4436 6752
rect 4488 6740 4494 6792
rect 6454 6740 6460 6792
rect 6512 6740 6518 6792
rect 7926 6780 7932 6792
rect 7887 6752 7932 6780
rect 7926 6740 7932 6752
rect 7984 6740 7990 6792
rect 4525 6715 4583 6721
rect 4525 6681 4537 6715
rect 4571 6712 4583 6715
rect 5353 6715 5411 6721
rect 5353 6712 5365 6715
rect 4571 6684 5365 6712
rect 4571 6681 4583 6684
rect 4525 6675 4583 6681
rect 5353 6681 5365 6684
rect 5399 6681 5411 6715
rect 5353 6675 5411 6681
rect 7466 6672 7472 6724
rect 7524 6712 7530 6724
rect 7834 6712 7840 6724
rect 7524 6684 7840 6712
rect 7524 6672 7530 6684
rect 7834 6672 7840 6684
rect 7892 6672 7898 6724
rect 4430 6604 4436 6656
rect 4488 6644 4494 6656
rect 6825 6647 6883 6653
rect 6825 6644 6837 6647
rect 4488 6616 6837 6644
rect 4488 6604 4494 6616
rect 6825 6613 6837 6616
rect 6871 6613 6883 6647
rect 6825 6607 6883 6613
rect 1104 6554 8832 6576
rect 1104 6502 3547 6554
rect 3599 6502 3611 6554
rect 3663 6502 3675 6554
rect 3727 6502 3739 6554
rect 3791 6502 3803 6554
rect 3855 6502 6144 6554
rect 6196 6502 6208 6554
rect 6260 6502 6272 6554
rect 6324 6502 6336 6554
rect 6388 6502 6400 6554
rect 6452 6502 8832 6554
rect 1104 6480 8832 6502
rect 5718 6400 5724 6452
rect 5776 6440 5782 6452
rect 5902 6440 5908 6452
rect 5776 6412 5908 6440
rect 5776 6400 5782 6412
rect 5902 6400 5908 6412
rect 5960 6400 5966 6452
rect 5629 6375 5687 6381
rect 5629 6341 5641 6375
rect 5675 6372 5687 6375
rect 7466 6372 7472 6384
rect 5675 6344 7472 6372
rect 5675 6341 5687 6344
rect 5629 6335 5687 6341
rect 7466 6332 7472 6344
rect 7524 6332 7530 6384
rect 5077 6307 5135 6313
rect 5077 6273 5089 6307
rect 5123 6304 5135 6307
rect 5902 6304 5908 6316
rect 5123 6276 5908 6304
rect 5123 6273 5135 6276
rect 5077 6267 5135 6273
rect 5902 6264 5908 6276
rect 5960 6264 5966 6316
rect 7098 6304 7104 6316
rect 6840 6276 7104 6304
rect 5813 6239 5871 6245
rect 5813 6205 5825 6239
rect 5859 6236 5871 6239
rect 6840 6236 6868 6276
rect 7098 6264 7104 6276
rect 7156 6304 7162 6316
rect 8113 6307 8171 6313
rect 8113 6304 8125 6307
rect 7156 6276 8125 6304
rect 7156 6264 7162 6276
rect 8113 6273 8125 6276
rect 8159 6273 8171 6307
rect 8113 6267 8171 6273
rect 5859 6208 6868 6236
rect 6917 6239 6975 6245
rect 5859 6205 5871 6208
rect 5813 6199 5871 6205
rect 6917 6205 6929 6239
rect 6963 6205 6975 6239
rect 6917 6199 6975 6205
rect 7469 6239 7527 6245
rect 7469 6205 7481 6239
rect 7515 6205 7527 6239
rect 7469 6199 7527 6205
rect 3881 6171 3939 6177
rect 3881 6137 3893 6171
rect 3927 6168 3939 6171
rect 4433 6171 4491 6177
rect 4433 6168 4445 6171
rect 3927 6140 4445 6168
rect 3927 6137 3939 6140
rect 3881 6131 3939 6137
rect 4433 6137 4445 6140
rect 4479 6168 4491 6171
rect 6932 6168 6960 6199
rect 4479 6140 6960 6168
rect 4479 6137 4491 6140
rect 4433 6131 4491 6137
rect 4985 6103 5043 6109
rect 4985 6069 4997 6103
rect 5031 6100 5043 6103
rect 5810 6100 5816 6112
rect 5031 6072 5816 6100
rect 5031 6069 5043 6072
rect 4985 6063 5043 6069
rect 5810 6060 5816 6072
rect 5868 6060 5874 6112
rect 5994 6060 6000 6112
rect 6052 6100 6058 6112
rect 6365 6103 6423 6109
rect 6365 6100 6377 6103
rect 6052 6072 6377 6100
rect 6052 6060 6058 6072
rect 6365 6069 6377 6072
rect 6411 6100 6423 6103
rect 6546 6100 6552 6112
rect 6411 6072 6552 6100
rect 6411 6069 6423 6072
rect 6365 6063 6423 6069
rect 6546 6060 6552 6072
rect 6604 6060 6610 6112
rect 6932 6100 6960 6140
rect 7006 6128 7012 6180
rect 7064 6168 7070 6180
rect 7377 6171 7435 6177
rect 7377 6168 7389 6171
rect 7064 6140 7389 6168
rect 7064 6128 7070 6140
rect 7377 6137 7389 6140
rect 7423 6137 7435 6171
rect 7484 6168 7512 6199
rect 7929 6171 7987 6177
rect 7929 6168 7941 6171
rect 7484 6140 7941 6168
rect 7377 6131 7435 6137
rect 7929 6137 7941 6140
rect 7975 6137 7987 6171
rect 7929 6131 7987 6137
rect 8110 6100 8116 6112
rect 6932 6072 8116 6100
rect 8110 6060 8116 6072
rect 8168 6060 8174 6112
rect 1104 6010 8832 6032
rect 1104 5958 2248 6010
rect 2300 5958 2312 6010
rect 2364 5958 2376 6010
rect 2428 5958 2440 6010
rect 2492 5958 2504 6010
rect 2556 5958 4846 6010
rect 4898 5958 4910 6010
rect 4962 5958 4974 6010
rect 5026 5958 5038 6010
rect 5090 5958 5102 6010
rect 5154 5958 7443 6010
rect 7495 5958 7507 6010
rect 7559 5958 7571 6010
rect 7623 5958 7635 6010
rect 7687 5958 7699 6010
rect 7751 5958 8832 6010
rect 1104 5936 8832 5958
rect 6362 5856 6368 5908
rect 6420 5896 6426 5908
rect 8018 5896 8024 5908
rect 6420 5868 8024 5896
rect 6420 5856 6426 5868
rect 8018 5856 8024 5868
rect 8076 5856 8082 5908
rect 7190 5828 7196 5840
rect 4540 5800 7196 5828
rect 4540 5701 4568 5800
rect 7190 5788 7196 5800
rect 7248 5788 7254 5840
rect 5261 5763 5319 5769
rect 5261 5729 5273 5763
rect 5307 5760 5319 5763
rect 6914 5760 6920 5772
rect 5307 5732 6920 5760
rect 5307 5729 5319 5732
rect 5261 5723 5319 5729
rect 6914 5720 6920 5732
rect 6972 5720 6978 5772
rect 4525 5695 4583 5701
rect 4525 5661 4537 5695
rect 4571 5661 4583 5695
rect 5718 5692 5724 5704
rect 4525 5655 4583 5661
rect 4632 5664 5724 5692
rect 3234 5624 3240 5636
rect 3147 5596 3240 5624
rect 3234 5584 3240 5596
rect 3292 5624 3298 5636
rect 4632 5624 4660 5664
rect 5718 5652 5724 5664
rect 5776 5692 5782 5704
rect 6362 5692 6368 5704
rect 5776 5664 6368 5692
rect 5776 5652 5782 5664
rect 6362 5652 6368 5664
rect 6420 5652 6426 5704
rect 6825 5695 6883 5701
rect 6825 5661 6837 5695
rect 6871 5692 6883 5695
rect 7098 5692 7104 5704
rect 6871 5664 7104 5692
rect 6871 5661 6883 5664
rect 6825 5655 6883 5661
rect 7098 5652 7104 5664
rect 7156 5652 7162 5704
rect 7745 5695 7803 5701
rect 7745 5661 7757 5695
rect 7791 5692 7803 5695
rect 8110 5692 8116 5704
rect 7791 5664 8116 5692
rect 7791 5661 7803 5664
rect 7745 5655 7803 5661
rect 8110 5652 8116 5664
rect 8168 5652 8174 5704
rect 5813 5627 5871 5633
rect 5813 5624 5825 5627
rect 3292 5596 4660 5624
rect 4724 5596 5825 5624
rect 3292 5584 3298 5596
rect 4062 5556 4068 5568
rect 4023 5528 4068 5556
rect 4062 5516 4068 5528
rect 4120 5516 4126 5568
rect 4724 5565 4752 5596
rect 5813 5593 5825 5596
rect 5859 5593 5871 5627
rect 5813 5587 5871 5593
rect 5902 5584 5908 5636
rect 5960 5624 5966 5636
rect 5960 5596 6005 5624
rect 5960 5584 5966 5596
rect 7006 5584 7012 5636
rect 7064 5624 7070 5636
rect 7064 5596 7157 5624
rect 7064 5584 7070 5596
rect 4709 5559 4767 5565
rect 4709 5525 4721 5559
rect 4755 5525 4767 5559
rect 4709 5519 4767 5525
rect 5353 5559 5411 5565
rect 5353 5525 5365 5559
rect 5399 5556 5411 5559
rect 7024 5556 7052 5584
rect 5399 5528 7052 5556
rect 5399 5525 5411 5528
rect 5353 5519 5411 5525
rect 1104 5466 8832 5488
rect 1104 5414 3547 5466
rect 3599 5414 3611 5466
rect 3663 5414 3675 5466
rect 3727 5414 3739 5466
rect 3791 5414 3803 5466
rect 3855 5414 6144 5466
rect 6196 5414 6208 5466
rect 6260 5414 6272 5466
rect 6324 5414 6336 5466
rect 6388 5414 6400 5466
rect 6452 5414 8832 5466
rect 1104 5392 8832 5414
rect 2593 5355 2651 5361
rect 2593 5321 2605 5355
rect 2639 5352 2651 5355
rect 3234 5352 3240 5364
rect 2639 5324 3240 5352
rect 2639 5321 2651 5324
rect 2593 5315 2651 5321
rect 3234 5312 3240 5324
rect 3292 5312 3298 5364
rect 5077 5355 5135 5361
rect 5077 5321 5089 5355
rect 5123 5352 5135 5355
rect 5534 5352 5540 5364
rect 5123 5324 5540 5352
rect 5123 5321 5135 5324
rect 5077 5315 5135 5321
rect 5534 5312 5540 5324
rect 5592 5312 5598 5364
rect 6549 5355 6607 5361
rect 6549 5321 6561 5355
rect 6595 5352 6607 5355
rect 7282 5352 7288 5364
rect 6595 5324 7288 5352
rect 6595 5321 6607 5324
rect 6549 5315 6607 5321
rect 7282 5312 7288 5324
rect 7340 5312 7346 5364
rect 5902 5244 5908 5296
rect 5960 5284 5966 5296
rect 7377 5287 7435 5293
rect 7377 5284 7389 5287
rect 5960 5256 7389 5284
rect 5960 5244 5966 5256
rect 7377 5253 7389 5256
rect 7423 5253 7435 5287
rect 7377 5247 7435 5253
rect 4341 5219 4399 5225
rect 4341 5216 4353 5219
rect 3620 5188 4353 5216
rect 2866 5040 2872 5092
rect 2924 5080 2930 5092
rect 3620 5089 3648 5188
rect 4341 5185 4353 5188
rect 4387 5185 4399 5219
rect 5166 5216 5172 5228
rect 5127 5188 5172 5216
rect 4341 5179 4399 5185
rect 5166 5176 5172 5188
rect 5224 5176 5230 5228
rect 6546 5176 6552 5228
rect 6604 5216 6610 5228
rect 6641 5219 6699 5225
rect 6641 5216 6653 5219
rect 6604 5188 6653 5216
rect 6604 5176 6610 5188
rect 6641 5185 6653 5188
rect 6687 5185 6699 5219
rect 7190 5216 7196 5228
rect 7151 5188 7196 5216
rect 6641 5179 6699 5185
rect 7190 5176 7196 5188
rect 7248 5176 7254 5228
rect 8018 5176 8024 5228
rect 8076 5216 8082 5228
rect 8113 5219 8171 5225
rect 8113 5216 8125 5219
rect 8076 5188 8125 5216
rect 8076 5176 8082 5188
rect 8113 5185 8125 5188
rect 8159 5185 8171 5219
rect 8113 5179 8171 5185
rect 4706 5108 4712 5160
rect 4764 5148 4770 5160
rect 4893 5151 4951 5157
rect 4893 5148 4905 5151
rect 4764 5120 4905 5148
rect 4764 5108 4770 5120
rect 4893 5117 4905 5120
rect 4939 5117 4951 5151
rect 4893 5111 4951 5117
rect 3605 5083 3663 5089
rect 3605 5080 3617 5083
rect 2924 5052 3617 5080
rect 2924 5040 2930 5052
rect 3605 5049 3617 5052
rect 3651 5049 3663 5083
rect 5537 5083 5595 5089
rect 3605 5043 3663 5049
rect 4172 5052 5488 5080
rect 3050 4972 3056 5024
rect 3108 5012 3114 5024
rect 3145 5015 3203 5021
rect 3145 5012 3157 5015
rect 3108 4984 3157 5012
rect 3108 4972 3114 4984
rect 3145 4981 3157 4984
rect 3191 5012 3203 5015
rect 4172 5012 4200 5052
rect 3191 4984 4200 5012
rect 4249 5015 4307 5021
rect 3191 4981 3203 4984
rect 3145 4975 3203 4981
rect 4249 4981 4261 5015
rect 4295 5012 4307 5015
rect 4338 5012 4344 5024
rect 4295 4984 4344 5012
rect 4295 4981 4307 4984
rect 4249 4975 4307 4981
rect 4338 4972 4344 4984
rect 4396 4972 4402 5024
rect 5460 5012 5488 5052
rect 5537 5049 5549 5083
rect 5583 5080 5595 5083
rect 6914 5080 6920 5092
rect 5583 5052 6920 5080
rect 5583 5049 5595 5052
rect 5537 5043 5595 5049
rect 6914 5040 6920 5052
rect 6972 5040 6978 5092
rect 8110 5012 8116 5024
rect 5460 4984 8116 5012
rect 8110 4972 8116 4984
rect 8168 4972 8174 5024
rect 1104 4922 8832 4944
rect 1104 4870 2248 4922
rect 2300 4870 2312 4922
rect 2364 4870 2376 4922
rect 2428 4870 2440 4922
rect 2492 4870 2504 4922
rect 2556 4870 4846 4922
rect 4898 4870 4910 4922
rect 4962 4870 4974 4922
rect 5026 4870 5038 4922
rect 5090 4870 5102 4922
rect 5154 4870 7443 4922
rect 7495 4870 7507 4922
rect 7559 4870 7571 4922
rect 7623 4870 7635 4922
rect 7687 4870 7699 4922
rect 7751 4870 8832 4922
rect 1104 4848 8832 4870
rect 4816 4780 7696 4808
rect 4816 4752 4844 4780
rect 4430 4700 4436 4752
rect 4488 4740 4494 4752
rect 4798 4740 4804 4752
rect 4488 4712 4804 4740
rect 4488 4700 4494 4712
rect 4798 4700 4804 4712
rect 4856 4700 4862 4752
rect 7024 4712 7604 4740
rect 4154 4632 4160 4684
rect 4212 4672 4218 4684
rect 4341 4675 4399 4681
rect 4341 4672 4353 4675
rect 4212 4644 4353 4672
rect 4212 4632 4218 4644
rect 4341 4641 4353 4644
rect 4387 4672 4399 4675
rect 4614 4672 4620 4684
rect 4387 4644 4620 4672
rect 4387 4641 4399 4644
rect 4341 4635 4399 4641
rect 4614 4632 4620 4644
rect 4672 4632 4678 4684
rect 5810 4632 5816 4684
rect 5868 4672 5874 4684
rect 7024 4672 7052 4712
rect 7576 4681 7604 4712
rect 5868 4644 7052 4672
rect 7561 4675 7619 4681
rect 5868 4632 5874 4644
rect 7561 4641 7573 4675
rect 7607 4641 7619 4675
rect 7561 4635 7619 4641
rect 4433 4607 4491 4613
rect 4433 4573 4445 4607
rect 4479 4573 4491 4607
rect 4433 4567 4491 4573
rect 4154 4536 4160 4548
rect 4115 4508 4160 4536
rect 4154 4496 4160 4508
rect 4212 4496 4218 4548
rect 4448 4536 4476 4567
rect 4522 4564 4528 4616
rect 4580 4604 4586 4616
rect 4709 4607 4767 4613
rect 4709 4604 4721 4607
rect 4580 4576 4721 4604
rect 4580 4564 4586 4576
rect 4709 4573 4721 4576
rect 4755 4573 4767 4607
rect 4709 4567 4767 4573
rect 7101 4607 7159 4613
rect 7101 4573 7113 4607
rect 7147 4604 7159 4607
rect 7668 4604 7696 4780
rect 8110 4604 8116 4616
rect 7147 4576 7696 4604
rect 8071 4576 8116 4604
rect 7147 4573 7159 4576
rect 7101 4567 7159 4573
rect 8110 4564 8116 4576
rect 8168 4564 8174 4616
rect 6822 4536 6828 4548
rect 4356 4508 4476 4536
rect 2682 4468 2688 4480
rect 2643 4440 2688 4468
rect 2682 4428 2688 4440
rect 2740 4428 2746 4480
rect 2866 4428 2872 4480
rect 2924 4468 2930 4480
rect 3145 4471 3203 4477
rect 3145 4468 3157 4471
rect 2924 4440 3157 4468
rect 2924 4428 2930 4440
rect 3145 4437 3157 4440
rect 3191 4468 3203 4471
rect 4356 4468 4384 4508
rect 6012 4480 6040 4522
rect 6783 4508 6828 4536
rect 6822 4496 6828 4508
rect 6880 4496 6886 4548
rect 7653 4539 7711 4545
rect 7653 4505 7665 4539
rect 7699 4505 7711 4539
rect 7653 4499 7711 4505
rect 3191 4440 4384 4468
rect 5353 4471 5411 4477
rect 3191 4437 3203 4440
rect 3145 4431 3203 4437
rect 5353 4437 5365 4471
rect 5399 4468 5411 4471
rect 5442 4468 5448 4480
rect 5399 4440 5448 4468
rect 5399 4437 5411 4440
rect 5353 4431 5411 4437
rect 5442 4428 5448 4440
rect 5500 4428 5506 4480
rect 5994 4428 6000 4480
rect 6052 4428 6058 4480
rect 6546 4428 6552 4480
rect 6604 4468 6610 4480
rect 7668 4468 7696 4499
rect 6604 4440 7696 4468
rect 6604 4428 6610 4440
rect 1104 4378 8832 4400
rect 1104 4326 3547 4378
rect 3599 4326 3611 4378
rect 3663 4326 3675 4378
rect 3727 4326 3739 4378
rect 3791 4326 3803 4378
rect 3855 4326 6144 4378
rect 6196 4326 6208 4378
rect 6260 4326 6272 4378
rect 6324 4326 6336 4378
rect 6388 4326 6400 4378
rect 6452 4326 8832 4378
rect 1104 4304 8832 4326
rect 3329 4267 3387 4273
rect 3329 4233 3341 4267
rect 3375 4264 3387 4267
rect 4430 4264 4436 4276
rect 3375 4236 4436 4264
rect 3375 4233 3387 4236
rect 3329 4227 3387 4233
rect 4430 4224 4436 4236
rect 4488 4224 4494 4276
rect 4617 4267 4675 4273
rect 4617 4233 4629 4267
rect 4663 4264 4675 4267
rect 5166 4264 5172 4276
rect 4663 4236 5172 4264
rect 4663 4233 4675 4236
rect 4617 4227 4675 4233
rect 5166 4224 5172 4236
rect 5224 4224 5230 4276
rect 5445 4267 5503 4273
rect 5445 4233 5457 4267
rect 5491 4264 5503 4267
rect 5534 4264 5540 4276
rect 5491 4236 5540 4264
rect 5491 4233 5503 4236
rect 5445 4227 5503 4233
rect 5534 4224 5540 4236
rect 5592 4224 5598 4276
rect 4154 4156 4160 4208
rect 4212 4156 4218 4208
rect 6546 4196 6552 4208
rect 6507 4168 6552 4196
rect 6546 4156 6552 4168
rect 6604 4156 6610 4208
rect 2777 4131 2835 4137
rect 2777 4128 2789 4131
rect 2240 4100 2789 4128
rect 934 3952 940 4004
rect 992 3992 998 4004
rect 2240 4001 2268 4100
rect 2777 4097 2789 4100
rect 2823 4097 2835 4131
rect 2777 4091 2835 4097
rect 3145 4131 3203 4137
rect 3145 4097 3157 4131
rect 3191 4128 3203 4131
rect 4172 4128 4200 4156
rect 3191 4100 3924 4128
rect 3191 4097 3203 4100
rect 3145 4091 3203 4097
rect 3237 4063 3295 4069
rect 3237 4029 3249 4063
rect 3283 4029 3295 4063
rect 3237 4023 3295 4029
rect 2225 3995 2283 4001
rect 2225 3992 2237 3995
rect 992 3964 2237 3992
rect 992 3952 998 3964
rect 2225 3961 2237 3964
rect 2271 3961 2283 3995
rect 2225 3955 2283 3961
rect 3252 3936 3280 4023
rect 3896 3992 3924 4100
rect 4080 4100 4200 4128
rect 4080 4069 4108 4100
rect 4246 4088 4252 4140
rect 4304 4128 4310 4140
rect 7190 4128 7196 4140
rect 4304 4100 4349 4128
rect 7151 4100 7196 4128
rect 4304 4088 4310 4100
rect 7190 4088 7196 4100
rect 7248 4088 7254 4140
rect 8110 4128 8116 4140
rect 8071 4100 8116 4128
rect 8110 4088 8116 4100
rect 8168 4088 8174 4140
rect 4065 4063 4123 4069
rect 4065 4029 4077 4063
rect 4111 4029 4123 4063
rect 4065 4023 4123 4029
rect 4157 4063 4215 4069
rect 4157 4029 4169 4063
rect 4203 4060 4215 4063
rect 4798 4060 4804 4072
rect 4203 4032 4804 4060
rect 4203 4029 4215 4032
rect 4157 4023 4215 4029
rect 4798 4020 4804 4032
rect 4856 4020 4862 4072
rect 5534 4060 5540 4072
rect 5495 4032 5540 4060
rect 5534 4020 5540 4032
rect 5592 4020 5598 4072
rect 5629 4063 5687 4069
rect 5629 4029 5641 4063
rect 5675 4029 5687 4063
rect 5629 4023 5687 4029
rect 4338 3992 4344 4004
rect 3896 3964 4344 3992
rect 4338 3952 4344 3964
rect 4396 3952 4402 4004
rect 5166 3952 5172 4004
rect 5224 3992 5230 4004
rect 5644 3992 5672 4023
rect 5224 3964 5672 3992
rect 5224 3952 5230 3964
rect 1765 3927 1823 3933
rect 1765 3893 1777 3927
rect 1811 3924 1823 3927
rect 3050 3924 3056 3936
rect 1811 3896 3056 3924
rect 1811 3893 1823 3896
rect 1765 3887 1823 3893
rect 3050 3884 3056 3896
rect 3108 3884 3114 3936
rect 3234 3924 3240 3936
rect 3147 3896 3240 3924
rect 3234 3884 3240 3896
rect 3292 3924 3298 3936
rect 4614 3924 4620 3936
rect 3292 3896 4620 3924
rect 3292 3884 3298 3896
rect 4614 3884 4620 3896
rect 4672 3884 4678 3936
rect 5077 3927 5135 3933
rect 5077 3893 5089 3927
rect 5123 3924 5135 3927
rect 5350 3924 5356 3936
rect 5123 3896 5356 3924
rect 5123 3893 5135 3896
rect 5077 3887 5135 3893
rect 5350 3884 5356 3896
rect 5408 3884 5414 3936
rect 1104 3834 8832 3856
rect 1104 3782 2248 3834
rect 2300 3782 2312 3834
rect 2364 3782 2376 3834
rect 2428 3782 2440 3834
rect 2492 3782 2504 3834
rect 2556 3782 4846 3834
rect 4898 3782 4910 3834
rect 4962 3782 4974 3834
rect 5026 3782 5038 3834
rect 5090 3782 5102 3834
rect 5154 3782 7443 3834
rect 7495 3782 7507 3834
rect 7559 3782 7571 3834
rect 7623 3782 7635 3834
rect 7687 3782 7699 3834
rect 7751 3782 8832 3834
rect 1104 3760 8832 3782
rect 5534 3680 5540 3732
rect 5592 3720 5598 3732
rect 6730 3720 6736 3732
rect 5592 3692 6736 3720
rect 5592 3680 5598 3692
rect 6730 3680 6736 3692
rect 6788 3720 6794 3732
rect 7193 3723 7251 3729
rect 7193 3720 7205 3723
rect 6788 3692 7205 3720
rect 6788 3680 6794 3692
rect 7193 3689 7205 3692
rect 7239 3689 7251 3723
rect 7193 3683 7251 3689
rect 2682 3652 2688 3664
rect 2595 3624 2688 3652
rect 2682 3612 2688 3624
rect 2740 3652 2746 3664
rect 3234 3652 3240 3664
rect 2740 3624 3240 3652
rect 2740 3612 2746 3624
rect 3234 3612 3240 3624
rect 3292 3612 3298 3664
rect 3160 3556 4660 3584
rect 2866 3340 2872 3392
rect 2924 3380 2930 3392
rect 3160 3389 3188 3556
rect 4632 3525 4660 3556
rect 4706 3544 4712 3596
rect 4764 3584 4770 3596
rect 4985 3587 5043 3593
rect 4985 3584 4997 3587
rect 4764 3556 4997 3584
rect 4764 3544 4770 3556
rect 4985 3553 4997 3556
rect 5031 3553 5043 3587
rect 5442 3584 5448 3596
rect 5403 3556 5448 3584
rect 4985 3547 5043 3553
rect 5442 3544 5448 3556
rect 5500 3544 5506 3596
rect 7190 3544 7196 3596
rect 7248 3584 7254 3596
rect 7837 3587 7895 3593
rect 7837 3584 7849 3587
rect 7248 3556 7849 3584
rect 7248 3544 7254 3556
rect 7837 3553 7849 3556
rect 7883 3553 7895 3587
rect 7837 3547 7895 3553
rect 4341 3519 4399 3525
rect 4341 3516 4353 3519
rect 3896 3488 4353 3516
rect 3896 3392 3924 3488
rect 4341 3485 4353 3488
rect 4387 3485 4399 3519
rect 4341 3479 4399 3485
rect 4617 3519 4675 3525
rect 4617 3485 4629 3519
rect 4663 3485 4675 3519
rect 4617 3479 4675 3485
rect 4801 3519 4859 3525
rect 4801 3485 4813 3519
rect 4847 3485 4859 3519
rect 4801 3479 4859 3485
rect 4706 3408 4712 3460
rect 4764 3448 4770 3460
rect 4816 3448 4844 3479
rect 5718 3448 5724 3460
rect 4764 3420 4844 3448
rect 5679 3420 5724 3448
rect 4764 3408 4770 3420
rect 5718 3408 5724 3420
rect 5776 3408 5782 3460
rect 8018 3448 8024 3460
rect 3145 3383 3203 3389
rect 3145 3380 3157 3383
rect 2924 3352 3157 3380
rect 2924 3340 2930 3352
rect 3145 3349 3157 3352
rect 3191 3349 3203 3383
rect 3878 3380 3884 3392
rect 3839 3352 3884 3380
rect 3145 3343 3203 3349
rect 3878 3340 3884 3352
rect 3936 3340 3942 3392
rect 5994 3340 6000 3392
rect 6052 3380 6058 3392
rect 6932 3380 6960 3434
rect 7979 3420 8024 3448
rect 8018 3408 8024 3420
rect 8076 3408 8082 3460
rect 8938 3380 8944 3392
rect 6052 3352 8944 3380
rect 6052 3340 6058 3352
rect 8938 3340 8944 3352
rect 8996 3340 9002 3392
rect 1104 3290 8832 3312
rect 1104 3238 3547 3290
rect 3599 3238 3611 3290
rect 3663 3238 3675 3290
rect 3727 3238 3739 3290
rect 3791 3238 3803 3290
rect 3855 3238 6144 3290
rect 6196 3238 6208 3290
rect 6260 3238 6272 3290
rect 6324 3238 6336 3290
rect 6388 3238 6400 3290
rect 6452 3238 8832 3290
rect 1104 3216 8832 3238
rect 4246 3136 4252 3188
rect 4304 3176 4310 3188
rect 4985 3179 5043 3185
rect 4985 3176 4997 3179
rect 4304 3148 4997 3176
rect 4304 3136 4310 3148
rect 4985 3145 4997 3148
rect 5031 3145 5043 3179
rect 5350 3176 5356 3188
rect 5311 3148 5356 3176
rect 4985 3139 5043 3145
rect 5350 3136 5356 3148
rect 5408 3136 5414 3188
rect 5442 3136 5448 3188
rect 5500 3176 5506 3188
rect 5500 3148 5545 3176
rect 5500 3136 5506 3148
rect 4341 3111 4399 3117
rect 4341 3077 4353 3111
rect 4387 3108 4399 3111
rect 4522 3108 4528 3120
rect 4387 3080 4528 3108
rect 4387 3077 4399 3080
rect 4341 3071 4399 3077
rect 4522 3068 4528 3080
rect 4580 3068 4586 3120
rect 4249 3043 4307 3049
rect 4249 3009 4261 3043
rect 4295 3009 4307 3043
rect 6546 3040 6552 3052
rect 6507 3012 6552 3040
rect 4249 3003 4307 3009
rect 934 2932 940 2984
rect 992 2972 998 2984
rect 3697 2975 3755 2981
rect 3697 2972 3709 2975
rect 992 2944 3709 2972
rect 992 2932 998 2944
rect 3697 2941 3709 2944
rect 3743 2972 3755 2975
rect 3878 2972 3884 2984
rect 3743 2944 3884 2972
rect 3743 2941 3755 2944
rect 3697 2935 3755 2941
rect 3878 2932 3884 2944
rect 3936 2972 3942 2984
rect 4264 2972 4292 3003
rect 6546 3000 6552 3012
rect 6604 3000 6610 3052
rect 7098 3000 7104 3052
rect 7156 3040 7162 3052
rect 7469 3043 7527 3049
rect 7469 3040 7481 3043
rect 7156 3012 7481 3040
rect 7156 3000 7162 3012
rect 7469 3009 7481 3012
rect 7515 3009 7527 3043
rect 7469 3003 7527 3009
rect 3936 2944 4292 2972
rect 3936 2932 3942 2944
rect 4430 2932 4436 2984
rect 4488 2972 4494 2984
rect 5537 2975 5595 2981
rect 5537 2972 5549 2975
rect 4488 2944 5549 2972
rect 4488 2932 4494 2944
rect 5537 2941 5549 2944
rect 5583 2941 5595 2975
rect 5537 2935 5595 2941
rect 3050 2864 3056 2916
rect 3108 2904 3114 2916
rect 6546 2904 6552 2916
rect 3108 2876 6552 2904
rect 3108 2864 3114 2876
rect 6546 2864 6552 2876
rect 6604 2864 6610 2916
rect 7190 2864 7196 2916
rect 7248 2904 7254 2916
rect 7837 2907 7895 2913
rect 7837 2904 7849 2907
rect 7248 2876 7849 2904
rect 7248 2864 7254 2876
rect 7837 2873 7849 2876
rect 7883 2904 7895 2907
rect 8018 2904 8024 2916
rect 7883 2876 8024 2904
rect 7883 2873 7895 2876
rect 7837 2867 7895 2873
rect 8018 2864 8024 2876
rect 8076 2864 8082 2916
rect 2685 2839 2743 2845
rect 2685 2805 2697 2839
rect 2731 2836 2743 2839
rect 3068 2836 3096 2864
rect 2731 2808 3096 2836
rect 3237 2839 3295 2845
rect 2731 2805 2743 2808
rect 2685 2799 2743 2805
rect 3237 2805 3249 2839
rect 3283 2836 3295 2839
rect 5994 2836 6000 2848
rect 3283 2808 6000 2836
rect 3283 2805 3295 2808
rect 3237 2799 3295 2805
rect 5994 2796 6000 2808
rect 6052 2796 6058 2848
rect 1104 2746 8832 2768
rect 1104 2694 2248 2746
rect 2300 2694 2312 2746
rect 2364 2694 2376 2746
rect 2428 2694 2440 2746
rect 2492 2694 2504 2746
rect 2556 2694 4846 2746
rect 4898 2694 4910 2746
rect 4962 2694 4974 2746
rect 5026 2694 5038 2746
rect 5090 2694 5102 2746
rect 5154 2694 7443 2746
rect 7495 2694 7507 2746
rect 7559 2694 7571 2746
rect 7623 2694 7635 2746
rect 7687 2694 7699 2746
rect 7751 2694 8832 2746
rect 1104 2672 8832 2694
rect 3050 2592 3056 2644
rect 3108 2632 3114 2644
rect 3145 2635 3203 2641
rect 3145 2632 3157 2635
rect 3108 2604 3157 2632
rect 3108 2592 3114 2604
rect 3145 2601 3157 2604
rect 3191 2601 3203 2635
rect 3145 2595 3203 2601
rect 5718 2592 5724 2644
rect 5776 2632 5782 2644
rect 6457 2635 6515 2641
rect 6457 2632 6469 2635
rect 5776 2604 6469 2632
rect 5776 2592 5782 2604
rect 6457 2601 6469 2604
rect 6503 2601 6515 2635
rect 6457 2595 6515 2601
rect 6546 2524 6552 2576
rect 6604 2564 6610 2576
rect 6604 2536 7696 2564
rect 6604 2524 6610 2536
rect 4246 2456 4252 2508
rect 4304 2496 4310 2508
rect 5166 2496 5172 2508
rect 4304 2468 4844 2496
rect 5127 2468 5172 2496
rect 4304 2456 4310 2468
rect 4522 2428 4528 2440
rect 4483 2400 4528 2428
rect 4522 2388 4528 2400
rect 4580 2388 4586 2440
rect 4816 2437 4844 2468
rect 5166 2456 5172 2468
rect 5224 2456 5230 2508
rect 5721 2499 5779 2505
rect 5721 2465 5733 2499
rect 5767 2496 5779 2499
rect 6822 2496 6828 2508
rect 5767 2468 6828 2496
rect 5767 2465 5779 2468
rect 5721 2459 5779 2465
rect 6822 2456 6828 2468
rect 6880 2456 6886 2508
rect 7190 2496 7196 2508
rect 7151 2468 7196 2496
rect 7190 2456 7196 2468
rect 7248 2456 7254 2508
rect 7668 2440 7696 2536
rect 4801 2431 4859 2437
rect 4801 2397 4813 2431
rect 4847 2397 4859 2431
rect 4801 2391 4859 2397
rect 4890 2388 4896 2440
rect 4948 2428 4954 2440
rect 4985 2431 5043 2437
rect 4985 2428 4997 2431
rect 4948 2400 4997 2428
rect 4948 2388 4954 2400
rect 4985 2397 4997 2400
rect 5031 2397 5043 2431
rect 4985 2391 5043 2397
rect 5442 2388 5448 2440
rect 5500 2428 5506 2440
rect 5629 2431 5687 2437
rect 5629 2428 5641 2431
rect 5500 2400 5641 2428
rect 5500 2388 5506 2400
rect 5629 2397 5641 2400
rect 5675 2397 5687 2431
rect 5629 2391 5687 2397
rect 6549 2431 6607 2437
rect 6549 2397 6561 2431
rect 6595 2428 6607 2431
rect 6730 2428 6736 2440
rect 6595 2400 6736 2428
rect 6595 2397 6607 2400
rect 6549 2391 6607 2397
rect 6730 2388 6736 2400
rect 6788 2388 6794 2440
rect 7006 2388 7012 2440
rect 7064 2428 7070 2440
rect 7101 2431 7159 2437
rect 7101 2428 7113 2431
rect 7064 2400 7113 2428
rect 7064 2388 7070 2400
rect 7101 2397 7113 2400
rect 7147 2397 7159 2431
rect 7650 2428 7656 2440
rect 7611 2400 7656 2428
rect 7101 2391 7159 2397
rect 7650 2388 7656 2400
rect 7708 2388 7714 2440
rect 4065 2363 4123 2369
rect 4065 2329 4077 2363
rect 4111 2360 4123 2363
rect 4706 2360 4712 2372
rect 4111 2332 4712 2360
rect 4111 2329 4123 2332
rect 4065 2323 4123 2329
rect 4706 2320 4712 2332
rect 4764 2360 4770 2372
rect 4908 2360 4936 2388
rect 4764 2332 4936 2360
rect 4764 2320 4770 2332
rect 1104 2202 8832 2224
rect 1104 2150 3547 2202
rect 3599 2150 3611 2202
rect 3663 2150 3675 2202
rect 3727 2150 3739 2202
rect 3791 2150 3803 2202
rect 3855 2150 6144 2202
rect 6196 2150 6208 2202
rect 6260 2150 6272 2202
rect 6324 2150 6336 2202
rect 6388 2150 6400 2202
rect 6452 2150 8832 2202
rect 1104 2128 8832 2150
<< via1 >>
rect 2248 27718 2300 27770
rect 2312 27718 2364 27770
rect 2376 27718 2428 27770
rect 2440 27718 2492 27770
rect 2504 27718 2556 27770
rect 4846 27718 4898 27770
rect 4910 27718 4962 27770
rect 4974 27718 5026 27770
rect 5038 27718 5090 27770
rect 5102 27718 5154 27770
rect 7443 27718 7495 27770
rect 7507 27718 7559 27770
rect 7571 27718 7623 27770
rect 7635 27718 7687 27770
rect 7699 27718 7751 27770
rect 7012 27480 7064 27532
rect 6552 27344 6604 27396
rect 5908 27276 5960 27328
rect 7840 27276 7892 27328
rect 3547 27174 3599 27226
rect 3611 27174 3663 27226
rect 3675 27174 3727 27226
rect 3739 27174 3791 27226
rect 3803 27174 3855 27226
rect 6144 27174 6196 27226
rect 6208 27174 6260 27226
rect 6272 27174 6324 27226
rect 6336 27174 6388 27226
rect 6400 27174 6452 27226
rect 6552 27115 6604 27124
rect 6552 27081 6561 27115
rect 6561 27081 6595 27115
rect 6595 27081 6604 27115
rect 6552 27072 6604 27081
rect 5908 27004 5960 27056
rect 6368 26979 6420 26988
rect 6368 26945 6377 26979
rect 6377 26945 6411 26979
rect 6411 26945 6420 26979
rect 6368 26936 6420 26945
rect 8116 26936 8168 26988
rect 5264 26868 5316 26920
rect 7104 26843 7156 26852
rect 7104 26809 7113 26843
rect 7113 26809 7147 26843
rect 7147 26809 7156 26843
rect 7104 26800 7156 26809
rect 2248 26630 2300 26682
rect 2312 26630 2364 26682
rect 2376 26630 2428 26682
rect 2440 26630 2492 26682
rect 2504 26630 2556 26682
rect 4846 26630 4898 26682
rect 4910 26630 4962 26682
rect 4974 26630 5026 26682
rect 5038 26630 5090 26682
rect 5102 26630 5154 26682
rect 7443 26630 7495 26682
rect 7507 26630 7559 26682
rect 7571 26630 7623 26682
rect 7635 26630 7687 26682
rect 7699 26630 7751 26682
rect 5264 26571 5316 26580
rect 5264 26537 5273 26571
rect 5273 26537 5307 26571
rect 5307 26537 5316 26571
rect 5264 26528 5316 26537
rect 7104 26460 7156 26512
rect 8024 26460 8076 26512
rect 7012 26392 7064 26444
rect 6368 26324 6420 26376
rect 6828 26367 6880 26376
rect 6828 26333 6837 26367
rect 6837 26333 6871 26367
rect 6871 26333 6880 26367
rect 6828 26324 6880 26333
rect 8116 26367 8168 26376
rect 8116 26333 8125 26367
rect 8125 26333 8159 26367
rect 8159 26333 8168 26367
rect 8116 26324 8168 26333
rect 6920 26188 6972 26240
rect 3547 26086 3599 26138
rect 3611 26086 3663 26138
rect 3675 26086 3727 26138
rect 3739 26086 3791 26138
rect 3803 26086 3855 26138
rect 6144 26086 6196 26138
rect 6208 26086 6260 26138
rect 6272 26086 6324 26138
rect 6336 26086 6388 26138
rect 6400 26086 6452 26138
rect 6828 25959 6880 25968
rect 6828 25925 6837 25959
rect 6837 25925 6871 25959
rect 6871 25925 6880 25959
rect 6828 25916 6880 25925
rect 7104 25959 7156 25968
rect 7104 25925 7113 25959
rect 7113 25925 7147 25959
rect 7147 25925 7156 25959
rect 7104 25916 7156 25925
rect 7840 25848 7892 25900
rect 2248 25542 2300 25594
rect 2312 25542 2364 25594
rect 2376 25542 2428 25594
rect 2440 25542 2492 25594
rect 2504 25542 2556 25594
rect 4846 25542 4898 25594
rect 4910 25542 4962 25594
rect 4974 25542 5026 25594
rect 5038 25542 5090 25594
rect 5102 25542 5154 25594
rect 7443 25542 7495 25594
rect 7507 25542 7559 25594
rect 7571 25542 7623 25594
rect 7635 25542 7687 25594
rect 7699 25542 7751 25594
rect 6920 25372 6972 25424
rect 7656 25372 7708 25424
rect 7196 25279 7248 25288
rect 7196 25245 7205 25279
rect 7205 25245 7239 25279
rect 7239 25245 7248 25279
rect 7196 25236 7248 25245
rect 6644 25100 6696 25152
rect 3547 24998 3599 25050
rect 3611 24998 3663 25050
rect 3675 24998 3727 25050
rect 3739 24998 3791 25050
rect 3803 24998 3855 25050
rect 6144 24998 6196 25050
rect 6208 24998 6260 25050
rect 6272 24998 6324 25050
rect 6336 24998 6388 25050
rect 6400 24998 6452 25050
rect 7656 24871 7708 24880
rect 7656 24837 7665 24871
rect 7665 24837 7699 24871
rect 7699 24837 7708 24871
rect 7656 24828 7708 24837
rect 7104 24803 7156 24812
rect 7104 24769 7113 24803
rect 7113 24769 7147 24803
rect 7147 24769 7156 24803
rect 7104 24760 7156 24769
rect 6644 24556 6696 24608
rect 2248 24454 2300 24506
rect 2312 24454 2364 24506
rect 2376 24454 2428 24506
rect 2440 24454 2492 24506
rect 2504 24454 2556 24506
rect 4846 24454 4898 24506
rect 4910 24454 4962 24506
rect 4974 24454 5026 24506
rect 5038 24454 5090 24506
rect 5102 24454 5154 24506
rect 7443 24454 7495 24506
rect 7507 24454 7559 24506
rect 7571 24454 7623 24506
rect 7635 24454 7687 24506
rect 7699 24454 7751 24506
rect 5816 24216 5868 24268
rect 7104 24148 7156 24200
rect 8116 24191 8168 24200
rect 8116 24157 8125 24191
rect 8125 24157 8159 24191
rect 8159 24157 8168 24191
rect 8116 24148 8168 24157
rect 7196 24123 7248 24132
rect 7196 24089 7205 24123
rect 7205 24089 7239 24123
rect 7239 24089 7248 24123
rect 7196 24080 7248 24089
rect 7564 24012 7616 24064
rect 3547 23910 3599 23962
rect 3611 23910 3663 23962
rect 3675 23910 3727 23962
rect 3739 23910 3791 23962
rect 3803 23910 3855 23962
rect 6144 23910 6196 23962
rect 6208 23910 6260 23962
rect 6272 23910 6324 23962
rect 6336 23910 6388 23962
rect 6400 23910 6452 23962
rect 5816 23851 5868 23860
rect 5816 23817 5825 23851
rect 5825 23817 5859 23851
rect 5859 23817 5868 23851
rect 5816 23808 5868 23817
rect 7196 23808 7248 23860
rect 7564 23783 7616 23792
rect 7564 23749 7573 23783
rect 7573 23749 7607 23783
rect 7607 23749 7616 23783
rect 7564 23740 7616 23749
rect 6552 23672 6604 23724
rect 7104 23672 7156 23724
rect 8116 23715 8168 23724
rect 8116 23681 8125 23715
rect 8125 23681 8159 23715
rect 8159 23681 8168 23715
rect 8116 23672 8168 23681
rect 2248 23366 2300 23418
rect 2312 23366 2364 23418
rect 2376 23366 2428 23418
rect 2440 23366 2492 23418
rect 2504 23366 2556 23418
rect 4846 23366 4898 23418
rect 4910 23366 4962 23418
rect 4974 23366 5026 23418
rect 5038 23366 5090 23418
rect 5102 23366 5154 23418
rect 7443 23366 7495 23418
rect 7507 23366 7559 23418
rect 7571 23366 7623 23418
rect 7635 23366 7687 23418
rect 7699 23366 7751 23418
rect 6736 23196 6788 23248
rect 7564 23060 7616 23112
rect 6920 23035 6972 23044
rect 6920 23001 6929 23035
rect 6929 23001 6963 23035
rect 6963 23001 6972 23035
rect 6920 22992 6972 23001
rect 6828 22924 6880 22976
rect 3547 22822 3599 22874
rect 3611 22822 3663 22874
rect 3675 22822 3727 22874
rect 3739 22822 3791 22874
rect 3803 22822 3855 22874
rect 6144 22822 6196 22874
rect 6208 22822 6260 22874
rect 6272 22822 6324 22874
rect 6336 22822 6388 22874
rect 6400 22822 6452 22874
rect 6828 22695 6880 22704
rect 6828 22661 6837 22695
rect 6837 22661 6871 22695
rect 6871 22661 6880 22695
rect 6828 22652 6880 22661
rect 6920 22695 6972 22704
rect 6920 22661 6929 22695
rect 6929 22661 6963 22695
rect 6963 22661 6972 22695
rect 6920 22652 6972 22661
rect 7564 22652 7616 22704
rect 7840 22695 7892 22704
rect 7840 22661 7849 22695
rect 7849 22661 7883 22695
rect 7883 22661 7892 22695
rect 7840 22652 7892 22661
rect 8024 22695 8076 22704
rect 8024 22661 8033 22695
rect 8033 22661 8067 22695
rect 8067 22661 8076 22695
rect 8024 22652 8076 22661
rect 6736 22516 6788 22568
rect 5724 22423 5776 22432
rect 5724 22389 5733 22423
rect 5733 22389 5767 22423
rect 5767 22389 5776 22423
rect 5724 22380 5776 22389
rect 2248 22278 2300 22330
rect 2312 22278 2364 22330
rect 2376 22278 2428 22330
rect 2440 22278 2492 22330
rect 2504 22278 2556 22330
rect 4846 22278 4898 22330
rect 4910 22278 4962 22330
rect 4974 22278 5026 22330
rect 5038 22278 5090 22330
rect 5102 22278 5154 22330
rect 7443 22278 7495 22330
rect 7507 22278 7559 22330
rect 7571 22278 7623 22330
rect 7635 22278 7687 22330
rect 7699 22278 7751 22330
rect 7840 22015 7892 22024
rect 7840 21981 7849 22015
rect 7849 21981 7883 22015
rect 7883 21981 7892 22015
rect 7840 21972 7892 21981
rect 7932 21947 7984 21956
rect 7932 21913 7941 21947
rect 7941 21913 7975 21947
rect 7975 21913 7984 21947
rect 7932 21904 7984 21913
rect 6000 21836 6052 21888
rect 3547 21734 3599 21786
rect 3611 21734 3663 21786
rect 3675 21734 3727 21786
rect 3739 21734 3791 21786
rect 3803 21734 3855 21786
rect 6144 21734 6196 21786
rect 6208 21734 6260 21786
rect 6272 21734 6324 21786
rect 6336 21734 6388 21786
rect 6400 21734 6452 21786
rect 5724 21564 5776 21616
rect 7932 21607 7984 21616
rect 7932 21573 7941 21607
rect 7941 21573 7975 21607
rect 7975 21573 7984 21607
rect 7932 21564 7984 21573
rect 5632 21539 5684 21548
rect 5632 21505 5641 21539
rect 5641 21505 5675 21539
rect 5675 21505 5684 21539
rect 5632 21496 5684 21505
rect 6000 21428 6052 21480
rect 8116 21403 8168 21412
rect 8116 21369 8125 21403
rect 8125 21369 8159 21403
rect 8159 21369 8168 21403
rect 8116 21360 8168 21369
rect 5172 21335 5224 21344
rect 5172 21301 5181 21335
rect 5181 21301 5215 21335
rect 5215 21301 5224 21335
rect 5172 21292 5224 21301
rect 6184 21292 6236 21344
rect 2248 21190 2300 21242
rect 2312 21190 2364 21242
rect 2376 21190 2428 21242
rect 2440 21190 2492 21242
rect 2504 21190 2556 21242
rect 4846 21190 4898 21242
rect 4910 21190 4962 21242
rect 4974 21190 5026 21242
rect 5038 21190 5090 21242
rect 5102 21190 5154 21242
rect 7443 21190 7495 21242
rect 7507 21190 7559 21242
rect 7571 21190 7623 21242
rect 7635 21190 7687 21242
rect 7699 21190 7751 21242
rect 6552 21020 6604 21072
rect 6184 20995 6236 21004
rect 6184 20961 6193 20995
rect 6193 20961 6227 20995
rect 6227 20961 6236 20995
rect 6184 20952 6236 20961
rect 5172 20927 5224 20936
rect 5172 20893 5181 20927
rect 5181 20893 5215 20927
rect 5215 20893 5224 20927
rect 5172 20884 5224 20893
rect 6644 20884 6696 20936
rect 8208 20884 8260 20936
rect 5632 20859 5684 20868
rect 5632 20825 5641 20859
rect 5641 20825 5675 20859
rect 5675 20825 5684 20859
rect 5632 20816 5684 20825
rect 5724 20859 5776 20868
rect 5724 20825 5733 20859
rect 5733 20825 5767 20859
rect 5767 20825 5776 20859
rect 7196 20859 7248 20868
rect 5724 20816 5776 20825
rect 7196 20825 7205 20859
rect 7205 20825 7239 20859
rect 7239 20825 7248 20859
rect 7196 20816 7248 20825
rect 5264 20748 5316 20800
rect 3547 20646 3599 20698
rect 3611 20646 3663 20698
rect 3675 20646 3727 20698
rect 3739 20646 3791 20698
rect 3803 20646 3855 20698
rect 6144 20646 6196 20698
rect 6208 20646 6260 20698
rect 6272 20646 6324 20698
rect 6336 20646 6388 20698
rect 6400 20646 6452 20698
rect 5172 20587 5224 20596
rect 5172 20553 5181 20587
rect 5181 20553 5215 20587
rect 5215 20553 5224 20587
rect 5172 20544 5224 20553
rect 5724 20544 5776 20596
rect 6552 20519 6604 20528
rect 6552 20485 6561 20519
rect 6561 20485 6595 20519
rect 6595 20485 6604 20519
rect 6552 20476 6604 20485
rect 6644 20476 6696 20528
rect 7196 20451 7248 20460
rect 7196 20417 7205 20451
rect 7205 20417 7239 20451
rect 7239 20417 7248 20451
rect 7196 20408 7248 20417
rect 8024 20408 8076 20460
rect 2248 20102 2300 20154
rect 2312 20102 2364 20154
rect 2376 20102 2428 20154
rect 2440 20102 2492 20154
rect 2504 20102 2556 20154
rect 4846 20102 4898 20154
rect 4910 20102 4962 20154
rect 4974 20102 5026 20154
rect 5038 20102 5090 20154
rect 5102 20102 5154 20154
rect 7443 20102 7495 20154
rect 7507 20102 7559 20154
rect 7571 20102 7623 20154
rect 7635 20102 7687 20154
rect 7699 20102 7751 20154
rect 5540 20000 5592 20052
rect 6736 19796 6788 19848
rect 8116 19839 8168 19848
rect 8116 19805 8125 19839
rect 8125 19805 8159 19839
rect 8159 19805 8168 19839
rect 8116 19796 8168 19805
rect 7196 19771 7248 19780
rect 7196 19737 7205 19771
rect 7205 19737 7239 19771
rect 7239 19737 7248 19771
rect 7196 19728 7248 19737
rect 5264 19660 5316 19712
rect 6644 19660 6696 19712
rect 7288 19660 7340 19712
rect 3547 19558 3599 19610
rect 3611 19558 3663 19610
rect 3675 19558 3727 19610
rect 3739 19558 3791 19610
rect 3803 19558 3855 19610
rect 6144 19558 6196 19610
rect 6208 19558 6260 19610
rect 6272 19558 6324 19610
rect 6336 19558 6388 19610
rect 6400 19558 6452 19610
rect 8024 19499 8076 19508
rect 8024 19465 8033 19499
rect 8033 19465 8067 19499
rect 8067 19465 8076 19499
rect 8024 19456 8076 19465
rect 7196 19431 7248 19440
rect 7196 19397 7205 19431
rect 7205 19397 7239 19431
rect 7239 19397 7248 19431
rect 7196 19388 7248 19397
rect 7288 19431 7340 19440
rect 7288 19397 7297 19431
rect 7297 19397 7331 19431
rect 7331 19397 7340 19431
rect 7288 19388 7340 19397
rect 6552 19320 6604 19372
rect 6736 19295 6788 19304
rect 6736 19261 6745 19295
rect 6745 19261 6779 19295
rect 6779 19261 6788 19295
rect 6736 19252 6788 19261
rect 5632 19116 5684 19168
rect 6828 19116 6880 19168
rect 2248 19014 2300 19066
rect 2312 19014 2364 19066
rect 2376 19014 2428 19066
rect 2440 19014 2492 19066
rect 2504 19014 2556 19066
rect 4846 19014 4898 19066
rect 4910 19014 4962 19066
rect 4974 19014 5026 19066
rect 5038 19014 5090 19066
rect 5102 19014 5154 19066
rect 7443 19014 7495 19066
rect 7507 19014 7559 19066
rect 7571 19014 7623 19066
rect 7635 19014 7687 19066
rect 7699 19014 7751 19066
rect 6736 18955 6788 18964
rect 6736 18921 6745 18955
rect 6745 18921 6779 18955
rect 6779 18921 6788 18955
rect 6736 18912 6788 18921
rect 7196 18751 7248 18760
rect 7196 18717 7205 18751
rect 7205 18717 7239 18751
rect 7239 18717 7248 18751
rect 7196 18708 7248 18717
rect 6736 18640 6788 18692
rect 7288 18615 7340 18624
rect 7288 18581 7297 18615
rect 7297 18581 7331 18615
rect 7331 18581 7340 18615
rect 7288 18572 7340 18581
rect 3547 18470 3599 18522
rect 3611 18470 3663 18522
rect 3675 18470 3727 18522
rect 3739 18470 3791 18522
rect 3803 18470 3855 18522
rect 6144 18470 6196 18522
rect 6208 18470 6260 18522
rect 6272 18470 6324 18522
rect 6336 18470 6388 18522
rect 6400 18470 6452 18522
rect 5724 18232 5776 18284
rect 6736 18232 6788 18284
rect 8116 18232 8168 18284
rect 7840 18139 7892 18148
rect 7840 18105 7849 18139
rect 7849 18105 7883 18139
rect 7883 18105 7892 18139
rect 7840 18096 7892 18105
rect 5724 18071 5776 18080
rect 5724 18037 5733 18071
rect 5733 18037 5767 18071
rect 5767 18037 5776 18071
rect 5724 18028 5776 18037
rect 2248 17926 2300 17978
rect 2312 17926 2364 17978
rect 2376 17926 2428 17978
rect 2440 17926 2492 17978
rect 2504 17926 2556 17978
rect 4846 17926 4898 17978
rect 4910 17926 4962 17978
rect 4974 17926 5026 17978
rect 5038 17926 5090 17978
rect 5102 17926 5154 17978
rect 7443 17926 7495 17978
rect 7507 17926 7559 17978
rect 7571 17926 7623 17978
rect 7635 17926 7687 17978
rect 7699 17926 7751 17978
rect 5540 17688 5592 17740
rect 5816 17731 5868 17740
rect 5816 17697 5825 17731
rect 5825 17697 5859 17731
rect 5859 17697 5868 17731
rect 5816 17688 5868 17697
rect 7104 17688 7156 17740
rect 7288 17688 7340 17740
rect 5724 17552 5776 17604
rect 7196 17620 7248 17672
rect 6920 17552 6972 17604
rect 7840 17552 7892 17604
rect 3547 17382 3599 17434
rect 3611 17382 3663 17434
rect 3675 17382 3727 17434
rect 3739 17382 3791 17434
rect 3803 17382 3855 17434
rect 6144 17382 6196 17434
rect 6208 17382 6260 17434
rect 6272 17382 6324 17434
rect 6336 17382 6388 17434
rect 6400 17382 6452 17434
rect 5908 17280 5960 17332
rect 6644 17280 6696 17332
rect 6552 17255 6604 17264
rect 6552 17221 6561 17255
rect 6561 17221 6595 17255
rect 6595 17221 6604 17255
rect 6552 17212 6604 17221
rect 7196 17187 7248 17196
rect 7196 17153 7205 17187
rect 7205 17153 7239 17187
rect 7239 17153 7248 17187
rect 7196 17144 7248 17153
rect 5816 16983 5868 16992
rect 5816 16949 5825 16983
rect 5825 16949 5859 16983
rect 5859 16949 5868 16983
rect 5816 16940 5868 16949
rect 2248 16838 2300 16890
rect 2312 16838 2364 16890
rect 2376 16838 2428 16890
rect 2440 16838 2492 16890
rect 2504 16838 2556 16890
rect 4846 16838 4898 16890
rect 4910 16838 4962 16890
rect 4974 16838 5026 16890
rect 5038 16838 5090 16890
rect 5102 16838 5154 16890
rect 7443 16838 7495 16890
rect 7507 16838 7559 16890
rect 7571 16838 7623 16890
rect 7635 16838 7687 16890
rect 7699 16838 7751 16890
rect 5540 16736 5592 16788
rect 6552 16668 6604 16720
rect 5816 16600 5868 16652
rect 7104 16532 7156 16584
rect 6736 16507 6788 16516
rect 6736 16473 6745 16507
rect 6745 16473 6779 16507
rect 6779 16473 6788 16507
rect 7196 16507 7248 16516
rect 6736 16464 6788 16473
rect 7196 16473 7205 16507
rect 7205 16473 7239 16507
rect 7239 16473 7248 16507
rect 7196 16464 7248 16473
rect 6552 16396 6604 16448
rect 3547 16294 3599 16346
rect 3611 16294 3663 16346
rect 3675 16294 3727 16346
rect 3739 16294 3791 16346
rect 3803 16294 3855 16346
rect 6144 16294 6196 16346
rect 6208 16294 6260 16346
rect 6272 16294 6324 16346
rect 6336 16294 6388 16346
rect 6400 16294 6452 16346
rect 6736 16192 6788 16244
rect 6920 16124 6972 16176
rect 7104 16124 7156 16176
rect 6736 16099 6788 16108
rect 6736 16065 6745 16099
rect 6745 16065 6779 16099
rect 6779 16065 6788 16099
rect 6736 16056 6788 16065
rect 7012 16056 7064 16108
rect 7840 16056 7892 16108
rect 5172 16031 5224 16040
rect 5172 15997 5181 16031
rect 5181 15997 5215 16031
rect 5215 15997 5224 16031
rect 5172 15988 5224 15997
rect 6460 15852 6512 15904
rect 2248 15750 2300 15802
rect 2312 15750 2364 15802
rect 2376 15750 2428 15802
rect 2440 15750 2492 15802
rect 2504 15750 2556 15802
rect 4846 15750 4898 15802
rect 4910 15750 4962 15802
rect 4974 15750 5026 15802
rect 5038 15750 5090 15802
rect 5102 15750 5154 15802
rect 7443 15750 7495 15802
rect 7507 15750 7559 15802
rect 7571 15750 7623 15802
rect 7635 15750 7687 15802
rect 7699 15750 7751 15802
rect 5172 15648 5224 15700
rect 5356 15648 5408 15700
rect 5356 15555 5408 15564
rect 5356 15521 5365 15555
rect 5365 15521 5399 15555
rect 5399 15521 5408 15555
rect 5356 15512 5408 15521
rect 6460 15555 6512 15564
rect 6460 15521 6469 15555
rect 6469 15521 6503 15555
rect 6503 15521 6512 15555
rect 6460 15512 6512 15521
rect 6736 15580 6788 15632
rect 7012 15555 7064 15564
rect 7012 15521 7021 15555
rect 7021 15521 7055 15555
rect 7055 15521 7064 15555
rect 7012 15512 7064 15521
rect 8116 15512 8168 15564
rect 7288 15444 7340 15496
rect 5816 15419 5868 15428
rect 5816 15385 5825 15419
rect 5825 15385 5859 15419
rect 5859 15385 5868 15419
rect 5816 15376 5868 15385
rect 7104 15376 7156 15428
rect 3547 15206 3599 15258
rect 3611 15206 3663 15258
rect 3675 15206 3727 15258
rect 3739 15206 3791 15258
rect 3803 15206 3855 15258
rect 6144 15206 6196 15258
rect 6208 15206 6260 15258
rect 6272 15206 6324 15258
rect 6336 15206 6388 15258
rect 6400 15206 6452 15258
rect 5356 15104 5408 15156
rect 7196 15104 7248 15156
rect 7840 15036 7892 15088
rect 6736 15011 6788 15020
rect 6736 14977 6745 15011
rect 6745 14977 6779 15011
rect 6779 14977 6788 15011
rect 6736 14968 6788 14977
rect 7012 14968 7064 15020
rect 7288 14968 7340 15020
rect 8116 15011 8168 15020
rect 8116 14977 8125 15011
rect 8125 14977 8159 15011
rect 8159 14977 8168 15011
rect 8116 14968 8168 14977
rect 5540 14832 5592 14884
rect 6552 14832 6604 14884
rect 6092 14764 6144 14816
rect 2248 14662 2300 14714
rect 2312 14662 2364 14714
rect 2376 14662 2428 14714
rect 2440 14662 2492 14714
rect 2504 14662 2556 14714
rect 4846 14662 4898 14714
rect 4910 14662 4962 14714
rect 4974 14662 5026 14714
rect 5038 14662 5090 14714
rect 5102 14662 5154 14714
rect 7443 14662 7495 14714
rect 7507 14662 7559 14714
rect 7571 14662 7623 14714
rect 7635 14662 7687 14714
rect 7699 14662 7751 14714
rect 7196 14492 7248 14544
rect 5816 14424 5868 14476
rect 5540 14356 5592 14408
rect 6736 14424 6788 14476
rect 6092 14399 6144 14408
rect 6092 14365 6101 14399
rect 6101 14365 6135 14399
rect 6135 14365 6144 14399
rect 6092 14356 6144 14365
rect 6920 14356 6972 14408
rect 6460 14288 6512 14340
rect 6736 14288 6788 14340
rect 3547 14118 3599 14170
rect 3611 14118 3663 14170
rect 3675 14118 3727 14170
rect 3739 14118 3791 14170
rect 3803 14118 3855 14170
rect 6144 14118 6196 14170
rect 6208 14118 6260 14170
rect 6272 14118 6324 14170
rect 6336 14118 6388 14170
rect 6400 14118 6452 14170
rect 6000 13880 6052 13932
rect 7012 13880 7064 13932
rect 7840 13787 7892 13796
rect 7840 13753 7849 13787
rect 7849 13753 7883 13787
rect 7883 13753 7892 13787
rect 7840 13744 7892 13753
rect 6000 13676 6052 13728
rect 2248 13574 2300 13626
rect 2312 13574 2364 13626
rect 2376 13574 2428 13626
rect 2440 13574 2492 13626
rect 2504 13574 2556 13626
rect 4846 13574 4898 13626
rect 4910 13574 4962 13626
rect 4974 13574 5026 13626
rect 5038 13574 5090 13626
rect 5102 13574 5154 13626
rect 7443 13574 7495 13626
rect 7507 13574 7559 13626
rect 7571 13574 7623 13626
rect 7635 13574 7687 13626
rect 7699 13574 7751 13626
rect 5540 13472 5592 13524
rect 7104 13515 7156 13524
rect 7104 13481 7113 13515
rect 7113 13481 7147 13515
rect 7147 13481 7156 13515
rect 7104 13472 7156 13481
rect 7840 13404 7892 13456
rect 7012 13268 7064 13320
rect 7288 13200 7340 13252
rect 6000 13132 6052 13184
rect 3547 13030 3599 13082
rect 3611 13030 3663 13082
rect 3675 13030 3727 13082
rect 3739 13030 3791 13082
rect 3803 13030 3855 13082
rect 6144 13030 6196 13082
rect 6208 13030 6260 13082
rect 6272 13030 6324 13082
rect 6336 13030 6388 13082
rect 6400 13030 6452 13082
rect 6828 12928 6880 12980
rect 7288 12971 7340 12980
rect 7288 12937 7297 12971
rect 7297 12937 7331 12971
rect 7331 12937 7340 12971
rect 7288 12928 7340 12937
rect 7380 12971 7432 12980
rect 7380 12937 7389 12971
rect 7389 12937 7423 12971
rect 7423 12937 7432 12971
rect 7380 12928 7432 12937
rect 8208 12860 8260 12912
rect 5540 12792 5592 12844
rect 6184 12792 6236 12844
rect 7196 12792 7248 12844
rect 6736 12767 6788 12776
rect 6736 12733 6745 12767
rect 6745 12733 6779 12767
rect 6779 12733 6788 12767
rect 6736 12724 6788 12733
rect 7840 12631 7892 12640
rect 7840 12597 7849 12631
rect 7849 12597 7883 12631
rect 7883 12597 7892 12631
rect 7840 12588 7892 12597
rect 2248 12486 2300 12538
rect 2312 12486 2364 12538
rect 2376 12486 2428 12538
rect 2440 12486 2492 12538
rect 2504 12486 2556 12538
rect 4846 12486 4898 12538
rect 4910 12486 4962 12538
rect 4974 12486 5026 12538
rect 5038 12486 5090 12538
rect 5102 12486 5154 12538
rect 7443 12486 7495 12538
rect 7507 12486 7559 12538
rect 7571 12486 7623 12538
rect 7635 12486 7687 12538
rect 7699 12486 7751 12538
rect 5264 12384 5316 12436
rect 5724 12384 5776 12436
rect 6736 12359 6788 12368
rect 6736 12325 6745 12359
rect 6745 12325 6779 12359
rect 6779 12325 6788 12359
rect 6736 12316 6788 12325
rect 6552 12248 6604 12300
rect 7840 12248 7892 12300
rect 5540 12180 5592 12232
rect 5816 12180 5868 12232
rect 5908 12180 5960 12232
rect 6184 12112 6236 12164
rect 7288 12112 7340 12164
rect 5816 12087 5868 12096
rect 5816 12053 5825 12087
rect 5825 12053 5859 12087
rect 5859 12053 5868 12087
rect 5816 12044 5868 12053
rect 6920 12044 6972 12096
rect 7104 12044 7156 12096
rect 3547 11942 3599 11994
rect 3611 11942 3663 11994
rect 3675 11942 3727 11994
rect 3739 11942 3791 11994
rect 3803 11942 3855 11994
rect 6144 11942 6196 11994
rect 6208 11942 6260 11994
rect 6272 11942 6324 11994
rect 6336 11942 6388 11994
rect 6400 11942 6452 11994
rect 7012 11815 7064 11824
rect 7012 11781 7021 11815
rect 7021 11781 7055 11815
rect 7055 11781 7064 11815
rect 7012 11772 7064 11781
rect 6828 11747 6880 11756
rect 6828 11713 6837 11747
rect 6837 11713 6871 11747
rect 6871 11713 6880 11747
rect 6828 11704 6880 11713
rect 6000 11636 6052 11688
rect 8300 11636 8352 11688
rect 5540 11500 5592 11552
rect 2248 11398 2300 11450
rect 2312 11398 2364 11450
rect 2376 11398 2428 11450
rect 2440 11398 2492 11450
rect 2504 11398 2556 11450
rect 4846 11398 4898 11450
rect 4910 11398 4962 11450
rect 4974 11398 5026 11450
rect 5038 11398 5090 11450
rect 5102 11398 5154 11450
rect 7443 11398 7495 11450
rect 7507 11398 7559 11450
rect 7571 11398 7623 11450
rect 7635 11398 7687 11450
rect 7699 11398 7751 11450
rect 5540 11296 5592 11348
rect 6000 11339 6052 11348
rect 6000 11305 6009 11339
rect 6009 11305 6043 11339
rect 6043 11305 6052 11339
rect 6000 11296 6052 11305
rect 6828 11271 6880 11280
rect 6828 11237 6837 11271
rect 6837 11237 6871 11271
rect 6871 11237 6880 11271
rect 6828 11228 6880 11237
rect 7196 11135 7248 11144
rect 7196 11101 7205 11135
rect 7205 11101 7239 11135
rect 7239 11101 7248 11135
rect 7196 11092 7248 11101
rect 8300 11092 8352 11144
rect 7288 11024 7340 11076
rect 3547 10854 3599 10906
rect 3611 10854 3663 10906
rect 3675 10854 3727 10906
rect 3739 10854 3791 10906
rect 3803 10854 3855 10906
rect 6144 10854 6196 10906
rect 6208 10854 6260 10906
rect 6272 10854 6324 10906
rect 6336 10854 6388 10906
rect 6400 10854 6452 10906
rect 6644 10752 6696 10804
rect 7932 10752 7984 10804
rect 7288 10727 7340 10736
rect 7288 10693 7297 10727
rect 7297 10693 7331 10727
rect 7331 10693 7340 10727
rect 7288 10684 7340 10693
rect 6552 10616 6604 10668
rect 7196 10616 7248 10668
rect 5816 10591 5868 10600
rect 5816 10557 5825 10591
rect 5825 10557 5859 10591
rect 5859 10557 5868 10591
rect 5816 10548 5868 10557
rect 2248 10310 2300 10362
rect 2312 10310 2364 10362
rect 2376 10310 2428 10362
rect 2440 10310 2492 10362
rect 2504 10310 2556 10362
rect 4846 10310 4898 10362
rect 4910 10310 4962 10362
rect 4974 10310 5026 10362
rect 5038 10310 5090 10362
rect 5102 10310 5154 10362
rect 7443 10310 7495 10362
rect 7507 10310 7559 10362
rect 7571 10310 7623 10362
rect 7635 10310 7687 10362
rect 7699 10310 7751 10362
rect 5540 10072 5592 10124
rect 7288 10004 7340 10056
rect 6920 9979 6972 9988
rect 6920 9945 6929 9979
rect 6929 9945 6963 9979
rect 6963 9945 6972 9979
rect 6920 9936 6972 9945
rect 8208 10004 8260 10056
rect 5448 9868 5500 9920
rect 5632 9868 5684 9920
rect 7932 9868 7984 9920
rect 3547 9766 3599 9818
rect 3611 9766 3663 9818
rect 3675 9766 3727 9818
rect 3739 9766 3791 9818
rect 3803 9766 3855 9818
rect 6144 9766 6196 9818
rect 6208 9766 6260 9818
rect 6272 9766 6324 9818
rect 6336 9766 6388 9818
rect 6400 9766 6452 9818
rect 5816 9571 5868 9580
rect 5816 9537 5825 9571
rect 5825 9537 5859 9571
rect 5859 9537 5868 9571
rect 5816 9528 5868 9537
rect 6644 9528 6696 9580
rect 7104 9571 7156 9580
rect 7104 9537 7113 9571
rect 7113 9537 7147 9571
rect 7147 9537 7156 9571
rect 7104 9528 7156 9537
rect 7840 9528 7892 9580
rect 7196 9324 7248 9376
rect 2248 9222 2300 9274
rect 2312 9222 2364 9274
rect 2376 9222 2428 9274
rect 2440 9222 2492 9274
rect 2504 9222 2556 9274
rect 4846 9222 4898 9274
rect 4910 9222 4962 9274
rect 4974 9222 5026 9274
rect 5038 9222 5090 9274
rect 5102 9222 5154 9274
rect 7443 9222 7495 9274
rect 7507 9222 7559 9274
rect 7571 9222 7623 9274
rect 7635 9222 7687 9274
rect 7699 9222 7751 9274
rect 5816 9120 5868 9172
rect 7104 9095 7156 9104
rect 7104 9061 7113 9095
rect 7113 9061 7147 9095
rect 7147 9061 7156 9095
rect 7104 9052 7156 9061
rect 6644 9027 6696 9036
rect 6644 8993 6653 9027
rect 6653 8993 6687 9027
rect 6687 8993 6696 9027
rect 6644 8984 6696 8993
rect 7196 9027 7248 9036
rect 7196 8993 7205 9027
rect 7205 8993 7239 9027
rect 7239 8993 7248 9027
rect 7196 8984 7248 8993
rect 7104 8848 7156 8900
rect 5816 8780 5868 8832
rect 6828 8780 6880 8832
rect 7840 8823 7892 8832
rect 7840 8789 7849 8823
rect 7849 8789 7883 8823
rect 7883 8789 7892 8823
rect 7840 8780 7892 8789
rect 3547 8678 3599 8730
rect 3611 8678 3663 8730
rect 3675 8678 3727 8730
rect 3739 8678 3791 8730
rect 3803 8678 3855 8730
rect 6144 8678 6196 8730
rect 6208 8678 6260 8730
rect 6272 8678 6324 8730
rect 6336 8678 6388 8730
rect 6400 8678 6452 8730
rect 5540 8576 5592 8628
rect 6920 8508 6972 8560
rect 7196 8483 7248 8492
rect 7196 8449 7205 8483
rect 7205 8449 7239 8483
rect 7239 8449 7248 8483
rect 7196 8440 7248 8449
rect 6552 8415 6604 8424
rect 6552 8381 6561 8415
rect 6561 8381 6595 8415
rect 6595 8381 6604 8415
rect 6552 8372 6604 8381
rect 5816 8304 5868 8356
rect 6460 8304 6512 8356
rect 2248 8134 2300 8186
rect 2312 8134 2364 8186
rect 2376 8134 2428 8186
rect 2440 8134 2492 8186
rect 2504 8134 2556 8186
rect 4846 8134 4898 8186
rect 4910 8134 4962 8186
rect 4974 8134 5026 8186
rect 5038 8134 5090 8186
rect 5102 8134 5154 8186
rect 7443 8134 7495 8186
rect 7507 8134 7559 8186
rect 7571 8134 7623 8186
rect 7635 8134 7687 8186
rect 7699 8134 7751 8186
rect 5908 8032 5960 8084
rect 5540 8007 5592 8016
rect 5540 7973 5549 8007
rect 5549 7973 5583 8007
rect 5583 7973 5592 8007
rect 5540 7964 5592 7973
rect 7932 7896 7984 7948
rect 5724 7871 5776 7880
rect 5724 7837 5733 7871
rect 5733 7837 5767 7871
rect 5767 7837 5776 7871
rect 5724 7828 5776 7837
rect 7288 7828 7340 7880
rect 5632 7760 5684 7812
rect 7196 7803 7248 7812
rect 7196 7769 7205 7803
rect 7205 7769 7239 7803
rect 7239 7769 7248 7803
rect 7196 7760 7248 7769
rect 7288 7692 7340 7744
rect 3547 7590 3599 7642
rect 3611 7590 3663 7642
rect 3675 7590 3727 7642
rect 3739 7590 3791 7642
rect 3803 7590 3855 7642
rect 6144 7590 6196 7642
rect 6208 7590 6260 7642
rect 6272 7590 6324 7642
rect 6336 7590 6388 7642
rect 6400 7590 6452 7642
rect 5724 7531 5776 7540
rect 5724 7497 5733 7531
rect 5733 7497 5767 7531
rect 5767 7497 5776 7531
rect 5724 7488 5776 7497
rect 7104 7420 7156 7472
rect 7840 7395 7892 7404
rect 7840 7361 7849 7395
rect 7849 7361 7883 7395
rect 7883 7361 7892 7395
rect 7840 7352 7892 7361
rect 7932 7284 7984 7336
rect 7840 7259 7892 7268
rect 7840 7225 7849 7259
rect 7849 7225 7883 7259
rect 7883 7225 7892 7259
rect 7840 7216 7892 7225
rect 5632 7148 5684 7200
rect 6460 7148 6512 7200
rect 2248 7046 2300 7098
rect 2312 7046 2364 7098
rect 2376 7046 2428 7098
rect 2440 7046 2492 7098
rect 2504 7046 2556 7098
rect 4846 7046 4898 7098
rect 4910 7046 4962 7098
rect 4974 7046 5026 7098
rect 5038 7046 5090 7098
rect 5102 7046 5154 7098
rect 7443 7046 7495 7098
rect 7507 7046 7559 7098
rect 7571 7046 7623 7098
rect 7635 7046 7687 7098
rect 7699 7046 7751 7098
rect 5448 6808 5500 6860
rect 6828 6808 6880 6860
rect 4436 6783 4488 6792
rect 4436 6749 4445 6783
rect 4445 6749 4479 6783
rect 4479 6749 4488 6783
rect 4436 6740 4488 6749
rect 6460 6740 6512 6792
rect 7932 6783 7984 6792
rect 7932 6749 7941 6783
rect 7941 6749 7975 6783
rect 7975 6749 7984 6783
rect 7932 6740 7984 6749
rect 7472 6715 7524 6724
rect 7472 6681 7481 6715
rect 7481 6681 7515 6715
rect 7515 6681 7524 6715
rect 7472 6672 7524 6681
rect 7840 6672 7892 6724
rect 4436 6604 4488 6656
rect 3547 6502 3599 6554
rect 3611 6502 3663 6554
rect 3675 6502 3727 6554
rect 3739 6502 3791 6554
rect 3803 6502 3855 6554
rect 6144 6502 6196 6554
rect 6208 6502 6260 6554
rect 6272 6502 6324 6554
rect 6336 6502 6388 6554
rect 6400 6502 6452 6554
rect 5724 6400 5776 6452
rect 5908 6400 5960 6452
rect 7472 6332 7524 6384
rect 5908 6264 5960 6316
rect 7104 6264 7156 6316
rect 5816 6060 5868 6112
rect 6000 6060 6052 6112
rect 6552 6060 6604 6112
rect 7012 6128 7064 6180
rect 8116 6060 8168 6112
rect 2248 5958 2300 6010
rect 2312 5958 2364 6010
rect 2376 5958 2428 6010
rect 2440 5958 2492 6010
rect 2504 5958 2556 6010
rect 4846 5958 4898 6010
rect 4910 5958 4962 6010
rect 4974 5958 5026 6010
rect 5038 5958 5090 6010
rect 5102 5958 5154 6010
rect 7443 5958 7495 6010
rect 7507 5958 7559 6010
rect 7571 5958 7623 6010
rect 7635 5958 7687 6010
rect 7699 5958 7751 6010
rect 6368 5856 6420 5908
rect 8024 5856 8076 5908
rect 7196 5788 7248 5840
rect 6920 5720 6972 5772
rect 3240 5627 3292 5636
rect 3240 5593 3249 5627
rect 3249 5593 3283 5627
rect 3283 5593 3292 5627
rect 5724 5652 5776 5704
rect 6368 5695 6420 5704
rect 6368 5661 6377 5695
rect 6377 5661 6411 5695
rect 6411 5661 6420 5695
rect 6368 5652 6420 5661
rect 7104 5652 7156 5704
rect 8116 5652 8168 5704
rect 3240 5584 3292 5593
rect 4068 5559 4120 5568
rect 4068 5525 4077 5559
rect 4077 5525 4111 5559
rect 4111 5525 4120 5559
rect 4068 5516 4120 5525
rect 5908 5627 5960 5636
rect 5908 5593 5917 5627
rect 5917 5593 5951 5627
rect 5951 5593 5960 5627
rect 5908 5584 5960 5593
rect 7012 5627 7064 5636
rect 7012 5593 7021 5627
rect 7021 5593 7055 5627
rect 7055 5593 7064 5627
rect 7012 5584 7064 5593
rect 3547 5414 3599 5466
rect 3611 5414 3663 5466
rect 3675 5414 3727 5466
rect 3739 5414 3791 5466
rect 3803 5414 3855 5466
rect 6144 5414 6196 5466
rect 6208 5414 6260 5466
rect 6272 5414 6324 5466
rect 6336 5414 6388 5466
rect 6400 5414 6452 5466
rect 3240 5312 3292 5364
rect 5540 5312 5592 5364
rect 7288 5312 7340 5364
rect 5908 5244 5960 5296
rect 2872 5040 2924 5092
rect 5172 5219 5224 5228
rect 5172 5185 5181 5219
rect 5181 5185 5215 5219
rect 5215 5185 5224 5219
rect 5172 5176 5224 5185
rect 6552 5176 6604 5228
rect 7196 5219 7248 5228
rect 7196 5185 7205 5219
rect 7205 5185 7239 5219
rect 7239 5185 7248 5219
rect 7196 5176 7248 5185
rect 8024 5176 8076 5228
rect 4712 5108 4764 5160
rect 3056 4972 3108 5024
rect 4344 4972 4396 5024
rect 6920 5040 6972 5092
rect 8116 4972 8168 5024
rect 2248 4870 2300 4922
rect 2312 4870 2364 4922
rect 2376 4870 2428 4922
rect 2440 4870 2492 4922
rect 2504 4870 2556 4922
rect 4846 4870 4898 4922
rect 4910 4870 4962 4922
rect 4974 4870 5026 4922
rect 5038 4870 5090 4922
rect 5102 4870 5154 4922
rect 7443 4870 7495 4922
rect 7507 4870 7559 4922
rect 7571 4870 7623 4922
rect 7635 4870 7687 4922
rect 7699 4870 7751 4922
rect 4436 4700 4488 4752
rect 4804 4700 4856 4752
rect 4160 4632 4212 4684
rect 4620 4632 4672 4684
rect 5816 4632 5868 4684
rect 4160 4539 4212 4548
rect 4160 4505 4169 4539
rect 4169 4505 4203 4539
rect 4203 4505 4212 4539
rect 4160 4496 4212 4505
rect 4528 4564 4580 4616
rect 8116 4607 8168 4616
rect 8116 4573 8125 4607
rect 8125 4573 8159 4607
rect 8159 4573 8168 4607
rect 8116 4564 8168 4573
rect 6828 4539 6880 4548
rect 2688 4471 2740 4480
rect 2688 4437 2697 4471
rect 2697 4437 2731 4471
rect 2731 4437 2740 4471
rect 2688 4428 2740 4437
rect 2872 4428 2924 4480
rect 6828 4505 6837 4539
rect 6837 4505 6871 4539
rect 6871 4505 6880 4539
rect 6828 4496 6880 4505
rect 5448 4428 5500 4480
rect 6000 4428 6052 4480
rect 6552 4428 6604 4480
rect 3547 4326 3599 4378
rect 3611 4326 3663 4378
rect 3675 4326 3727 4378
rect 3739 4326 3791 4378
rect 3803 4326 3855 4378
rect 6144 4326 6196 4378
rect 6208 4326 6260 4378
rect 6272 4326 6324 4378
rect 6336 4326 6388 4378
rect 6400 4326 6452 4378
rect 4436 4224 4488 4276
rect 5172 4224 5224 4276
rect 5540 4224 5592 4276
rect 4160 4156 4212 4208
rect 6552 4199 6604 4208
rect 6552 4165 6561 4199
rect 6561 4165 6595 4199
rect 6595 4165 6604 4199
rect 6552 4156 6604 4165
rect 940 3952 992 4004
rect 4252 4131 4304 4140
rect 4252 4097 4261 4131
rect 4261 4097 4295 4131
rect 4295 4097 4304 4131
rect 7196 4131 7248 4140
rect 4252 4088 4304 4097
rect 7196 4097 7205 4131
rect 7205 4097 7239 4131
rect 7239 4097 7248 4131
rect 7196 4088 7248 4097
rect 8116 4131 8168 4140
rect 8116 4097 8125 4131
rect 8125 4097 8159 4131
rect 8159 4097 8168 4131
rect 8116 4088 8168 4097
rect 4804 4020 4856 4072
rect 5540 4063 5592 4072
rect 5540 4029 5549 4063
rect 5549 4029 5583 4063
rect 5583 4029 5592 4063
rect 5540 4020 5592 4029
rect 4344 3952 4396 4004
rect 5172 3952 5224 4004
rect 3056 3884 3108 3936
rect 3240 3884 3292 3936
rect 4620 3884 4672 3936
rect 5356 3884 5408 3936
rect 2248 3782 2300 3834
rect 2312 3782 2364 3834
rect 2376 3782 2428 3834
rect 2440 3782 2492 3834
rect 2504 3782 2556 3834
rect 4846 3782 4898 3834
rect 4910 3782 4962 3834
rect 4974 3782 5026 3834
rect 5038 3782 5090 3834
rect 5102 3782 5154 3834
rect 7443 3782 7495 3834
rect 7507 3782 7559 3834
rect 7571 3782 7623 3834
rect 7635 3782 7687 3834
rect 7699 3782 7751 3834
rect 5540 3680 5592 3732
rect 6736 3680 6788 3732
rect 2688 3655 2740 3664
rect 2688 3621 2697 3655
rect 2697 3621 2731 3655
rect 2731 3621 2740 3655
rect 2688 3612 2740 3621
rect 3240 3612 3292 3664
rect 2872 3340 2924 3392
rect 4712 3544 4764 3596
rect 5448 3587 5500 3596
rect 5448 3553 5457 3587
rect 5457 3553 5491 3587
rect 5491 3553 5500 3587
rect 5448 3544 5500 3553
rect 7196 3544 7248 3596
rect 4712 3408 4764 3460
rect 5724 3451 5776 3460
rect 5724 3417 5733 3451
rect 5733 3417 5767 3451
rect 5767 3417 5776 3451
rect 5724 3408 5776 3417
rect 8024 3451 8076 3460
rect 3884 3383 3936 3392
rect 3884 3349 3893 3383
rect 3893 3349 3927 3383
rect 3927 3349 3936 3383
rect 3884 3340 3936 3349
rect 6000 3340 6052 3392
rect 8024 3417 8033 3451
rect 8033 3417 8067 3451
rect 8067 3417 8076 3451
rect 8024 3408 8076 3417
rect 8944 3340 8996 3392
rect 3547 3238 3599 3290
rect 3611 3238 3663 3290
rect 3675 3238 3727 3290
rect 3739 3238 3791 3290
rect 3803 3238 3855 3290
rect 6144 3238 6196 3290
rect 6208 3238 6260 3290
rect 6272 3238 6324 3290
rect 6336 3238 6388 3290
rect 6400 3238 6452 3290
rect 4252 3136 4304 3188
rect 5356 3179 5408 3188
rect 5356 3145 5365 3179
rect 5365 3145 5399 3179
rect 5399 3145 5408 3179
rect 5356 3136 5408 3145
rect 5448 3179 5500 3188
rect 5448 3145 5457 3179
rect 5457 3145 5491 3179
rect 5491 3145 5500 3179
rect 5448 3136 5500 3145
rect 4528 3068 4580 3120
rect 6552 3043 6604 3052
rect 940 2932 992 2984
rect 3884 2932 3936 2984
rect 6552 3009 6561 3043
rect 6561 3009 6595 3043
rect 6595 3009 6604 3043
rect 6552 3000 6604 3009
rect 7104 3000 7156 3052
rect 4436 2932 4488 2984
rect 3056 2864 3108 2916
rect 6552 2864 6604 2916
rect 7196 2864 7248 2916
rect 8024 2864 8076 2916
rect 6000 2796 6052 2848
rect 2248 2694 2300 2746
rect 2312 2694 2364 2746
rect 2376 2694 2428 2746
rect 2440 2694 2492 2746
rect 2504 2694 2556 2746
rect 4846 2694 4898 2746
rect 4910 2694 4962 2746
rect 4974 2694 5026 2746
rect 5038 2694 5090 2746
rect 5102 2694 5154 2746
rect 7443 2694 7495 2746
rect 7507 2694 7559 2746
rect 7571 2694 7623 2746
rect 7635 2694 7687 2746
rect 7699 2694 7751 2746
rect 3056 2592 3108 2644
rect 5724 2592 5776 2644
rect 6552 2524 6604 2576
rect 4252 2456 4304 2508
rect 5172 2499 5224 2508
rect 4528 2431 4580 2440
rect 4528 2397 4537 2431
rect 4537 2397 4571 2431
rect 4571 2397 4580 2431
rect 4528 2388 4580 2397
rect 5172 2465 5181 2499
rect 5181 2465 5215 2499
rect 5215 2465 5224 2499
rect 5172 2456 5224 2465
rect 6828 2456 6880 2508
rect 7196 2499 7248 2508
rect 7196 2465 7205 2499
rect 7205 2465 7239 2499
rect 7239 2465 7248 2499
rect 7196 2456 7248 2465
rect 4896 2388 4948 2440
rect 5448 2388 5500 2440
rect 6736 2388 6788 2440
rect 7012 2388 7064 2440
rect 7656 2431 7708 2440
rect 7656 2397 7665 2431
rect 7665 2397 7699 2431
rect 7699 2397 7708 2431
rect 7656 2388 7708 2397
rect 4712 2320 4764 2372
rect 3547 2150 3599 2202
rect 3611 2150 3663 2202
rect 3675 2150 3727 2202
rect 3739 2150 3791 2202
rect 3803 2150 3855 2202
rect 6144 2150 6196 2202
rect 6208 2150 6260 2202
rect 6272 2150 6324 2202
rect 6336 2150 6388 2202
rect 6400 2150 6452 2202
<< metal2 >>
rect 8206 29472 8262 29481
rect 8206 29407 8262 29416
rect 5538 28384 5594 28393
rect 5538 28319 5594 28328
rect 2248 27772 2556 27792
rect 2248 27770 2254 27772
rect 2310 27770 2334 27772
rect 2390 27770 2414 27772
rect 2470 27770 2494 27772
rect 2550 27770 2556 27772
rect 2310 27718 2312 27770
rect 2492 27718 2494 27770
rect 2248 27716 2254 27718
rect 2310 27716 2334 27718
rect 2390 27716 2414 27718
rect 2470 27716 2494 27718
rect 2550 27716 2556 27718
rect 2248 27696 2556 27716
rect 4846 27772 5154 27792
rect 4846 27770 4852 27772
rect 4908 27770 4932 27772
rect 4988 27770 5012 27772
rect 5068 27770 5092 27772
rect 5148 27770 5154 27772
rect 4908 27718 4910 27770
rect 5090 27718 5092 27770
rect 4846 27716 4852 27718
rect 4908 27716 4932 27718
rect 4988 27716 5012 27718
rect 5068 27716 5092 27718
rect 5148 27716 5154 27718
rect 4846 27696 5154 27716
rect 3547 27228 3855 27248
rect 3547 27226 3553 27228
rect 3609 27226 3633 27228
rect 3689 27226 3713 27228
rect 3769 27226 3793 27228
rect 3849 27226 3855 27228
rect 3609 27174 3611 27226
rect 3791 27174 3793 27226
rect 3547 27172 3553 27174
rect 3609 27172 3633 27174
rect 3689 27172 3713 27174
rect 3769 27172 3793 27174
rect 3849 27172 3855 27174
rect 3547 27152 3855 27172
rect 5264 26920 5316 26926
rect 5264 26862 5316 26868
rect 2248 26684 2556 26704
rect 2248 26682 2254 26684
rect 2310 26682 2334 26684
rect 2390 26682 2414 26684
rect 2470 26682 2494 26684
rect 2550 26682 2556 26684
rect 2310 26630 2312 26682
rect 2492 26630 2494 26682
rect 2248 26628 2254 26630
rect 2310 26628 2334 26630
rect 2390 26628 2414 26630
rect 2470 26628 2494 26630
rect 2550 26628 2556 26630
rect 2248 26608 2556 26628
rect 4846 26684 5154 26704
rect 4846 26682 4852 26684
rect 4908 26682 4932 26684
rect 4988 26682 5012 26684
rect 5068 26682 5092 26684
rect 5148 26682 5154 26684
rect 4908 26630 4910 26682
rect 5090 26630 5092 26682
rect 4846 26628 4852 26630
rect 4908 26628 4932 26630
rect 4988 26628 5012 26630
rect 5068 26628 5092 26630
rect 5148 26628 5154 26630
rect 4846 26608 5154 26628
rect 5276 26586 5304 26862
rect 5264 26580 5316 26586
rect 5264 26522 5316 26528
rect 3547 26140 3855 26160
rect 3547 26138 3553 26140
rect 3609 26138 3633 26140
rect 3689 26138 3713 26140
rect 3769 26138 3793 26140
rect 3849 26138 3855 26140
rect 3609 26086 3611 26138
rect 3791 26086 3793 26138
rect 3547 26084 3553 26086
rect 3609 26084 3633 26086
rect 3689 26084 3713 26086
rect 3769 26084 3793 26086
rect 3849 26084 3855 26086
rect 3547 26064 3855 26084
rect 2248 25596 2556 25616
rect 2248 25594 2254 25596
rect 2310 25594 2334 25596
rect 2390 25594 2414 25596
rect 2470 25594 2494 25596
rect 2550 25594 2556 25596
rect 2310 25542 2312 25594
rect 2492 25542 2494 25594
rect 2248 25540 2254 25542
rect 2310 25540 2334 25542
rect 2390 25540 2414 25542
rect 2470 25540 2494 25542
rect 2550 25540 2556 25542
rect 2248 25520 2556 25540
rect 4846 25596 5154 25616
rect 4846 25594 4852 25596
rect 4908 25594 4932 25596
rect 4988 25594 5012 25596
rect 5068 25594 5092 25596
rect 5148 25594 5154 25596
rect 4908 25542 4910 25594
rect 5090 25542 5092 25594
rect 4846 25540 4852 25542
rect 4908 25540 4932 25542
rect 4988 25540 5012 25542
rect 5068 25540 5092 25542
rect 5148 25540 5154 25542
rect 4846 25520 5154 25540
rect 3547 25052 3855 25072
rect 3547 25050 3553 25052
rect 3609 25050 3633 25052
rect 3689 25050 3713 25052
rect 3769 25050 3793 25052
rect 3849 25050 3855 25052
rect 3609 24998 3611 25050
rect 3791 24998 3793 25050
rect 3547 24996 3553 24998
rect 3609 24996 3633 24998
rect 3689 24996 3713 24998
rect 3769 24996 3793 24998
rect 3849 24996 3855 24998
rect 3547 24976 3855 24996
rect 2248 24508 2556 24528
rect 2248 24506 2254 24508
rect 2310 24506 2334 24508
rect 2390 24506 2414 24508
rect 2470 24506 2494 24508
rect 2550 24506 2556 24508
rect 2310 24454 2312 24506
rect 2492 24454 2494 24506
rect 2248 24452 2254 24454
rect 2310 24452 2334 24454
rect 2390 24452 2414 24454
rect 2470 24452 2494 24454
rect 2550 24452 2556 24454
rect 2248 24432 2556 24452
rect 4846 24508 5154 24528
rect 4846 24506 4852 24508
rect 4908 24506 4932 24508
rect 4988 24506 5012 24508
rect 5068 24506 5092 24508
rect 5148 24506 5154 24508
rect 4908 24454 4910 24506
rect 5090 24454 5092 24506
rect 4846 24452 4852 24454
rect 4908 24452 4932 24454
rect 4988 24452 5012 24454
rect 5068 24452 5092 24454
rect 5148 24452 5154 24454
rect 4846 24432 5154 24452
rect 3547 23964 3855 23984
rect 3547 23962 3553 23964
rect 3609 23962 3633 23964
rect 3689 23962 3713 23964
rect 3769 23962 3793 23964
rect 3849 23962 3855 23964
rect 3609 23910 3611 23962
rect 3791 23910 3793 23962
rect 3547 23908 3553 23910
rect 3609 23908 3633 23910
rect 3689 23908 3713 23910
rect 3769 23908 3793 23910
rect 3849 23908 3855 23910
rect 3547 23888 3855 23908
rect 2248 23420 2556 23440
rect 2248 23418 2254 23420
rect 2310 23418 2334 23420
rect 2390 23418 2414 23420
rect 2470 23418 2494 23420
rect 2550 23418 2556 23420
rect 2310 23366 2312 23418
rect 2492 23366 2494 23418
rect 2248 23364 2254 23366
rect 2310 23364 2334 23366
rect 2390 23364 2414 23366
rect 2470 23364 2494 23366
rect 2550 23364 2556 23366
rect 2248 23344 2556 23364
rect 4846 23420 5154 23440
rect 4846 23418 4852 23420
rect 4908 23418 4932 23420
rect 4988 23418 5012 23420
rect 5068 23418 5092 23420
rect 5148 23418 5154 23420
rect 4908 23366 4910 23418
rect 5090 23366 5092 23418
rect 4846 23364 4852 23366
rect 4908 23364 4932 23366
rect 4988 23364 5012 23366
rect 5068 23364 5092 23366
rect 5148 23364 5154 23366
rect 4846 23344 5154 23364
rect 3547 22876 3855 22896
rect 3547 22874 3553 22876
rect 3609 22874 3633 22876
rect 3689 22874 3713 22876
rect 3769 22874 3793 22876
rect 3849 22874 3855 22876
rect 3609 22822 3611 22874
rect 3791 22822 3793 22874
rect 3547 22820 3553 22822
rect 3609 22820 3633 22822
rect 3689 22820 3713 22822
rect 3769 22820 3793 22822
rect 3849 22820 3855 22822
rect 3547 22800 3855 22820
rect 2248 22332 2556 22352
rect 2248 22330 2254 22332
rect 2310 22330 2334 22332
rect 2390 22330 2414 22332
rect 2470 22330 2494 22332
rect 2550 22330 2556 22332
rect 2310 22278 2312 22330
rect 2492 22278 2494 22330
rect 2248 22276 2254 22278
rect 2310 22276 2334 22278
rect 2390 22276 2414 22278
rect 2470 22276 2494 22278
rect 2550 22276 2556 22278
rect 2248 22256 2556 22276
rect 4846 22332 5154 22352
rect 4846 22330 4852 22332
rect 4908 22330 4932 22332
rect 4988 22330 5012 22332
rect 5068 22330 5092 22332
rect 5148 22330 5154 22332
rect 4908 22278 4910 22330
rect 5090 22278 5092 22330
rect 4846 22276 4852 22278
rect 4908 22276 4932 22278
rect 4988 22276 5012 22278
rect 5068 22276 5092 22278
rect 5148 22276 5154 22278
rect 4846 22256 5154 22276
rect 3547 21788 3855 21808
rect 3547 21786 3553 21788
rect 3609 21786 3633 21788
rect 3689 21786 3713 21788
rect 3769 21786 3793 21788
rect 3849 21786 3855 21788
rect 3609 21734 3611 21786
rect 3791 21734 3793 21786
rect 3547 21732 3553 21734
rect 3609 21732 3633 21734
rect 3689 21732 3713 21734
rect 3769 21732 3793 21734
rect 3849 21732 3855 21734
rect 3547 21712 3855 21732
rect 5354 21448 5410 21457
rect 5354 21383 5410 21392
rect 5172 21344 5224 21350
rect 5172 21286 5224 21292
rect 2248 21244 2556 21264
rect 2248 21242 2254 21244
rect 2310 21242 2334 21244
rect 2390 21242 2414 21244
rect 2470 21242 2494 21244
rect 2550 21242 2556 21244
rect 2310 21190 2312 21242
rect 2492 21190 2494 21242
rect 2248 21188 2254 21190
rect 2310 21188 2334 21190
rect 2390 21188 2414 21190
rect 2470 21188 2494 21190
rect 2550 21188 2556 21190
rect 2248 21168 2556 21188
rect 4846 21244 5154 21264
rect 4846 21242 4852 21244
rect 4908 21242 4932 21244
rect 4988 21242 5012 21244
rect 5068 21242 5092 21244
rect 5148 21242 5154 21244
rect 4908 21190 4910 21242
rect 5090 21190 5092 21242
rect 4846 21188 4852 21190
rect 4908 21188 4932 21190
rect 4988 21188 5012 21190
rect 5068 21188 5092 21190
rect 5148 21188 5154 21190
rect 4846 21168 5154 21188
rect 5184 20942 5212 21286
rect 5172 20936 5224 20942
rect 5172 20878 5224 20884
rect 3547 20700 3855 20720
rect 3547 20698 3553 20700
rect 3609 20698 3633 20700
rect 3689 20698 3713 20700
rect 3769 20698 3793 20700
rect 3849 20698 3855 20700
rect 3609 20646 3611 20698
rect 3791 20646 3793 20698
rect 3547 20644 3553 20646
rect 3609 20644 3633 20646
rect 3689 20644 3713 20646
rect 3769 20644 3793 20646
rect 3849 20644 3855 20646
rect 3547 20624 3855 20644
rect 5184 20602 5212 20878
rect 5264 20800 5316 20806
rect 5264 20742 5316 20748
rect 5172 20596 5224 20602
rect 5172 20538 5224 20544
rect 2248 20156 2556 20176
rect 2248 20154 2254 20156
rect 2310 20154 2334 20156
rect 2390 20154 2414 20156
rect 2470 20154 2494 20156
rect 2550 20154 2556 20156
rect 2310 20102 2312 20154
rect 2492 20102 2494 20154
rect 2248 20100 2254 20102
rect 2310 20100 2334 20102
rect 2390 20100 2414 20102
rect 2470 20100 2494 20102
rect 2550 20100 2556 20102
rect 2248 20080 2556 20100
rect 4846 20156 5154 20176
rect 4846 20154 4852 20156
rect 4908 20154 4932 20156
rect 4988 20154 5012 20156
rect 5068 20154 5092 20156
rect 5148 20154 5154 20156
rect 4908 20102 4910 20154
rect 5090 20102 5092 20154
rect 4846 20100 4852 20102
rect 4908 20100 4932 20102
rect 4988 20100 5012 20102
rect 5068 20100 5092 20102
rect 5148 20100 5154 20102
rect 4846 20080 5154 20100
rect 5276 19718 5304 20742
rect 5264 19712 5316 19718
rect 5264 19654 5316 19660
rect 3547 19612 3855 19632
rect 3547 19610 3553 19612
rect 3609 19610 3633 19612
rect 3689 19610 3713 19612
rect 3769 19610 3793 19612
rect 3849 19610 3855 19612
rect 3609 19558 3611 19610
rect 3791 19558 3793 19610
rect 3547 19556 3553 19558
rect 3609 19556 3633 19558
rect 3689 19556 3713 19558
rect 3769 19556 3793 19558
rect 3849 19556 3855 19558
rect 3547 19536 3855 19556
rect 2248 19068 2556 19088
rect 2248 19066 2254 19068
rect 2310 19066 2334 19068
rect 2390 19066 2414 19068
rect 2470 19066 2494 19068
rect 2550 19066 2556 19068
rect 2310 19014 2312 19066
rect 2492 19014 2494 19066
rect 2248 19012 2254 19014
rect 2310 19012 2334 19014
rect 2390 19012 2414 19014
rect 2470 19012 2494 19014
rect 2550 19012 2556 19014
rect 2248 18992 2556 19012
rect 4846 19068 5154 19088
rect 4846 19066 4852 19068
rect 4908 19066 4932 19068
rect 4988 19066 5012 19068
rect 5068 19066 5092 19068
rect 5148 19066 5154 19068
rect 4908 19014 4910 19066
rect 5090 19014 5092 19066
rect 4846 19012 4852 19014
rect 4908 19012 4932 19014
rect 4988 19012 5012 19014
rect 5068 19012 5092 19014
rect 5148 19012 5154 19014
rect 4846 18992 5154 19012
rect 3547 18524 3855 18544
rect 3547 18522 3553 18524
rect 3609 18522 3633 18524
rect 3689 18522 3713 18524
rect 3769 18522 3793 18524
rect 3849 18522 3855 18524
rect 3609 18470 3611 18522
rect 3791 18470 3793 18522
rect 3547 18468 3553 18470
rect 3609 18468 3633 18470
rect 3689 18468 3713 18470
rect 3769 18468 3793 18470
rect 3849 18468 3855 18470
rect 3547 18448 3855 18468
rect 2248 17980 2556 18000
rect 2248 17978 2254 17980
rect 2310 17978 2334 17980
rect 2390 17978 2414 17980
rect 2470 17978 2494 17980
rect 2550 17978 2556 17980
rect 2310 17926 2312 17978
rect 2492 17926 2494 17978
rect 2248 17924 2254 17926
rect 2310 17924 2334 17926
rect 2390 17924 2414 17926
rect 2470 17924 2494 17926
rect 2550 17924 2556 17926
rect 2248 17904 2556 17924
rect 4846 17980 5154 18000
rect 4846 17978 4852 17980
rect 4908 17978 4932 17980
rect 4988 17978 5012 17980
rect 5068 17978 5092 17980
rect 5148 17978 5154 17980
rect 4908 17926 4910 17978
rect 5090 17926 5092 17978
rect 4846 17924 4852 17926
rect 4908 17924 4932 17926
rect 4988 17924 5012 17926
rect 5068 17924 5092 17926
rect 5148 17924 5154 17926
rect 4846 17904 5154 17924
rect 3547 17436 3855 17456
rect 3547 17434 3553 17436
rect 3609 17434 3633 17436
rect 3689 17434 3713 17436
rect 3769 17434 3793 17436
rect 3849 17434 3855 17436
rect 3609 17382 3611 17434
rect 3791 17382 3793 17434
rect 3547 17380 3553 17382
rect 3609 17380 3633 17382
rect 3689 17380 3713 17382
rect 3769 17380 3793 17382
rect 3849 17380 3855 17382
rect 3547 17360 3855 17380
rect 2248 16892 2556 16912
rect 2248 16890 2254 16892
rect 2310 16890 2334 16892
rect 2390 16890 2414 16892
rect 2470 16890 2494 16892
rect 2550 16890 2556 16892
rect 2310 16838 2312 16890
rect 2492 16838 2494 16890
rect 2248 16836 2254 16838
rect 2310 16836 2334 16838
rect 2390 16836 2414 16838
rect 2470 16836 2494 16838
rect 2550 16836 2556 16838
rect 2248 16816 2556 16836
rect 4846 16892 5154 16912
rect 4846 16890 4852 16892
rect 4908 16890 4932 16892
rect 4988 16890 5012 16892
rect 5068 16890 5092 16892
rect 5148 16890 5154 16892
rect 4908 16838 4910 16890
rect 5090 16838 5092 16890
rect 4846 16836 4852 16838
rect 4908 16836 4932 16838
rect 4988 16836 5012 16838
rect 5068 16836 5092 16838
rect 5148 16836 5154 16838
rect 4846 16816 5154 16836
rect 3547 16348 3855 16368
rect 3547 16346 3553 16348
rect 3609 16346 3633 16348
rect 3689 16346 3713 16348
rect 3769 16346 3793 16348
rect 3849 16346 3855 16348
rect 3609 16294 3611 16346
rect 3791 16294 3793 16346
rect 3547 16292 3553 16294
rect 3609 16292 3633 16294
rect 3689 16292 3713 16294
rect 3769 16292 3793 16294
rect 3849 16292 3855 16294
rect 3547 16272 3855 16292
rect 5172 16040 5224 16046
rect 5172 15982 5224 15988
rect 2248 15804 2556 15824
rect 2248 15802 2254 15804
rect 2310 15802 2334 15804
rect 2390 15802 2414 15804
rect 2470 15802 2494 15804
rect 2550 15802 2556 15804
rect 2310 15750 2312 15802
rect 2492 15750 2494 15802
rect 2248 15748 2254 15750
rect 2310 15748 2334 15750
rect 2390 15748 2414 15750
rect 2470 15748 2494 15750
rect 2550 15748 2556 15750
rect 2248 15728 2556 15748
rect 4846 15804 5154 15824
rect 4846 15802 4852 15804
rect 4908 15802 4932 15804
rect 4988 15802 5012 15804
rect 5068 15802 5092 15804
rect 5148 15802 5154 15804
rect 4908 15750 4910 15802
rect 5090 15750 5092 15802
rect 4846 15748 4852 15750
rect 4908 15748 4932 15750
rect 4988 15748 5012 15750
rect 5068 15748 5092 15750
rect 5148 15748 5154 15750
rect 4846 15728 5154 15748
rect 5184 15706 5212 15982
rect 5172 15700 5224 15706
rect 5172 15642 5224 15648
rect 3547 15260 3855 15280
rect 3547 15258 3553 15260
rect 3609 15258 3633 15260
rect 3689 15258 3713 15260
rect 3769 15258 3793 15260
rect 3849 15258 3855 15260
rect 3609 15206 3611 15258
rect 3791 15206 3793 15258
rect 3547 15204 3553 15206
rect 3609 15204 3633 15206
rect 3689 15204 3713 15206
rect 3769 15204 3793 15206
rect 3849 15204 3855 15206
rect 3547 15184 3855 15204
rect 2248 14716 2556 14736
rect 2248 14714 2254 14716
rect 2310 14714 2334 14716
rect 2390 14714 2414 14716
rect 2470 14714 2494 14716
rect 2550 14714 2556 14716
rect 2310 14662 2312 14714
rect 2492 14662 2494 14714
rect 2248 14660 2254 14662
rect 2310 14660 2334 14662
rect 2390 14660 2414 14662
rect 2470 14660 2494 14662
rect 2550 14660 2556 14662
rect 2248 14640 2556 14660
rect 4846 14716 5154 14736
rect 4846 14714 4852 14716
rect 4908 14714 4932 14716
rect 4988 14714 5012 14716
rect 5068 14714 5092 14716
rect 5148 14714 5154 14716
rect 4908 14662 4910 14714
rect 5090 14662 5092 14714
rect 4846 14660 4852 14662
rect 4908 14660 4932 14662
rect 4988 14660 5012 14662
rect 5068 14660 5092 14662
rect 5148 14660 5154 14662
rect 4846 14640 5154 14660
rect 3547 14172 3855 14192
rect 3547 14170 3553 14172
rect 3609 14170 3633 14172
rect 3689 14170 3713 14172
rect 3769 14170 3793 14172
rect 3849 14170 3855 14172
rect 3609 14118 3611 14170
rect 3791 14118 3793 14170
rect 3547 14116 3553 14118
rect 3609 14116 3633 14118
rect 3689 14116 3713 14118
rect 3769 14116 3793 14118
rect 3849 14116 3855 14118
rect 3547 14096 3855 14116
rect 2248 13628 2556 13648
rect 2248 13626 2254 13628
rect 2310 13626 2334 13628
rect 2390 13626 2414 13628
rect 2470 13626 2494 13628
rect 2550 13626 2556 13628
rect 2310 13574 2312 13626
rect 2492 13574 2494 13626
rect 2248 13572 2254 13574
rect 2310 13572 2334 13574
rect 2390 13572 2414 13574
rect 2470 13572 2494 13574
rect 2550 13572 2556 13574
rect 2248 13552 2556 13572
rect 4846 13628 5154 13648
rect 4846 13626 4852 13628
rect 4908 13626 4932 13628
rect 4988 13626 5012 13628
rect 5068 13626 5092 13628
rect 5148 13626 5154 13628
rect 4908 13574 4910 13626
rect 5090 13574 5092 13626
rect 4846 13572 4852 13574
rect 4908 13572 4932 13574
rect 4988 13572 5012 13574
rect 5068 13572 5092 13574
rect 5148 13572 5154 13574
rect 4846 13552 5154 13572
rect 3547 13084 3855 13104
rect 3547 13082 3553 13084
rect 3609 13082 3633 13084
rect 3689 13082 3713 13084
rect 3769 13082 3793 13084
rect 3849 13082 3855 13084
rect 3609 13030 3611 13082
rect 3791 13030 3793 13082
rect 3547 13028 3553 13030
rect 3609 13028 3633 13030
rect 3689 13028 3713 13030
rect 3769 13028 3793 13030
rect 3849 13028 3855 13030
rect 3547 13008 3855 13028
rect 2248 12540 2556 12560
rect 2248 12538 2254 12540
rect 2310 12538 2334 12540
rect 2390 12538 2414 12540
rect 2470 12538 2494 12540
rect 2550 12538 2556 12540
rect 2310 12486 2312 12538
rect 2492 12486 2494 12538
rect 2248 12484 2254 12486
rect 2310 12484 2334 12486
rect 2390 12484 2414 12486
rect 2470 12484 2494 12486
rect 2550 12484 2556 12486
rect 2248 12464 2556 12484
rect 4846 12540 5154 12560
rect 4846 12538 4852 12540
rect 4908 12538 4932 12540
rect 4988 12538 5012 12540
rect 5068 12538 5092 12540
rect 5148 12538 5154 12540
rect 4908 12486 4910 12538
rect 5090 12486 5092 12538
rect 4846 12484 4852 12486
rect 4908 12484 4932 12486
rect 4988 12484 5012 12486
rect 5068 12484 5092 12486
rect 5148 12484 5154 12486
rect 4846 12464 5154 12484
rect 5276 12442 5304 19654
rect 5368 15706 5396 21383
rect 5552 20058 5580 28319
rect 7443 27772 7751 27792
rect 7443 27770 7449 27772
rect 7505 27770 7529 27772
rect 7585 27770 7609 27772
rect 7665 27770 7689 27772
rect 7745 27770 7751 27772
rect 7505 27718 7507 27770
rect 7687 27718 7689 27770
rect 7443 27716 7449 27718
rect 7505 27716 7529 27718
rect 7585 27716 7609 27718
rect 7665 27716 7689 27718
rect 7745 27716 7751 27718
rect 7443 27696 7751 27716
rect 7012 27532 7064 27538
rect 7012 27474 7064 27480
rect 6552 27396 6604 27402
rect 6552 27338 6604 27344
rect 5908 27328 5960 27334
rect 5908 27270 5960 27276
rect 5920 27062 5948 27270
rect 6144 27228 6452 27248
rect 6144 27226 6150 27228
rect 6206 27226 6230 27228
rect 6286 27226 6310 27228
rect 6366 27226 6390 27228
rect 6446 27226 6452 27228
rect 6206 27174 6208 27226
rect 6388 27174 6390 27226
rect 6144 27172 6150 27174
rect 6206 27172 6230 27174
rect 6286 27172 6310 27174
rect 6366 27172 6390 27174
rect 6446 27172 6452 27174
rect 6144 27152 6452 27172
rect 6564 27130 6592 27338
rect 6734 27160 6790 27169
rect 6552 27124 6604 27130
rect 6734 27095 6790 27104
rect 6552 27066 6604 27072
rect 5908 27056 5960 27062
rect 5908 26998 5960 27004
rect 5816 24268 5868 24274
rect 5816 24210 5868 24216
rect 5828 23866 5856 24210
rect 5816 23860 5868 23866
rect 5816 23802 5868 23808
rect 5814 22536 5870 22545
rect 5814 22471 5870 22480
rect 5724 22432 5776 22438
rect 5724 22374 5776 22380
rect 5736 21622 5764 22374
rect 5724 21616 5776 21622
rect 5724 21558 5776 21564
rect 5632 21548 5684 21554
rect 5632 21490 5684 21496
rect 5644 20874 5672 21490
rect 5632 20868 5684 20874
rect 5632 20810 5684 20816
rect 5724 20868 5776 20874
rect 5724 20810 5776 20816
rect 5736 20602 5764 20810
rect 5724 20596 5776 20602
rect 5724 20538 5776 20544
rect 5540 20052 5592 20058
rect 5540 19994 5592 20000
rect 5538 19952 5594 19961
rect 5538 19887 5594 19896
rect 5552 17898 5580 19887
rect 5632 19168 5684 19174
rect 5632 19110 5684 19116
rect 5460 17870 5580 17898
rect 5460 16674 5488 17870
rect 5540 17740 5592 17746
rect 5540 17682 5592 17688
rect 5552 16794 5580 17682
rect 5540 16788 5592 16794
rect 5540 16730 5592 16736
rect 5460 16646 5580 16674
rect 5356 15700 5408 15706
rect 5356 15642 5408 15648
rect 5368 15570 5396 15642
rect 5356 15564 5408 15570
rect 5356 15506 5408 15512
rect 5368 15162 5396 15506
rect 5356 15156 5408 15162
rect 5356 15098 5408 15104
rect 5552 15042 5580 16646
rect 5460 15014 5580 15042
rect 5460 13410 5488 15014
rect 5540 14884 5592 14890
rect 5540 14826 5592 14832
rect 5552 14414 5580 14826
rect 5540 14408 5592 14414
rect 5540 14350 5592 14356
rect 5552 13530 5580 14350
rect 5540 13524 5592 13530
rect 5540 13466 5592 13472
rect 5460 13382 5580 13410
rect 5552 12850 5580 13382
rect 5540 12844 5592 12850
rect 5540 12786 5592 12792
rect 5264 12436 5316 12442
rect 5264 12378 5316 12384
rect 5540 12232 5592 12238
rect 5540 12174 5592 12180
rect 3547 11996 3855 12016
rect 3547 11994 3553 11996
rect 3609 11994 3633 11996
rect 3689 11994 3713 11996
rect 3769 11994 3793 11996
rect 3849 11994 3855 11996
rect 3609 11942 3611 11994
rect 3791 11942 3793 11994
rect 3547 11940 3553 11942
rect 3609 11940 3633 11942
rect 3689 11940 3713 11942
rect 3769 11940 3793 11942
rect 3849 11940 3855 11942
rect 3547 11920 3855 11940
rect 5552 11642 5580 12174
rect 5460 11614 5580 11642
rect 2248 11452 2556 11472
rect 2248 11450 2254 11452
rect 2310 11450 2334 11452
rect 2390 11450 2414 11452
rect 2470 11450 2494 11452
rect 2550 11450 2556 11452
rect 2310 11398 2312 11450
rect 2492 11398 2494 11450
rect 2248 11396 2254 11398
rect 2310 11396 2334 11398
rect 2390 11396 2414 11398
rect 2470 11396 2494 11398
rect 2550 11396 2556 11398
rect 2248 11376 2556 11396
rect 4846 11452 5154 11472
rect 4846 11450 4852 11452
rect 4908 11450 4932 11452
rect 4988 11450 5012 11452
rect 5068 11450 5092 11452
rect 5148 11450 5154 11452
rect 4908 11398 4910 11450
rect 5090 11398 5092 11450
rect 4846 11396 4852 11398
rect 4908 11396 4932 11398
rect 4988 11396 5012 11398
rect 5068 11396 5092 11398
rect 5148 11396 5154 11398
rect 4846 11376 5154 11396
rect 5460 11098 5488 11614
rect 5540 11552 5592 11558
rect 5540 11494 5592 11500
rect 5552 11354 5580 11494
rect 5540 11348 5592 11354
rect 5540 11290 5592 11296
rect 5460 11070 5580 11098
rect 3547 10908 3855 10928
rect 3547 10906 3553 10908
rect 3609 10906 3633 10908
rect 3689 10906 3713 10908
rect 3769 10906 3793 10908
rect 3849 10906 3855 10908
rect 3609 10854 3611 10906
rect 3791 10854 3793 10906
rect 3547 10852 3553 10854
rect 3609 10852 3633 10854
rect 3689 10852 3713 10854
rect 3769 10852 3793 10854
rect 3849 10852 3855 10854
rect 3547 10832 3855 10852
rect 2248 10364 2556 10384
rect 2248 10362 2254 10364
rect 2310 10362 2334 10364
rect 2390 10362 2414 10364
rect 2470 10362 2494 10364
rect 2550 10362 2556 10364
rect 2310 10310 2312 10362
rect 2492 10310 2494 10362
rect 2248 10308 2254 10310
rect 2310 10308 2334 10310
rect 2390 10308 2414 10310
rect 2470 10308 2494 10310
rect 2550 10308 2556 10310
rect 2248 10288 2556 10308
rect 4846 10364 5154 10384
rect 4846 10362 4852 10364
rect 4908 10362 4932 10364
rect 4988 10362 5012 10364
rect 5068 10362 5092 10364
rect 5148 10362 5154 10364
rect 4908 10310 4910 10362
rect 5090 10310 5092 10362
rect 4846 10308 4852 10310
rect 4908 10308 4932 10310
rect 4988 10308 5012 10310
rect 5068 10308 5092 10310
rect 5148 10308 5154 10310
rect 4846 10288 5154 10308
rect 5552 10282 5580 11070
rect 5460 10254 5580 10282
rect 5460 9926 5488 10254
rect 5540 10124 5592 10130
rect 5540 10066 5592 10072
rect 5448 9920 5500 9926
rect 5448 9862 5500 9868
rect 3547 9820 3855 9840
rect 3547 9818 3553 9820
rect 3609 9818 3633 9820
rect 3689 9818 3713 9820
rect 3769 9818 3793 9820
rect 3849 9818 3855 9820
rect 3609 9766 3611 9818
rect 3791 9766 3793 9818
rect 3547 9764 3553 9766
rect 3609 9764 3633 9766
rect 3689 9764 3713 9766
rect 3769 9764 3793 9766
rect 3849 9764 3855 9766
rect 3547 9744 3855 9764
rect 2248 9276 2556 9296
rect 2248 9274 2254 9276
rect 2310 9274 2334 9276
rect 2390 9274 2414 9276
rect 2470 9274 2494 9276
rect 2550 9274 2556 9276
rect 2310 9222 2312 9274
rect 2492 9222 2494 9274
rect 2248 9220 2254 9222
rect 2310 9220 2334 9222
rect 2390 9220 2414 9222
rect 2470 9220 2494 9222
rect 2550 9220 2556 9222
rect 2248 9200 2556 9220
rect 4846 9276 5154 9296
rect 4846 9274 4852 9276
rect 4908 9274 4932 9276
rect 4988 9274 5012 9276
rect 5068 9274 5092 9276
rect 5148 9274 5154 9276
rect 4908 9222 4910 9274
rect 5090 9222 5092 9274
rect 4846 9220 4852 9222
rect 4908 9220 4932 9222
rect 4988 9220 5012 9222
rect 5068 9220 5092 9222
rect 5148 9220 5154 9222
rect 4846 9200 5154 9220
rect 3547 8732 3855 8752
rect 3547 8730 3553 8732
rect 3609 8730 3633 8732
rect 3689 8730 3713 8732
rect 3769 8730 3793 8732
rect 3849 8730 3855 8732
rect 3609 8678 3611 8730
rect 3791 8678 3793 8730
rect 3547 8676 3553 8678
rect 3609 8676 3633 8678
rect 3689 8676 3713 8678
rect 3769 8676 3793 8678
rect 3849 8676 3855 8678
rect 3547 8656 3855 8676
rect 5552 8634 5580 10066
rect 5644 10033 5672 19110
rect 5724 18284 5776 18290
rect 5724 18226 5776 18232
rect 5736 18086 5764 18226
rect 5724 18080 5776 18086
rect 5724 18022 5776 18028
rect 5736 17610 5764 18022
rect 5828 17746 5856 22471
rect 5816 17740 5868 17746
rect 5816 17682 5868 17688
rect 5724 17604 5776 17610
rect 5724 17546 5776 17552
rect 5736 13297 5764 17546
rect 5920 17338 5948 26998
rect 6368 26988 6420 26994
rect 6368 26930 6420 26936
rect 6380 26382 6408 26930
rect 6368 26376 6420 26382
rect 6368 26318 6420 26324
rect 6144 26140 6452 26160
rect 6144 26138 6150 26140
rect 6206 26138 6230 26140
rect 6286 26138 6310 26140
rect 6366 26138 6390 26140
rect 6446 26138 6452 26140
rect 6206 26086 6208 26138
rect 6388 26086 6390 26138
rect 6144 26084 6150 26086
rect 6206 26084 6230 26086
rect 6286 26084 6310 26086
rect 6366 26084 6390 26086
rect 6446 26084 6452 26086
rect 6144 26064 6452 26084
rect 6644 25152 6696 25158
rect 6644 25094 6696 25100
rect 6144 25052 6452 25072
rect 6144 25050 6150 25052
rect 6206 25050 6230 25052
rect 6286 25050 6310 25052
rect 6366 25050 6390 25052
rect 6446 25050 6452 25052
rect 6206 24998 6208 25050
rect 6388 24998 6390 25050
rect 6144 24996 6150 24998
rect 6206 24996 6230 24998
rect 6286 24996 6310 24998
rect 6366 24996 6390 24998
rect 6446 24996 6452 24998
rect 6144 24976 6452 24996
rect 6656 24614 6684 25094
rect 6644 24608 6696 24614
rect 6644 24550 6696 24556
rect 6144 23964 6452 23984
rect 6144 23962 6150 23964
rect 6206 23962 6230 23964
rect 6286 23962 6310 23964
rect 6366 23962 6390 23964
rect 6446 23962 6452 23964
rect 6206 23910 6208 23962
rect 6388 23910 6390 23962
rect 6144 23908 6150 23910
rect 6206 23908 6230 23910
rect 6286 23908 6310 23910
rect 6366 23908 6390 23910
rect 6446 23908 6452 23910
rect 6144 23888 6452 23908
rect 6552 23724 6604 23730
rect 6552 23666 6604 23672
rect 6144 22876 6452 22896
rect 6144 22874 6150 22876
rect 6206 22874 6230 22876
rect 6286 22874 6310 22876
rect 6366 22874 6390 22876
rect 6446 22874 6452 22876
rect 6206 22822 6208 22874
rect 6388 22822 6390 22874
rect 6144 22820 6150 22822
rect 6206 22820 6230 22822
rect 6286 22820 6310 22822
rect 6366 22820 6390 22822
rect 6446 22820 6452 22822
rect 6144 22800 6452 22820
rect 6000 21888 6052 21894
rect 6000 21830 6052 21836
rect 6012 21486 6040 21830
rect 6144 21788 6452 21808
rect 6144 21786 6150 21788
rect 6206 21786 6230 21788
rect 6286 21786 6310 21788
rect 6366 21786 6390 21788
rect 6446 21786 6452 21788
rect 6206 21734 6208 21786
rect 6388 21734 6390 21786
rect 6144 21732 6150 21734
rect 6206 21732 6230 21734
rect 6286 21732 6310 21734
rect 6366 21732 6390 21734
rect 6446 21732 6452 21734
rect 6144 21712 6452 21732
rect 6000 21480 6052 21486
rect 6000 21422 6052 21428
rect 6012 17921 6040 21422
rect 6184 21344 6236 21350
rect 6184 21286 6236 21292
rect 6196 21010 6224 21286
rect 6564 21078 6592 23666
rect 6656 22386 6684 24550
rect 6748 23254 6776 27095
rect 7024 26450 7052 27474
rect 7840 27328 7892 27334
rect 7840 27270 7892 27276
rect 7104 26852 7156 26858
rect 7104 26794 7156 26800
rect 7116 26518 7144 26794
rect 7443 26684 7751 26704
rect 7443 26682 7449 26684
rect 7505 26682 7529 26684
rect 7585 26682 7609 26684
rect 7665 26682 7689 26684
rect 7745 26682 7751 26684
rect 7505 26630 7507 26682
rect 7687 26630 7689 26682
rect 7443 26628 7449 26630
rect 7505 26628 7529 26630
rect 7585 26628 7609 26630
rect 7665 26628 7689 26630
rect 7745 26628 7751 26630
rect 7443 26608 7751 26628
rect 7104 26512 7156 26518
rect 7104 26454 7156 26460
rect 7012 26444 7064 26450
rect 7012 26386 7064 26392
rect 6828 26376 6880 26382
rect 6828 26318 6880 26324
rect 6840 25974 6868 26318
rect 6920 26240 6972 26246
rect 7024 26234 7052 26386
rect 7024 26206 7144 26234
rect 6920 26182 6972 26188
rect 6828 25968 6880 25974
rect 6828 25910 6880 25916
rect 6932 25430 6960 26182
rect 7116 25974 7144 26206
rect 7852 26081 7880 27270
rect 8116 26988 8168 26994
rect 8116 26930 8168 26936
rect 8024 26512 8076 26518
rect 8024 26454 8076 26460
rect 7838 26072 7894 26081
rect 7838 26007 7894 26016
rect 7104 25968 7156 25974
rect 7104 25910 7156 25916
rect 7852 25906 7880 26007
rect 7840 25900 7892 25906
rect 7840 25842 7892 25848
rect 7443 25596 7751 25616
rect 7443 25594 7449 25596
rect 7505 25594 7529 25596
rect 7585 25594 7609 25596
rect 7665 25594 7689 25596
rect 7745 25594 7751 25596
rect 7505 25542 7507 25594
rect 7687 25542 7689 25594
rect 7443 25540 7449 25542
rect 7505 25540 7529 25542
rect 7585 25540 7609 25542
rect 7665 25540 7689 25542
rect 7745 25540 7751 25542
rect 7443 25520 7751 25540
rect 6920 25424 6972 25430
rect 6920 25366 6972 25372
rect 7656 25424 7708 25430
rect 7656 25366 7708 25372
rect 7196 25288 7248 25294
rect 7196 25230 7248 25236
rect 7104 24812 7156 24818
rect 7104 24754 7156 24760
rect 7116 24206 7144 24754
rect 7104 24200 7156 24206
rect 7104 24142 7156 24148
rect 7116 23730 7144 24142
rect 7208 24138 7236 25230
rect 7668 24886 7696 25366
rect 7656 24880 7708 24886
rect 7656 24822 7708 24828
rect 7443 24508 7751 24528
rect 7443 24506 7449 24508
rect 7505 24506 7529 24508
rect 7585 24506 7609 24508
rect 7665 24506 7689 24508
rect 7745 24506 7751 24508
rect 7505 24454 7507 24506
rect 7687 24454 7689 24506
rect 7443 24452 7449 24454
rect 7505 24452 7529 24454
rect 7585 24452 7609 24454
rect 7665 24452 7689 24454
rect 7745 24452 7751 24454
rect 7443 24432 7751 24452
rect 7196 24132 7248 24138
rect 7196 24074 7248 24080
rect 7208 23866 7236 24074
rect 7564 24064 7616 24070
rect 7564 24006 7616 24012
rect 7196 23860 7248 23866
rect 7196 23802 7248 23808
rect 7576 23798 7604 24006
rect 7564 23792 7616 23798
rect 7564 23734 7616 23740
rect 7104 23724 7156 23730
rect 7104 23666 7156 23672
rect 7443 23420 7751 23440
rect 7443 23418 7449 23420
rect 7505 23418 7529 23420
rect 7585 23418 7609 23420
rect 7665 23418 7689 23420
rect 7745 23418 7751 23420
rect 7505 23366 7507 23418
rect 7687 23366 7689 23418
rect 7443 23364 7449 23366
rect 7505 23364 7529 23366
rect 7585 23364 7609 23366
rect 7665 23364 7689 23366
rect 7745 23364 7751 23366
rect 7443 23344 7751 23364
rect 6736 23248 6788 23254
rect 6736 23190 6788 23196
rect 6748 22574 6776 23190
rect 7564 23112 7616 23118
rect 7564 23054 7616 23060
rect 6920 23044 6972 23050
rect 6920 22986 6972 22992
rect 6828 22976 6880 22982
rect 6828 22918 6880 22924
rect 6840 22710 6868 22918
rect 6932 22710 6960 22986
rect 7576 22710 7604 23054
rect 8036 22710 8064 26454
rect 8128 26382 8156 26930
rect 8116 26376 8168 26382
rect 8116 26318 8168 26324
rect 8114 24848 8170 24857
rect 8114 24783 8170 24792
rect 8128 24206 8156 24783
rect 8116 24200 8168 24206
rect 8116 24142 8168 24148
rect 8128 23730 8156 24142
rect 8116 23724 8168 23730
rect 8116 23666 8168 23672
rect 6828 22704 6880 22710
rect 6828 22646 6880 22652
rect 6920 22704 6972 22710
rect 6920 22646 6972 22652
rect 7564 22704 7616 22710
rect 7564 22646 7616 22652
rect 7840 22704 7892 22710
rect 7840 22646 7892 22652
rect 8024 22704 8076 22710
rect 8024 22646 8076 22652
rect 6736 22568 6788 22574
rect 6736 22510 6788 22516
rect 6656 22358 6868 22386
rect 6552 21072 6604 21078
rect 6552 21014 6604 21020
rect 6184 21004 6236 21010
rect 6184 20946 6236 20952
rect 6144 20700 6452 20720
rect 6144 20698 6150 20700
rect 6206 20698 6230 20700
rect 6286 20698 6310 20700
rect 6366 20698 6390 20700
rect 6446 20698 6452 20700
rect 6206 20646 6208 20698
rect 6388 20646 6390 20698
rect 6144 20644 6150 20646
rect 6206 20644 6230 20646
rect 6286 20644 6310 20646
rect 6366 20644 6390 20646
rect 6446 20644 6452 20646
rect 6144 20624 6452 20644
rect 6564 20534 6592 21014
rect 6644 20936 6696 20942
rect 6644 20878 6696 20884
rect 6656 20534 6684 20878
rect 6552 20528 6604 20534
rect 6552 20470 6604 20476
rect 6644 20528 6696 20534
rect 6644 20470 6696 20476
rect 6656 19718 6684 20470
rect 6736 19848 6788 19854
rect 6736 19790 6788 19796
rect 6644 19712 6696 19718
rect 6644 19654 6696 19660
rect 6144 19612 6452 19632
rect 6144 19610 6150 19612
rect 6206 19610 6230 19612
rect 6286 19610 6310 19612
rect 6366 19610 6390 19612
rect 6446 19610 6452 19612
rect 6206 19558 6208 19610
rect 6388 19558 6390 19610
rect 6144 19556 6150 19558
rect 6206 19556 6230 19558
rect 6286 19556 6310 19558
rect 6366 19556 6390 19558
rect 6446 19556 6452 19558
rect 6144 19536 6452 19556
rect 6552 19372 6604 19378
rect 6552 19314 6604 19320
rect 6144 18524 6452 18544
rect 6144 18522 6150 18524
rect 6206 18522 6230 18524
rect 6286 18522 6310 18524
rect 6366 18522 6390 18524
rect 6446 18522 6452 18524
rect 6206 18470 6208 18522
rect 6388 18470 6390 18522
rect 6144 18468 6150 18470
rect 6206 18468 6230 18470
rect 6286 18468 6310 18470
rect 6366 18468 6390 18470
rect 6446 18468 6452 18470
rect 6144 18448 6452 18468
rect 5998 17912 6054 17921
rect 5998 17847 6054 17856
rect 5998 17776 6054 17785
rect 5998 17711 6054 17720
rect 5908 17332 5960 17338
rect 5908 17274 5960 17280
rect 5816 16992 5868 16998
rect 5816 16934 5868 16940
rect 5828 16658 5856 16934
rect 6012 16674 6040 17711
rect 6144 17436 6452 17456
rect 6144 17434 6150 17436
rect 6206 17434 6230 17436
rect 6286 17434 6310 17436
rect 6366 17434 6390 17436
rect 6446 17434 6452 17436
rect 6206 17382 6208 17434
rect 6388 17382 6390 17434
rect 6144 17380 6150 17382
rect 6206 17380 6230 17382
rect 6286 17380 6310 17382
rect 6366 17380 6390 17382
rect 6446 17380 6452 17382
rect 6144 17360 6452 17380
rect 6564 17270 6592 19314
rect 6748 19310 6776 19790
rect 6736 19304 6788 19310
rect 6736 19246 6788 19252
rect 6748 18970 6776 19246
rect 6840 19174 6868 22358
rect 7443 22332 7751 22352
rect 7443 22330 7449 22332
rect 7505 22330 7529 22332
rect 7585 22330 7609 22332
rect 7665 22330 7689 22332
rect 7745 22330 7751 22332
rect 7505 22278 7507 22330
rect 7687 22278 7689 22330
rect 7443 22276 7449 22278
rect 7505 22276 7529 22278
rect 7585 22276 7609 22278
rect 7665 22276 7689 22278
rect 7745 22276 7751 22278
rect 7443 22256 7751 22276
rect 7852 22030 7880 22646
rect 8220 22094 8248 29407
rect 8298 23760 8354 23769
rect 8298 23695 8354 23704
rect 8036 22066 8248 22094
rect 7840 22024 7892 22030
rect 7840 21966 7892 21972
rect 7932 21956 7984 21962
rect 7932 21898 7984 21904
rect 7944 21622 7972 21898
rect 7932 21616 7984 21622
rect 7932 21558 7984 21564
rect 7443 21244 7751 21264
rect 7443 21242 7449 21244
rect 7505 21242 7529 21244
rect 7585 21242 7609 21244
rect 7665 21242 7689 21244
rect 7745 21242 7751 21244
rect 7505 21190 7507 21242
rect 7687 21190 7689 21242
rect 7443 21188 7449 21190
rect 7505 21188 7529 21190
rect 7585 21188 7609 21190
rect 7665 21188 7689 21190
rect 7745 21188 7751 21190
rect 7443 21168 7751 21188
rect 7196 20868 7248 20874
rect 7196 20810 7248 20816
rect 7208 20466 7236 20810
rect 8036 20618 8064 22066
rect 8116 21412 8168 21418
rect 8116 21354 8168 21360
rect 7944 20590 8064 20618
rect 7196 20460 7248 20466
rect 7196 20402 7248 20408
rect 7443 20156 7751 20176
rect 7443 20154 7449 20156
rect 7505 20154 7529 20156
rect 7585 20154 7609 20156
rect 7665 20154 7689 20156
rect 7745 20154 7751 20156
rect 7505 20102 7507 20154
rect 7687 20102 7689 20154
rect 7443 20100 7449 20102
rect 7505 20100 7529 20102
rect 7585 20100 7609 20102
rect 7665 20100 7689 20102
rect 7745 20100 7751 20102
rect 7443 20080 7751 20100
rect 7196 19780 7248 19786
rect 7196 19722 7248 19728
rect 7208 19446 7236 19722
rect 7288 19712 7340 19718
rect 7288 19654 7340 19660
rect 7300 19446 7328 19654
rect 7196 19440 7248 19446
rect 7196 19382 7248 19388
rect 7288 19440 7340 19446
rect 7288 19382 7340 19388
rect 6828 19168 6880 19174
rect 6828 19110 6880 19116
rect 6736 18964 6788 18970
rect 6736 18906 6788 18912
rect 6826 18864 6882 18873
rect 6826 18799 6882 18808
rect 6736 18692 6788 18698
rect 6736 18634 6788 18640
rect 6748 18290 6776 18634
rect 6736 18284 6788 18290
rect 6736 18226 6788 18232
rect 6644 17332 6696 17338
rect 6644 17274 6696 17280
rect 6552 17264 6604 17270
rect 6552 17206 6604 17212
rect 6564 16726 6592 17206
rect 5816 16652 5868 16658
rect 5816 16594 5868 16600
rect 5920 16646 6040 16674
rect 6552 16720 6604 16726
rect 6552 16662 6604 16668
rect 5816 15428 5868 15434
rect 5816 15370 5868 15376
rect 5828 14482 5856 15370
rect 5816 14476 5868 14482
rect 5816 14418 5868 14424
rect 5920 14362 5948 16646
rect 6552 16448 6604 16454
rect 6552 16390 6604 16396
rect 6144 16348 6452 16368
rect 6144 16346 6150 16348
rect 6206 16346 6230 16348
rect 6286 16346 6310 16348
rect 6366 16346 6390 16348
rect 6446 16346 6452 16348
rect 6206 16294 6208 16346
rect 6388 16294 6390 16346
rect 6144 16292 6150 16294
rect 6206 16292 6230 16294
rect 6286 16292 6310 16294
rect 6366 16292 6390 16294
rect 6446 16292 6452 16294
rect 6144 16272 6452 16292
rect 6460 15904 6512 15910
rect 6460 15846 6512 15852
rect 6472 15570 6500 15846
rect 6460 15564 6512 15570
rect 6460 15506 6512 15512
rect 6144 15260 6452 15280
rect 6144 15258 6150 15260
rect 6206 15258 6230 15260
rect 6286 15258 6310 15260
rect 6366 15258 6390 15260
rect 6446 15258 6452 15260
rect 6206 15206 6208 15258
rect 6388 15206 6390 15258
rect 6144 15204 6150 15206
rect 6206 15204 6230 15206
rect 6286 15204 6310 15206
rect 6366 15204 6390 15206
rect 6446 15204 6452 15206
rect 6144 15184 6452 15204
rect 6564 15042 6592 16390
rect 6472 15014 6592 15042
rect 6092 14816 6144 14822
rect 6092 14758 6144 14764
rect 6104 14414 6132 14758
rect 5828 14334 5948 14362
rect 6092 14408 6144 14414
rect 6092 14350 6144 14356
rect 6472 14346 6500 15014
rect 6552 14884 6604 14890
rect 6552 14826 6604 14832
rect 6460 14340 6512 14346
rect 5722 13288 5778 13297
rect 5722 13223 5778 13232
rect 5724 12436 5776 12442
rect 5724 12378 5776 12384
rect 5630 10024 5686 10033
rect 5630 9959 5686 9968
rect 5632 9920 5684 9926
rect 5632 9862 5684 9868
rect 5540 8628 5592 8634
rect 5540 8570 5592 8576
rect 2248 8188 2556 8208
rect 2248 8186 2254 8188
rect 2310 8186 2334 8188
rect 2390 8186 2414 8188
rect 2470 8186 2494 8188
rect 2550 8186 2556 8188
rect 2310 8134 2312 8186
rect 2492 8134 2494 8186
rect 2248 8132 2254 8134
rect 2310 8132 2334 8134
rect 2390 8132 2414 8134
rect 2470 8132 2494 8134
rect 2550 8132 2556 8134
rect 2248 8112 2556 8132
rect 4846 8188 5154 8208
rect 4846 8186 4852 8188
rect 4908 8186 4932 8188
rect 4988 8186 5012 8188
rect 5068 8186 5092 8188
rect 5148 8186 5154 8188
rect 4908 8134 4910 8186
rect 5090 8134 5092 8186
rect 4846 8132 4852 8134
rect 4908 8132 4932 8134
rect 4988 8132 5012 8134
rect 5068 8132 5092 8134
rect 5148 8132 5154 8134
rect 4846 8112 5154 8132
rect 5540 8016 5592 8022
rect 5540 7958 5592 7964
rect 5644 7970 5672 9862
rect 5736 8945 5764 12378
rect 5828 12238 5856 14334
rect 6460 14282 6512 14288
rect 6144 14172 6452 14192
rect 6144 14170 6150 14172
rect 6206 14170 6230 14172
rect 6286 14170 6310 14172
rect 6366 14170 6390 14172
rect 6446 14170 6452 14172
rect 6206 14118 6208 14170
rect 6388 14118 6390 14170
rect 6144 14116 6150 14118
rect 6206 14116 6230 14118
rect 6286 14116 6310 14118
rect 6366 14116 6390 14118
rect 6446 14116 6452 14118
rect 6144 14096 6452 14116
rect 6000 13932 6052 13938
rect 6000 13874 6052 13880
rect 6012 13734 6040 13874
rect 6000 13728 6052 13734
rect 6000 13670 6052 13676
rect 6012 13190 6040 13670
rect 6000 13184 6052 13190
rect 6000 13126 6052 13132
rect 6012 12866 6040 13126
rect 6144 13084 6452 13104
rect 6144 13082 6150 13084
rect 6206 13082 6230 13084
rect 6286 13082 6310 13084
rect 6366 13082 6390 13084
rect 6446 13082 6452 13084
rect 6206 13030 6208 13082
rect 6388 13030 6390 13082
rect 6144 13028 6150 13030
rect 6206 13028 6230 13030
rect 6286 13028 6310 13030
rect 6366 13028 6390 13030
rect 6446 13028 6452 13030
rect 6144 13008 6452 13028
rect 6012 12838 6132 12866
rect 5998 12744 6054 12753
rect 5998 12679 6054 12688
rect 6012 12345 6040 12679
rect 5998 12336 6054 12345
rect 5998 12271 6054 12280
rect 5816 12232 5868 12238
rect 5816 12174 5868 12180
rect 5908 12232 5960 12238
rect 6104 12186 6132 12838
rect 6184 12844 6236 12850
rect 6184 12786 6236 12792
rect 5908 12174 5960 12180
rect 5816 12096 5868 12102
rect 5816 12038 5868 12044
rect 5828 10606 5856 12038
rect 5816 10600 5868 10606
rect 5816 10542 5868 10548
rect 5816 9580 5868 9586
rect 5816 9522 5868 9528
rect 5828 9178 5856 9522
rect 5816 9172 5868 9178
rect 5816 9114 5868 9120
rect 5722 8936 5778 8945
rect 5722 8871 5778 8880
rect 5816 8832 5868 8838
rect 5816 8774 5868 8780
rect 5828 8362 5856 8774
rect 5816 8356 5868 8362
rect 5816 8298 5868 8304
rect 5920 8090 5948 12174
rect 6012 12158 6132 12186
rect 6196 12170 6224 12786
rect 6564 12306 6592 14826
rect 6552 12300 6604 12306
rect 6552 12242 6604 12248
rect 6184 12164 6236 12170
rect 6012 11778 6040 12158
rect 6184 12106 6236 12112
rect 6144 11996 6452 12016
rect 6144 11994 6150 11996
rect 6206 11994 6230 11996
rect 6286 11994 6310 11996
rect 6366 11994 6390 11996
rect 6446 11994 6452 11996
rect 6206 11942 6208 11994
rect 6388 11942 6390 11994
rect 6144 11940 6150 11942
rect 6206 11940 6230 11942
rect 6286 11940 6310 11942
rect 6366 11940 6390 11942
rect 6446 11940 6452 11942
rect 6144 11920 6452 11940
rect 6012 11750 6132 11778
rect 6000 11688 6052 11694
rect 6000 11630 6052 11636
rect 6012 11354 6040 11630
rect 6000 11348 6052 11354
rect 6000 11290 6052 11296
rect 6104 11098 6132 11750
rect 6012 11070 6132 11098
rect 5908 8084 5960 8090
rect 5908 8026 5960 8032
rect 3547 7644 3855 7664
rect 3547 7642 3553 7644
rect 3609 7642 3633 7644
rect 3689 7642 3713 7644
rect 3769 7642 3793 7644
rect 3849 7642 3855 7644
rect 3609 7590 3611 7642
rect 3791 7590 3793 7642
rect 3547 7588 3553 7590
rect 3609 7588 3633 7590
rect 3689 7588 3713 7590
rect 3769 7588 3793 7590
rect 3849 7588 3855 7590
rect 3547 7568 3855 7588
rect 2248 7100 2556 7120
rect 2248 7098 2254 7100
rect 2310 7098 2334 7100
rect 2390 7098 2414 7100
rect 2470 7098 2494 7100
rect 2550 7098 2556 7100
rect 2310 7046 2312 7098
rect 2492 7046 2494 7098
rect 2248 7044 2254 7046
rect 2310 7044 2334 7046
rect 2390 7044 2414 7046
rect 2470 7044 2494 7046
rect 2550 7044 2556 7046
rect 2248 7024 2556 7044
rect 4846 7100 5154 7120
rect 4846 7098 4852 7100
rect 4908 7098 4932 7100
rect 4988 7098 5012 7100
rect 5068 7098 5092 7100
rect 5148 7098 5154 7100
rect 4908 7046 4910 7098
rect 5090 7046 5092 7098
rect 4846 7044 4852 7046
rect 4908 7044 4932 7046
rect 4988 7044 5012 7046
rect 5068 7044 5092 7046
rect 5148 7044 5154 7046
rect 4846 7024 5154 7044
rect 5552 6882 5580 7958
rect 5644 7942 5948 7970
rect 5724 7880 5776 7886
rect 5724 7822 5776 7828
rect 5632 7812 5684 7818
rect 5632 7754 5684 7760
rect 5644 7206 5672 7754
rect 5736 7546 5764 7822
rect 5724 7540 5776 7546
rect 5724 7482 5776 7488
rect 5632 7200 5684 7206
rect 5632 7142 5684 7148
rect 5460 6866 5580 6882
rect 5448 6860 5580 6866
rect 5500 6854 5580 6860
rect 5448 6802 5500 6808
rect 4436 6792 4488 6798
rect 4436 6734 4488 6740
rect 4448 6662 4476 6734
rect 4436 6656 4488 6662
rect 4436 6598 4488 6604
rect 3547 6556 3855 6576
rect 3547 6554 3553 6556
rect 3609 6554 3633 6556
rect 3689 6554 3713 6556
rect 3769 6554 3793 6556
rect 3849 6554 3855 6556
rect 3609 6502 3611 6554
rect 3791 6502 3793 6554
rect 3547 6500 3553 6502
rect 3609 6500 3633 6502
rect 3689 6500 3713 6502
rect 3769 6500 3793 6502
rect 3849 6500 3855 6502
rect 3547 6480 3855 6500
rect 2248 6012 2556 6032
rect 2248 6010 2254 6012
rect 2310 6010 2334 6012
rect 2390 6010 2414 6012
rect 2470 6010 2494 6012
rect 2550 6010 2556 6012
rect 2310 5958 2312 6010
rect 2492 5958 2494 6010
rect 2248 5956 2254 5958
rect 2310 5956 2334 5958
rect 2390 5956 2414 5958
rect 2470 5956 2494 5958
rect 2550 5956 2556 5958
rect 2248 5936 2556 5956
rect 3240 5636 3292 5642
rect 3240 5578 3292 5584
rect 3252 5370 3280 5578
rect 4068 5568 4120 5574
rect 4120 5516 4200 5522
rect 4068 5510 4200 5516
rect 4080 5494 4200 5510
rect 3547 5468 3855 5488
rect 3547 5466 3553 5468
rect 3609 5466 3633 5468
rect 3689 5466 3713 5468
rect 3769 5466 3793 5468
rect 3849 5466 3855 5468
rect 3609 5414 3611 5466
rect 3791 5414 3793 5466
rect 3547 5412 3553 5414
rect 3609 5412 3633 5414
rect 3689 5412 3713 5414
rect 3769 5412 3793 5414
rect 3849 5412 3855 5414
rect 3547 5392 3855 5412
rect 3240 5364 3292 5370
rect 3240 5306 3292 5312
rect 2872 5092 2924 5098
rect 2872 5034 2924 5040
rect 2248 4924 2556 4944
rect 2248 4922 2254 4924
rect 2310 4922 2334 4924
rect 2390 4922 2414 4924
rect 2470 4922 2494 4924
rect 2550 4922 2556 4924
rect 2310 4870 2312 4922
rect 2492 4870 2494 4922
rect 2248 4868 2254 4870
rect 2310 4868 2334 4870
rect 2390 4868 2414 4870
rect 2470 4868 2494 4870
rect 2550 4868 2556 4870
rect 2248 4848 2556 4868
rect 2884 4486 2912 5034
rect 3056 5024 3108 5030
rect 3056 4966 3108 4972
rect 2688 4480 2740 4486
rect 2688 4422 2740 4428
rect 2872 4480 2924 4486
rect 2872 4422 2924 4428
rect 940 4004 992 4010
rect 940 3946 992 3952
rect 952 2990 980 3946
rect 2248 3836 2556 3856
rect 2248 3834 2254 3836
rect 2310 3834 2334 3836
rect 2390 3834 2414 3836
rect 2470 3834 2494 3836
rect 2550 3834 2556 3836
rect 2310 3782 2312 3834
rect 2492 3782 2494 3834
rect 2248 3780 2254 3782
rect 2310 3780 2334 3782
rect 2390 3780 2414 3782
rect 2470 3780 2494 3782
rect 2550 3780 2556 3782
rect 2248 3760 2556 3780
rect 2700 3670 2728 4422
rect 2688 3664 2740 3670
rect 2688 3606 2740 3612
rect 2884 3398 2912 4422
rect 3068 3942 3096 4966
rect 4172 4690 4200 5494
rect 4344 5024 4396 5030
rect 4344 4966 4396 4972
rect 4160 4684 4212 4690
rect 4160 4626 4212 4632
rect 4160 4548 4212 4554
rect 4160 4490 4212 4496
rect 3547 4380 3855 4400
rect 3547 4378 3553 4380
rect 3609 4378 3633 4380
rect 3689 4378 3713 4380
rect 3769 4378 3793 4380
rect 3849 4378 3855 4380
rect 3609 4326 3611 4378
rect 3791 4326 3793 4378
rect 3547 4324 3553 4326
rect 3609 4324 3633 4326
rect 3689 4324 3713 4326
rect 3769 4324 3793 4326
rect 3849 4324 3855 4326
rect 3547 4304 3855 4324
rect 4172 4214 4200 4490
rect 4160 4208 4212 4214
rect 4160 4150 4212 4156
rect 4252 4140 4304 4146
rect 4252 4082 4304 4088
rect 3056 3936 3108 3942
rect 3056 3878 3108 3884
rect 3240 3936 3292 3942
rect 3240 3878 3292 3884
rect 3252 3670 3280 3878
rect 3240 3664 3292 3670
rect 3240 3606 3292 3612
rect 2872 3392 2924 3398
rect 2872 3334 2924 3340
rect 3884 3392 3936 3398
rect 3884 3334 3936 3340
rect 940 2984 992 2990
rect 940 2926 992 2932
rect 952 800 980 2926
rect 2248 2748 2556 2768
rect 2248 2746 2254 2748
rect 2310 2746 2334 2748
rect 2390 2746 2414 2748
rect 2470 2746 2494 2748
rect 2550 2746 2556 2748
rect 2310 2694 2312 2746
rect 2492 2694 2494 2746
rect 2248 2692 2254 2694
rect 2310 2692 2334 2694
rect 2390 2692 2414 2694
rect 2470 2692 2494 2694
rect 2550 2692 2556 2694
rect 2248 2672 2556 2692
rect 2884 800 2912 3334
rect 3547 3292 3855 3312
rect 3547 3290 3553 3292
rect 3609 3290 3633 3292
rect 3689 3290 3713 3292
rect 3769 3290 3793 3292
rect 3849 3290 3855 3292
rect 3609 3238 3611 3290
rect 3791 3238 3793 3290
rect 3547 3236 3553 3238
rect 3609 3236 3633 3238
rect 3689 3236 3713 3238
rect 3769 3236 3793 3238
rect 3849 3236 3855 3238
rect 3547 3216 3855 3236
rect 3896 2990 3924 3334
rect 4264 3194 4292 4082
rect 4356 4010 4384 4966
rect 4448 4758 4476 6598
rect 4846 6012 5154 6032
rect 4846 6010 4852 6012
rect 4908 6010 4932 6012
rect 4988 6010 5012 6012
rect 5068 6010 5092 6012
rect 5148 6010 5154 6012
rect 4908 5958 4910 6010
rect 5090 5958 5092 6010
rect 4846 5956 4852 5958
rect 4908 5956 4932 5958
rect 4988 5956 5012 5958
rect 5068 5956 5092 5958
rect 5148 5956 5154 5958
rect 4846 5936 5154 5956
rect 5552 5370 5580 6854
rect 5920 6458 5948 7942
rect 5724 6452 5776 6458
rect 5724 6394 5776 6400
rect 5908 6452 5960 6458
rect 5908 6394 5960 6400
rect 5736 5710 5764 6394
rect 6012 6361 6040 11070
rect 6656 10985 6684 17274
rect 6736 16516 6788 16522
rect 6736 16458 6788 16464
rect 6748 16250 6776 16458
rect 6736 16244 6788 16250
rect 6736 16186 6788 16192
rect 6736 16108 6788 16114
rect 6736 16050 6788 16056
rect 6748 15638 6776 16050
rect 6736 15632 6788 15638
rect 6736 15574 6788 15580
rect 6736 15020 6788 15026
rect 6736 14962 6788 14968
rect 6748 14521 6776 14962
rect 6734 14512 6790 14521
rect 6734 14447 6736 14456
rect 6788 14447 6790 14456
rect 6736 14418 6788 14424
rect 6748 14387 6776 14418
rect 6736 14340 6788 14346
rect 6736 14282 6788 14288
rect 6748 12866 6776 14282
rect 6840 12986 6868 18799
rect 7208 18766 7236 19382
rect 7443 19068 7751 19088
rect 7443 19066 7449 19068
rect 7505 19066 7529 19068
rect 7585 19066 7609 19068
rect 7665 19066 7689 19068
rect 7745 19066 7751 19068
rect 7505 19014 7507 19066
rect 7687 19014 7689 19066
rect 7443 19012 7449 19014
rect 7505 19012 7529 19014
rect 7585 19012 7609 19014
rect 7665 19012 7689 19014
rect 7745 19012 7751 19014
rect 7443 18992 7751 19012
rect 7196 18760 7248 18766
rect 7196 18702 7248 18708
rect 7288 18624 7340 18630
rect 7288 18566 7340 18572
rect 7300 17746 7328 18566
rect 7840 18148 7892 18154
rect 7840 18090 7892 18096
rect 7443 17980 7751 18000
rect 7443 17978 7449 17980
rect 7505 17978 7529 17980
rect 7585 17978 7609 17980
rect 7665 17978 7689 17980
rect 7745 17978 7751 17980
rect 7505 17926 7507 17978
rect 7687 17926 7689 17978
rect 7443 17924 7449 17926
rect 7505 17924 7529 17926
rect 7585 17924 7609 17926
rect 7665 17924 7689 17926
rect 7745 17924 7751 17926
rect 7443 17904 7751 17924
rect 7104 17740 7156 17746
rect 7104 17682 7156 17688
rect 7288 17740 7340 17746
rect 7288 17682 7340 17688
rect 6920 17604 6972 17610
rect 6920 17546 6972 17552
rect 6932 16182 6960 17546
rect 7116 16590 7144 17682
rect 7196 17672 7248 17678
rect 7196 17614 7248 17620
rect 7208 17202 7236 17614
rect 7852 17610 7880 18090
rect 7840 17604 7892 17610
rect 7840 17546 7892 17552
rect 7196 17196 7248 17202
rect 7196 17138 7248 17144
rect 7104 16584 7156 16590
rect 7104 16526 7156 16532
rect 7116 16182 7144 16526
rect 7208 16522 7236 17138
rect 7443 16892 7751 16912
rect 7443 16890 7449 16892
rect 7505 16890 7529 16892
rect 7585 16890 7609 16892
rect 7665 16890 7689 16892
rect 7745 16890 7751 16892
rect 7505 16838 7507 16890
rect 7687 16838 7689 16890
rect 7443 16836 7449 16838
rect 7505 16836 7529 16838
rect 7585 16836 7609 16838
rect 7665 16836 7689 16838
rect 7745 16836 7751 16838
rect 7443 16816 7751 16836
rect 7196 16516 7248 16522
rect 7196 16458 7248 16464
rect 6920 16176 6972 16182
rect 6920 16118 6972 16124
rect 7104 16176 7156 16182
rect 7104 16118 7156 16124
rect 6932 14414 6960 16118
rect 7012 16108 7064 16114
rect 7012 16050 7064 16056
rect 7024 15570 7052 16050
rect 7012 15564 7064 15570
rect 7012 15506 7064 15512
rect 7104 15428 7156 15434
rect 7104 15370 7156 15376
rect 7012 15020 7064 15026
rect 7012 14962 7064 14968
rect 6920 14408 6972 14414
rect 6920 14350 6972 14356
rect 7024 13938 7052 14962
rect 7012 13932 7064 13938
rect 7012 13874 7064 13880
rect 7024 13326 7052 13874
rect 7116 13530 7144 15370
rect 7208 15162 7236 16458
rect 7944 16130 7972 20590
rect 8024 20460 8076 20466
rect 8024 20402 8076 20408
rect 8036 19514 8064 20402
rect 8128 19854 8156 21354
rect 8312 21026 8340 23695
rect 8220 20998 8340 21026
rect 8220 20942 8248 20998
rect 8208 20936 8260 20942
rect 8208 20878 8260 20884
rect 8116 19848 8168 19854
rect 8116 19790 8168 19796
rect 8024 19508 8076 19514
rect 8024 19450 8076 19456
rect 8128 18290 8156 19790
rect 8116 18284 8168 18290
rect 8116 18226 8168 18232
rect 8022 16824 8078 16833
rect 8022 16759 8078 16768
rect 7852 16114 7972 16130
rect 7840 16108 7972 16114
rect 7892 16102 7972 16108
rect 7840 16050 7892 16056
rect 7443 15804 7751 15824
rect 7443 15802 7449 15804
rect 7505 15802 7529 15804
rect 7585 15802 7609 15804
rect 7665 15802 7689 15804
rect 7745 15802 7751 15804
rect 7505 15750 7507 15802
rect 7687 15750 7689 15802
rect 7443 15748 7449 15750
rect 7505 15748 7529 15750
rect 7585 15748 7609 15750
rect 7665 15748 7689 15750
rect 7745 15748 7751 15750
rect 7443 15728 7751 15748
rect 7930 15600 7986 15609
rect 7930 15535 7986 15544
rect 7288 15496 7340 15502
rect 7288 15438 7340 15444
rect 7196 15156 7248 15162
rect 7196 15098 7248 15104
rect 7300 15026 7328 15438
rect 7840 15088 7892 15094
rect 7840 15030 7892 15036
rect 7288 15020 7340 15026
rect 7288 14962 7340 14968
rect 7196 14544 7248 14550
rect 7196 14486 7248 14492
rect 7104 13524 7156 13530
rect 7104 13466 7156 13472
rect 7208 13410 7236 14486
rect 7116 13382 7236 13410
rect 7300 13410 7328 14962
rect 7443 14716 7751 14736
rect 7443 14714 7449 14716
rect 7505 14714 7529 14716
rect 7585 14714 7609 14716
rect 7665 14714 7689 14716
rect 7745 14714 7751 14716
rect 7505 14662 7507 14714
rect 7687 14662 7689 14714
rect 7443 14660 7449 14662
rect 7505 14660 7529 14662
rect 7585 14660 7609 14662
rect 7665 14660 7689 14662
rect 7745 14660 7751 14662
rect 7443 14640 7751 14660
rect 7852 13802 7880 15030
rect 7840 13796 7892 13802
rect 7840 13738 7892 13744
rect 7443 13628 7751 13648
rect 7443 13626 7449 13628
rect 7505 13626 7529 13628
rect 7585 13626 7609 13628
rect 7665 13626 7689 13628
rect 7745 13626 7751 13628
rect 7505 13574 7507 13626
rect 7687 13574 7689 13626
rect 7443 13572 7449 13574
rect 7505 13572 7529 13574
rect 7585 13572 7609 13574
rect 7665 13572 7689 13574
rect 7745 13572 7751 13574
rect 7443 13552 7751 13572
rect 7852 13462 7880 13738
rect 7840 13456 7892 13462
rect 7300 13382 7420 13410
rect 7840 13398 7892 13404
rect 7012 13320 7064 13326
rect 7012 13262 7064 13268
rect 6828 12980 6880 12986
rect 6828 12922 6880 12928
rect 6748 12838 6868 12866
rect 6736 12776 6788 12782
rect 6736 12718 6788 12724
rect 6748 12374 6776 12718
rect 6736 12368 6788 12374
rect 6736 12310 6788 12316
rect 6840 11914 6868 12838
rect 6920 12096 6972 12102
rect 6920 12038 6972 12044
rect 6748 11886 6868 11914
rect 6642 10976 6698 10985
rect 6144 10908 6452 10928
rect 6642 10911 6698 10920
rect 6144 10906 6150 10908
rect 6206 10906 6230 10908
rect 6286 10906 6310 10908
rect 6366 10906 6390 10908
rect 6446 10906 6452 10908
rect 6206 10854 6208 10906
rect 6388 10854 6390 10906
rect 6144 10852 6150 10854
rect 6206 10852 6230 10854
rect 6286 10852 6310 10854
rect 6366 10852 6390 10854
rect 6446 10852 6452 10854
rect 6144 10832 6452 10852
rect 6644 10804 6696 10810
rect 6644 10746 6696 10752
rect 6552 10668 6604 10674
rect 6552 10610 6604 10616
rect 6144 9820 6452 9840
rect 6144 9818 6150 9820
rect 6206 9818 6230 9820
rect 6286 9818 6310 9820
rect 6366 9818 6390 9820
rect 6446 9818 6452 9820
rect 6206 9766 6208 9818
rect 6388 9766 6390 9818
rect 6144 9764 6150 9766
rect 6206 9764 6230 9766
rect 6286 9764 6310 9766
rect 6366 9764 6390 9766
rect 6446 9764 6452 9766
rect 6144 9744 6452 9764
rect 6144 8732 6452 8752
rect 6144 8730 6150 8732
rect 6206 8730 6230 8732
rect 6286 8730 6310 8732
rect 6366 8730 6390 8732
rect 6446 8730 6452 8732
rect 6206 8678 6208 8730
rect 6388 8678 6390 8730
rect 6144 8676 6150 8678
rect 6206 8676 6230 8678
rect 6286 8676 6310 8678
rect 6366 8676 6390 8678
rect 6446 8676 6452 8678
rect 6144 8656 6452 8676
rect 6564 8430 6592 10610
rect 6656 9586 6684 10746
rect 6644 9580 6696 9586
rect 6644 9522 6696 9528
rect 6656 9042 6684 9522
rect 6644 9036 6696 9042
rect 6644 8978 6696 8984
rect 6552 8424 6604 8430
rect 6552 8366 6604 8372
rect 6460 8356 6512 8362
rect 6460 8298 6512 8304
rect 6472 8242 6500 8298
rect 6472 8214 6592 8242
rect 6144 7644 6452 7664
rect 6144 7642 6150 7644
rect 6206 7642 6230 7644
rect 6286 7642 6310 7644
rect 6366 7642 6390 7644
rect 6446 7642 6452 7644
rect 6206 7590 6208 7642
rect 6388 7590 6390 7642
rect 6144 7588 6150 7590
rect 6206 7588 6230 7590
rect 6286 7588 6310 7590
rect 6366 7588 6390 7590
rect 6446 7588 6452 7590
rect 6144 7568 6452 7588
rect 6564 7290 6592 8214
rect 6748 7585 6776 11886
rect 6828 11756 6880 11762
rect 6828 11698 6880 11704
rect 6840 11286 6868 11698
rect 6932 11642 6960 12038
rect 7024 11830 7052 13262
rect 7116 12102 7144 13382
rect 7288 13252 7340 13258
rect 7288 13194 7340 13200
rect 7300 12986 7328 13194
rect 7392 12986 7420 13382
rect 7288 12980 7340 12986
rect 7288 12922 7340 12928
rect 7380 12980 7432 12986
rect 7380 12922 7432 12928
rect 7196 12844 7248 12850
rect 7196 12786 7248 12792
rect 7104 12096 7156 12102
rect 7104 12038 7156 12044
rect 7012 11824 7064 11830
rect 7012 11766 7064 11772
rect 6932 11614 7052 11642
rect 6828 11280 6880 11286
rect 6828 11222 6880 11228
rect 6920 9988 6972 9994
rect 6920 9930 6972 9936
rect 6828 8832 6880 8838
rect 6828 8774 6880 8780
rect 6734 7576 6790 7585
rect 6734 7511 6790 7520
rect 6564 7262 6776 7290
rect 6460 7200 6512 7206
rect 6460 7142 6512 7148
rect 6472 6798 6500 7142
rect 6460 6792 6512 6798
rect 6512 6740 6592 6746
rect 6460 6734 6592 6740
rect 6472 6718 6592 6734
rect 6144 6556 6452 6576
rect 6144 6554 6150 6556
rect 6206 6554 6230 6556
rect 6286 6554 6310 6556
rect 6366 6554 6390 6556
rect 6446 6554 6452 6556
rect 6206 6502 6208 6554
rect 6388 6502 6390 6554
rect 6144 6500 6150 6502
rect 6206 6500 6230 6502
rect 6286 6500 6310 6502
rect 6366 6500 6390 6502
rect 6446 6500 6452 6502
rect 6144 6480 6452 6500
rect 5998 6352 6054 6361
rect 5908 6316 5960 6322
rect 5998 6287 6054 6296
rect 5908 6258 5960 6264
rect 5816 6112 5868 6118
rect 5816 6054 5868 6060
rect 5724 5704 5776 5710
rect 5724 5646 5776 5652
rect 5540 5364 5592 5370
rect 5540 5306 5592 5312
rect 5172 5228 5224 5234
rect 5172 5170 5224 5176
rect 4712 5160 4764 5166
rect 4712 5102 4764 5108
rect 4436 4752 4488 4758
rect 4436 4694 4488 4700
rect 4620 4684 4672 4690
rect 4620 4626 4672 4632
rect 4528 4616 4580 4622
rect 4528 4558 4580 4564
rect 4436 4276 4488 4282
rect 4436 4218 4488 4224
rect 4344 4004 4396 4010
rect 4344 3946 4396 3952
rect 4252 3188 4304 3194
rect 4252 3130 4304 3136
rect 3884 2984 3936 2990
rect 3884 2926 3936 2932
rect 3056 2916 3108 2922
rect 3056 2858 3108 2864
rect 3068 2650 3096 2858
rect 4356 2774 4384 3946
rect 4448 2990 4476 4218
rect 4540 3126 4568 4558
rect 4632 3942 4660 4626
rect 4620 3936 4672 3942
rect 4620 3878 4672 3884
rect 4632 3482 4660 3878
rect 4724 3602 4752 5102
rect 4846 4924 5154 4944
rect 4846 4922 4852 4924
rect 4908 4922 4932 4924
rect 4988 4922 5012 4924
rect 5068 4922 5092 4924
rect 5148 4922 5154 4924
rect 4908 4870 4910 4922
rect 5090 4870 5092 4922
rect 4846 4868 4852 4870
rect 4908 4868 4932 4870
rect 4988 4868 5012 4870
rect 5068 4868 5092 4870
rect 5148 4868 5154 4870
rect 4846 4848 5154 4868
rect 4804 4752 4856 4758
rect 4804 4694 4856 4700
rect 4816 4078 4844 4694
rect 5184 4282 5212 5170
rect 5448 4480 5500 4486
rect 5448 4422 5500 4428
rect 5172 4276 5224 4282
rect 5172 4218 5224 4224
rect 4804 4072 4856 4078
rect 4804 4014 4856 4020
rect 5172 4004 5224 4010
rect 5172 3946 5224 3952
rect 4846 3836 5154 3856
rect 4846 3834 4852 3836
rect 4908 3834 4932 3836
rect 4988 3834 5012 3836
rect 5068 3834 5092 3836
rect 5148 3834 5154 3836
rect 4908 3782 4910 3834
rect 5090 3782 5092 3834
rect 4846 3780 4852 3782
rect 4908 3780 4932 3782
rect 4988 3780 5012 3782
rect 5068 3780 5092 3782
rect 5148 3780 5154 3782
rect 4846 3760 5154 3780
rect 4712 3596 4764 3602
rect 4712 3538 4764 3544
rect 4632 3466 4752 3482
rect 4632 3460 4764 3466
rect 4632 3454 4712 3460
rect 4712 3402 4764 3408
rect 4528 3120 4580 3126
rect 4528 3062 4580 3068
rect 4436 2984 4488 2990
rect 4436 2926 4488 2932
rect 4264 2746 4384 2774
rect 3056 2644 3108 2650
rect 3056 2586 3108 2592
rect 4264 2514 4292 2746
rect 4252 2508 4304 2514
rect 4252 2450 4304 2456
rect 4540 2446 4568 3062
rect 4528 2440 4580 2446
rect 4528 2382 4580 2388
rect 4724 2378 4752 3402
rect 4846 2748 5154 2768
rect 4846 2746 4852 2748
rect 4908 2746 4932 2748
rect 4988 2746 5012 2748
rect 5068 2746 5092 2748
rect 5148 2746 5154 2748
rect 4908 2694 4910 2746
rect 5090 2694 5092 2746
rect 4846 2692 4852 2694
rect 4908 2692 4932 2694
rect 4988 2692 5012 2694
rect 5068 2692 5092 2694
rect 5148 2692 5154 2694
rect 4846 2672 5154 2692
rect 5184 2514 5212 3946
rect 5356 3936 5408 3942
rect 5356 3878 5408 3884
rect 5368 3194 5396 3878
rect 5460 3602 5488 4422
rect 5552 4282 5580 5306
rect 5828 4690 5856 6054
rect 5920 5642 5948 6258
rect 6564 6118 6592 6718
rect 6000 6112 6052 6118
rect 6000 6054 6052 6060
rect 6552 6112 6604 6118
rect 6552 6054 6604 6060
rect 5908 5636 5960 5642
rect 5908 5578 5960 5584
rect 5920 5302 5948 5578
rect 5908 5296 5960 5302
rect 5908 5238 5960 5244
rect 5816 4684 5868 4690
rect 5816 4626 5868 4632
rect 6012 4486 6040 6054
rect 6368 5908 6420 5914
rect 6368 5850 6420 5856
rect 6380 5710 6408 5850
rect 6368 5704 6420 5710
rect 6368 5646 6420 5652
rect 6144 5468 6452 5488
rect 6144 5466 6150 5468
rect 6206 5466 6230 5468
rect 6286 5466 6310 5468
rect 6366 5466 6390 5468
rect 6446 5466 6452 5468
rect 6206 5414 6208 5466
rect 6388 5414 6390 5466
rect 6144 5412 6150 5414
rect 6206 5412 6230 5414
rect 6286 5412 6310 5414
rect 6366 5412 6390 5414
rect 6446 5412 6452 5414
rect 6144 5392 6452 5412
rect 6552 5228 6604 5234
rect 6552 5170 6604 5176
rect 6564 4486 6592 5170
rect 6000 4480 6052 4486
rect 6000 4422 6052 4428
rect 6552 4480 6604 4486
rect 6552 4422 6604 4428
rect 5540 4276 5592 4282
rect 5540 4218 5592 4224
rect 5540 4072 5592 4078
rect 5540 4014 5592 4020
rect 5552 3738 5580 4014
rect 5540 3732 5592 3738
rect 5540 3674 5592 3680
rect 5448 3596 5500 3602
rect 5448 3538 5500 3544
rect 5460 3194 5488 3538
rect 5724 3460 5776 3466
rect 5724 3402 5776 3408
rect 5356 3188 5408 3194
rect 5356 3130 5408 3136
rect 5448 3188 5500 3194
rect 5448 3130 5500 3136
rect 5172 2508 5224 2514
rect 5172 2450 5224 2456
rect 5460 2446 5488 3130
rect 5736 2650 5764 3402
rect 6012 3398 6040 4422
rect 6144 4380 6452 4400
rect 6144 4378 6150 4380
rect 6206 4378 6230 4380
rect 6286 4378 6310 4380
rect 6366 4378 6390 4380
rect 6446 4378 6452 4380
rect 6206 4326 6208 4378
rect 6388 4326 6390 4378
rect 6144 4324 6150 4326
rect 6206 4324 6230 4326
rect 6286 4324 6310 4326
rect 6366 4324 6390 4326
rect 6446 4324 6452 4326
rect 6144 4304 6452 4324
rect 6564 4214 6592 4422
rect 6552 4208 6604 4214
rect 6552 4150 6604 4156
rect 6748 4049 6776 7262
rect 6840 6866 6868 8774
rect 6932 8566 6960 9930
rect 7024 8922 7052 11614
rect 7208 11150 7236 12786
rect 7840 12640 7892 12646
rect 7840 12582 7892 12588
rect 7443 12540 7751 12560
rect 7443 12538 7449 12540
rect 7505 12538 7529 12540
rect 7585 12538 7609 12540
rect 7665 12538 7689 12540
rect 7745 12538 7751 12540
rect 7505 12486 7507 12538
rect 7687 12486 7689 12538
rect 7443 12484 7449 12486
rect 7505 12484 7529 12486
rect 7585 12484 7609 12486
rect 7665 12484 7689 12486
rect 7745 12484 7751 12486
rect 7443 12464 7751 12484
rect 7852 12306 7880 12582
rect 7840 12300 7892 12306
rect 7840 12242 7892 12248
rect 7288 12164 7340 12170
rect 7288 12106 7340 12112
rect 7196 11144 7248 11150
rect 7196 11086 7248 11092
rect 7208 10674 7236 11086
rect 7300 11082 7328 12106
rect 7443 11452 7751 11472
rect 7443 11450 7449 11452
rect 7505 11450 7529 11452
rect 7585 11450 7609 11452
rect 7665 11450 7689 11452
rect 7745 11450 7751 11452
rect 7505 11398 7507 11450
rect 7687 11398 7689 11450
rect 7443 11396 7449 11398
rect 7505 11396 7529 11398
rect 7585 11396 7609 11398
rect 7665 11396 7689 11398
rect 7745 11396 7751 11398
rect 7443 11376 7751 11396
rect 7288 11076 7340 11082
rect 7288 11018 7340 11024
rect 7300 10742 7328 11018
rect 7944 10810 7972 15535
rect 8036 12434 8064 16759
rect 8116 15564 8168 15570
rect 8116 15506 8168 15512
rect 8128 15026 8156 15506
rect 8116 15020 8168 15026
rect 8116 14962 8168 14968
rect 8208 12912 8260 12918
rect 8208 12854 8260 12860
rect 8036 12406 8156 12434
rect 7932 10804 7984 10810
rect 7932 10746 7984 10752
rect 7288 10736 7340 10742
rect 7288 10678 7340 10684
rect 7196 10668 7248 10674
rect 7196 10610 7248 10616
rect 7443 10364 7751 10384
rect 7443 10362 7449 10364
rect 7505 10362 7529 10364
rect 7585 10362 7609 10364
rect 7665 10362 7689 10364
rect 7745 10362 7751 10364
rect 7505 10310 7507 10362
rect 7687 10310 7689 10362
rect 7443 10308 7449 10310
rect 7505 10308 7529 10310
rect 7585 10308 7609 10310
rect 7665 10308 7689 10310
rect 7745 10308 7751 10310
rect 7443 10288 7751 10308
rect 7288 10056 7340 10062
rect 7288 9998 7340 10004
rect 7104 9580 7156 9586
rect 7104 9522 7156 9528
rect 7116 9110 7144 9522
rect 7196 9376 7248 9382
rect 7196 9318 7248 9324
rect 7104 9104 7156 9110
rect 7104 9046 7156 9052
rect 7208 9042 7236 9318
rect 7196 9036 7248 9042
rect 7196 8978 7248 8984
rect 7024 8906 7144 8922
rect 7024 8900 7156 8906
rect 7024 8894 7104 8900
rect 7104 8842 7156 8848
rect 6920 8560 6972 8566
rect 6920 8502 6972 8508
rect 7116 7478 7144 8842
rect 7196 8492 7248 8498
rect 7196 8434 7248 8440
rect 7208 7818 7236 8434
rect 7300 7886 7328 9998
rect 7932 9920 7984 9926
rect 7932 9862 7984 9868
rect 7840 9580 7892 9586
rect 7840 9522 7892 9528
rect 7443 9276 7751 9296
rect 7443 9274 7449 9276
rect 7505 9274 7529 9276
rect 7585 9274 7609 9276
rect 7665 9274 7689 9276
rect 7745 9274 7751 9276
rect 7505 9222 7507 9274
rect 7687 9222 7689 9274
rect 7443 9220 7449 9222
rect 7505 9220 7529 9222
rect 7585 9220 7609 9222
rect 7665 9220 7689 9222
rect 7745 9220 7751 9222
rect 7443 9200 7751 9220
rect 7852 8838 7880 9522
rect 7840 8832 7892 8838
rect 7840 8774 7892 8780
rect 7443 8188 7751 8208
rect 7443 8186 7449 8188
rect 7505 8186 7529 8188
rect 7585 8186 7609 8188
rect 7665 8186 7689 8188
rect 7745 8186 7751 8188
rect 7505 8134 7507 8186
rect 7687 8134 7689 8186
rect 7443 8132 7449 8134
rect 7505 8132 7529 8134
rect 7585 8132 7609 8134
rect 7665 8132 7689 8134
rect 7745 8132 7751 8134
rect 7443 8112 7751 8132
rect 7288 7880 7340 7886
rect 7288 7822 7340 7828
rect 7196 7812 7248 7818
rect 7196 7754 7248 7760
rect 7288 7744 7340 7750
rect 7288 7686 7340 7692
rect 7104 7472 7156 7478
rect 7104 7414 7156 7420
rect 6828 6860 6880 6866
rect 6828 6802 6880 6808
rect 7104 6316 7156 6322
rect 7104 6258 7156 6264
rect 7012 6180 7064 6186
rect 7012 6122 7064 6128
rect 6920 5772 6972 5778
rect 6920 5714 6972 5720
rect 6932 5250 6960 5714
rect 7024 5642 7052 6122
rect 7116 5710 7144 6258
rect 7196 5840 7248 5846
rect 7196 5782 7248 5788
rect 7104 5704 7156 5710
rect 7104 5646 7156 5652
rect 7012 5636 7064 5642
rect 7012 5578 7064 5584
rect 6932 5222 7052 5250
rect 6920 5092 6972 5098
rect 6920 5034 6972 5040
rect 6828 4548 6880 4554
rect 6828 4490 6880 4496
rect 6734 4040 6790 4049
rect 6734 3975 6790 3984
rect 6736 3732 6788 3738
rect 6736 3674 6788 3680
rect 6000 3392 6052 3398
rect 6000 3334 6052 3340
rect 6012 2854 6040 3334
rect 6144 3292 6452 3312
rect 6144 3290 6150 3292
rect 6206 3290 6230 3292
rect 6286 3290 6310 3292
rect 6366 3290 6390 3292
rect 6446 3290 6452 3292
rect 6206 3238 6208 3290
rect 6388 3238 6390 3290
rect 6144 3236 6150 3238
rect 6206 3236 6230 3238
rect 6286 3236 6310 3238
rect 6366 3236 6390 3238
rect 6446 3236 6452 3238
rect 6144 3216 6452 3236
rect 6552 3052 6604 3058
rect 6552 2994 6604 3000
rect 6564 2922 6592 2994
rect 6552 2916 6604 2922
rect 6552 2858 6604 2864
rect 6000 2848 6052 2854
rect 6000 2790 6052 2796
rect 5724 2644 5776 2650
rect 5724 2586 5776 2592
rect 6564 2582 6592 2858
rect 6552 2576 6604 2582
rect 6552 2518 6604 2524
rect 6748 2446 6776 3674
rect 6840 2514 6868 4490
rect 6828 2508 6880 2514
rect 6828 2450 6880 2456
rect 4896 2440 4948 2446
rect 4896 2382 4948 2388
rect 5448 2440 5500 2446
rect 5448 2382 5500 2388
rect 6736 2440 6788 2446
rect 6736 2382 6788 2388
rect 4712 2372 4764 2378
rect 4712 2314 4764 2320
rect 3547 2204 3855 2224
rect 3547 2202 3553 2204
rect 3609 2202 3633 2204
rect 3689 2202 3713 2204
rect 3769 2202 3793 2204
rect 3849 2202 3855 2204
rect 3609 2150 3611 2202
rect 3791 2150 3793 2202
rect 3547 2148 3553 2150
rect 3609 2148 3633 2150
rect 3689 2148 3713 2150
rect 3769 2148 3793 2150
rect 3849 2148 3855 2150
rect 3547 2128 3855 2148
rect 4908 800 4936 2382
rect 6144 2204 6452 2224
rect 6144 2202 6150 2204
rect 6206 2202 6230 2204
rect 6286 2202 6310 2204
rect 6366 2202 6390 2204
rect 6446 2202 6452 2204
rect 6206 2150 6208 2202
rect 6388 2150 6390 2202
rect 6144 2148 6150 2150
rect 6206 2148 6230 2150
rect 6286 2148 6310 2150
rect 6366 2148 6390 2150
rect 6446 2148 6452 2150
rect 6144 2128 6452 2148
rect 6932 800 6960 5034
rect 7024 2446 7052 5222
rect 7116 3058 7144 5646
rect 7208 5234 7236 5782
rect 7300 5370 7328 7686
rect 7852 7410 7880 8774
rect 7944 7954 7972 9862
rect 7932 7948 7984 7954
rect 7932 7890 7984 7896
rect 7840 7404 7892 7410
rect 7840 7346 7892 7352
rect 7932 7336 7984 7342
rect 7932 7278 7984 7284
rect 7840 7268 7892 7274
rect 7840 7210 7892 7216
rect 7443 7100 7751 7120
rect 7443 7098 7449 7100
rect 7505 7098 7529 7100
rect 7585 7098 7609 7100
rect 7665 7098 7689 7100
rect 7745 7098 7751 7100
rect 7505 7046 7507 7098
rect 7687 7046 7689 7098
rect 7443 7044 7449 7046
rect 7505 7044 7529 7046
rect 7585 7044 7609 7046
rect 7665 7044 7689 7046
rect 7745 7044 7751 7046
rect 7443 7024 7751 7044
rect 7852 6730 7880 7210
rect 7944 6798 7972 7278
rect 7932 6792 7984 6798
rect 7932 6734 7984 6740
rect 7472 6724 7524 6730
rect 7472 6666 7524 6672
rect 7840 6724 7892 6730
rect 7840 6666 7892 6672
rect 7484 6390 7512 6666
rect 7472 6384 7524 6390
rect 7472 6326 7524 6332
rect 7443 6012 7751 6032
rect 7443 6010 7449 6012
rect 7505 6010 7529 6012
rect 7585 6010 7609 6012
rect 7665 6010 7689 6012
rect 7745 6010 7751 6012
rect 7505 5958 7507 6010
rect 7687 5958 7689 6010
rect 7443 5956 7449 5958
rect 7505 5956 7529 5958
rect 7585 5956 7609 5958
rect 7665 5956 7689 5958
rect 7745 5956 7751 5958
rect 7443 5936 7751 5956
rect 7288 5364 7340 5370
rect 7288 5306 7340 5312
rect 7196 5228 7248 5234
rect 7196 5170 7248 5176
rect 7208 4146 7236 5170
rect 7443 4924 7751 4944
rect 7443 4922 7449 4924
rect 7505 4922 7529 4924
rect 7585 4922 7609 4924
rect 7665 4922 7689 4924
rect 7745 4922 7751 4924
rect 7505 4870 7507 4922
rect 7687 4870 7689 4922
rect 7443 4868 7449 4870
rect 7505 4868 7529 4870
rect 7585 4868 7609 4870
rect 7665 4868 7689 4870
rect 7745 4868 7751 4870
rect 7443 4848 7751 4868
rect 7196 4140 7248 4146
rect 7196 4082 7248 4088
rect 7208 3602 7236 4082
rect 7443 3836 7751 3856
rect 7443 3834 7449 3836
rect 7505 3834 7529 3836
rect 7585 3834 7609 3836
rect 7665 3834 7689 3836
rect 7745 3834 7751 3836
rect 7505 3782 7507 3834
rect 7687 3782 7689 3834
rect 7443 3780 7449 3782
rect 7505 3780 7529 3782
rect 7585 3780 7609 3782
rect 7665 3780 7689 3782
rect 7745 3780 7751 3782
rect 7443 3760 7751 3780
rect 7196 3596 7248 3602
rect 7196 3538 7248 3544
rect 7104 3052 7156 3058
rect 7104 2994 7156 3000
rect 7196 2916 7248 2922
rect 7196 2858 7248 2864
rect 7208 2514 7236 2858
rect 7443 2748 7751 2768
rect 7443 2746 7449 2748
rect 7505 2746 7529 2748
rect 7585 2746 7609 2748
rect 7665 2746 7689 2748
rect 7745 2746 7751 2748
rect 7505 2694 7507 2746
rect 7687 2694 7689 2746
rect 7443 2692 7449 2694
rect 7505 2692 7529 2694
rect 7585 2692 7609 2694
rect 7665 2692 7689 2694
rect 7745 2692 7751 2694
rect 7443 2672 7751 2692
rect 7196 2508 7248 2514
rect 7196 2450 7248 2456
rect 7012 2440 7064 2446
rect 7012 2382 7064 2388
rect 7656 2440 7708 2446
rect 7656 2382 7708 2388
rect 7668 1737 7696 2382
rect 7654 1728 7710 1737
rect 7654 1663 7710 1672
rect 938 0 994 800
rect 2870 0 2926 800
rect 4894 0 4950 800
rect 6918 0 6974 800
rect 7944 649 7972 6734
rect 8128 6118 8156 12406
rect 8220 10062 8248 12854
rect 8300 11688 8352 11694
rect 8300 11630 8352 11636
rect 8312 11150 8340 11630
rect 8300 11144 8352 11150
rect 8300 11086 8352 11092
rect 8208 10056 8260 10062
rect 8208 9998 8260 10004
rect 8116 6112 8168 6118
rect 8116 6054 8168 6060
rect 8024 5908 8076 5914
rect 8024 5850 8076 5856
rect 8036 5234 8064 5850
rect 8128 5710 8156 6054
rect 8116 5704 8168 5710
rect 8116 5646 8168 5652
rect 8312 5273 8340 11086
rect 8298 5264 8354 5273
rect 8024 5228 8076 5234
rect 8298 5199 8354 5208
rect 8024 5170 8076 5176
rect 8116 5024 8168 5030
rect 8116 4966 8168 4972
rect 8128 4622 8156 4966
rect 8116 4616 8168 4622
rect 8116 4558 8168 4564
rect 8128 4146 8156 4558
rect 8116 4140 8168 4146
rect 8116 4082 8168 4088
rect 8024 3460 8076 3466
rect 8024 3402 8076 3408
rect 8036 2922 8064 3402
rect 8128 2961 8156 4082
rect 8944 3392 8996 3398
rect 8944 3334 8996 3340
rect 8114 2952 8170 2961
rect 8024 2916 8076 2922
rect 8114 2887 8170 2896
rect 8024 2858 8076 2864
rect 8956 800 8984 3334
rect 7930 640 7986 649
rect 7930 575 7986 584
rect 8942 0 8998 800
<< via2 >>
rect 8206 29416 8262 29472
rect 5538 28328 5594 28384
rect 2254 27770 2310 27772
rect 2334 27770 2390 27772
rect 2414 27770 2470 27772
rect 2494 27770 2550 27772
rect 2254 27718 2300 27770
rect 2300 27718 2310 27770
rect 2334 27718 2364 27770
rect 2364 27718 2376 27770
rect 2376 27718 2390 27770
rect 2414 27718 2428 27770
rect 2428 27718 2440 27770
rect 2440 27718 2470 27770
rect 2494 27718 2504 27770
rect 2504 27718 2550 27770
rect 2254 27716 2310 27718
rect 2334 27716 2390 27718
rect 2414 27716 2470 27718
rect 2494 27716 2550 27718
rect 4852 27770 4908 27772
rect 4932 27770 4988 27772
rect 5012 27770 5068 27772
rect 5092 27770 5148 27772
rect 4852 27718 4898 27770
rect 4898 27718 4908 27770
rect 4932 27718 4962 27770
rect 4962 27718 4974 27770
rect 4974 27718 4988 27770
rect 5012 27718 5026 27770
rect 5026 27718 5038 27770
rect 5038 27718 5068 27770
rect 5092 27718 5102 27770
rect 5102 27718 5148 27770
rect 4852 27716 4908 27718
rect 4932 27716 4988 27718
rect 5012 27716 5068 27718
rect 5092 27716 5148 27718
rect 3553 27226 3609 27228
rect 3633 27226 3689 27228
rect 3713 27226 3769 27228
rect 3793 27226 3849 27228
rect 3553 27174 3599 27226
rect 3599 27174 3609 27226
rect 3633 27174 3663 27226
rect 3663 27174 3675 27226
rect 3675 27174 3689 27226
rect 3713 27174 3727 27226
rect 3727 27174 3739 27226
rect 3739 27174 3769 27226
rect 3793 27174 3803 27226
rect 3803 27174 3849 27226
rect 3553 27172 3609 27174
rect 3633 27172 3689 27174
rect 3713 27172 3769 27174
rect 3793 27172 3849 27174
rect 2254 26682 2310 26684
rect 2334 26682 2390 26684
rect 2414 26682 2470 26684
rect 2494 26682 2550 26684
rect 2254 26630 2300 26682
rect 2300 26630 2310 26682
rect 2334 26630 2364 26682
rect 2364 26630 2376 26682
rect 2376 26630 2390 26682
rect 2414 26630 2428 26682
rect 2428 26630 2440 26682
rect 2440 26630 2470 26682
rect 2494 26630 2504 26682
rect 2504 26630 2550 26682
rect 2254 26628 2310 26630
rect 2334 26628 2390 26630
rect 2414 26628 2470 26630
rect 2494 26628 2550 26630
rect 4852 26682 4908 26684
rect 4932 26682 4988 26684
rect 5012 26682 5068 26684
rect 5092 26682 5148 26684
rect 4852 26630 4898 26682
rect 4898 26630 4908 26682
rect 4932 26630 4962 26682
rect 4962 26630 4974 26682
rect 4974 26630 4988 26682
rect 5012 26630 5026 26682
rect 5026 26630 5038 26682
rect 5038 26630 5068 26682
rect 5092 26630 5102 26682
rect 5102 26630 5148 26682
rect 4852 26628 4908 26630
rect 4932 26628 4988 26630
rect 5012 26628 5068 26630
rect 5092 26628 5148 26630
rect 3553 26138 3609 26140
rect 3633 26138 3689 26140
rect 3713 26138 3769 26140
rect 3793 26138 3849 26140
rect 3553 26086 3599 26138
rect 3599 26086 3609 26138
rect 3633 26086 3663 26138
rect 3663 26086 3675 26138
rect 3675 26086 3689 26138
rect 3713 26086 3727 26138
rect 3727 26086 3739 26138
rect 3739 26086 3769 26138
rect 3793 26086 3803 26138
rect 3803 26086 3849 26138
rect 3553 26084 3609 26086
rect 3633 26084 3689 26086
rect 3713 26084 3769 26086
rect 3793 26084 3849 26086
rect 2254 25594 2310 25596
rect 2334 25594 2390 25596
rect 2414 25594 2470 25596
rect 2494 25594 2550 25596
rect 2254 25542 2300 25594
rect 2300 25542 2310 25594
rect 2334 25542 2364 25594
rect 2364 25542 2376 25594
rect 2376 25542 2390 25594
rect 2414 25542 2428 25594
rect 2428 25542 2440 25594
rect 2440 25542 2470 25594
rect 2494 25542 2504 25594
rect 2504 25542 2550 25594
rect 2254 25540 2310 25542
rect 2334 25540 2390 25542
rect 2414 25540 2470 25542
rect 2494 25540 2550 25542
rect 4852 25594 4908 25596
rect 4932 25594 4988 25596
rect 5012 25594 5068 25596
rect 5092 25594 5148 25596
rect 4852 25542 4898 25594
rect 4898 25542 4908 25594
rect 4932 25542 4962 25594
rect 4962 25542 4974 25594
rect 4974 25542 4988 25594
rect 5012 25542 5026 25594
rect 5026 25542 5038 25594
rect 5038 25542 5068 25594
rect 5092 25542 5102 25594
rect 5102 25542 5148 25594
rect 4852 25540 4908 25542
rect 4932 25540 4988 25542
rect 5012 25540 5068 25542
rect 5092 25540 5148 25542
rect 3553 25050 3609 25052
rect 3633 25050 3689 25052
rect 3713 25050 3769 25052
rect 3793 25050 3849 25052
rect 3553 24998 3599 25050
rect 3599 24998 3609 25050
rect 3633 24998 3663 25050
rect 3663 24998 3675 25050
rect 3675 24998 3689 25050
rect 3713 24998 3727 25050
rect 3727 24998 3739 25050
rect 3739 24998 3769 25050
rect 3793 24998 3803 25050
rect 3803 24998 3849 25050
rect 3553 24996 3609 24998
rect 3633 24996 3689 24998
rect 3713 24996 3769 24998
rect 3793 24996 3849 24998
rect 2254 24506 2310 24508
rect 2334 24506 2390 24508
rect 2414 24506 2470 24508
rect 2494 24506 2550 24508
rect 2254 24454 2300 24506
rect 2300 24454 2310 24506
rect 2334 24454 2364 24506
rect 2364 24454 2376 24506
rect 2376 24454 2390 24506
rect 2414 24454 2428 24506
rect 2428 24454 2440 24506
rect 2440 24454 2470 24506
rect 2494 24454 2504 24506
rect 2504 24454 2550 24506
rect 2254 24452 2310 24454
rect 2334 24452 2390 24454
rect 2414 24452 2470 24454
rect 2494 24452 2550 24454
rect 4852 24506 4908 24508
rect 4932 24506 4988 24508
rect 5012 24506 5068 24508
rect 5092 24506 5148 24508
rect 4852 24454 4898 24506
rect 4898 24454 4908 24506
rect 4932 24454 4962 24506
rect 4962 24454 4974 24506
rect 4974 24454 4988 24506
rect 5012 24454 5026 24506
rect 5026 24454 5038 24506
rect 5038 24454 5068 24506
rect 5092 24454 5102 24506
rect 5102 24454 5148 24506
rect 4852 24452 4908 24454
rect 4932 24452 4988 24454
rect 5012 24452 5068 24454
rect 5092 24452 5148 24454
rect 3553 23962 3609 23964
rect 3633 23962 3689 23964
rect 3713 23962 3769 23964
rect 3793 23962 3849 23964
rect 3553 23910 3599 23962
rect 3599 23910 3609 23962
rect 3633 23910 3663 23962
rect 3663 23910 3675 23962
rect 3675 23910 3689 23962
rect 3713 23910 3727 23962
rect 3727 23910 3739 23962
rect 3739 23910 3769 23962
rect 3793 23910 3803 23962
rect 3803 23910 3849 23962
rect 3553 23908 3609 23910
rect 3633 23908 3689 23910
rect 3713 23908 3769 23910
rect 3793 23908 3849 23910
rect 2254 23418 2310 23420
rect 2334 23418 2390 23420
rect 2414 23418 2470 23420
rect 2494 23418 2550 23420
rect 2254 23366 2300 23418
rect 2300 23366 2310 23418
rect 2334 23366 2364 23418
rect 2364 23366 2376 23418
rect 2376 23366 2390 23418
rect 2414 23366 2428 23418
rect 2428 23366 2440 23418
rect 2440 23366 2470 23418
rect 2494 23366 2504 23418
rect 2504 23366 2550 23418
rect 2254 23364 2310 23366
rect 2334 23364 2390 23366
rect 2414 23364 2470 23366
rect 2494 23364 2550 23366
rect 4852 23418 4908 23420
rect 4932 23418 4988 23420
rect 5012 23418 5068 23420
rect 5092 23418 5148 23420
rect 4852 23366 4898 23418
rect 4898 23366 4908 23418
rect 4932 23366 4962 23418
rect 4962 23366 4974 23418
rect 4974 23366 4988 23418
rect 5012 23366 5026 23418
rect 5026 23366 5038 23418
rect 5038 23366 5068 23418
rect 5092 23366 5102 23418
rect 5102 23366 5148 23418
rect 4852 23364 4908 23366
rect 4932 23364 4988 23366
rect 5012 23364 5068 23366
rect 5092 23364 5148 23366
rect 3553 22874 3609 22876
rect 3633 22874 3689 22876
rect 3713 22874 3769 22876
rect 3793 22874 3849 22876
rect 3553 22822 3599 22874
rect 3599 22822 3609 22874
rect 3633 22822 3663 22874
rect 3663 22822 3675 22874
rect 3675 22822 3689 22874
rect 3713 22822 3727 22874
rect 3727 22822 3739 22874
rect 3739 22822 3769 22874
rect 3793 22822 3803 22874
rect 3803 22822 3849 22874
rect 3553 22820 3609 22822
rect 3633 22820 3689 22822
rect 3713 22820 3769 22822
rect 3793 22820 3849 22822
rect 2254 22330 2310 22332
rect 2334 22330 2390 22332
rect 2414 22330 2470 22332
rect 2494 22330 2550 22332
rect 2254 22278 2300 22330
rect 2300 22278 2310 22330
rect 2334 22278 2364 22330
rect 2364 22278 2376 22330
rect 2376 22278 2390 22330
rect 2414 22278 2428 22330
rect 2428 22278 2440 22330
rect 2440 22278 2470 22330
rect 2494 22278 2504 22330
rect 2504 22278 2550 22330
rect 2254 22276 2310 22278
rect 2334 22276 2390 22278
rect 2414 22276 2470 22278
rect 2494 22276 2550 22278
rect 4852 22330 4908 22332
rect 4932 22330 4988 22332
rect 5012 22330 5068 22332
rect 5092 22330 5148 22332
rect 4852 22278 4898 22330
rect 4898 22278 4908 22330
rect 4932 22278 4962 22330
rect 4962 22278 4974 22330
rect 4974 22278 4988 22330
rect 5012 22278 5026 22330
rect 5026 22278 5038 22330
rect 5038 22278 5068 22330
rect 5092 22278 5102 22330
rect 5102 22278 5148 22330
rect 4852 22276 4908 22278
rect 4932 22276 4988 22278
rect 5012 22276 5068 22278
rect 5092 22276 5148 22278
rect 3553 21786 3609 21788
rect 3633 21786 3689 21788
rect 3713 21786 3769 21788
rect 3793 21786 3849 21788
rect 3553 21734 3599 21786
rect 3599 21734 3609 21786
rect 3633 21734 3663 21786
rect 3663 21734 3675 21786
rect 3675 21734 3689 21786
rect 3713 21734 3727 21786
rect 3727 21734 3739 21786
rect 3739 21734 3769 21786
rect 3793 21734 3803 21786
rect 3803 21734 3849 21786
rect 3553 21732 3609 21734
rect 3633 21732 3689 21734
rect 3713 21732 3769 21734
rect 3793 21732 3849 21734
rect 5354 21392 5410 21448
rect 2254 21242 2310 21244
rect 2334 21242 2390 21244
rect 2414 21242 2470 21244
rect 2494 21242 2550 21244
rect 2254 21190 2300 21242
rect 2300 21190 2310 21242
rect 2334 21190 2364 21242
rect 2364 21190 2376 21242
rect 2376 21190 2390 21242
rect 2414 21190 2428 21242
rect 2428 21190 2440 21242
rect 2440 21190 2470 21242
rect 2494 21190 2504 21242
rect 2504 21190 2550 21242
rect 2254 21188 2310 21190
rect 2334 21188 2390 21190
rect 2414 21188 2470 21190
rect 2494 21188 2550 21190
rect 4852 21242 4908 21244
rect 4932 21242 4988 21244
rect 5012 21242 5068 21244
rect 5092 21242 5148 21244
rect 4852 21190 4898 21242
rect 4898 21190 4908 21242
rect 4932 21190 4962 21242
rect 4962 21190 4974 21242
rect 4974 21190 4988 21242
rect 5012 21190 5026 21242
rect 5026 21190 5038 21242
rect 5038 21190 5068 21242
rect 5092 21190 5102 21242
rect 5102 21190 5148 21242
rect 4852 21188 4908 21190
rect 4932 21188 4988 21190
rect 5012 21188 5068 21190
rect 5092 21188 5148 21190
rect 3553 20698 3609 20700
rect 3633 20698 3689 20700
rect 3713 20698 3769 20700
rect 3793 20698 3849 20700
rect 3553 20646 3599 20698
rect 3599 20646 3609 20698
rect 3633 20646 3663 20698
rect 3663 20646 3675 20698
rect 3675 20646 3689 20698
rect 3713 20646 3727 20698
rect 3727 20646 3739 20698
rect 3739 20646 3769 20698
rect 3793 20646 3803 20698
rect 3803 20646 3849 20698
rect 3553 20644 3609 20646
rect 3633 20644 3689 20646
rect 3713 20644 3769 20646
rect 3793 20644 3849 20646
rect 2254 20154 2310 20156
rect 2334 20154 2390 20156
rect 2414 20154 2470 20156
rect 2494 20154 2550 20156
rect 2254 20102 2300 20154
rect 2300 20102 2310 20154
rect 2334 20102 2364 20154
rect 2364 20102 2376 20154
rect 2376 20102 2390 20154
rect 2414 20102 2428 20154
rect 2428 20102 2440 20154
rect 2440 20102 2470 20154
rect 2494 20102 2504 20154
rect 2504 20102 2550 20154
rect 2254 20100 2310 20102
rect 2334 20100 2390 20102
rect 2414 20100 2470 20102
rect 2494 20100 2550 20102
rect 4852 20154 4908 20156
rect 4932 20154 4988 20156
rect 5012 20154 5068 20156
rect 5092 20154 5148 20156
rect 4852 20102 4898 20154
rect 4898 20102 4908 20154
rect 4932 20102 4962 20154
rect 4962 20102 4974 20154
rect 4974 20102 4988 20154
rect 5012 20102 5026 20154
rect 5026 20102 5038 20154
rect 5038 20102 5068 20154
rect 5092 20102 5102 20154
rect 5102 20102 5148 20154
rect 4852 20100 4908 20102
rect 4932 20100 4988 20102
rect 5012 20100 5068 20102
rect 5092 20100 5148 20102
rect 3553 19610 3609 19612
rect 3633 19610 3689 19612
rect 3713 19610 3769 19612
rect 3793 19610 3849 19612
rect 3553 19558 3599 19610
rect 3599 19558 3609 19610
rect 3633 19558 3663 19610
rect 3663 19558 3675 19610
rect 3675 19558 3689 19610
rect 3713 19558 3727 19610
rect 3727 19558 3739 19610
rect 3739 19558 3769 19610
rect 3793 19558 3803 19610
rect 3803 19558 3849 19610
rect 3553 19556 3609 19558
rect 3633 19556 3689 19558
rect 3713 19556 3769 19558
rect 3793 19556 3849 19558
rect 2254 19066 2310 19068
rect 2334 19066 2390 19068
rect 2414 19066 2470 19068
rect 2494 19066 2550 19068
rect 2254 19014 2300 19066
rect 2300 19014 2310 19066
rect 2334 19014 2364 19066
rect 2364 19014 2376 19066
rect 2376 19014 2390 19066
rect 2414 19014 2428 19066
rect 2428 19014 2440 19066
rect 2440 19014 2470 19066
rect 2494 19014 2504 19066
rect 2504 19014 2550 19066
rect 2254 19012 2310 19014
rect 2334 19012 2390 19014
rect 2414 19012 2470 19014
rect 2494 19012 2550 19014
rect 4852 19066 4908 19068
rect 4932 19066 4988 19068
rect 5012 19066 5068 19068
rect 5092 19066 5148 19068
rect 4852 19014 4898 19066
rect 4898 19014 4908 19066
rect 4932 19014 4962 19066
rect 4962 19014 4974 19066
rect 4974 19014 4988 19066
rect 5012 19014 5026 19066
rect 5026 19014 5038 19066
rect 5038 19014 5068 19066
rect 5092 19014 5102 19066
rect 5102 19014 5148 19066
rect 4852 19012 4908 19014
rect 4932 19012 4988 19014
rect 5012 19012 5068 19014
rect 5092 19012 5148 19014
rect 3553 18522 3609 18524
rect 3633 18522 3689 18524
rect 3713 18522 3769 18524
rect 3793 18522 3849 18524
rect 3553 18470 3599 18522
rect 3599 18470 3609 18522
rect 3633 18470 3663 18522
rect 3663 18470 3675 18522
rect 3675 18470 3689 18522
rect 3713 18470 3727 18522
rect 3727 18470 3739 18522
rect 3739 18470 3769 18522
rect 3793 18470 3803 18522
rect 3803 18470 3849 18522
rect 3553 18468 3609 18470
rect 3633 18468 3689 18470
rect 3713 18468 3769 18470
rect 3793 18468 3849 18470
rect 2254 17978 2310 17980
rect 2334 17978 2390 17980
rect 2414 17978 2470 17980
rect 2494 17978 2550 17980
rect 2254 17926 2300 17978
rect 2300 17926 2310 17978
rect 2334 17926 2364 17978
rect 2364 17926 2376 17978
rect 2376 17926 2390 17978
rect 2414 17926 2428 17978
rect 2428 17926 2440 17978
rect 2440 17926 2470 17978
rect 2494 17926 2504 17978
rect 2504 17926 2550 17978
rect 2254 17924 2310 17926
rect 2334 17924 2390 17926
rect 2414 17924 2470 17926
rect 2494 17924 2550 17926
rect 4852 17978 4908 17980
rect 4932 17978 4988 17980
rect 5012 17978 5068 17980
rect 5092 17978 5148 17980
rect 4852 17926 4898 17978
rect 4898 17926 4908 17978
rect 4932 17926 4962 17978
rect 4962 17926 4974 17978
rect 4974 17926 4988 17978
rect 5012 17926 5026 17978
rect 5026 17926 5038 17978
rect 5038 17926 5068 17978
rect 5092 17926 5102 17978
rect 5102 17926 5148 17978
rect 4852 17924 4908 17926
rect 4932 17924 4988 17926
rect 5012 17924 5068 17926
rect 5092 17924 5148 17926
rect 3553 17434 3609 17436
rect 3633 17434 3689 17436
rect 3713 17434 3769 17436
rect 3793 17434 3849 17436
rect 3553 17382 3599 17434
rect 3599 17382 3609 17434
rect 3633 17382 3663 17434
rect 3663 17382 3675 17434
rect 3675 17382 3689 17434
rect 3713 17382 3727 17434
rect 3727 17382 3739 17434
rect 3739 17382 3769 17434
rect 3793 17382 3803 17434
rect 3803 17382 3849 17434
rect 3553 17380 3609 17382
rect 3633 17380 3689 17382
rect 3713 17380 3769 17382
rect 3793 17380 3849 17382
rect 2254 16890 2310 16892
rect 2334 16890 2390 16892
rect 2414 16890 2470 16892
rect 2494 16890 2550 16892
rect 2254 16838 2300 16890
rect 2300 16838 2310 16890
rect 2334 16838 2364 16890
rect 2364 16838 2376 16890
rect 2376 16838 2390 16890
rect 2414 16838 2428 16890
rect 2428 16838 2440 16890
rect 2440 16838 2470 16890
rect 2494 16838 2504 16890
rect 2504 16838 2550 16890
rect 2254 16836 2310 16838
rect 2334 16836 2390 16838
rect 2414 16836 2470 16838
rect 2494 16836 2550 16838
rect 4852 16890 4908 16892
rect 4932 16890 4988 16892
rect 5012 16890 5068 16892
rect 5092 16890 5148 16892
rect 4852 16838 4898 16890
rect 4898 16838 4908 16890
rect 4932 16838 4962 16890
rect 4962 16838 4974 16890
rect 4974 16838 4988 16890
rect 5012 16838 5026 16890
rect 5026 16838 5038 16890
rect 5038 16838 5068 16890
rect 5092 16838 5102 16890
rect 5102 16838 5148 16890
rect 4852 16836 4908 16838
rect 4932 16836 4988 16838
rect 5012 16836 5068 16838
rect 5092 16836 5148 16838
rect 3553 16346 3609 16348
rect 3633 16346 3689 16348
rect 3713 16346 3769 16348
rect 3793 16346 3849 16348
rect 3553 16294 3599 16346
rect 3599 16294 3609 16346
rect 3633 16294 3663 16346
rect 3663 16294 3675 16346
rect 3675 16294 3689 16346
rect 3713 16294 3727 16346
rect 3727 16294 3739 16346
rect 3739 16294 3769 16346
rect 3793 16294 3803 16346
rect 3803 16294 3849 16346
rect 3553 16292 3609 16294
rect 3633 16292 3689 16294
rect 3713 16292 3769 16294
rect 3793 16292 3849 16294
rect 2254 15802 2310 15804
rect 2334 15802 2390 15804
rect 2414 15802 2470 15804
rect 2494 15802 2550 15804
rect 2254 15750 2300 15802
rect 2300 15750 2310 15802
rect 2334 15750 2364 15802
rect 2364 15750 2376 15802
rect 2376 15750 2390 15802
rect 2414 15750 2428 15802
rect 2428 15750 2440 15802
rect 2440 15750 2470 15802
rect 2494 15750 2504 15802
rect 2504 15750 2550 15802
rect 2254 15748 2310 15750
rect 2334 15748 2390 15750
rect 2414 15748 2470 15750
rect 2494 15748 2550 15750
rect 4852 15802 4908 15804
rect 4932 15802 4988 15804
rect 5012 15802 5068 15804
rect 5092 15802 5148 15804
rect 4852 15750 4898 15802
rect 4898 15750 4908 15802
rect 4932 15750 4962 15802
rect 4962 15750 4974 15802
rect 4974 15750 4988 15802
rect 5012 15750 5026 15802
rect 5026 15750 5038 15802
rect 5038 15750 5068 15802
rect 5092 15750 5102 15802
rect 5102 15750 5148 15802
rect 4852 15748 4908 15750
rect 4932 15748 4988 15750
rect 5012 15748 5068 15750
rect 5092 15748 5148 15750
rect 3553 15258 3609 15260
rect 3633 15258 3689 15260
rect 3713 15258 3769 15260
rect 3793 15258 3849 15260
rect 3553 15206 3599 15258
rect 3599 15206 3609 15258
rect 3633 15206 3663 15258
rect 3663 15206 3675 15258
rect 3675 15206 3689 15258
rect 3713 15206 3727 15258
rect 3727 15206 3739 15258
rect 3739 15206 3769 15258
rect 3793 15206 3803 15258
rect 3803 15206 3849 15258
rect 3553 15204 3609 15206
rect 3633 15204 3689 15206
rect 3713 15204 3769 15206
rect 3793 15204 3849 15206
rect 2254 14714 2310 14716
rect 2334 14714 2390 14716
rect 2414 14714 2470 14716
rect 2494 14714 2550 14716
rect 2254 14662 2300 14714
rect 2300 14662 2310 14714
rect 2334 14662 2364 14714
rect 2364 14662 2376 14714
rect 2376 14662 2390 14714
rect 2414 14662 2428 14714
rect 2428 14662 2440 14714
rect 2440 14662 2470 14714
rect 2494 14662 2504 14714
rect 2504 14662 2550 14714
rect 2254 14660 2310 14662
rect 2334 14660 2390 14662
rect 2414 14660 2470 14662
rect 2494 14660 2550 14662
rect 4852 14714 4908 14716
rect 4932 14714 4988 14716
rect 5012 14714 5068 14716
rect 5092 14714 5148 14716
rect 4852 14662 4898 14714
rect 4898 14662 4908 14714
rect 4932 14662 4962 14714
rect 4962 14662 4974 14714
rect 4974 14662 4988 14714
rect 5012 14662 5026 14714
rect 5026 14662 5038 14714
rect 5038 14662 5068 14714
rect 5092 14662 5102 14714
rect 5102 14662 5148 14714
rect 4852 14660 4908 14662
rect 4932 14660 4988 14662
rect 5012 14660 5068 14662
rect 5092 14660 5148 14662
rect 3553 14170 3609 14172
rect 3633 14170 3689 14172
rect 3713 14170 3769 14172
rect 3793 14170 3849 14172
rect 3553 14118 3599 14170
rect 3599 14118 3609 14170
rect 3633 14118 3663 14170
rect 3663 14118 3675 14170
rect 3675 14118 3689 14170
rect 3713 14118 3727 14170
rect 3727 14118 3739 14170
rect 3739 14118 3769 14170
rect 3793 14118 3803 14170
rect 3803 14118 3849 14170
rect 3553 14116 3609 14118
rect 3633 14116 3689 14118
rect 3713 14116 3769 14118
rect 3793 14116 3849 14118
rect 2254 13626 2310 13628
rect 2334 13626 2390 13628
rect 2414 13626 2470 13628
rect 2494 13626 2550 13628
rect 2254 13574 2300 13626
rect 2300 13574 2310 13626
rect 2334 13574 2364 13626
rect 2364 13574 2376 13626
rect 2376 13574 2390 13626
rect 2414 13574 2428 13626
rect 2428 13574 2440 13626
rect 2440 13574 2470 13626
rect 2494 13574 2504 13626
rect 2504 13574 2550 13626
rect 2254 13572 2310 13574
rect 2334 13572 2390 13574
rect 2414 13572 2470 13574
rect 2494 13572 2550 13574
rect 4852 13626 4908 13628
rect 4932 13626 4988 13628
rect 5012 13626 5068 13628
rect 5092 13626 5148 13628
rect 4852 13574 4898 13626
rect 4898 13574 4908 13626
rect 4932 13574 4962 13626
rect 4962 13574 4974 13626
rect 4974 13574 4988 13626
rect 5012 13574 5026 13626
rect 5026 13574 5038 13626
rect 5038 13574 5068 13626
rect 5092 13574 5102 13626
rect 5102 13574 5148 13626
rect 4852 13572 4908 13574
rect 4932 13572 4988 13574
rect 5012 13572 5068 13574
rect 5092 13572 5148 13574
rect 3553 13082 3609 13084
rect 3633 13082 3689 13084
rect 3713 13082 3769 13084
rect 3793 13082 3849 13084
rect 3553 13030 3599 13082
rect 3599 13030 3609 13082
rect 3633 13030 3663 13082
rect 3663 13030 3675 13082
rect 3675 13030 3689 13082
rect 3713 13030 3727 13082
rect 3727 13030 3739 13082
rect 3739 13030 3769 13082
rect 3793 13030 3803 13082
rect 3803 13030 3849 13082
rect 3553 13028 3609 13030
rect 3633 13028 3689 13030
rect 3713 13028 3769 13030
rect 3793 13028 3849 13030
rect 2254 12538 2310 12540
rect 2334 12538 2390 12540
rect 2414 12538 2470 12540
rect 2494 12538 2550 12540
rect 2254 12486 2300 12538
rect 2300 12486 2310 12538
rect 2334 12486 2364 12538
rect 2364 12486 2376 12538
rect 2376 12486 2390 12538
rect 2414 12486 2428 12538
rect 2428 12486 2440 12538
rect 2440 12486 2470 12538
rect 2494 12486 2504 12538
rect 2504 12486 2550 12538
rect 2254 12484 2310 12486
rect 2334 12484 2390 12486
rect 2414 12484 2470 12486
rect 2494 12484 2550 12486
rect 4852 12538 4908 12540
rect 4932 12538 4988 12540
rect 5012 12538 5068 12540
rect 5092 12538 5148 12540
rect 4852 12486 4898 12538
rect 4898 12486 4908 12538
rect 4932 12486 4962 12538
rect 4962 12486 4974 12538
rect 4974 12486 4988 12538
rect 5012 12486 5026 12538
rect 5026 12486 5038 12538
rect 5038 12486 5068 12538
rect 5092 12486 5102 12538
rect 5102 12486 5148 12538
rect 4852 12484 4908 12486
rect 4932 12484 4988 12486
rect 5012 12484 5068 12486
rect 5092 12484 5148 12486
rect 7449 27770 7505 27772
rect 7529 27770 7585 27772
rect 7609 27770 7665 27772
rect 7689 27770 7745 27772
rect 7449 27718 7495 27770
rect 7495 27718 7505 27770
rect 7529 27718 7559 27770
rect 7559 27718 7571 27770
rect 7571 27718 7585 27770
rect 7609 27718 7623 27770
rect 7623 27718 7635 27770
rect 7635 27718 7665 27770
rect 7689 27718 7699 27770
rect 7699 27718 7745 27770
rect 7449 27716 7505 27718
rect 7529 27716 7585 27718
rect 7609 27716 7665 27718
rect 7689 27716 7745 27718
rect 6150 27226 6206 27228
rect 6230 27226 6286 27228
rect 6310 27226 6366 27228
rect 6390 27226 6446 27228
rect 6150 27174 6196 27226
rect 6196 27174 6206 27226
rect 6230 27174 6260 27226
rect 6260 27174 6272 27226
rect 6272 27174 6286 27226
rect 6310 27174 6324 27226
rect 6324 27174 6336 27226
rect 6336 27174 6366 27226
rect 6390 27174 6400 27226
rect 6400 27174 6446 27226
rect 6150 27172 6206 27174
rect 6230 27172 6286 27174
rect 6310 27172 6366 27174
rect 6390 27172 6446 27174
rect 6734 27104 6790 27160
rect 5814 22480 5870 22536
rect 5538 19896 5594 19952
rect 3553 11994 3609 11996
rect 3633 11994 3689 11996
rect 3713 11994 3769 11996
rect 3793 11994 3849 11996
rect 3553 11942 3599 11994
rect 3599 11942 3609 11994
rect 3633 11942 3663 11994
rect 3663 11942 3675 11994
rect 3675 11942 3689 11994
rect 3713 11942 3727 11994
rect 3727 11942 3739 11994
rect 3739 11942 3769 11994
rect 3793 11942 3803 11994
rect 3803 11942 3849 11994
rect 3553 11940 3609 11942
rect 3633 11940 3689 11942
rect 3713 11940 3769 11942
rect 3793 11940 3849 11942
rect 2254 11450 2310 11452
rect 2334 11450 2390 11452
rect 2414 11450 2470 11452
rect 2494 11450 2550 11452
rect 2254 11398 2300 11450
rect 2300 11398 2310 11450
rect 2334 11398 2364 11450
rect 2364 11398 2376 11450
rect 2376 11398 2390 11450
rect 2414 11398 2428 11450
rect 2428 11398 2440 11450
rect 2440 11398 2470 11450
rect 2494 11398 2504 11450
rect 2504 11398 2550 11450
rect 2254 11396 2310 11398
rect 2334 11396 2390 11398
rect 2414 11396 2470 11398
rect 2494 11396 2550 11398
rect 4852 11450 4908 11452
rect 4932 11450 4988 11452
rect 5012 11450 5068 11452
rect 5092 11450 5148 11452
rect 4852 11398 4898 11450
rect 4898 11398 4908 11450
rect 4932 11398 4962 11450
rect 4962 11398 4974 11450
rect 4974 11398 4988 11450
rect 5012 11398 5026 11450
rect 5026 11398 5038 11450
rect 5038 11398 5068 11450
rect 5092 11398 5102 11450
rect 5102 11398 5148 11450
rect 4852 11396 4908 11398
rect 4932 11396 4988 11398
rect 5012 11396 5068 11398
rect 5092 11396 5148 11398
rect 3553 10906 3609 10908
rect 3633 10906 3689 10908
rect 3713 10906 3769 10908
rect 3793 10906 3849 10908
rect 3553 10854 3599 10906
rect 3599 10854 3609 10906
rect 3633 10854 3663 10906
rect 3663 10854 3675 10906
rect 3675 10854 3689 10906
rect 3713 10854 3727 10906
rect 3727 10854 3739 10906
rect 3739 10854 3769 10906
rect 3793 10854 3803 10906
rect 3803 10854 3849 10906
rect 3553 10852 3609 10854
rect 3633 10852 3689 10854
rect 3713 10852 3769 10854
rect 3793 10852 3849 10854
rect 2254 10362 2310 10364
rect 2334 10362 2390 10364
rect 2414 10362 2470 10364
rect 2494 10362 2550 10364
rect 2254 10310 2300 10362
rect 2300 10310 2310 10362
rect 2334 10310 2364 10362
rect 2364 10310 2376 10362
rect 2376 10310 2390 10362
rect 2414 10310 2428 10362
rect 2428 10310 2440 10362
rect 2440 10310 2470 10362
rect 2494 10310 2504 10362
rect 2504 10310 2550 10362
rect 2254 10308 2310 10310
rect 2334 10308 2390 10310
rect 2414 10308 2470 10310
rect 2494 10308 2550 10310
rect 4852 10362 4908 10364
rect 4932 10362 4988 10364
rect 5012 10362 5068 10364
rect 5092 10362 5148 10364
rect 4852 10310 4898 10362
rect 4898 10310 4908 10362
rect 4932 10310 4962 10362
rect 4962 10310 4974 10362
rect 4974 10310 4988 10362
rect 5012 10310 5026 10362
rect 5026 10310 5038 10362
rect 5038 10310 5068 10362
rect 5092 10310 5102 10362
rect 5102 10310 5148 10362
rect 4852 10308 4908 10310
rect 4932 10308 4988 10310
rect 5012 10308 5068 10310
rect 5092 10308 5148 10310
rect 3553 9818 3609 9820
rect 3633 9818 3689 9820
rect 3713 9818 3769 9820
rect 3793 9818 3849 9820
rect 3553 9766 3599 9818
rect 3599 9766 3609 9818
rect 3633 9766 3663 9818
rect 3663 9766 3675 9818
rect 3675 9766 3689 9818
rect 3713 9766 3727 9818
rect 3727 9766 3739 9818
rect 3739 9766 3769 9818
rect 3793 9766 3803 9818
rect 3803 9766 3849 9818
rect 3553 9764 3609 9766
rect 3633 9764 3689 9766
rect 3713 9764 3769 9766
rect 3793 9764 3849 9766
rect 2254 9274 2310 9276
rect 2334 9274 2390 9276
rect 2414 9274 2470 9276
rect 2494 9274 2550 9276
rect 2254 9222 2300 9274
rect 2300 9222 2310 9274
rect 2334 9222 2364 9274
rect 2364 9222 2376 9274
rect 2376 9222 2390 9274
rect 2414 9222 2428 9274
rect 2428 9222 2440 9274
rect 2440 9222 2470 9274
rect 2494 9222 2504 9274
rect 2504 9222 2550 9274
rect 2254 9220 2310 9222
rect 2334 9220 2390 9222
rect 2414 9220 2470 9222
rect 2494 9220 2550 9222
rect 4852 9274 4908 9276
rect 4932 9274 4988 9276
rect 5012 9274 5068 9276
rect 5092 9274 5148 9276
rect 4852 9222 4898 9274
rect 4898 9222 4908 9274
rect 4932 9222 4962 9274
rect 4962 9222 4974 9274
rect 4974 9222 4988 9274
rect 5012 9222 5026 9274
rect 5026 9222 5038 9274
rect 5038 9222 5068 9274
rect 5092 9222 5102 9274
rect 5102 9222 5148 9274
rect 4852 9220 4908 9222
rect 4932 9220 4988 9222
rect 5012 9220 5068 9222
rect 5092 9220 5148 9222
rect 3553 8730 3609 8732
rect 3633 8730 3689 8732
rect 3713 8730 3769 8732
rect 3793 8730 3849 8732
rect 3553 8678 3599 8730
rect 3599 8678 3609 8730
rect 3633 8678 3663 8730
rect 3663 8678 3675 8730
rect 3675 8678 3689 8730
rect 3713 8678 3727 8730
rect 3727 8678 3739 8730
rect 3739 8678 3769 8730
rect 3793 8678 3803 8730
rect 3803 8678 3849 8730
rect 3553 8676 3609 8678
rect 3633 8676 3689 8678
rect 3713 8676 3769 8678
rect 3793 8676 3849 8678
rect 6150 26138 6206 26140
rect 6230 26138 6286 26140
rect 6310 26138 6366 26140
rect 6390 26138 6446 26140
rect 6150 26086 6196 26138
rect 6196 26086 6206 26138
rect 6230 26086 6260 26138
rect 6260 26086 6272 26138
rect 6272 26086 6286 26138
rect 6310 26086 6324 26138
rect 6324 26086 6336 26138
rect 6336 26086 6366 26138
rect 6390 26086 6400 26138
rect 6400 26086 6446 26138
rect 6150 26084 6206 26086
rect 6230 26084 6286 26086
rect 6310 26084 6366 26086
rect 6390 26084 6446 26086
rect 6150 25050 6206 25052
rect 6230 25050 6286 25052
rect 6310 25050 6366 25052
rect 6390 25050 6446 25052
rect 6150 24998 6196 25050
rect 6196 24998 6206 25050
rect 6230 24998 6260 25050
rect 6260 24998 6272 25050
rect 6272 24998 6286 25050
rect 6310 24998 6324 25050
rect 6324 24998 6336 25050
rect 6336 24998 6366 25050
rect 6390 24998 6400 25050
rect 6400 24998 6446 25050
rect 6150 24996 6206 24998
rect 6230 24996 6286 24998
rect 6310 24996 6366 24998
rect 6390 24996 6446 24998
rect 6150 23962 6206 23964
rect 6230 23962 6286 23964
rect 6310 23962 6366 23964
rect 6390 23962 6446 23964
rect 6150 23910 6196 23962
rect 6196 23910 6206 23962
rect 6230 23910 6260 23962
rect 6260 23910 6272 23962
rect 6272 23910 6286 23962
rect 6310 23910 6324 23962
rect 6324 23910 6336 23962
rect 6336 23910 6366 23962
rect 6390 23910 6400 23962
rect 6400 23910 6446 23962
rect 6150 23908 6206 23910
rect 6230 23908 6286 23910
rect 6310 23908 6366 23910
rect 6390 23908 6446 23910
rect 6150 22874 6206 22876
rect 6230 22874 6286 22876
rect 6310 22874 6366 22876
rect 6390 22874 6446 22876
rect 6150 22822 6196 22874
rect 6196 22822 6206 22874
rect 6230 22822 6260 22874
rect 6260 22822 6272 22874
rect 6272 22822 6286 22874
rect 6310 22822 6324 22874
rect 6324 22822 6336 22874
rect 6336 22822 6366 22874
rect 6390 22822 6400 22874
rect 6400 22822 6446 22874
rect 6150 22820 6206 22822
rect 6230 22820 6286 22822
rect 6310 22820 6366 22822
rect 6390 22820 6446 22822
rect 6150 21786 6206 21788
rect 6230 21786 6286 21788
rect 6310 21786 6366 21788
rect 6390 21786 6446 21788
rect 6150 21734 6196 21786
rect 6196 21734 6206 21786
rect 6230 21734 6260 21786
rect 6260 21734 6272 21786
rect 6272 21734 6286 21786
rect 6310 21734 6324 21786
rect 6324 21734 6336 21786
rect 6336 21734 6366 21786
rect 6390 21734 6400 21786
rect 6400 21734 6446 21786
rect 6150 21732 6206 21734
rect 6230 21732 6286 21734
rect 6310 21732 6366 21734
rect 6390 21732 6446 21734
rect 7449 26682 7505 26684
rect 7529 26682 7585 26684
rect 7609 26682 7665 26684
rect 7689 26682 7745 26684
rect 7449 26630 7495 26682
rect 7495 26630 7505 26682
rect 7529 26630 7559 26682
rect 7559 26630 7571 26682
rect 7571 26630 7585 26682
rect 7609 26630 7623 26682
rect 7623 26630 7635 26682
rect 7635 26630 7665 26682
rect 7689 26630 7699 26682
rect 7699 26630 7745 26682
rect 7449 26628 7505 26630
rect 7529 26628 7585 26630
rect 7609 26628 7665 26630
rect 7689 26628 7745 26630
rect 7838 26016 7894 26072
rect 7449 25594 7505 25596
rect 7529 25594 7585 25596
rect 7609 25594 7665 25596
rect 7689 25594 7745 25596
rect 7449 25542 7495 25594
rect 7495 25542 7505 25594
rect 7529 25542 7559 25594
rect 7559 25542 7571 25594
rect 7571 25542 7585 25594
rect 7609 25542 7623 25594
rect 7623 25542 7635 25594
rect 7635 25542 7665 25594
rect 7689 25542 7699 25594
rect 7699 25542 7745 25594
rect 7449 25540 7505 25542
rect 7529 25540 7585 25542
rect 7609 25540 7665 25542
rect 7689 25540 7745 25542
rect 7449 24506 7505 24508
rect 7529 24506 7585 24508
rect 7609 24506 7665 24508
rect 7689 24506 7745 24508
rect 7449 24454 7495 24506
rect 7495 24454 7505 24506
rect 7529 24454 7559 24506
rect 7559 24454 7571 24506
rect 7571 24454 7585 24506
rect 7609 24454 7623 24506
rect 7623 24454 7635 24506
rect 7635 24454 7665 24506
rect 7689 24454 7699 24506
rect 7699 24454 7745 24506
rect 7449 24452 7505 24454
rect 7529 24452 7585 24454
rect 7609 24452 7665 24454
rect 7689 24452 7745 24454
rect 7449 23418 7505 23420
rect 7529 23418 7585 23420
rect 7609 23418 7665 23420
rect 7689 23418 7745 23420
rect 7449 23366 7495 23418
rect 7495 23366 7505 23418
rect 7529 23366 7559 23418
rect 7559 23366 7571 23418
rect 7571 23366 7585 23418
rect 7609 23366 7623 23418
rect 7623 23366 7635 23418
rect 7635 23366 7665 23418
rect 7689 23366 7699 23418
rect 7699 23366 7745 23418
rect 7449 23364 7505 23366
rect 7529 23364 7585 23366
rect 7609 23364 7665 23366
rect 7689 23364 7745 23366
rect 8114 24792 8170 24848
rect 6150 20698 6206 20700
rect 6230 20698 6286 20700
rect 6310 20698 6366 20700
rect 6390 20698 6446 20700
rect 6150 20646 6196 20698
rect 6196 20646 6206 20698
rect 6230 20646 6260 20698
rect 6260 20646 6272 20698
rect 6272 20646 6286 20698
rect 6310 20646 6324 20698
rect 6324 20646 6336 20698
rect 6336 20646 6366 20698
rect 6390 20646 6400 20698
rect 6400 20646 6446 20698
rect 6150 20644 6206 20646
rect 6230 20644 6286 20646
rect 6310 20644 6366 20646
rect 6390 20644 6446 20646
rect 6150 19610 6206 19612
rect 6230 19610 6286 19612
rect 6310 19610 6366 19612
rect 6390 19610 6446 19612
rect 6150 19558 6196 19610
rect 6196 19558 6206 19610
rect 6230 19558 6260 19610
rect 6260 19558 6272 19610
rect 6272 19558 6286 19610
rect 6310 19558 6324 19610
rect 6324 19558 6336 19610
rect 6336 19558 6366 19610
rect 6390 19558 6400 19610
rect 6400 19558 6446 19610
rect 6150 19556 6206 19558
rect 6230 19556 6286 19558
rect 6310 19556 6366 19558
rect 6390 19556 6446 19558
rect 6150 18522 6206 18524
rect 6230 18522 6286 18524
rect 6310 18522 6366 18524
rect 6390 18522 6446 18524
rect 6150 18470 6196 18522
rect 6196 18470 6206 18522
rect 6230 18470 6260 18522
rect 6260 18470 6272 18522
rect 6272 18470 6286 18522
rect 6310 18470 6324 18522
rect 6324 18470 6336 18522
rect 6336 18470 6366 18522
rect 6390 18470 6400 18522
rect 6400 18470 6446 18522
rect 6150 18468 6206 18470
rect 6230 18468 6286 18470
rect 6310 18468 6366 18470
rect 6390 18468 6446 18470
rect 5998 17856 6054 17912
rect 5998 17720 6054 17776
rect 6150 17434 6206 17436
rect 6230 17434 6286 17436
rect 6310 17434 6366 17436
rect 6390 17434 6446 17436
rect 6150 17382 6196 17434
rect 6196 17382 6206 17434
rect 6230 17382 6260 17434
rect 6260 17382 6272 17434
rect 6272 17382 6286 17434
rect 6310 17382 6324 17434
rect 6324 17382 6336 17434
rect 6336 17382 6366 17434
rect 6390 17382 6400 17434
rect 6400 17382 6446 17434
rect 6150 17380 6206 17382
rect 6230 17380 6286 17382
rect 6310 17380 6366 17382
rect 6390 17380 6446 17382
rect 7449 22330 7505 22332
rect 7529 22330 7585 22332
rect 7609 22330 7665 22332
rect 7689 22330 7745 22332
rect 7449 22278 7495 22330
rect 7495 22278 7505 22330
rect 7529 22278 7559 22330
rect 7559 22278 7571 22330
rect 7571 22278 7585 22330
rect 7609 22278 7623 22330
rect 7623 22278 7635 22330
rect 7635 22278 7665 22330
rect 7689 22278 7699 22330
rect 7699 22278 7745 22330
rect 7449 22276 7505 22278
rect 7529 22276 7585 22278
rect 7609 22276 7665 22278
rect 7689 22276 7745 22278
rect 8298 23704 8354 23760
rect 7449 21242 7505 21244
rect 7529 21242 7585 21244
rect 7609 21242 7665 21244
rect 7689 21242 7745 21244
rect 7449 21190 7495 21242
rect 7495 21190 7505 21242
rect 7529 21190 7559 21242
rect 7559 21190 7571 21242
rect 7571 21190 7585 21242
rect 7609 21190 7623 21242
rect 7623 21190 7635 21242
rect 7635 21190 7665 21242
rect 7689 21190 7699 21242
rect 7699 21190 7745 21242
rect 7449 21188 7505 21190
rect 7529 21188 7585 21190
rect 7609 21188 7665 21190
rect 7689 21188 7745 21190
rect 7449 20154 7505 20156
rect 7529 20154 7585 20156
rect 7609 20154 7665 20156
rect 7689 20154 7745 20156
rect 7449 20102 7495 20154
rect 7495 20102 7505 20154
rect 7529 20102 7559 20154
rect 7559 20102 7571 20154
rect 7571 20102 7585 20154
rect 7609 20102 7623 20154
rect 7623 20102 7635 20154
rect 7635 20102 7665 20154
rect 7689 20102 7699 20154
rect 7699 20102 7745 20154
rect 7449 20100 7505 20102
rect 7529 20100 7585 20102
rect 7609 20100 7665 20102
rect 7689 20100 7745 20102
rect 6826 18808 6882 18864
rect 6150 16346 6206 16348
rect 6230 16346 6286 16348
rect 6310 16346 6366 16348
rect 6390 16346 6446 16348
rect 6150 16294 6196 16346
rect 6196 16294 6206 16346
rect 6230 16294 6260 16346
rect 6260 16294 6272 16346
rect 6272 16294 6286 16346
rect 6310 16294 6324 16346
rect 6324 16294 6336 16346
rect 6336 16294 6366 16346
rect 6390 16294 6400 16346
rect 6400 16294 6446 16346
rect 6150 16292 6206 16294
rect 6230 16292 6286 16294
rect 6310 16292 6366 16294
rect 6390 16292 6446 16294
rect 6150 15258 6206 15260
rect 6230 15258 6286 15260
rect 6310 15258 6366 15260
rect 6390 15258 6446 15260
rect 6150 15206 6196 15258
rect 6196 15206 6206 15258
rect 6230 15206 6260 15258
rect 6260 15206 6272 15258
rect 6272 15206 6286 15258
rect 6310 15206 6324 15258
rect 6324 15206 6336 15258
rect 6336 15206 6366 15258
rect 6390 15206 6400 15258
rect 6400 15206 6446 15258
rect 6150 15204 6206 15206
rect 6230 15204 6286 15206
rect 6310 15204 6366 15206
rect 6390 15204 6446 15206
rect 5722 13232 5778 13288
rect 5630 9968 5686 10024
rect 2254 8186 2310 8188
rect 2334 8186 2390 8188
rect 2414 8186 2470 8188
rect 2494 8186 2550 8188
rect 2254 8134 2300 8186
rect 2300 8134 2310 8186
rect 2334 8134 2364 8186
rect 2364 8134 2376 8186
rect 2376 8134 2390 8186
rect 2414 8134 2428 8186
rect 2428 8134 2440 8186
rect 2440 8134 2470 8186
rect 2494 8134 2504 8186
rect 2504 8134 2550 8186
rect 2254 8132 2310 8134
rect 2334 8132 2390 8134
rect 2414 8132 2470 8134
rect 2494 8132 2550 8134
rect 4852 8186 4908 8188
rect 4932 8186 4988 8188
rect 5012 8186 5068 8188
rect 5092 8186 5148 8188
rect 4852 8134 4898 8186
rect 4898 8134 4908 8186
rect 4932 8134 4962 8186
rect 4962 8134 4974 8186
rect 4974 8134 4988 8186
rect 5012 8134 5026 8186
rect 5026 8134 5038 8186
rect 5038 8134 5068 8186
rect 5092 8134 5102 8186
rect 5102 8134 5148 8186
rect 4852 8132 4908 8134
rect 4932 8132 4988 8134
rect 5012 8132 5068 8134
rect 5092 8132 5148 8134
rect 6150 14170 6206 14172
rect 6230 14170 6286 14172
rect 6310 14170 6366 14172
rect 6390 14170 6446 14172
rect 6150 14118 6196 14170
rect 6196 14118 6206 14170
rect 6230 14118 6260 14170
rect 6260 14118 6272 14170
rect 6272 14118 6286 14170
rect 6310 14118 6324 14170
rect 6324 14118 6336 14170
rect 6336 14118 6366 14170
rect 6390 14118 6400 14170
rect 6400 14118 6446 14170
rect 6150 14116 6206 14118
rect 6230 14116 6286 14118
rect 6310 14116 6366 14118
rect 6390 14116 6446 14118
rect 6150 13082 6206 13084
rect 6230 13082 6286 13084
rect 6310 13082 6366 13084
rect 6390 13082 6446 13084
rect 6150 13030 6196 13082
rect 6196 13030 6206 13082
rect 6230 13030 6260 13082
rect 6260 13030 6272 13082
rect 6272 13030 6286 13082
rect 6310 13030 6324 13082
rect 6324 13030 6336 13082
rect 6336 13030 6366 13082
rect 6390 13030 6400 13082
rect 6400 13030 6446 13082
rect 6150 13028 6206 13030
rect 6230 13028 6286 13030
rect 6310 13028 6366 13030
rect 6390 13028 6446 13030
rect 5998 12688 6054 12744
rect 5998 12280 6054 12336
rect 5722 8880 5778 8936
rect 6150 11994 6206 11996
rect 6230 11994 6286 11996
rect 6310 11994 6366 11996
rect 6390 11994 6446 11996
rect 6150 11942 6196 11994
rect 6196 11942 6206 11994
rect 6230 11942 6260 11994
rect 6260 11942 6272 11994
rect 6272 11942 6286 11994
rect 6310 11942 6324 11994
rect 6324 11942 6336 11994
rect 6336 11942 6366 11994
rect 6390 11942 6400 11994
rect 6400 11942 6446 11994
rect 6150 11940 6206 11942
rect 6230 11940 6286 11942
rect 6310 11940 6366 11942
rect 6390 11940 6446 11942
rect 3553 7642 3609 7644
rect 3633 7642 3689 7644
rect 3713 7642 3769 7644
rect 3793 7642 3849 7644
rect 3553 7590 3599 7642
rect 3599 7590 3609 7642
rect 3633 7590 3663 7642
rect 3663 7590 3675 7642
rect 3675 7590 3689 7642
rect 3713 7590 3727 7642
rect 3727 7590 3739 7642
rect 3739 7590 3769 7642
rect 3793 7590 3803 7642
rect 3803 7590 3849 7642
rect 3553 7588 3609 7590
rect 3633 7588 3689 7590
rect 3713 7588 3769 7590
rect 3793 7588 3849 7590
rect 2254 7098 2310 7100
rect 2334 7098 2390 7100
rect 2414 7098 2470 7100
rect 2494 7098 2550 7100
rect 2254 7046 2300 7098
rect 2300 7046 2310 7098
rect 2334 7046 2364 7098
rect 2364 7046 2376 7098
rect 2376 7046 2390 7098
rect 2414 7046 2428 7098
rect 2428 7046 2440 7098
rect 2440 7046 2470 7098
rect 2494 7046 2504 7098
rect 2504 7046 2550 7098
rect 2254 7044 2310 7046
rect 2334 7044 2390 7046
rect 2414 7044 2470 7046
rect 2494 7044 2550 7046
rect 4852 7098 4908 7100
rect 4932 7098 4988 7100
rect 5012 7098 5068 7100
rect 5092 7098 5148 7100
rect 4852 7046 4898 7098
rect 4898 7046 4908 7098
rect 4932 7046 4962 7098
rect 4962 7046 4974 7098
rect 4974 7046 4988 7098
rect 5012 7046 5026 7098
rect 5026 7046 5038 7098
rect 5038 7046 5068 7098
rect 5092 7046 5102 7098
rect 5102 7046 5148 7098
rect 4852 7044 4908 7046
rect 4932 7044 4988 7046
rect 5012 7044 5068 7046
rect 5092 7044 5148 7046
rect 3553 6554 3609 6556
rect 3633 6554 3689 6556
rect 3713 6554 3769 6556
rect 3793 6554 3849 6556
rect 3553 6502 3599 6554
rect 3599 6502 3609 6554
rect 3633 6502 3663 6554
rect 3663 6502 3675 6554
rect 3675 6502 3689 6554
rect 3713 6502 3727 6554
rect 3727 6502 3739 6554
rect 3739 6502 3769 6554
rect 3793 6502 3803 6554
rect 3803 6502 3849 6554
rect 3553 6500 3609 6502
rect 3633 6500 3689 6502
rect 3713 6500 3769 6502
rect 3793 6500 3849 6502
rect 2254 6010 2310 6012
rect 2334 6010 2390 6012
rect 2414 6010 2470 6012
rect 2494 6010 2550 6012
rect 2254 5958 2300 6010
rect 2300 5958 2310 6010
rect 2334 5958 2364 6010
rect 2364 5958 2376 6010
rect 2376 5958 2390 6010
rect 2414 5958 2428 6010
rect 2428 5958 2440 6010
rect 2440 5958 2470 6010
rect 2494 5958 2504 6010
rect 2504 5958 2550 6010
rect 2254 5956 2310 5958
rect 2334 5956 2390 5958
rect 2414 5956 2470 5958
rect 2494 5956 2550 5958
rect 3553 5466 3609 5468
rect 3633 5466 3689 5468
rect 3713 5466 3769 5468
rect 3793 5466 3849 5468
rect 3553 5414 3599 5466
rect 3599 5414 3609 5466
rect 3633 5414 3663 5466
rect 3663 5414 3675 5466
rect 3675 5414 3689 5466
rect 3713 5414 3727 5466
rect 3727 5414 3739 5466
rect 3739 5414 3769 5466
rect 3793 5414 3803 5466
rect 3803 5414 3849 5466
rect 3553 5412 3609 5414
rect 3633 5412 3689 5414
rect 3713 5412 3769 5414
rect 3793 5412 3849 5414
rect 2254 4922 2310 4924
rect 2334 4922 2390 4924
rect 2414 4922 2470 4924
rect 2494 4922 2550 4924
rect 2254 4870 2300 4922
rect 2300 4870 2310 4922
rect 2334 4870 2364 4922
rect 2364 4870 2376 4922
rect 2376 4870 2390 4922
rect 2414 4870 2428 4922
rect 2428 4870 2440 4922
rect 2440 4870 2470 4922
rect 2494 4870 2504 4922
rect 2504 4870 2550 4922
rect 2254 4868 2310 4870
rect 2334 4868 2390 4870
rect 2414 4868 2470 4870
rect 2494 4868 2550 4870
rect 2254 3834 2310 3836
rect 2334 3834 2390 3836
rect 2414 3834 2470 3836
rect 2494 3834 2550 3836
rect 2254 3782 2300 3834
rect 2300 3782 2310 3834
rect 2334 3782 2364 3834
rect 2364 3782 2376 3834
rect 2376 3782 2390 3834
rect 2414 3782 2428 3834
rect 2428 3782 2440 3834
rect 2440 3782 2470 3834
rect 2494 3782 2504 3834
rect 2504 3782 2550 3834
rect 2254 3780 2310 3782
rect 2334 3780 2390 3782
rect 2414 3780 2470 3782
rect 2494 3780 2550 3782
rect 3553 4378 3609 4380
rect 3633 4378 3689 4380
rect 3713 4378 3769 4380
rect 3793 4378 3849 4380
rect 3553 4326 3599 4378
rect 3599 4326 3609 4378
rect 3633 4326 3663 4378
rect 3663 4326 3675 4378
rect 3675 4326 3689 4378
rect 3713 4326 3727 4378
rect 3727 4326 3739 4378
rect 3739 4326 3769 4378
rect 3793 4326 3803 4378
rect 3803 4326 3849 4378
rect 3553 4324 3609 4326
rect 3633 4324 3689 4326
rect 3713 4324 3769 4326
rect 3793 4324 3849 4326
rect 2254 2746 2310 2748
rect 2334 2746 2390 2748
rect 2414 2746 2470 2748
rect 2494 2746 2550 2748
rect 2254 2694 2300 2746
rect 2300 2694 2310 2746
rect 2334 2694 2364 2746
rect 2364 2694 2376 2746
rect 2376 2694 2390 2746
rect 2414 2694 2428 2746
rect 2428 2694 2440 2746
rect 2440 2694 2470 2746
rect 2494 2694 2504 2746
rect 2504 2694 2550 2746
rect 2254 2692 2310 2694
rect 2334 2692 2390 2694
rect 2414 2692 2470 2694
rect 2494 2692 2550 2694
rect 3553 3290 3609 3292
rect 3633 3290 3689 3292
rect 3713 3290 3769 3292
rect 3793 3290 3849 3292
rect 3553 3238 3599 3290
rect 3599 3238 3609 3290
rect 3633 3238 3663 3290
rect 3663 3238 3675 3290
rect 3675 3238 3689 3290
rect 3713 3238 3727 3290
rect 3727 3238 3739 3290
rect 3739 3238 3769 3290
rect 3793 3238 3803 3290
rect 3803 3238 3849 3290
rect 3553 3236 3609 3238
rect 3633 3236 3689 3238
rect 3713 3236 3769 3238
rect 3793 3236 3849 3238
rect 4852 6010 4908 6012
rect 4932 6010 4988 6012
rect 5012 6010 5068 6012
rect 5092 6010 5148 6012
rect 4852 5958 4898 6010
rect 4898 5958 4908 6010
rect 4932 5958 4962 6010
rect 4962 5958 4974 6010
rect 4974 5958 4988 6010
rect 5012 5958 5026 6010
rect 5026 5958 5038 6010
rect 5038 5958 5068 6010
rect 5092 5958 5102 6010
rect 5102 5958 5148 6010
rect 4852 5956 4908 5958
rect 4932 5956 4988 5958
rect 5012 5956 5068 5958
rect 5092 5956 5148 5958
rect 6734 14476 6790 14512
rect 6734 14456 6736 14476
rect 6736 14456 6788 14476
rect 6788 14456 6790 14476
rect 7449 19066 7505 19068
rect 7529 19066 7585 19068
rect 7609 19066 7665 19068
rect 7689 19066 7745 19068
rect 7449 19014 7495 19066
rect 7495 19014 7505 19066
rect 7529 19014 7559 19066
rect 7559 19014 7571 19066
rect 7571 19014 7585 19066
rect 7609 19014 7623 19066
rect 7623 19014 7635 19066
rect 7635 19014 7665 19066
rect 7689 19014 7699 19066
rect 7699 19014 7745 19066
rect 7449 19012 7505 19014
rect 7529 19012 7585 19014
rect 7609 19012 7665 19014
rect 7689 19012 7745 19014
rect 7449 17978 7505 17980
rect 7529 17978 7585 17980
rect 7609 17978 7665 17980
rect 7689 17978 7745 17980
rect 7449 17926 7495 17978
rect 7495 17926 7505 17978
rect 7529 17926 7559 17978
rect 7559 17926 7571 17978
rect 7571 17926 7585 17978
rect 7609 17926 7623 17978
rect 7623 17926 7635 17978
rect 7635 17926 7665 17978
rect 7689 17926 7699 17978
rect 7699 17926 7745 17978
rect 7449 17924 7505 17926
rect 7529 17924 7585 17926
rect 7609 17924 7665 17926
rect 7689 17924 7745 17926
rect 7449 16890 7505 16892
rect 7529 16890 7585 16892
rect 7609 16890 7665 16892
rect 7689 16890 7745 16892
rect 7449 16838 7495 16890
rect 7495 16838 7505 16890
rect 7529 16838 7559 16890
rect 7559 16838 7571 16890
rect 7571 16838 7585 16890
rect 7609 16838 7623 16890
rect 7623 16838 7635 16890
rect 7635 16838 7665 16890
rect 7689 16838 7699 16890
rect 7699 16838 7745 16890
rect 7449 16836 7505 16838
rect 7529 16836 7585 16838
rect 7609 16836 7665 16838
rect 7689 16836 7745 16838
rect 8022 16768 8078 16824
rect 7449 15802 7505 15804
rect 7529 15802 7585 15804
rect 7609 15802 7665 15804
rect 7689 15802 7745 15804
rect 7449 15750 7495 15802
rect 7495 15750 7505 15802
rect 7529 15750 7559 15802
rect 7559 15750 7571 15802
rect 7571 15750 7585 15802
rect 7609 15750 7623 15802
rect 7623 15750 7635 15802
rect 7635 15750 7665 15802
rect 7689 15750 7699 15802
rect 7699 15750 7745 15802
rect 7449 15748 7505 15750
rect 7529 15748 7585 15750
rect 7609 15748 7665 15750
rect 7689 15748 7745 15750
rect 7930 15544 7986 15600
rect 7449 14714 7505 14716
rect 7529 14714 7585 14716
rect 7609 14714 7665 14716
rect 7689 14714 7745 14716
rect 7449 14662 7495 14714
rect 7495 14662 7505 14714
rect 7529 14662 7559 14714
rect 7559 14662 7571 14714
rect 7571 14662 7585 14714
rect 7609 14662 7623 14714
rect 7623 14662 7635 14714
rect 7635 14662 7665 14714
rect 7689 14662 7699 14714
rect 7699 14662 7745 14714
rect 7449 14660 7505 14662
rect 7529 14660 7585 14662
rect 7609 14660 7665 14662
rect 7689 14660 7745 14662
rect 7449 13626 7505 13628
rect 7529 13626 7585 13628
rect 7609 13626 7665 13628
rect 7689 13626 7745 13628
rect 7449 13574 7495 13626
rect 7495 13574 7505 13626
rect 7529 13574 7559 13626
rect 7559 13574 7571 13626
rect 7571 13574 7585 13626
rect 7609 13574 7623 13626
rect 7623 13574 7635 13626
rect 7635 13574 7665 13626
rect 7689 13574 7699 13626
rect 7699 13574 7745 13626
rect 7449 13572 7505 13574
rect 7529 13572 7585 13574
rect 7609 13572 7665 13574
rect 7689 13572 7745 13574
rect 6642 10920 6698 10976
rect 6150 10906 6206 10908
rect 6230 10906 6286 10908
rect 6310 10906 6366 10908
rect 6390 10906 6446 10908
rect 6150 10854 6196 10906
rect 6196 10854 6206 10906
rect 6230 10854 6260 10906
rect 6260 10854 6272 10906
rect 6272 10854 6286 10906
rect 6310 10854 6324 10906
rect 6324 10854 6336 10906
rect 6336 10854 6366 10906
rect 6390 10854 6400 10906
rect 6400 10854 6446 10906
rect 6150 10852 6206 10854
rect 6230 10852 6286 10854
rect 6310 10852 6366 10854
rect 6390 10852 6446 10854
rect 6150 9818 6206 9820
rect 6230 9818 6286 9820
rect 6310 9818 6366 9820
rect 6390 9818 6446 9820
rect 6150 9766 6196 9818
rect 6196 9766 6206 9818
rect 6230 9766 6260 9818
rect 6260 9766 6272 9818
rect 6272 9766 6286 9818
rect 6310 9766 6324 9818
rect 6324 9766 6336 9818
rect 6336 9766 6366 9818
rect 6390 9766 6400 9818
rect 6400 9766 6446 9818
rect 6150 9764 6206 9766
rect 6230 9764 6286 9766
rect 6310 9764 6366 9766
rect 6390 9764 6446 9766
rect 6150 8730 6206 8732
rect 6230 8730 6286 8732
rect 6310 8730 6366 8732
rect 6390 8730 6446 8732
rect 6150 8678 6196 8730
rect 6196 8678 6206 8730
rect 6230 8678 6260 8730
rect 6260 8678 6272 8730
rect 6272 8678 6286 8730
rect 6310 8678 6324 8730
rect 6324 8678 6336 8730
rect 6336 8678 6366 8730
rect 6390 8678 6400 8730
rect 6400 8678 6446 8730
rect 6150 8676 6206 8678
rect 6230 8676 6286 8678
rect 6310 8676 6366 8678
rect 6390 8676 6446 8678
rect 6150 7642 6206 7644
rect 6230 7642 6286 7644
rect 6310 7642 6366 7644
rect 6390 7642 6446 7644
rect 6150 7590 6196 7642
rect 6196 7590 6206 7642
rect 6230 7590 6260 7642
rect 6260 7590 6272 7642
rect 6272 7590 6286 7642
rect 6310 7590 6324 7642
rect 6324 7590 6336 7642
rect 6336 7590 6366 7642
rect 6390 7590 6400 7642
rect 6400 7590 6446 7642
rect 6150 7588 6206 7590
rect 6230 7588 6286 7590
rect 6310 7588 6366 7590
rect 6390 7588 6446 7590
rect 6734 7520 6790 7576
rect 6150 6554 6206 6556
rect 6230 6554 6286 6556
rect 6310 6554 6366 6556
rect 6390 6554 6446 6556
rect 6150 6502 6196 6554
rect 6196 6502 6206 6554
rect 6230 6502 6260 6554
rect 6260 6502 6272 6554
rect 6272 6502 6286 6554
rect 6310 6502 6324 6554
rect 6324 6502 6336 6554
rect 6336 6502 6366 6554
rect 6390 6502 6400 6554
rect 6400 6502 6446 6554
rect 6150 6500 6206 6502
rect 6230 6500 6286 6502
rect 6310 6500 6366 6502
rect 6390 6500 6446 6502
rect 5998 6296 6054 6352
rect 4852 4922 4908 4924
rect 4932 4922 4988 4924
rect 5012 4922 5068 4924
rect 5092 4922 5148 4924
rect 4852 4870 4898 4922
rect 4898 4870 4908 4922
rect 4932 4870 4962 4922
rect 4962 4870 4974 4922
rect 4974 4870 4988 4922
rect 5012 4870 5026 4922
rect 5026 4870 5038 4922
rect 5038 4870 5068 4922
rect 5092 4870 5102 4922
rect 5102 4870 5148 4922
rect 4852 4868 4908 4870
rect 4932 4868 4988 4870
rect 5012 4868 5068 4870
rect 5092 4868 5148 4870
rect 4852 3834 4908 3836
rect 4932 3834 4988 3836
rect 5012 3834 5068 3836
rect 5092 3834 5148 3836
rect 4852 3782 4898 3834
rect 4898 3782 4908 3834
rect 4932 3782 4962 3834
rect 4962 3782 4974 3834
rect 4974 3782 4988 3834
rect 5012 3782 5026 3834
rect 5026 3782 5038 3834
rect 5038 3782 5068 3834
rect 5092 3782 5102 3834
rect 5102 3782 5148 3834
rect 4852 3780 4908 3782
rect 4932 3780 4988 3782
rect 5012 3780 5068 3782
rect 5092 3780 5148 3782
rect 4852 2746 4908 2748
rect 4932 2746 4988 2748
rect 5012 2746 5068 2748
rect 5092 2746 5148 2748
rect 4852 2694 4898 2746
rect 4898 2694 4908 2746
rect 4932 2694 4962 2746
rect 4962 2694 4974 2746
rect 4974 2694 4988 2746
rect 5012 2694 5026 2746
rect 5026 2694 5038 2746
rect 5038 2694 5068 2746
rect 5092 2694 5102 2746
rect 5102 2694 5148 2746
rect 4852 2692 4908 2694
rect 4932 2692 4988 2694
rect 5012 2692 5068 2694
rect 5092 2692 5148 2694
rect 6150 5466 6206 5468
rect 6230 5466 6286 5468
rect 6310 5466 6366 5468
rect 6390 5466 6446 5468
rect 6150 5414 6196 5466
rect 6196 5414 6206 5466
rect 6230 5414 6260 5466
rect 6260 5414 6272 5466
rect 6272 5414 6286 5466
rect 6310 5414 6324 5466
rect 6324 5414 6336 5466
rect 6336 5414 6366 5466
rect 6390 5414 6400 5466
rect 6400 5414 6446 5466
rect 6150 5412 6206 5414
rect 6230 5412 6286 5414
rect 6310 5412 6366 5414
rect 6390 5412 6446 5414
rect 6150 4378 6206 4380
rect 6230 4378 6286 4380
rect 6310 4378 6366 4380
rect 6390 4378 6446 4380
rect 6150 4326 6196 4378
rect 6196 4326 6206 4378
rect 6230 4326 6260 4378
rect 6260 4326 6272 4378
rect 6272 4326 6286 4378
rect 6310 4326 6324 4378
rect 6324 4326 6336 4378
rect 6336 4326 6366 4378
rect 6390 4326 6400 4378
rect 6400 4326 6446 4378
rect 6150 4324 6206 4326
rect 6230 4324 6286 4326
rect 6310 4324 6366 4326
rect 6390 4324 6446 4326
rect 7449 12538 7505 12540
rect 7529 12538 7585 12540
rect 7609 12538 7665 12540
rect 7689 12538 7745 12540
rect 7449 12486 7495 12538
rect 7495 12486 7505 12538
rect 7529 12486 7559 12538
rect 7559 12486 7571 12538
rect 7571 12486 7585 12538
rect 7609 12486 7623 12538
rect 7623 12486 7635 12538
rect 7635 12486 7665 12538
rect 7689 12486 7699 12538
rect 7699 12486 7745 12538
rect 7449 12484 7505 12486
rect 7529 12484 7585 12486
rect 7609 12484 7665 12486
rect 7689 12484 7745 12486
rect 7449 11450 7505 11452
rect 7529 11450 7585 11452
rect 7609 11450 7665 11452
rect 7689 11450 7745 11452
rect 7449 11398 7495 11450
rect 7495 11398 7505 11450
rect 7529 11398 7559 11450
rect 7559 11398 7571 11450
rect 7571 11398 7585 11450
rect 7609 11398 7623 11450
rect 7623 11398 7635 11450
rect 7635 11398 7665 11450
rect 7689 11398 7699 11450
rect 7699 11398 7745 11450
rect 7449 11396 7505 11398
rect 7529 11396 7585 11398
rect 7609 11396 7665 11398
rect 7689 11396 7745 11398
rect 7449 10362 7505 10364
rect 7529 10362 7585 10364
rect 7609 10362 7665 10364
rect 7689 10362 7745 10364
rect 7449 10310 7495 10362
rect 7495 10310 7505 10362
rect 7529 10310 7559 10362
rect 7559 10310 7571 10362
rect 7571 10310 7585 10362
rect 7609 10310 7623 10362
rect 7623 10310 7635 10362
rect 7635 10310 7665 10362
rect 7689 10310 7699 10362
rect 7699 10310 7745 10362
rect 7449 10308 7505 10310
rect 7529 10308 7585 10310
rect 7609 10308 7665 10310
rect 7689 10308 7745 10310
rect 7449 9274 7505 9276
rect 7529 9274 7585 9276
rect 7609 9274 7665 9276
rect 7689 9274 7745 9276
rect 7449 9222 7495 9274
rect 7495 9222 7505 9274
rect 7529 9222 7559 9274
rect 7559 9222 7571 9274
rect 7571 9222 7585 9274
rect 7609 9222 7623 9274
rect 7623 9222 7635 9274
rect 7635 9222 7665 9274
rect 7689 9222 7699 9274
rect 7699 9222 7745 9274
rect 7449 9220 7505 9222
rect 7529 9220 7585 9222
rect 7609 9220 7665 9222
rect 7689 9220 7745 9222
rect 7449 8186 7505 8188
rect 7529 8186 7585 8188
rect 7609 8186 7665 8188
rect 7689 8186 7745 8188
rect 7449 8134 7495 8186
rect 7495 8134 7505 8186
rect 7529 8134 7559 8186
rect 7559 8134 7571 8186
rect 7571 8134 7585 8186
rect 7609 8134 7623 8186
rect 7623 8134 7635 8186
rect 7635 8134 7665 8186
rect 7689 8134 7699 8186
rect 7699 8134 7745 8186
rect 7449 8132 7505 8134
rect 7529 8132 7585 8134
rect 7609 8132 7665 8134
rect 7689 8132 7745 8134
rect 6734 3984 6790 4040
rect 6150 3290 6206 3292
rect 6230 3290 6286 3292
rect 6310 3290 6366 3292
rect 6390 3290 6446 3292
rect 6150 3238 6196 3290
rect 6196 3238 6206 3290
rect 6230 3238 6260 3290
rect 6260 3238 6272 3290
rect 6272 3238 6286 3290
rect 6310 3238 6324 3290
rect 6324 3238 6336 3290
rect 6336 3238 6366 3290
rect 6390 3238 6400 3290
rect 6400 3238 6446 3290
rect 6150 3236 6206 3238
rect 6230 3236 6286 3238
rect 6310 3236 6366 3238
rect 6390 3236 6446 3238
rect 3553 2202 3609 2204
rect 3633 2202 3689 2204
rect 3713 2202 3769 2204
rect 3793 2202 3849 2204
rect 3553 2150 3599 2202
rect 3599 2150 3609 2202
rect 3633 2150 3663 2202
rect 3663 2150 3675 2202
rect 3675 2150 3689 2202
rect 3713 2150 3727 2202
rect 3727 2150 3739 2202
rect 3739 2150 3769 2202
rect 3793 2150 3803 2202
rect 3803 2150 3849 2202
rect 3553 2148 3609 2150
rect 3633 2148 3689 2150
rect 3713 2148 3769 2150
rect 3793 2148 3849 2150
rect 6150 2202 6206 2204
rect 6230 2202 6286 2204
rect 6310 2202 6366 2204
rect 6390 2202 6446 2204
rect 6150 2150 6196 2202
rect 6196 2150 6206 2202
rect 6230 2150 6260 2202
rect 6260 2150 6272 2202
rect 6272 2150 6286 2202
rect 6310 2150 6324 2202
rect 6324 2150 6336 2202
rect 6336 2150 6366 2202
rect 6390 2150 6400 2202
rect 6400 2150 6446 2202
rect 6150 2148 6206 2150
rect 6230 2148 6286 2150
rect 6310 2148 6366 2150
rect 6390 2148 6446 2150
rect 7449 7098 7505 7100
rect 7529 7098 7585 7100
rect 7609 7098 7665 7100
rect 7689 7098 7745 7100
rect 7449 7046 7495 7098
rect 7495 7046 7505 7098
rect 7529 7046 7559 7098
rect 7559 7046 7571 7098
rect 7571 7046 7585 7098
rect 7609 7046 7623 7098
rect 7623 7046 7635 7098
rect 7635 7046 7665 7098
rect 7689 7046 7699 7098
rect 7699 7046 7745 7098
rect 7449 7044 7505 7046
rect 7529 7044 7585 7046
rect 7609 7044 7665 7046
rect 7689 7044 7745 7046
rect 7449 6010 7505 6012
rect 7529 6010 7585 6012
rect 7609 6010 7665 6012
rect 7689 6010 7745 6012
rect 7449 5958 7495 6010
rect 7495 5958 7505 6010
rect 7529 5958 7559 6010
rect 7559 5958 7571 6010
rect 7571 5958 7585 6010
rect 7609 5958 7623 6010
rect 7623 5958 7635 6010
rect 7635 5958 7665 6010
rect 7689 5958 7699 6010
rect 7699 5958 7745 6010
rect 7449 5956 7505 5958
rect 7529 5956 7585 5958
rect 7609 5956 7665 5958
rect 7689 5956 7745 5958
rect 7449 4922 7505 4924
rect 7529 4922 7585 4924
rect 7609 4922 7665 4924
rect 7689 4922 7745 4924
rect 7449 4870 7495 4922
rect 7495 4870 7505 4922
rect 7529 4870 7559 4922
rect 7559 4870 7571 4922
rect 7571 4870 7585 4922
rect 7609 4870 7623 4922
rect 7623 4870 7635 4922
rect 7635 4870 7665 4922
rect 7689 4870 7699 4922
rect 7699 4870 7745 4922
rect 7449 4868 7505 4870
rect 7529 4868 7585 4870
rect 7609 4868 7665 4870
rect 7689 4868 7745 4870
rect 7449 3834 7505 3836
rect 7529 3834 7585 3836
rect 7609 3834 7665 3836
rect 7689 3834 7745 3836
rect 7449 3782 7495 3834
rect 7495 3782 7505 3834
rect 7529 3782 7559 3834
rect 7559 3782 7571 3834
rect 7571 3782 7585 3834
rect 7609 3782 7623 3834
rect 7623 3782 7635 3834
rect 7635 3782 7665 3834
rect 7689 3782 7699 3834
rect 7699 3782 7745 3834
rect 7449 3780 7505 3782
rect 7529 3780 7585 3782
rect 7609 3780 7665 3782
rect 7689 3780 7745 3782
rect 7449 2746 7505 2748
rect 7529 2746 7585 2748
rect 7609 2746 7665 2748
rect 7689 2746 7745 2748
rect 7449 2694 7495 2746
rect 7495 2694 7505 2746
rect 7529 2694 7559 2746
rect 7559 2694 7571 2746
rect 7571 2694 7585 2746
rect 7609 2694 7623 2746
rect 7623 2694 7635 2746
rect 7635 2694 7665 2746
rect 7689 2694 7699 2746
rect 7699 2694 7745 2746
rect 7449 2692 7505 2694
rect 7529 2692 7585 2694
rect 7609 2692 7665 2694
rect 7689 2692 7745 2694
rect 7654 1672 7710 1728
rect 8298 5208 8354 5264
rect 8114 2896 8170 2952
rect 7930 584 7986 640
<< metal3 >>
rect 8201 29474 8267 29477
rect 9200 29474 10000 29504
rect 8201 29472 10000 29474
rect 8201 29416 8206 29472
rect 8262 29416 10000 29472
rect 8201 29414 10000 29416
rect 8201 29411 8267 29414
rect 9200 29384 10000 29414
rect 5533 28386 5599 28389
rect 9200 28386 10000 28416
rect 5533 28384 10000 28386
rect 5533 28328 5538 28384
rect 5594 28328 10000 28384
rect 5533 28326 10000 28328
rect 5533 28323 5599 28326
rect 9200 28296 10000 28326
rect 2242 27776 2562 27777
rect 2242 27712 2250 27776
rect 2314 27712 2330 27776
rect 2394 27712 2410 27776
rect 2474 27712 2490 27776
rect 2554 27712 2562 27776
rect 2242 27711 2562 27712
rect 4840 27776 5160 27777
rect 4840 27712 4848 27776
rect 4912 27712 4928 27776
rect 4992 27712 5008 27776
rect 5072 27712 5088 27776
rect 5152 27712 5160 27776
rect 4840 27711 5160 27712
rect 7437 27776 7757 27777
rect 7437 27712 7445 27776
rect 7509 27712 7525 27776
rect 7589 27712 7605 27776
rect 7669 27712 7685 27776
rect 7749 27712 7757 27776
rect 7437 27711 7757 27712
rect 3541 27232 3861 27233
rect 3541 27168 3549 27232
rect 3613 27168 3629 27232
rect 3693 27168 3709 27232
rect 3773 27168 3789 27232
rect 3853 27168 3861 27232
rect 3541 27167 3861 27168
rect 6138 27232 6458 27233
rect 6138 27168 6146 27232
rect 6210 27168 6226 27232
rect 6290 27168 6306 27232
rect 6370 27168 6386 27232
rect 6450 27168 6458 27232
rect 6138 27167 6458 27168
rect 6729 27162 6795 27165
rect 9200 27162 10000 27192
rect 6729 27160 10000 27162
rect 6729 27104 6734 27160
rect 6790 27104 10000 27160
rect 6729 27102 10000 27104
rect 6729 27099 6795 27102
rect 9200 27072 10000 27102
rect 2242 26688 2562 26689
rect 2242 26624 2250 26688
rect 2314 26624 2330 26688
rect 2394 26624 2410 26688
rect 2474 26624 2490 26688
rect 2554 26624 2562 26688
rect 2242 26623 2562 26624
rect 4840 26688 5160 26689
rect 4840 26624 4848 26688
rect 4912 26624 4928 26688
rect 4992 26624 5008 26688
rect 5072 26624 5088 26688
rect 5152 26624 5160 26688
rect 4840 26623 5160 26624
rect 7437 26688 7757 26689
rect 7437 26624 7445 26688
rect 7509 26624 7525 26688
rect 7589 26624 7605 26688
rect 7669 26624 7685 26688
rect 7749 26624 7757 26688
rect 7437 26623 7757 26624
rect 3541 26144 3861 26145
rect 3541 26080 3549 26144
rect 3613 26080 3629 26144
rect 3693 26080 3709 26144
rect 3773 26080 3789 26144
rect 3853 26080 3861 26144
rect 3541 26079 3861 26080
rect 6138 26144 6458 26145
rect 6138 26080 6146 26144
rect 6210 26080 6226 26144
rect 6290 26080 6306 26144
rect 6370 26080 6386 26144
rect 6450 26080 6458 26144
rect 6138 26079 6458 26080
rect 7833 26074 7899 26077
rect 9200 26074 10000 26104
rect 7833 26072 10000 26074
rect 7833 26016 7838 26072
rect 7894 26016 10000 26072
rect 7833 26014 10000 26016
rect 7833 26011 7899 26014
rect 9200 25984 10000 26014
rect 2242 25600 2562 25601
rect 2242 25536 2250 25600
rect 2314 25536 2330 25600
rect 2394 25536 2410 25600
rect 2474 25536 2490 25600
rect 2554 25536 2562 25600
rect 2242 25535 2562 25536
rect 4840 25600 5160 25601
rect 4840 25536 4848 25600
rect 4912 25536 4928 25600
rect 4992 25536 5008 25600
rect 5072 25536 5088 25600
rect 5152 25536 5160 25600
rect 4840 25535 5160 25536
rect 7437 25600 7757 25601
rect 7437 25536 7445 25600
rect 7509 25536 7525 25600
rect 7589 25536 7605 25600
rect 7669 25536 7685 25600
rect 7749 25536 7757 25600
rect 7437 25535 7757 25536
rect 3541 25056 3861 25057
rect 3541 24992 3549 25056
rect 3613 24992 3629 25056
rect 3693 24992 3709 25056
rect 3773 24992 3789 25056
rect 3853 24992 3861 25056
rect 3541 24991 3861 24992
rect 6138 25056 6458 25057
rect 6138 24992 6146 25056
rect 6210 24992 6226 25056
rect 6290 24992 6306 25056
rect 6370 24992 6386 25056
rect 6450 24992 6458 25056
rect 6138 24991 6458 24992
rect 8109 24850 8175 24853
rect 9200 24850 10000 24880
rect 8109 24848 10000 24850
rect 8109 24792 8114 24848
rect 8170 24792 10000 24848
rect 8109 24790 10000 24792
rect 8109 24787 8175 24790
rect 9200 24760 10000 24790
rect 2242 24512 2562 24513
rect 2242 24448 2250 24512
rect 2314 24448 2330 24512
rect 2394 24448 2410 24512
rect 2474 24448 2490 24512
rect 2554 24448 2562 24512
rect 2242 24447 2562 24448
rect 4840 24512 5160 24513
rect 4840 24448 4848 24512
rect 4912 24448 4928 24512
rect 4992 24448 5008 24512
rect 5072 24448 5088 24512
rect 5152 24448 5160 24512
rect 4840 24447 5160 24448
rect 7437 24512 7757 24513
rect 7437 24448 7445 24512
rect 7509 24448 7525 24512
rect 7589 24448 7605 24512
rect 7669 24448 7685 24512
rect 7749 24448 7757 24512
rect 7437 24447 7757 24448
rect 3541 23968 3861 23969
rect 3541 23904 3549 23968
rect 3613 23904 3629 23968
rect 3693 23904 3709 23968
rect 3773 23904 3789 23968
rect 3853 23904 3861 23968
rect 3541 23903 3861 23904
rect 6138 23968 6458 23969
rect 6138 23904 6146 23968
rect 6210 23904 6226 23968
rect 6290 23904 6306 23968
rect 6370 23904 6386 23968
rect 6450 23904 6458 23968
rect 6138 23903 6458 23904
rect 8293 23762 8359 23765
rect 9200 23762 10000 23792
rect 8293 23760 10000 23762
rect 8293 23704 8298 23760
rect 8354 23704 10000 23760
rect 8293 23702 10000 23704
rect 8293 23699 8359 23702
rect 9200 23672 10000 23702
rect 2242 23424 2562 23425
rect 2242 23360 2250 23424
rect 2314 23360 2330 23424
rect 2394 23360 2410 23424
rect 2474 23360 2490 23424
rect 2554 23360 2562 23424
rect 2242 23359 2562 23360
rect 4840 23424 5160 23425
rect 4840 23360 4848 23424
rect 4912 23360 4928 23424
rect 4992 23360 5008 23424
rect 5072 23360 5088 23424
rect 5152 23360 5160 23424
rect 4840 23359 5160 23360
rect 7437 23424 7757 23425
rect 7437 23360 7445 23424
rect 7509 23360 7525 23424
rect 7589 23360 7605 23424
rect 7669 23360 7685 23424
rect 7749 23360 7757 23424
rect 7437 23359 7757 23360
rect 3541 22880 3861 22881
rect 3541 22816 3549 22880
rect 3613 22816 3629 22880
rect 3693 22816 3709 22880
rect 3773 22816 3789 22880
rect 3853 22816 3861 22880
rect 3541 22815 3861 22816
rect 6138 22880 6458 22881
rect 6138 22816 6146 22880
rect 6210 22816 6226 22880
rect 6290 22816 6306 22880
rect 6370 22816 6386 22880
rect 6450 22816 6458 22880
rect 6138 22815 6458 22816
rect 5809 22538 5875 22541
rect 9200 22538 10000 22568
rect 5809 22536 10000 22538
rect 5809 22480 5814 22536
rect 5870 22480 10000 22536
rect 5809 22478 10000 22480
rect 5809 22475 5875 22478
rect 9200 22448 10000 22478
rect 2242 22336 2562 22337
rect 2242 22272 2250 22336
rect 2314 22272 2330 22336
rect 2394 22272 2410 22336
rect 2474 22272 2490 22336
rect 2554 22272 2562 22336
rect 2242 22271 2562 22272
rect 4840 22336 5160 22337
rect 4840 22272 4848 22336
rect 4912 22272 4928 22336
rect 4992 22272 5008 22336
rect 5072 22272 5088 22336
rect 5152 22272 5160 22336
rect 4840 22271 5160 22272
rect 7437 22336 7757 22337
rect 7437 22272 7445 22336
rect 7509 22272 7525 22336
rect 7589 22272 7605 22336
rect 7669 22272 7685 22336
rect 7749 22272 7757 22336
rect 7437 22271 7757 22272
rect 3541 21792 3861 21793
rect 3541 21728 3549 21792
rect 3613 21728 3629 21792
rect 3693 21728 3709 21792
rect 3773 21728 3789 21792
rect 3853 21728 3861 21792
rect 3541 21727 3861 21728
rect 6138 21792 6458 21793
rect 6138 21728 6146 21792
rect 6210 21728 6226 21792
rect 6290 21728 6306 21792
rect 6370 21728 6386 21792
rect 6450 21728 6458 21792
rect 6138 21727 6458 21728
rect 5349 21450 5415 21453
rect 9200 21450 10000 21480
rect 5349 21448 10000 21450
rect 5349 21392 5354 21448
rect 5410 21392 10000 21448
rect 5349 21390 10000 21392
rect 5349 21387 5415 21390
rect 9200 21360 10000 21390
rect 2242 21248 2562 21249
rect 2242 21184 2250 21248
rect 2314 21184 2330 21248
rect 2394 21184 2410 21248
rect 2474 21184 2490 21248
rect 2554 21184 2562 21248
rect 2242 21183 2562 21184
rect 4840 21248 5160 21249
rect 4840 21184 4848 21248
rect 4912 21184 4928 21248
rect 4992 21184 5008 21248
rect 5072 21184 5088 21248
rect 5152 21184 5160 21248
rect 4840 21183 5160 21184
rect 7437 21248 7757 21249
rect 7437 21184 7445 21248
rect 7509 21184 7525 21248
rect 7589 21184 7605 21248
rect 7669 21184 7685 21248
rect 7749 21184 7757 21248
rect 7437 21183 7757 21184
rect 3541 20704 3861 20705
rect 3541 20640 3549 20704
rect 3613 20640 3629 20704
rect 3693 20640 3709 20704
rect 3773 20640 3789 20704
rect 3853 20640 3861 20704
rect 3541 20639 3861 20640
rect 6138 20704 6458 20705
rect 6138 20640 6146 20704
rect 6210 20640 6226 20704
rect 6290 20640 6306 20704
rect 6370 20640 6386 20704
rect 6450 20640 6458 20704
rect 6138 20639 6458 20640
rect 9200 20226 10000 20256
rect 7974 20166 10000 20226
rect 2242 20160 2562 20161
rect 2242 20096 2250 20160
rect 2314 20096 2330 20160
rect 2394 20096 2410 20160
rect 2474 20096 2490 20160
rect 2554 20096 2562 20160
rect 2242 20095 2562 20096
rect 4840 20160 5160 20161
rect 4840 20096 4848 20160
rect 4912 20096 4928 20160
rect 4992 20096 5008 20160
rect 5072 20096 5088 20160
rect 5152 20096 5160 20160
rect 4840 20095 5160 20096
rect 7437 20160 7757 20161
rect 7437 20096 7445 20160
rect 7509 20096 7525 20160
rect 7589 20096 7605 20160
rect 7669 20096 7685 20160
rect 7749 20096 7757 20160
rect 7437 20095 7757 20096
rect 5533 19954 5599 19957
rect 7974 19954 8034 20166
rect 9200 20136 10000 20166
rect 5533 19952 8034 19954
rect 5533 19896 5538 19952
rect 5594 19896 8034 19952
rect 5533 19894 8034 19896
rect 5533 19891 5599 19894
rect 3541 19616 3861 19617
rect 3541 19552 3549 19616
rect 3613 19552 3629 19616
rect 3693 19552 3709 19616
rect 3773 19552 3789 19616
rect 3853 19552 3861 19616
rect 3541 19551 3861 19552
rect 6138 19616 6458 19617
rect 6138 19552 6146 19616
rect 6210 19552 6226 19616
rect 6290 19552 6306 19616
rect 6370 19552 6386 19616
rect 6450 19552 6458 19616
rect 6138 19551 6458 19552
rect 9200 19138 10000 19168
rect 7974 19078 10000 19138
rect 2242 19072 2562 19073
rect 2242 19008 2250 19072
rect 2314 19008 2330 19072
rect 2394 19008 2410 19072
rect 2474 19008 2490 19072
rect 2554 19008 2562 19072
rect 2242 19007 2562 19008
rect 4840 19072 5160 19073
rect 4840 19008 4848 19072
rect 4912 19008 4928 19072
rect 4992 19008 5008 19072
rect 5072 19008 5088 19072
rect 5152 19008 5160 19072
rect 4840 19007 5160 19008
rect 7437 19072 7757 19073
rect 7437 19008 7445 19072
rect 7509 19008 7525 19072
rect 7589 19008 7605 19072
rect 7669 19008 7685 19072
rect 7749 19008 7757 19072
rect 7437 19007 7757 19008
rect 6821 18866 6887 18869
rect 7974 18866 8034 19078
rect 9200 19048 10000 19078
rect 6821 18864 8034 18866
rect 6821 18808 6826 18864
rect 6882 18808 8034 18864
rect 6821 18806 8034 18808
rect 6821 18803 6887 18806
rect 3541 18528 3861 18529
rect 3541 18464 3549 18528
rect 3613 18464 3629 18528
rect 3693 18464 3709 18528
rect 3773 18464 3789 18528
rect 3853 18464 3861 18528
rect 3541 18463 3861 18464
rect 6138 18528 6458 18529
rect 6138 18464 6146 18528
rect 6210 18464 6226 18528
rect 6290 18464 6306 18528
rect 6370 18464 6386 18528
rect 6450 18464 6458 18528
rect 6138 18463 6458 18464
rect 2242 17984 2562 17985
rect 2242 17920 2250 17984
rect 2314 17920 2330 17984
rect 2394 17920 2410 17984
rect 2474 17920 2490 17984
rect 2554 17920 2562 17984
rect 2242 17919 2562 17920
rect 4840 17984 5160 17985
rect 4840 17920 4848 17984
rect 4912 17920 4928 17984
rect 4992 17920 5008 17984
rect 5072 17920 5088 17984
rect 5152 17920 5160 17984
rect 4840 17919 5160 17920
rect 7437 17984 7757 17985
rect 7437 17920 7445 17984
rect 7509 17920 7525 17984
rect 7589 17920 7605 17984
rect 7669 17920 7685 17984
rect 7749 17920 7757 17984
rect 7437 17919 7757 17920
rect 5993 17916 6059 17917
rect 5942 17852 5948 17916
rect 6012 17914 6059 17916
rect 9200 17914 10000 17944
rect 6012 17912 6104 17914
rect 6054 17856 6104 17912
rect 6012 17854 6104 17856
rect 7974 17854 10000 17914
rect 6012 17852 6059 17854
rect 5993 17851 6059 17852
rect 5993 17778 6059 17781
rect 7974 17778 8034 17854
rect 9200 17824 10000 17854
rect 5993 17776 8034 17778
rect 5993 17720 5998 17776
rect 6054 17720 8034 17776
rect 5993 17718 8034 17720
rect 5993 17715 6059 17718
rect 3541 17440 3861 17441
rect 3541 17376 3549 17440
rect 3613 17376 3629 17440
rect 3693 17376 3709 17440
rect 3773 17376 3789 17440
rect 3853 17376 3861 17440
rect 3541 17375 3861 17376
rect 6138 17440 6458 17441
rect 6138 17376 6146 17440
rect 6210 17376 6226 17440
rect 6290 17376 6306 17440
rect 6370 17376 6386 17440
rect 6450 17376 6458 17440
rect 6138 17375 6458 17376
rect 2242 16896 2562 16897
rect 2242 16832 2250 16896
rect 2314 16832 2330 16896
rect 2394 16832 2410 16896
rect 2474 16832 2490 16896
rect 2554 16832 2562 16896
rect 2242 16831 2562 16832
rect 4840 16896 5160 16897
rect 4840 16832 4848 16896
rect 4912 16832 4928 16896
rect 4992 16832 5008 16896
rect 5072 16832 5088 16896
rect 5152 16832 5160 16896
rect 4840 16831 5160 16832
rect 7437 16896 7757 16897
rect 7437 16832 7445 16896
rect 7509 16832 7525 16896
rect 7589 16832 7605 16896
rect 7669 16832 7685 16896
rect 7749 16832 7757 16896
rect 7437 16831 7757 16832
rect 8017 16826 8083 16829
rect 9200 16826 10000 16856
rect 8017 16824 10000 16826
rect 8017 16768 8022 16824
rect 8078 16768 10000 16824
rect 8017 16766 10000 16768
rect 8017 16763 8083 16766
rect 9200 16736 10000 16766
rect 3541 16352 3861 16353
rect 3541 16288 3549 16352
rect 3613 16288 3629 16352
rect 3693 16288 3709 16352
rect 3773 16288 3789 16352
rect 3853 16288 3861 16352
rect 3541 16287 3861 16288
rect 6138 16352 6458 16353
rect 6138 16288 6146 16352
rect 6210 16288 6226 16352
rect 6290 16288 6306 16352
rect 6370 16288 6386 16352
rect 6450 16288 6458 16352
rect 6138 16287 6458 16288
rect 2242 15808 2562 15809
rect 2242 15744 2250 15808
rect 2314 15744 2330 15808
rect 2394 15744 2410 15808
rect 2474 15744 2490 15808
rect 2554 15744 2562 15808
rect 2242 15743 2562 15744
rect 4840 15808 5160 15809
rect 4840 15744 4848 15808
rect 4912 15744 4928 15808
rect 4992 15744 5008 15808
rect 5072 15744 5088 15808
rect 5152 15744 5160 15808
rect 4840 15743 5160 15744
rect 7437 15808 7757 15809
rect 7437 15744 7445 15808
rect 7509 15744 7525 15808
rect 7589 15744 7605 15808
rect 7669 15744 7685 15808
rect 7749 15744 7757 15808
rect 7437 15743 7757 15744
rect 7925 15602 7991 15605
rect 9200 15602 10000 15632
rect 7925 15600 10000 15602
rect 7925 15544 7930 15600
rect 7986 15544 10000 15600
rect 7925 15542 10000 15544
rect 7925 15539 7991 15542
rect 9200 15512 10000 15542
rect 3541 15264 3861 15265
rect 3541 15200 3549 15264
rect 3613 15200 3629 15264
rect 3693 15200 3709 15264
rect 3773 15200 3789 15264
rect 3853 15200 3861 15264
rect 3541 15199 3861 15200
rect 6138 15264 6458 15265
rect 6138 15200 6146 15264
rect 6210 15200 6226 15264
rect 6290 15200 6306 15264
rect 6370 15200 6386 15264
rect 6450 15200 6458 15264
rect 6138 15199 6458 15200
rect 2242 14720 2562 14721
rect 2242 14656 2250 14720
rect 2314 14656 2330 14720
rect 2394 14656 2410 14720
rect 2474 14656 2490 14720
rect 2554 14656 2562 14720
rect 2242 14655 2562 14656
rect 4840 14720 5160 14721
rect 4840 14656 4848 14720
rect 4912 14656 4928 14720
rect 4992 14656 5008 14720
rect 5072 14656 5088 14720
rect 5152 14656 5160 14720
rect 4840 14655 5160 14656
rect 7437 14720 7757 14721
rect 7437 14656 7445 14720
rect 7509 14656 7525 14720
rect 7589 14656 7605 14720
rect 7669 14656 7685 14720
rect 7749 14656 7757 14720
rect 7437 14655 7757 14656
rect 6729 14514 6795 14517
rect 9200 14514 10000 14544
rect 6729 14512 10000 14514
rect 6729 14456 6734 14512
rect 6790 14456 10000 14512
rect 6729 14454 10000 14456
rect 6729 14451 6795 14454
rect 9200 14424 10000 14454
rect 3541 14176 3861 14177
rect 3541 14112 3549 14176
rect 3613 14112 3629 14176
rect 3693 14112 3709 14176
rect 3773 14112 3789 14176
rect 3853 14112 3861 14176
rect 3541 14111 3861 14112
rect 6138 14176 6458 14177
rect 6138 14112 6146 14176
rect 6210 14112 6226 14176
rect 6290 14112 6306 14176
rect 6370 14112 6386 14176
rect 6450 14112 6458 14176
rect 6138 14111 6458 14112
rect 2242 13632 2562 13633
rect 2242 13568 2250 13632
rect 2314 13568 2330 13632
rect 2394 13568 2410 13632
rect 2474 13568 2490 13632
rect 2554 13568 2562 13632
rect 2242 13567 2562 13568
rect 4840 13632 5160 13633
rect 4840 13568 4848 13632
rect 4912 13568 4928 13632
rect 4992 13568 5008 13632
rect 5072 13568 5088 13632
rect 5152 13568 5160 13632
rect 4840 13567 5160 13568
rect 7437 13632 7757 13633
rect 7437 13568 7445 13632
rect 7509 13568 7525 13632
rect 7589 13568 7605 13632
rect 7669 13568 7685 13632
rect 7749 13568 7757 13632
rect 7437 13567 7757 13568
rect 5717 13290 5783 13293
rect 9200 13290 10000 13320
rect 5717 13288 10000 13290
rect 5717 13232 5722 13288
rect 5778 13232 10000 13288
rect 5717 13230 10000 13232
rect 5717 13227 5783 13230
rect 9200 13200 10000 13230
rect 3541 13088 3861 13089
rect 3541 13024 3549 13088
rect 3613 13024 3629 13088
rect 3693 13024 3709 13088
rect 3773 13024 3789 13088
rect 3853 13024 3861 13088
rect 3541 13023 3861 13024
rect 6138 13088 6458 13089
rect 6138 13024 6146 13088
rect 6210 13024 6226 13088
rect 6290 13024 6306 13088
rect 6370 13024 6386 13088
rect 6450 13024 6458 13088
rect 6138 13023 6458 13024
rect 5993 12748 6059 12749
rect 5942 12746 5948 12748
rect 5902 12686 5948 12746
rect 6012 12744 6059 12748
rect 6054 12688 6059 12744
rect 5942 12684 5948 12686
rect 6012 12684 6059 12688
rect 5993 12683 6059 12684
rect 2242 12544 2562 12545
rect 2242 12480 2250 12544
rect 2314 12480 2330 12544
rect 2394 12480 2410 12544
rect 2474 12480 2490 12544
rect 2554 12480 2562 12544
rect 2242 12479 2562 12480
rect 4840 12544 5160 12545
rect 4840 12480 4848 12544
rect 4912 12480 4928 12544
rect 4992 12480 5008 12544
rect 5072 12480 5088 12544
rect 5152 12480 5160 12544
rect 4840 12479 5160 12480
rect 7437 12544 7757 12545
rect 7437 12480 7445 12544
rect 7509 12480 7525 12544
rect 7589 12480 7605 12544
rect 7669 12480 7685 12544
rect 7749 12480 7757 12544
rect 7437 12479 7757 12480
rect 5993 12336 6059 12341
rect 5993 12280 5998 12336
rect 6054 12280 6059 12336
rect 5993 12275 6059 12280
rect 5996 12202 6056 12275
rect 9200 12202 10000 12232
rect 5996 12142 10000 12202
rect 9200 12112 10000 12142
rect 3541 12000 3861 12001
rect 3541 11936 3549 12000
rect 3613 11936 3629 12000
rect 3693 11936 3709 12000
rect 3773 11936 3789 12000
rect 3853 11936 3861 12000
rect 3541 11935 3861 11936
rect 6138 12000 6458 12001
rect 6138 11936 6146 12000
rect 6210 11936 6226 12000
rect 6290 11936 6306 12000
rect 6370 11936 6386 12000
rect 6450 11936 6458 12000
rect 6138 11935 6458 11936
rect 2242 11456 2562 11457
rect 2242 11392 2250 11456
rect 2314 11392 2330 11456
rect 2394 11392 2410 11456
rect 2474 11392 2490 11456
rect 2554 11392 2562 11456
rect 2242 11391 2562 11392
rect 4840 11456 5160 11457
rect 4840 11392 4848 11456
rect 4912 11392 4928 11456
rect 4992 11392 5008 11456
rect 5072 11392 5088 11456
rect 5152 11392 5160 11456
rect 4840 11391 5160 11392
rect 7437 11456 7757 11457
rect 7437 11392 7445 11456
rect 7509 11392 7525 11456
rect 7589 11392 7605 11456
rect 7669 11392 7685 11456
rect 7749 11392 7757 11456
rect 7437 11391 7757 11392
rect 6637 10978 6703 10981
rect 9200 10978 10000 11008
rect 6637 10976 10000 10978
rect 6637 10920 6642 10976
rect 6698 10920 10000 10976
rect 6637 10918 10000 10920
rect 6637 10915 6703 10918
rect 3541 10912 3861 10913
rect 3541 10848 3549 10912
rect 3613 10848 3629 10912
rect 3693 10848 3709 10912
rect 3773 10848 3789 10912
rect 3853 10848 3861 10912
rect 3541 10847 3861 10848
rect 6138 10912 6458 10913
rect 6138 10848 6146 10912
rect 6210 10848 6226 10912
rect 6290 10848 6306 10912
rect 6370 10848 6386 10912
rect 6450 10848 6458 10912
rect 9200 10888 10000 10918
rect 6138 10847 6458 10848
rect 2242 10368 2562 10369
rect 2242 10304 2250 10368
rect 2314 10304 2330 10368
rect 2394 10304 2410 10368
rect 2474 10304 2490 10368
rect 2554 10304 2562 10368
rect 2242 10303 2562 10304
rect 4840 10368 5160 10369
rect 4840 10304 4848 10368
rect 4912 10304 4928 10368
rect 4992 10304 5008 10368
rect 5072 10304 5088 10368
rect 5152 10304 5160 10368
rect 4840 10303 5160 10304
rect 7437 10368 7757 10369
rect 7437 10304 7445 10368
rect 7509 10304 7525 10368
rect 7589 10304 7605 10368
rect 7669 10304 7685 10368
rect 7749 10304 7757 10368
rect 7437 10303 7757 10304
rect 5625 10026 5691 10029
rect 5625 10024 6746 10026
rect 5625 9968 5630 10024
rect 5686 9968 6746 10024
rect 5625 9966 6746 9968
rect 5625 9963 5691 9966
rect 6686 9890 6746 9966
rect 9200 9890 10000 9920
rect 6686 9830 10000 9890
rect 3541 9824 3861 9825
rect 3541 9760 3549 9824
rect 3613 9760 3629 9824
rect 3693 9760 3709 9824
rect 3773 9760 3789 9824
rect 3853 9760 3861 9824
rect 3541 9759 3861 9760
rect 6138 9824 6458 9825
rect 6138 9760 6146 9824
rect 6210 9760 6226 9824
rect 6290 9760 6306 9824
rect 6370 9760 6386 9824
rect 6450 9760 6458 9824
rect 9200 9800 10000 9830
rect 6138 9759 6458 9760
rect 2242 9280 2562 9281
rect 2242 9216 2250 9280
rect 2314 9216 2330 9280
rect 2394 9216 2410 9280
rect 2474 9216 2490 9280
rect 2554 9216 2562 9280
rect 2242 9215 2562 9216
rect 4840 9280 5160 9281
rect 4840 9216 4848 9280
rect 4912 9216 4928 9280
rect 4992 9216 5008 9280
rect 5072 9216 5088 9280
rect 5152 9216 5160 9280
rect 4840 9215 5160 9216
rect 7437 9280 7757 9281
rect 7437 9216 7445 9280
rect 7509 9216 7525 9280
rect 7589 9216 7605 9280
rect 7669 9216 7685 9280
rect 7749 9216 7757 9280
rect 7437 9215 7757 9216
rect 5717 8938 5783 8941
rect 5717 8936 6746 8938
rect 5717 8880 5722 8936
rect 5778 8880 6746 8936
rect 5717 8878 6746 8880
rect 5717 8875 5783 8878
rect 3541 8736 3861 8737
rect 3541 8672 3549 8736
rect 3613 8672 3629 8736
rect 3693 8672 3709 8736
rect 3773 8672 3789 8736
rect 3853 8672 3861 8736
rect 3541 8671 3861 8672
rect 6138 8736 6458 8737
rect 6138 8672 6146 8736
rect 6210 8672 6226 8736
rect 6290 8672 6306 8736
rect 6370 8672 6386 8736
rect 6450 8672 6458 8736
rect 6138 8671 6458 8672
rect 6686 8666 6746 8878
rect 9200 8666 10000 8696
rect 6686 8606 10000 8666
rect 9200 8576 10000 8606
rect 2242 8192 2562 8193
rect 2242 8128 2250 8192
rect 2314 8128 2330 8192
rect 2394 8128 2410 8192
rect 2474 8128 2490 8192
rect 2554 8128 2562 8192
rect 2242 8127 2562 8128
rect 4840 8192 5160 8193
rect 4840 8128 4848 8192
rect 4912 8128 4928 8192
rect 4992 8128 5008 8192
rect 5072 8128 5088 8192
rect 5152 8128 5160 8192
rect 4840 8127 5160 8128
rect 7437 8192 7757 8193
rect 7437 8128 7445 8192
rect 7509 8128 7525 8192
rect 7589 8128 7605 8192
rect 7669 8128 7685 8192
rect 7749 8128 7757 8192
rect 7437 8127 7757 8128
rect 3541 7648 3861 7649
rect 3541 7584 3549 7648
rect 3613 7584 3629 7648
rect 3693 7584 3709 7648
rect 3773 7584 3789 7648
rect 3853 7584 3861 7648
rect 3541 7583 3861 7584
rect 6138 7648 6458 7649
rect 6138 7584 6146 7648
rect 6210 7584 6226 7648
rect 6290 7584 6306 7648
rect 6370 7584 6386 7648
rect 6450 7584 6458 7648
rect 6138 7583 6458 7584
rect 6729 7578 6795 7581
rect 9200 7578 10000 7608
rect 6729 7576 10000 7578
rect 6729 7520 6734 7576
rect 6790 7520 10000 7576
rect 6729 7518 10000 7520
rect 6729 7515 6795 7518
rect 9200 7488 10000 7518
rect 2242 7104 2562 7105
rect 2242 7040 2250 7104
rect 2314 7040 2330 7104
rect 2394 7040 2410 7104
rect 2474 7040 2490 7104
rect 2554 7040 2562 7104
rect 2242 7039 2562 7040
rect 4840 7104 5160 7105
rect 4840 7040 4848 7104
rect 4912 7040 4928 7104
rect 4992 7040 5008 7104
rect 5072 7040 5088 7104
rect 5152 7040 5160 7104
rect 4840 7039 5160 7040
rect 7437 7104 7757 7105
rect 7437 7040 7445 7104
rect 7509 7040 7525 7104
rect 7589 7040 7605 7104
rect 7669 7040 7685 7104
rect 7749 7040 7757 7104
rect 7437 7039 7757 7040
rect 3541 6560 3861 6561
rect 3541 6496 3549 6560
rect 3613 6496 3629 6560
rect 3693 6496 3709 6560
rect 3773 6496 3789 6560
rect 3853 6496 3861 6560
rect 3541 6495 3861 6496
rect 6138 6560 6458 6561
rect 6138 6496 6146 6560
rect 6210 6496 6226 6560
rect 6290 6496 6306 6560
rect 6370 6496 6386 6560
rect 6450 6496 6458 6560
rect 6138 6495 6458 6496
rect 5993 6354 6059 6357
rect 9200 6354 10000 6384
rect 5993 6352 10000 6354
rect 5993 6296 5998 6352
rect 6054 6296 10000 6352
rect 5993 6294 10000 6296
rect 5993 6291 6059 6294
rect 9200 6264 10000 6294
rect 2242 6016 2562 6017
rect 2242 5952 2250 6016
rect 2314 5952 2330 6016
rect 2394 5952 2410 6016
rect 2474 5952 2490 6016
rect 2554 5952 2562 6016
rect 2242 5951 2562 5952
rect 4840 6016 5160 6017
rect 4840 5952 4848 6016
rect 4912 5952 4928 6016
rect 4992 5952 5008 6016
rect 5072 5952 5088 6016
rect 5152 5952 5160 6016
rect 4840 5951 5160 5952
rect 7437 6016 7757 6017
rect 7437 5952 7445 6016
rect 7509 5952 7525 6016
rect 7589 5952 7605 6016
rect 7669 5952 7685 6016
rect 7749 5952 7757 6016
rect 7437 5951 7757 5952
rect 3541 5472 3861 5473
rect 3541 5408 3549 5472
rect 3613 5408 3629 5472
rect 3693 5408 3709 5472
rect 3773 5408 3789 5472
rect 3853 5408 3861 5472
rect 3541 5407 3861 5408
rect 6138 5472 6458 5473
rect 6138 5408 6146 5472
rect 6210 5408 6226 5472
rect 6290 5408 6306 5472
rect 6370 5408 6386 5472
rect 6450 5408 6458 5472
rect 6138 5407 6458 5408
rect 8293 5266 8359 5269
rect 9200 5266 10000 5296
rect 8293 5264 10000 5266
rect 8293 5208 8298 5264
rect 8354 5208 10000 5264
rect 8293 5206 10000 5208
rect 8293 5203 8359 5206
rect 9200 5176 10000 5206
rect 2242 4928 2562 4929
rect 2242 4864 2250 4928
rect 2314 4864 2330 4928
rect 2394 4864 2410 4928
rect 2474 4864 2490 4928
rect 2554 4864 2562 4928
rect 2242 4863 2562 4864
rect 4840 4928 5160 4929
rect 4840 4864 4848 4928
rect 4912 4864 4928 4928
rect 4992 4864 5008 4928
rect 5072 4864 5088 4928
rect 5152 4864 5160 4928
rect 4840 4863 5160 4864
rect 7437 4928 7757 4929
rect 7437 4864 7445 4928
rect 7509 4864 7525 4928
rect 7589 4864 7605 4928
rect 7669 4864 7685 4928
rect 7749 4864 7757 4928
rect 7437 4863 7757 4864
rect 3541 4384 3861 4385
rect 3541 4320 3549 4384
rect 3613 4320 3629 4384
rect 3693 4320 3709 4384
rect 3773 4320 3789 4384
rect 3853 4320 3861 4384
rect 3541 4319 3861 4320
rect 6138 4384 6458 4385
rect 6138 4320 6146 4384
rect 6210 4320 6226 4384
rect 6290 4320 6306 4384
rect 6370 4320 6386 4384
rect 6450 4320 6458 4384
rect 6138 4319 6458 4320
rect 6729 4042 6795 4045
rect 9200 4042 10000 4072
rect 6729 4040 10000 4042
rect 6729 3984 6734 4040
rect 6790 3984 10000 4040
rect 6729 3982 10000 3984
rect 6729 3979 6795 3982
rect 9200 3952 10000 3982
rect 2242 3840 2562 3841
rect 2242 3776 2250 3840
rect 2314 3776 2330 3840
rect 2394 3776 2410 3840
rect 2474 3776 2490 3840
rect 2554 3776 2562 3840
rect 2242 3775 2562 3776
rect 4840 3840 5160 3841
rect 4840 3776 4848 3840
rect 4912 3776 4928 3840
rect 4992 3776 5008 3840
rect 5072 3776 5088 3840
rect 5152 3776 5160 3840
rect 4840 3775 5160 3776
rect 7437 3840 7757 3841
rect 7437 3776 7445 3840
rect 7509 3776 7525 3840
rect 7589 3776 7605 3840
rect 7669 3776 7685 3840
rect 7749 3776 7757 3840
rect 7437 3775 7757 3776
rect 3541 3296 3861 3297
rect 3541 3232 3549 3296
rect 3613 3232 3629 3296
rect 3693 3232 3709 3296
rect 3773 3232 3789 3296
rect 3853 3232 3861 3296
rect 3541 3231 3861 3232
rect 6138 3296 6458 3297
rect 6138 3232 6146 3296
rect 6210 3232 6226 3296
rect 6290 3232 6306 3296
rect 6370 3232 6386 3296
rect 6450 3232 6458 3296
rect 6138 3231 6458 3232
rect 8109 2954 8175 2957
rect 9200 2954 10000 2984
rect 8109 2952 10000 2954
rect 8109 2896 8114 2952
rect 8170 2896 10000 2952
rect 8109 2894 10000 2896
rect 8109 2891 8175 2894
rect 9200 2864 10000 2894
rect 2242 2752 2562 2753
rect 2242 2688 2250 2752
rect 2314 2688 2330 2752
rect 2394 2688 2410 2752
rect 2474 2688 2490 2752
rect 2554 2688 2562 2752
rect 2242 2687 2562 2688
rect 4840 2752 5160 2753
rect 4840 2688 4848 2752
rect 4912 2688 4928 2752
rect 4992 2688 5008 2752
rect 5072 2688 5088 2752
rect 5152 2688 5160 2752
rect 4840 2687 5160 2688
rect 7437 2752 7757 2753
rect 7437 2688 7445 2752
rect 7509 2688 7525 2752
rect 7589 2688 7605 2752
rect 7669 2688 7685 2752
rect 7749 2688 7757 2752
rect 7437 2687 7757 2688
rect 3541 2208 3861 2209
rect 3541 2144 3549 2208
rect 3613 2144 3629 2208
rect 3693 2144 3709 2208
rect 3773 2144 3789 2208
rect 3853 2144 3861 2208
rect 3541 2143 3861 2144
rect 6138 2208 6458 2209
rect 6138 2144 6146 2208
rect 6210 2144 6226 2208
rect 6290 2144 6306 2208
rect 6370 2144 6386 2208
rect 6450 2144 6458 2208
rect 6138 2143 6458 2144
rect 7649 1730 7715 1733
rect 9200 1730 10000 1760
rect 7649 1728 10000 1730
rect 7649 1672 7654 1728
rect 7710 1672 10000 1728
rect 7649 1670 10000 1672
rect 7649 1667 7715 1670
rect 9200 1640 10000 1670
rect 7925 642 7991 645
rect 9200 642 10000 672
rect 7925 640 10000 642
rect 7925 584 7930 640
rect 7986 584 10000 640
rect 7925 582 10000 584
rect 7925 579 7991 582
rect 9200 552 10000 582
<< via3 >>
rect 2250 27772 2314 27776
rect 2250 27716 2254 27772
rect 2254 27716 2310 27772
rect 2310 27716 2314 27772
rect 2250 27712 2314 27716
rect 2330 27772 2394 27776
rect 2330 27716 2334 27772
rect 2334 27716 2390 27772
rect 2390 27716 2394 27772
rect 2330 27712 2394 27716
rect 2410 27772 2474 27776
rect 2410 27716 2414 27772
rect 2414 27716 2470 27772
rect 2470 27716 2474 27772
rect 2410 27712 2474 27716
rect 2490 27772 2554 27776
rect 2490 27716 2494 27772
rect 2494 27716 2550 27772
rect 2550 27716 2554 27772
rect 2490 27712 2554 27716
rect 4848 27772 4912 27776
rect 4848 27716 4852 27772
rect 4852 27716 4908 27772
rect 4908 27716 4912 27772
rect 4848 27712 4912 27716
rect 4928 27772 4992 27776
rect 4928 27716 4932 27772
rect 4932 27716 4988 27772
rect 4988 27716 4992 27772
rect 4928 27712 4992 27716
rect 5008 27772 5072 27776
rect 5008 27716 5012 27772
rect 5012 27716 5068 27772
rect 5068 27716 5072 27772
rect 5008 27712 5072 27716
rect 5088 27772 5152 27776
rect 5088 27716 5092 27772
rect 5092 27716 5148 27772
rect 5148 27716 5152 27772
rect 5088 27712 5152 27716
rect 7445 27772 7509 27776
rect 7445 27716 7449 27772
rect 7449 27716 7505 27772
rect 7505 27716 7509 27772
rect 7445 27712 7509 27716
rect 7525 27772 7589 27776
rect 7525 27716 7529 27772
rect 7529 27716 7585 27772
rect 7585 27716 7589 27772
rect 7525 27712 7589 27716
rect 7605 27772 7669 27776
rect 7605 27716 7609 27772
rect 7609 27716 7665 27772
rect 7665 27716 7669 27772
rect 7605 27712 7669 27716
rect 7685 27772 7749 27776
rect 7685 27716 7689 27772
rect 7689 27716 7745 27772
rect 7745 27716 7749 27772
rect 7685 27712 7749 27716
rect 3549 27228 3613 27232
rect 3549 27172 3553 27228
rect 3553 27172 3609 27228
rect 3609 27172 3613 27228
rect 3549 27168 3613 27172
rect 3629 27228 3693 27232
rect 3629 27172 3633 27228
rect 3633 27172 3689 27228
rect 3689 27172 3693 27228
rect 3629 27168 3693 27172
rect 3709 27228 3773 27232
rect 3709 27172 3713 27228
rect 3713 27172 3769 27228
rect 3769 27172 3773 27228
rect 3709 27168 3773 27172
rect 3789 27228 3853 27232
rect 3789 27172 3793 27228
rect 3793 27172 3849 27228
rect 3849 27172 3853 27228
rect 3789 27168 3853 27172
rect 6146 27228 6210 27232
rect 6146 27172 6150 27228
rect 6150 27172 6206 27228
rect 6206 27172 6210 27228
rect 6146 27168 6210 27172
rect 6226 27228 6290 27232
rect 6226 27172 6230 27228
rect 6230 27172 6286 27228
rect 6286 27172 6290 27228
rect 6226 27168 6290 27172
rect 6306 27228 6370 27232
rect 6306 27172 6310 27228
rect 6310 27172 6366 27228
rect 6366 27172 6370 27228
rect 6306 27168 6370 27172
rect 6386 27228 6450 27232
rect 6386 27172 6390 27228
rect 6390 27172 6446 27228
rect 6446 27172 6450 27228
rect 6386 27168 6450 27172
rect 2250 26684 2314 26688
rect 2250 26628 2254 26684
rect 2254 26628 2310 26684
rect 2310 26628 2314 26684
rect 2250 26624 2314 26628
rect 2330 26684 2394 26688
rect 2330 26628 2334 26684
rect 2334 26628 2390 26684
rect 2390 26628 2394 26684
rect 2330 26624 2394 26628
rect 2410 26684 2474 26688
rect 2410 26628 2414 26684
rect 2414 26628 2470 26684
rect 2470 26628 2474 26684
rect 2410 26624 2474 26628
rect 2490 26684 2554 26688
rect 2490 26628 2494 26684
rect 2494 26628 2550 26684
rect 2550 26628 2554 26684
rect 2490 26624 2554 26628
rect 4848 26684 4912 26688
rect 4848 26628 4852 26684
rect 4852 26628 4908 26684
rect 4908 26628 4912 26684
rect 4848 26624 4912 26628
rect 4928 26684 4992 26688
rect 4928 26628 4932 26684
rect 4932 26628 4988 26684
rect 4988 26628 4992 26684
rect 4928 26624 4992 26628
rect 5008 26684 5072 26688
rect 5008 26628 5012 26684
rect 5012 26628 5068 26684
rect 5068 26628 5072 26684
rect 5008 26624 5072 26628
rect 5088 26684 5152 26688
rect 5088 26628 5092 26684
rect 5092 26628 5148 26684
rect 5148 26628 5152 26684
rect 5088 26624 5152 26628
rect 7445 26684 7509 26688
rect 7445 26628 7449 26684
rect 7449 26628 7505 26684
rect 7505 26628 7509 26684
rect 7445 26624 7509 26628
rect 7525 26684 7589 26688
rect 7525 26628 7529 26684
rect 7529 26628 7585 26684
rect 7585 26628 7589 26684
rect 7525 26624 7589 26628
rect 7605 26684 7669 26688
rect 7605 26628 7609 26684
rect 7609 26628 7665 26684
rect 7665 26628 7669 26684
rect 7605 26624 7669 26628
rect 7685 26684 7749 26688
rect 7685 26628 7689 26684
rect 7689 26628 7745 26684
rect 7745 26628 7749 26684
rect 7685 26624 7749 26628
rect 3549 26140 3613 26144
rect 3549 26084 3553 26140
rect 3553 26084 3609 26140
rect 3609 26084 3613 26140
rect 3549 26080 3613 26084
rect 3629 26140 3693 26144
rect 3629 26084 3633 26140
rect 3633 26084 3689 26140
rect 3689 26084 3693 26140
rect 3629 26080 3693 26084
rect 3709 26140 3773 26144
rect 3709 26084 3713 26140
rect 3713 26084 3769 26140
rect 3769 26084 3773 26140
rect 3709 26080 3773 26084
rect 3789 26140 3853 26144
rect 3789 26084 3793 26140
rect 3793 26084 3849 26140
rect 3849 26084 3853 26140
rect 3789 26080 3853 26084
rect 6146 26140 6210 26144
rect 6146 26084 6150 26140
rect 6150 26084 6206 26140
rect 6206 26084 6210 26140
rect 6146 26080 6210 26084
rect 6226 26140 6290 26144
rect 6226 26084 6230 26140
rect 6230 26084 6286 26140
rect 6286 26084 6290 26140
rect 6226 26080 6290 26084
rect 6306 26140 6370 26144
rect 6306 26084 6310 26140
rect 6310 26084 6366 26140
rect 6366 26084 6370 26140
rect 6306 26080 6370 26084
rect 6386 26140 6450 26144
rect 6386 26084 6390 26140
rect 6390 26084 6446 26140
rect 6446 26084 6450 26140
rect 6386 26080 6450 26084
rect 2250 25596 2314 25600
rect 2250 25540 2254 25596
rect 2254 25540 2310 25596
rect 2310 25540 2314 25596
rect 2250 25536 2314 25540
rect 2330 25596 2394 25600
rect 2330 25540 2334 25596
rect 2334 25540 2390 25596
rect 2390 25540 2394 25596
rect 2330 25536 2394 25540
rect 2410 25596 2474 25600
rect 2410 25540 2414 25596
rect 2414 25540 2470 25596
rect 2470 25540 2474 25596
rect 2410 25536 2474 25540
rect 2490 25596 2554 25600
rect 2490 25540 2494 25596
rect 2494 25540 2550 25596
rect 2550 25540 2554 25596
rect 2490 25536 2554 25540
rect 4848 25596 4912 25600
rect 4848 25540 4852 25596
rect 4852 25540 4908 25596
rect 4908 25540 4912 25596
rect 4848 25536 4912 25540
rect 4928 25596 4992 25600
rect 4928 25540 4932 25596
rect 4932 25540 4988 25596
rect 4988 25540 4992 25596
rect 4928 25536 4992 25540
rect 5008 25596 5072 25600
rect 5008 25540 5012 25596
rect 5012 25540 5068 25596
rect 5068 25540 5072 25596
rect 5008 25536 5072 25540
rect 5088 25596 5152 25600
rect 5088 25540 5092 25596
rect 5092 25540 5148 25596
rect 5148 25540 5152 25596
rect 5088 25536 5152 25540
rect 7445 25596 7509 25600
rect 7445 25540 7449 25596
rect 7449 25540 7505 25596
rect 7505 25540 7509 25596
rect 7445 25536 7509 25540
rect 7525 25596 7589 25600
rect 7525 25540 7529 25596
rect 7529 25540 7585 25596
rect 7585 25540 7589 25596
rect 7525 25536 7589 25540
rect 7605 25596 7669 25600
rect 7605 25540 7609 25596
rect 7609 25540 7665 25596
rect 7665 25540 7669 25596
rect 7605 25536 7669 25540
rect 7685 25596 7749 25600
rect 7685 25540 7689 25596
rect 7689 25540 7745 25596
rect 7745 25540 7749 25596
rect 7685 25536 7749 25540
rect 3549 25052 3613 25056
rect 3549 24996 3553 25052
rect 3553 24996 3609 25052
rect 3609 24996 3613 25052
rect 3549 24992 3613 24996
rect 3629 25052 3693 25056
rect 3629 24996 3633 25052
rect 3633 24996 3689 25052
rect 3689 24996 3693 25052
rect 3629 24992 3693 24996
rect 3709 25052 3773 25056
rect 3709 24996 3713 25052
rect 3713 24996 3769 25052
rect 3769 24996 3773 25052
rect 3709 24992 3773 24996
rect 3789 25052 3853 25056
rect 3789 24996 3793 25052
rect 3793 24996 3849 25052
rect 3849 24996 3853 25052
rect 3789 24992 3853 24996
rect 6146 25052 6210 25056
rect 6146 24996 6150 25052
rect 6150 24996 6206 25052
rect 6206 24996 6210 25052
rect 6146 24992 6210 24996
rect 6226 25052 6290 25056
rect 6226 24996 6230 25052
rect 6230 24996 6286 25052
rect 6286 24996 6290 25052
rect 6226 24992 6290 24996
rect 6306 25052 6370 25056
rect 6306 24996 6310 25052
rect 6310 24996 6366 25052
rect 6366 24996 6370 25052
rect 6306 24992 6370 24996
rect 6386 25052 6450 25056
rect 6386 24996 6390 25052
rect 6390 24996 6446 25052
rect 6446 24996 6450 25052
rect 6386 24992 6450 24996
rect 2250 24508 2314 24512
rect 2250 24452 2254 24508
rect 2254 24452 2310 24508
rect 2310 24452 2314 24508
rect 2250 24448 2314 24452
rect 2330 24508 2394 24512
rect 2330 24452 2334 24508
rect 2334 24452 2390 24508
rect 2390 24452 2394 24508
rect 2330 24448 2394 24452
rect 2410 24508 2474 24512
rect 2410 24452 2414 24508
rect 2414 24452 2470 24508
rect 2470 24452 2474 24508
rect 2410 24448 2474 24452
rect 2490 24508 2554 24512
rect 2490 24452 2494 24508
rect 2494 24452 2550 24508
rect 2550 24452 2554 24508
rect 2490 24448 2554 24452
rect 4848 24508 4912 24512
rect 4848 24452 4852 24508
rect 4852 24452 4908 24508
rect 4908 24452 4912 24508
rect 4848 24448 4912 24452
rect 4928 24508 4992 24512
rect 4928 24452 4932 24508
rect 4932 24452 4988 24508
rect 4988 24452 4992 24508
rect 4928 24448 4992 24452
rect 5008 24508 5072 24512
rect 5008 24452 5012 24508
rect 5012 24452 5068 24508
rect 5068 24452 5072 24508
rect 5008 24448 5072 24452
rect 5088 24508 5152 24512
rect 5088 24452 5092 24508
rect 5092 24452 5148 24508
rect 5148 24452 5152 24508
rect 5088 24448 5152 24452
rect 7445 24508 7509 24512
rect 7445 24452 7449 24508
rect 7449 24452 7505 24508
rect 7505 24452 7509 24508
rect 7445 24448 7509 24452
rect 7525 24508 7589 24512
rect 7525 24452 7529 24508
rect 7529 24452 7585 24508
rect 7585 24452 7589 24508
rect 7525 24448 7589 24452
rect 7605 24508 7669 24512
rect 7605 24452 7609 24508
rect 7609 24452 7665 24508
rect 7665 24452 7669 24508
rect 7605 24448 7669 24452
rect 7685 24508 7749 24512
rect 7685 24452 7689 24508
rect 7689 24452 7745 24508
rect 7745 24452 7749 24508
rect 7685 24448 7749 24452
rect 3549 23964 3613 23968
rect 3549 23908 3553 23964
rect 3553 23908 3609 23964
rect 3609 23908 3613 23964
rect 3549 23904 3613 23908
rect 3629 23964 3693 23968
rect 3629 23908 3633 23964
rect 3633 23908 3689 23964
rect 3689 23908 3693 23964
rect 3629 23904 3693 23908
rect 3709 23964 3773 23968
rect 3709 23908 3713 23964
rect 3713 23908 3769 23964
rect 3769 23908 3773 23964
rect 3709 23904 3773 23908
rect 3789 23964 3853 23968
rect 3789 23908 3793 23964
rect 3793 23908 3849 23964
rect 3849 23908 3853 23964
rect 3789 23904 3853 23908
rect 6146 23964 6210 23968
rect 6146 23908 6150 23964
rect 6150 23908 6206 23964
rect 6206 23908 6210 23964
rect 6146 23904 6210 23908
rect 6226 23964 6290 23968
rect 6226 23908 6230 23964
rect 6230 23908 6286 23964
rect 6286 23908 6290 23964
rect 6226 23904 6290 23908
rect 6306 23964 6370 23968
rect 6306 23908 6310 23964
rect 6310 23908 6366 23964
rect 6366 23908 6370 23964
rect 6306 23904 6370 23908
rect 6386 23964 6450 23968
rect 6386 23908 6390 23964
rect 6390 23908 6446 23964
rect 6446 23908 6450 23964
rect 6386 23904 6450 23908
rect 2250 23420 2314 23424
rect 2250 23364 2254 23420
rect 2254 23364 2310 23420
rect 2310 23364 2314 23420
rect 2250 23360 2314 23364
rect 2330 23420 2394 23424
rect 2330 23364 2334 23420
rect 2334 23364 2390 23420
rect 2390 23364 2394 23420
rect 2330 23360 2394 23364
rect 2410 23420 2474 23424
rect 2410 23364 2414 23420
rect 2414 23364 2470 23420
rect 2470 23364 2474 23420
rect 2410 23360 2474 23364
rect 2490 23420 2554 23424
rect 2490 23364 2494 23420
rect 2494 23364 2550 23420
rect 2550 23364 2554 23420
rect 2490 23360 2554 23364
rect 4848 23420 4912 23424
rect 4848 23364 4852 23420
rect 4852 23364 4908 23420
rect 4908 23364 4912 23420
rect 4848 23360 4912 23364
rect 4928 23420 4992 23424
rect 4928 23364 4932 23420
rect 4932 23364 4988 23420
rect 4988 23364 4992 23420
rect 4928 23360 4992 23364
rect 5008 23420 5072 23424
rect 5008 23364 5012 23420
rect 5012 23364 5068 23420
rect 5068 23364 5072 23420
rect 5008 23360 5072 23364
rect 5088 23420 5152 23424
rect 5088 23364 5092 23420
rect 5092 23364 5148 23420
rect 5148 23364 5152 23420
rect 5088 23360 5152 23364
rect 7445 23420 7509 23424
rect 7445 23364 7449 23420
rect 7449 23364 7505 23420
rect 7505 23364 7509 23420
rect 7445 23360 7509 23364
rect 7525 23420 7589 23424
rect 7525 23364 7529 23420
rect 7529 23364 7585 23420
rect 7585 23364 7589 23420
rect 7525 23360 7589 23364
rect 7605 23420 7669 23424
rect 7605 23364 7609 23420
rect 7609 23364 7665 23420
rect 7665 23364 7669 23420
rect 7605 23360 7669 23364
rect 7685 23420 7749 23424
rect 7685 23364 7689 23420
rect 7689 23364 7745 23420
rect 7745 23364 7749 23420
rect 7685 23360 7749 23364
rect 3549 22876 3613 22880
rect 3549 22820 3553 22876
rect 3553 22820 3609 22876
rect 3609 22820 3613 22876
rect 3549 22816 3613 22820
rect 3629 22876 3693 22880
rect 3629 22820 3633 22876
rect 3633 22820 3689 22876
rect 3689 22820 3693 22876
rect 3629 22816 3693 22820
rect 3709 22876 3773 22880
rect 3709 22820 3713 22876
rect 3713 22820 3769 22876
rect 3769 22820 3773 22876
rect 3709 22816 3773 22820
rect 3789 22876 3853 22880
rect 3789 22820 3793 22876
rect 3793 22820 3849 22876
rect 3849 22820 3853 22876
rect 3789 22816 3853 22820
rect 6146 22876 6210 22880
rect 6146 22820 6150 22876
rect 6150 22820 6206 22876
rect 6206 22820 6210 22876
rect 6146 22816 6210 22820
rect 6226 22876 6290 22880
rect 6226 22820 6230 22876
rect 6230 22820 6286 22876
rect 6286 22820 6290 22876
rect 6226 22816 6290 22820
rect 6306 22876 6370 22880
rect 6306 22820 6310 22876
rect 6310 22820 6366 22876
rect 6366 22820 6370 22876
rect 6306 22816 6370 22820
rect 6386 22876 6450 22880
rect 6386 22820 6390 22876
rect 6390 22820 6446 22876
rect 6446 22820 6450 22876
rect 6386 22816 6450 22820
rect 2250 22332 2314 22336
rect 2250 22276 2254 22332
rect 2254 22276 2310 22332
rect 2310 22276 2314 22332
rect 2250 22272 2314 22276
rect 2330 22332 2394 22336
rect 2330 22276 2334 22332
rect 2334 22276 2390 22332
rect 2390 22276 2394 22332
rect 2330 22272 2394 22276
rect 2410 22332 2474 22336
rect 2410 22276 2414 22332
rect 2414 22276 2470 22332
rect 2470 22276 2474 22332
rect 2410 22272 2474 22276
rect 2490 22332 2554 22336
rect 2490 22276 2494 22332
rect 2494 22276 2550 22332
rect 2550 22276 2554 22332
rect 2490 22272 2554 22276
rect 4848 22332 4912 22336
rect 4848 22276 4852 22332
rect 4852 22276 4908 22332
rect 4908 22276 4912 22332
rect 4848 22272 4912 22276
rect 4928 22332 4992 22336
rect 4928 22276 4932 22332
rect 4932 22276 4988 22332
rect 4988 22276 4992 22332
rect 4928 22272 4992 22276
rect 5008 22332 5072 22336
rect 5008 22276 5012 22332
rect 5012 22276 5068 22332
rect 5068 22276 5072 22332
rect 5008 22272 5072 22276
rect 5088 22332 5152 22336
rect 5088 22276 5092 22332
rect 5092 22276 5148 22332
rect 5148 22276 5152 22332
rect 5088 22272 5152 22276
rect 7445 22332 7509 22336
rect 7445 22276 7449 22332
rect 7449 22276 7505 22332
rect 7505 22276 7509 22332
rect 7445 22272 7509 22276
rect 7525 22332 7589 22336
rect 7525 22276 7529 22332
rect 7529 22276 7585 22332
rect 7585 22276 7589 22332
rect 7525 22272 7589 22276
rect 7605 22332 7669 22336
rect 7605 22276 7609 22332
rect 7609 22276 7665 22332
rect 7665 22276 7669 22332
rect 7605 22272 7669 22276
rect 7685 22332 7749 22336
rect 7685 22276 7689 22332
rect 7689 22276 7745 22332
rect 7745 22276 7749 22332
rect 7685 22272 7749 22276
rect 3549 21788 3613 21792
rect 3549 21732 3553 21788
rect 3553 21732 3609 21788
rect 3609 21732 3613 21788
rect 3549 21728 3613 21732
rect 3629 21788 3693 21792
rect 3629 21732 3633 21788
rect 3633 21732 3689 21788
rect 3689 21732 3693 21788
rect 3629 21728 3693 21732
rect 3709 21788 3773 21792
rect 3709 21732 3713 21788
rect 3713 21732 3769 21788
rect 3769 21732 3773 21788
rect 3709 21728 3773 21732
rect 3789 21788 3853 21792
rect 3789 21732 3793 21788
rect 3793 21732 3849 21788
rect 3849 21732 3853 21788
rect 3789 21728 3853 21732
rect 6146 21788 6210 21792
rect 6146 21732 6150 21788
rect 6150 21732 6206 21788
rect 6206 21732 6210 21788
rect 6146 21728 6210 21732
rect 6226 21788 6290 21792
rect 6226 21732 6230 21788
rect 6230 21732 6286 21788
rect 6286 21732 6290 21788
rect 6226 21728 6290 21732
rect 6306 21788 6370 21792
rect 6306 21732 6310 21788
rect 6310 21732 6366 21788
rect 6366 21732 6370 21788
rect 6306 21728 6370 21732
rect 6386 21788 6450 21792
rect 6386 21732 6390 21788
rect 6390 21732 6446 21788
rect 6446 21732 6450 21788
rect 6386 21728 6450 21732
rect 2250 21244 2314 21248
rect 2250 21188 2254 21244
rect 2254 21188 2310 21244
rect 2310 21188 2314 21244
rect 2250 21184 2314 21188
rect 2330 21244 2394 21248
rect 2330 21188 2334 21244
rect 2334 21188 2390 21244
rect 2390 21188 2394 21244
rect 2330 21184 2394 21188
rect 2410 21244 2474 21248
rect 2410 21188 2414 21244
rect 2414 21188 2470 21244
rect 2470 21188 2474 21244
rect 2410 21184 2474 21188
rect 2490 21244 2554 21248
rect 2490 21188 2494 21244
rect 2494 21188 2550 21244
rect 2550 21188 2554 21244
rect 2490 21184 2554 21188
rect 4848 21244 4912 21248
rect 4848 21188 4852 21244
rect 4852 21188 4908 21244
rect 4908 21188 4912 21244
rect 4848 21184 4912 21188
rect 4928 21244 4992 21248
rect 4928 21188 4932 21244
rect 4932 21188 4988 21244
rect 4988 21188 4992 21244
rect 4928 21184 4992 21188
rect 5008 21244 5072 21248
rect 5008 21188 5012 21244
rect 5012 21188 5068 21244
rect 5068 21188 5072 21244
rect 5008 21184 5072 21188
rect 5088 21244 5152 21248
rect 5088 21188 5092 21244
rect 5092 21188 5148 21244
rect 5148 21188 5152 21244
rect 5088 21184 5152 21188
rect 7445 21244 7509 21248
rect 7445 21188 7449 21244
rect 7449 21188 7505 21244
rect 7505 21188 7509 21244
rect 7445 21184 7509 21188
rect 7525 21244 7589 21248
rect 7525 21188 7529 21244
rect 7529 21188 7585 21244
rect 7585 21188 7589 21244
rect 7525 21184 7589 21188
rect 7605 21244 7669 21248
rect 7605 21188 7609 21244
rect 7609 21188 7665 21244
rect 7665 21188 7669 21244
rect 7605 21184 7669 21188
rect 7685 21244 7749 21248
rect 7685 21188 7689 21244
rect 7689 21188 7745 21244
rect 7745 21188 7749 21244
rect 7685 21184 7749 21188
rect 3549 20700 3613 20704
rect 3549 20644 3553 20700
rect 3553 20644 3609 20700
rect 3609 20644 3613 20700
rect 3549 20640 3613 20644
rect 3629 20700 3693 20704
rect 3629 20644 3633 20700
rect 3633 20644 3689 20700
rect 3689 20644 3693 20700
rect 3629 20640 3693 20644
rect 3709 20700 3773 20704
rect 3709 20644 3713 20700
rect 3713 20644 3769 20700
rect 3769 20644 3773 20700
rect 3709 20640 3773 20644
rect 3789 20700 3853 20704
rect 3789 20644 3793 20700
rect 3793 20644 3849 20700
rect 3849 20644 3853 20700
rect 3789 20640 3853 20644
rect 6146 20700 6210 20704
rect 6146 20644 6150 20700
rect 6150 20644 6206 20700
rect 6206 20644 6210 20700
rect 6146 20640 6210 20644
rect 6226 20700 6290 20704
rect 6226 20644 6230 20700
rect 6230 20644 6286 20700
rect 6286 20644 6290 20700
rect 6226 20640 6290 20644
rect 6306 20700 6370 20704
rect 6306 20644 6310 20700
rect 6310 20644 6366 20700
rect 6366 20644 6370 20700
rect 6306 20640 6370 20644
rect 6386 20700 6450 20704
rect 6386 20644 6390 20700
rect 6390 20644 6446 20700
rect 6446 20644 6450 20700
rect 6386 20640 6450 20644
rect 2250 20156 2314 20160
rect 2250 20100 2254 20156
rect 2254 20100 2310 20156
rect 2310 20100 2314 20156
rect 2250 20096 2314 20100
rect 2330 20156 2394 20160
rect 2330 20100 2334 20156
rect 2334 20100 2390 20156
rect 2390 20100 2394 20156
rect 2330 20096 2394 20100
rect 2410 20156 2474 20160
rect 2410 20100 2414 20156
rect 2414 20100 2470 20156
rect 2470 20100 2474 20156
rect 2410 20096 2474 20100
rect 2490 20156 2554 20160
rect 2490 20100 2494 20156
rect 2494 20100 2550 20156
rect 2550 20100 2554 20156
rect 2490 20096 2554 20100
rect 4848 20156 4912 20160
rect 4848 20100 4852 20156
rect 4852 20100 4908 20156
rect 4908 20100 4912 20156
rect 4848 20096 4912 20100
rect 4928 20156 4992 20160
rect 4928 20100 4932 20156
rect 4932 20100 4988 20156
rect 4988 20100 4992 20156
rect 4928 20096 4992 20100
rect 5008 20156 5072 20160
rect 5008 20100 5012 20156
rect 5012 20100 5068 20156
rect 5068 20100 5072 20156
rect 5008 20096 5072 20100
rect 5088 20156 5152 20160
rect 5088 20100 5092 20156
rect 5092 20100 5148 20156
rect 5148 20100 5152 20156
rect 5088 20096 5152 20100
rect 7445 20156 7509 20160
rect 7445 20100 7449 20156
rect 7449 20100 7505 20156
rect 7505 20100 7509 20156
rect 7445 20096 7509 20100
rect 7525 20156 7589 20160
rect 7525 20100 7529 20156
rect 7529 20100 7585 20156
rect 7585 20100 7589 20156
rect 7525 20096 7589 20100
rect 7605 20156 7669 20160
rect 7605 20100 7609 20156
rect 7609 20100 7665 20156
rect 7665 20100 7669 20156
rect 7605 20096 7669 20100
rect 7685 20156 7749 20160
rect 7685 20100 7689 20156
rect 7689 20100 7745 20156
rect 7745 20100 7749 20156
rect 7685 20096 7749 20100
rect 3549 19612 3613 19616
rect 3549 19556 3553 19612
rect 3553 19556 3609 19612
rect 3609 19556 3613 19612
rect 3549 19552 3613 19556
rect 3629 19612 3693 19616
rect 3629 19556 3633 19612
rect 3633 19556 3689 19612
rect 3689 19556 3693 19612
rect 3629 19552 3693 19556
rect 3709 19612 3773 19616
rect 3709 19556 3713 19612
rect 3713 19556 3769 19612
rect 3769 19556 3773 19612
rect 3709 19552 3773 19556
rect 3789 19612 3853 19616
rect 3789 19556 3793 19612
rect 3793 19556 3849 19612
rect 3849 19556 3853 19612
rect 3789 19552 3853 19556
rect 6146 19612 6210 19616
rect 6146 19556 6150 19612
rect 6150 19556 6206 19612
rect 6206 19556 6210 19612
rect 6146 19552 6210 19556
rect 6226 19612 6290 19616
rect 6226 19556 6230 19612
rect 6230 19556 6286 19612
rect 6286 19556 6290 19612
rect 6226 19552 6290 19556
rect 6306 19612 6370 19616
rect 6306 19556 6310 19612
rect 6310 19556 6366 19612
rect 6366 19556 6370 19612
rect 6306 19552 6370 19556
rect 6386 19612 6450 19616
rect 6386 19556 6390 19612
rect 6390 19556 6446 19612
rect 6446 19556 6450 19612
rect 6386 19552 6450 19556
rect 2250 19068 2314 19072
rect 2250 19012 2254 19068
rect 2254 19012 2310 19068
rect 2310 19012 2314 19068
rect 2250 19008 2314 19012
rect 2330 19068 2394 19072
rect 2330 19012 2334 19068
rect 2334 19012 2390 19068
rect 2390 19012 2394 19068
rect 2330 19008 2394 19012
rect 2410 19068 2474 19072
rect 2410 19012 2414 19068
rect 2414 19012 2470 19068
rect 2470 19012 2474 19068
rect 2410 19008 2474 19012
rect 2490 19068 2554 19072
rect 2490 19012 2494 19068
rect 2494 19012 2550 19068
rect 2550 19012 2554 19068
rect 2490 19008 2554 19012
rect 4848 19068 4912 19072
rect 4848 19012 4852 19068
rect 4852 19012 4908 19068
rect 4908 19012 4912 19068
rect 4848 19008 4912 19012
rect 4928 19068 4992 19072
rect 4928 19012 4932 19068
rect 4932 19012 4988 19068
rect 4988 19012 4992 19068
rect 4928 19008 4992 19012
rect 5008 19068 5072 19072
rect 5008 19012 5012 19068
rect 5012 19012 5068 19068
rect 5068 19012 5072 19068
rect 5008 19008 5072 19012
rect 5088 19068 5152 19072
rect 5088 19012 5092 19068
rect 5092 19012 5148 19068
rect 5148 19012 5152 19068
rect 5088 19008 5152 19012
rect 7445 19068 7509 19072
rect 7445 19012 7449 19068
rect 7449 19012 7505 19068
rect 7505 19012 7509 19068
rect 7445 19008 7509 19012
rect 7525 19068 7589 19072
rect 7525 19012 7529 19068
rect 7529 19012 7585 19068
rect 7585 19012 7589 19068
rect 7525 19008 7589 19012
rect 7605 19068 7669 19072
rect 7605 19012 7609 19068
rect 7609 19012 7665 19068
rect 7665 19012 7669 19068
rect 7605 19008 7669 19012
rect 7685 19068 7749 19072
rect 7685 19012 7689 19068
rect 7689 19012 7745 19068
rect 7745 19012 7749 19068
rect 7685 19008 7749 19012
rect 3549 18524 3613 18528
rect 3549 18468 3553 18524
rect 3553 18468 3609 18524
rect 3609 18468 3613 18524
rect 3549 18464 3613 18468
rect 3629 18524 3693 18528
rect 3629 18468 3633 18524
rect 3633 18468 3689 18524
rect 3689 18468 3693 18524
rect 3629 18464 3693 18468
rect 3709 18524 3773 18528
rect 3709 18468 3713 18524
rect 3713 18468 3769 18524
rect 3769 18468 3773 18524
rect 3709 18464 3773 18468
rect 3789 18524 3853 18528
rect 3789 18468 3793 18524
rect 3793 18468 3849 18524
rect 3849 18468 3853 18524
rect 3789 18464 3853 18468
rect 6146 18524 6210 18528
rect 6146 18468 6150 18524
rect 6150 18468 6206 18524
rect 6206 18468 6210 18524
rect 6146 18464 6210 18468
rect 6226 18524 6290 18528
rect 6226 18468 6230 18524
rect 6230 18468 6286 18524
rect 6286 18468 6290 18524
rect 6226 18464 6290 18468
rect 6306 18524 6370 18528
rect 6306 18468 6310 18524
rect 6310 18468 6366 18524
rect 6366 18468 6370 18524
rect 6306 18464 6370 18468
rect 6386 18524 6450 18528
rect 6386 18468 6390 18524
rect 6390 18468 6446 18524
rect 6446 18468 6450 18524
rect 6386 18464 6450 18468
rect 2250 17980 2314 17984
rect 2250 17924 2254 17980
rect 2254 17924 2310 17980
rect 2310 17924 2314 17980
rect 2250 17920 2314 17924
rect 2330 17980 2394 17984
rect 2330 17924 2334 17980
rect 2334 17924 2390 17980
rect 2390 17924 2394 17980
rect 2330 17920 2394 17924
rect 2410 17980 2474 17984
rect 2410 17924 2414 17980
rect 2414 17924 2470 17980
rect 2470 17924 2474 17980
rect 2410 17920 2474 17924
rect 2490 17980 2554 17984
rect 2490 17924 2494 17980
rect 2494 17924 2550 17980
rect 2550 17924 2554 17980
rect 2490 17920 2554 17924
rect 4848 17980 4912 17984
rect 4848 17924 4852 17980
rect 4852 17924 4908 17980
rect 4908 17924 4912 17980
rect 4848 17920 4912 17924
rect 4928 17980 4992 17984
rect 4928 17924 4932 17980
rect 4932 17924 4988 17980
rect 4988 17924 4992 17980
rect 4928 17920 4992 17924
rect 5008 17980 5072 17984
rect 5008 17924 5012 17980
rect 5012 17924 5068 17980
rect 5068 17924 5072 17980
rect 5008 17920 5072 17924
rect 5088 17980 5152 17984
rect 5088 17924 5092 17980
rect 5092 17924 5148 17980
rect 5148 17924 5152 17980
rect 5088 17920 5152 17924
rect 7445 17980 7509 17984
rect 7445 17924 7449 17980
rect 7449 17924 7505 17980
rect 7505 17924 7509 17980
rect 7445 17920 7509 17924
rect 7525 17980 7589 17984
rect 7525 17924 7529 17980
rect 7529 17924 7585 17980
rect 7585 17924 7589 17980
rect 7525 17920 7589 17924
rect 7605 17980 7669 17984
rect 7605 17924 7609 17980
rect 7609 17924 7665 17980
rect 7665 17924 7669 17980
rect 7605 17920 7669 17924
rect 7685 17980 7749 17984
rect 7685 17924 7689 17980
rect 7689 17924 7745 17980
rect 7745 17924 7749 17980
rect 7685 17920 7749 17924
rect 5948 17912 6012 17916
rect 5948 17856 5998 17912
rect 5998 17856 6012 17912
rect 5948 17852 6012 17856
rect 3549 17436 3613 17440
rect 3549 17380 3553 17436
rect 3553 17380 3609 17436
rect 3609 17380 3613 17436
rect 3549 17376 3613 17380
rect 3629 17436 3693 17440
rect 3629 17380 3633 17436
rect 3633 17380 3689 17436
rect 3689 17380 3693 17436
rect 3629 17376 3693 17380
rect 3709 17436 3773 17440
rect 3709 17380 3713 17436
rect 3713 17380 3769 17436
rect 3769 17380 3773 17436
rect 3709 17376 3773 17380
rect 3789 17436 3853 17440
rect 3789 17380 3793 17436
rect 3793 17380 3849 17436
rect 3849 17380 3853 17436
rect 3789 17376 3853 17380
rect 6146 17436 6210 17440
rect 6146 17380 6150 17436
rect 6150 17380 6206 17436
rect 6206 17380 6210 17436
rect 6146 17376 6210 17380
rect 6226 17436 6290 17440
rect 6226 17380 6230 17436
rect 6230 17380 6286 17436
rect 6286 17380 6290 17436
rect 6226 17376 6290 17380
rect 6306 17436 6370 17440
rect 6306 17380 6310 17436
rect 6310 17380 6366 17436
rect 6366 17380 6370 17436
rect 6306 17376 6370 17380
rect 6386 17436 6450 17440
rect 6386 17380 6390 17436
rect 6390 17380 6446 17436
rect 6446 17380 6450 17436
rect 6386 17376 6450 17380
rect 2250 16892 2314 16896
rect 2250 16836 2254 16892
rect 2254 16836 2310 16892
rect 2310 16836 2314 16892
rect 2250 16832 2314 16836
rect 2330 16892 2394 16896
rect 2330 16836 2334 16892
rect 2334 16836 2390 16892
rect 2390 16836 2394 16892
rect 2330 16832 2394 16836
rect 2410 16892 2474 16896
rect 2410 16836 2414 16892
rect 2414 16836 2470 16892
rect 2470 16836 2474 16892
rect 2410 16832 2474 16836
rect 2490 16892 2554 16896
rect 2490 16836 2494 16892
rect 2494 16836 2550 16892
rect 2550 16836 2554 16892
rect 2490 16832 2554 16836
rect 4848 16892 4912 16896
rect 4848 16836 4852 16892
rect 4852 16836 4908 16892
rect 4908 16836 4912 16892
rect 4848 16832 4912 16836
rect 4928 16892 4992 16896
rect 4928 16836 4932 16892
rect 4932 16836 4988 16892
rect 4988 16836 4992 16892
rect 4928 16832 4992 16836
rect 5008 16892 5072 16896
rect 5008 16836 5012 16892
rect 5012 16836 5068 16892
rect 5068 16836 5072 16892
rect 5008 16832 5072 16836
rect 5088 16892 5152 16896
rect 5088 16836 5092 16892
rect 5092 16836 5148 16892
rect 5148 16836 5152 16892
rect 5088 16832 5152 16836
rect 7445 16892 7509 16896
rect 7445 16836 7449 16892
rect 7449 16836 7505 16892
rect 7505 16836 7509 16892
rect 7445 16832 7509 16836
rect 7525 16892 7589 16896
rect 7525 16836 7529 16892
rect 7529 16836 7585 16892
rect 7585 16836 7589 16892
rect 7525 16832 7589 16836
rect 7605 16892 7669 16896
rect 7605 16836 7609 16892
rect 7609 16836 7665 16892
rect 7665 16836 7669 16892
rect 7605 16832 7669 16836
rect 7685 16892 7749 16896
rect 7685 16836 7689 16892
rect 7689 16836 7745 16892
rect 7745 16836 7749 16892
rect 7685 16832 7749 16836
rect 3549 16348 3613 16352
rect 3549 16292 3553 16348
rect 3553 16292 3609 16348
rect 3609 16292 3613 16348
rect 3549 16288 3613 16292
rect 3629 16348 3693 16352
rect 3629 16292 3633 16348
rect 3633 16292 3689 16348
rect 3689 16292 3693 16348
rect 3629 16288 3693 16292
rect 3709 16348 3773 16352
rect 3709 16292 3713 16348
rect 3713 16292 3769 16348
rect 3769 16292 3773 16348
rect 3709 16288 3773 16292
rect 3789 16348 3853 16352
rect 3789 16292 3793 16348
rect 3793 16292 3849 16348
rect 3849 16292 3853 16348
rect 3789 16288 3853 16292
rect 6146 16348 6210 16352
rect 6146 16292 6150 16348
rect 6150 16292 6206 16348
rect 6206 16292 6210 16348
rect 6146 16288 6210 16292
rect 6226 16348 6290 16352
rect 6226 16292 6230 16348
rect 6230 16292 6286 16348
rect 6286 16292 6290 16348
rect 6226 16288 6290 16292
rect 6306 16348 6370 16352
rect 6306 16292 6310 16348
rect 6310 16292 6366 16348
rect 6366 16292 6370 16348
rect 6306 16288 6370 16292
rect 6386 16348 6450 16352
rect 6386 16292 6390 16348
rect 6390 16292 6446 16348
rect 6446 16292 6450 16348
rect 6386 16288 6450 16292
rect 2250 15804 2314 15808
rect 2250 15748 2254 15804
rect 2254 15748 2310 15804
rect 2310 15748 2314 15804
rect 2250 15744 2314 15748
rect 2330 15804 2394 15808
rect 2330 15748 2334 15804
rect 2334 15748 2390 15804
rect 2390 15748 2394 15804
rect 2330 15744 2394 15748
rect 2410 15804 2474 15808
rect 2410 15748 2414 15804
rect 2414 15748 2470 15804
rect 2470 15748 2474 15804
rect 2410 15744 2474 15748
rect 2490 15804 2554 15808
rect 2490 15748 2494 15804
rect 2494 15748 2550 15804
rect 2550 15748 2554 15804
rect 2490 15744 2554 15748
rect 4848 15804 4912 15808
rect 4848 15748 4852 15804
rect 4852 15748 4908 15804
rect 4908 15748 4912 15804
rect 4848 15744 4912 15748
rect 4928 15804 4992 15808
rect 4928 15748 4932 15804
rect 4932 15748 4988 15804
rect 4988 15748 4992 15804
rect 4928 15744 4992 15748
rect 5008 15804 5072 15808
rect 5008 15748 5012 15804
rect 5012 15748 5068 15804
rect 5068 15748 5072 15804
rect 5008 15744 5072 15748
rect 5088 15804 5152 15808
rect 5088 15748 5092 15804
rect 5092 15748 5148 15804
rect 5148 15748 5152 15804
rect 5088 15744 5152 15748
rect 7445 15804 7509 15808
rect 7445 15748 7449 15804
rect 7449 15748 7505 15804
rect 7505 15748 7509 15804
rect 7445 15744 7509 15748
rect 7525 15804 7589 15808
rect 7525 15748 7529 15804
rect 7529 15748 7585 15804
rect 7585 15748 7589 15804
rect 7525 15744 7589 15748
rect 7605 15804 7669 15808
rect 7605 15748 7609 15804
rect 7609 15748 7665 15804
rect 7665 15748 7669 15804
rect 7605 15744 7669 15748
rect 7685 15804 7749 15808
rect 7685 15748 7689 15804
rect 7689 15748 7745 15804
rect 7745 15748 7749 15804
rect 7685 15744 7749 15748
rect 3549 15260 3613 15264
rect 3549 15204 3553 15260
rect 3553 15204 3609 15260
rect 3609 15204 3613 15260
rect 3549 15200 3613 15204
rect 3629 15260 3693 15264
rect 3629 15204 3633 15260
rect 3633 15204 3689 15260
rect 3689 15204 3693 15260
rect 3629 15200 3693 15204
rect 3709 15260 3773 15264
rect 3709 15204 3713 15260
rect 3713 15204 3769 15260
rect 3769 15204 3773 15260
rect 3709 15200 3773 15204
rect 3789 15260 3853 15264
rect 3789 15204 3793 15260
rect 3793 15204 3849 15260
rect 3849 15204 3853 15260
rect 3789 15200 3853 15204
rect 6146 15260 6210 15264
rect 6146 15204 6150 15260
rect 6150 15204 6206 15260
rect 6206 15204 6210 15260
rect 6146 15200 6210 15204
rect 6226 15260 6290 15264
rect 6226 15204 6230 15260
rect 6230 15204 6286 15260
rect 6286 15204 6290 15260
rect 6226 15200 6290 15204
rect 6306 15260 6370 15264
rect 6306 15204 6310 15260
rect 6310 15204 6366 15260
rect 6366 15204 6370 15260
rect 6306 15200 6370 15204
rect 6386 15260 6450 15264
rect 6386 15204 6390 15260
rect 6390 15204 6446 15260
rect 6446 15204 6450 15260
rect 6386 15200 6450 15204
rect 2250 14716 2314 14720
rect 2250 14660 2254 14716
rect 2254 14660 2310 14716
rect 2310 14660 2314 14716
rect 2250 14656 2314 14660
rect 2330 14716 2394 14720
rect 2330 14660 2334 14716
rect 2334 14660 2390 14716
rect 2390 14660 2394 14716
rect 2330 14656 2394 14660
rect 2410 14716 2474 14720
rect 2410 14660 2414 14716
rect 2414 14660 2470 14716
rect 2470 14660 2474 14716
rect 2410 14656 2474 14660
rect 2490 14716 2554 14720
rect 2490 14660 2494 14716
rect 2494 14660 2550 14716
rect 2550 14660 2554 14716
rect 2490 14656 2554 14660
rect 4848 14716 4912 14720
rect 4848 14660 4852 14716
rect 4852 14660 4908 14716
rect 4908 14660 4912 14716
rect 4848 14656 4912 14660
rect 4928 14716 4992 14720
rect 4928 14660 4932 14716
rect 4932 14660 4988 14716
rect 4988 14660 4992 14716
rect 4928 14656 4992 14660
rect 5008 14716 5072 14720
rect 5008 14660 5012 14716
rect 5012 14660 5068 14716
rect 5068 14660 5072 14716
rect 5008 14656 5072 14660
rect 5088 14716 5152 14720
rect 5088 14660 5092 14716
rect 5092 14660 5148 14716
rect 5148 14660 5152 14716
rect 5088 14656 5152 14660
rect 7445 14716 7509 14720
rect 7445 14660 7449 14716
rect 7449 14660 7505 14716
rect 7505 14660 7509 14716
rect 7445 14656 7509 14660
rect 7525 14716 7589 14720
rect 7525 14660 7529 14716
rect 7529 14660 7585 14716
rect 7585 14660 7589 14716
rect 7525 14656 7589 14660
rect 7605 14716 7669 14720
rect 7605 14660 7609 14716
rect 7609 14660 7665 14716
rect 7665 14660 7669 14716
rect 7605 14656 7669 14660
rect 7685 14716 7749 14720
rect 7685 14660 7689 14716
rect 7689 14660 7745 14716
rect 7745 14660 7749 14716
rect 7685 14656 7749 14660
rect 3549 14172 3613 14176
rect 3549 14116 3553 14172
rect 3553 14116 3609 14172
rect 3609 14116 3613 14172
rect 3549 14112 3613 14116
rect 3629 14172 3693 14176
rect 3629 14116 3633 14172
rect 3633 14116 3689 14172
rect 3689 14116 3693 14172
rect 3629 14112 3693 14116
rect 3709 14172 3773 14176
rect 3709 14116 3713 14172
rect 3713 14116 3769 14172
rect 3769 14116 3773 14172
rect 3709 14112 3773 14116
rect 3789 14172 3853 14176
rect 3789 14116 3793 14172
rect 3793 14116 3849 14172
rect 3849 14116 3853 14172
rect 3789 14112 3853 14116
rect 6146 14172 6210 14176
rect 6146 14116 6150 14172
rect 6150 14116 6206 14172
rect 6206 14116 6210 14172
rect 6146 14112 6210 14116
rect 6226 14172 6290 14176
rect 6226 14116 6230 14172
rect 6230 14116 6286 14172
rect 6286 14116 6290 14172
rect 6226 14112 6290 14116
rect 6306 14172 6370 14176
rect 6306 14116 6310 14172
rect 6310 14116 6366 14172
rect 6366 14116 6370 14172
rect 6306 14112 6370 14116
rect 6386 14172 6450 14176
rect 6386 14116 6390 14172
rect 6390 14116 6446 14172
rect 6446 14116 6450 14172
rect 6386 14112 6450 14116
rect 2250 13628 2314 13632
rect 2250 13572 2254 13628
rect 2254 13572 2310 13628
rect 2310 13572 2314 13628
rect 2250 13568 2314 13572
rect 2330 13628 2394 13632
rect 2330 13572 2334 13628
rect 2334 13572 2390 13628
rect 2390 13572 2394 13628
rect 2330 13568 2394 13572
rect 2410 13628 2474 13632
rect 2410 13572 2414 13628
rect 2414 13572 2470 13628
rect 2470 13572 2474 13628
rect 2410 13568 2474 13572
rect 2490 13628 2554 13632
rect 2490 13572 2494 13628
rect 2494 13572 2550 13628
rect 2550 13572 2554 13628
rect 2490 13568 2554 13572
rect 4848 13628 4912 13632
rect 4848 13572 4852 13628
rect 4852 13572 4908 13628
rect 4908 13572 4912 13628
rect 4848 13568 4912 13572
rect 4928 13628 4992 13632
rect 4928 13572 4932 13628
rect 4932 13572 4988 13628
rect 4988 13572 4992 13628
rect 4928 13568 4992 13572
rect 5008 13628 5072 13632
rect 5008 13572 5012 13628
rect 5012 13572 5068 13628
rect 5068 13572 5072 13628
rect 5008 13568 5072 13572
rect 5088 13628 5152 13632
rect 5088 13572 5092 13628
rect 5092 13572 5148 13628
rect 5148 13572 5152 13628
rect 5088 13568 5152 13572
rect 7445 13628 7509 13632
rect 7445 13572 7449 13628
rect 7449 13572 7505 13628
rect 7505 13572 7509 13628
rect 7445 13568 7509 13572
rect 7525 13628 7589 13632
rect 7525 13572 7529 13628
rect 7529 13572 7585 13628
rect 7585 13572 7589 13628
rect 7525 13568 7589 13572
rect 7605 13628 7669 13632
rect 7605 13572 7609 13628
rect 7609 13572 7665 13628
rect 7665 13572 7669 13628
rect 7605 13568 7669 13572
rect 7685 13628 7749 13632
rect 7685 13572 7689 13628
rect 7689 13572 7745 13628
rect 7745 13572 7749 13628
rect 7685 13568 7749 13572
rect 3549 13084 3613 13088
rect 3549 13028 3553 13084
rect 3553 13028 3609 13084
rect 3609 13028 3613 13084
rect 3549 13024 3613 13028
rect 3629 13084 3693 13088
rect 3629 13028 3633 13084
rect 3633 13028 3689 13084
rect 3689 13028 3693 13084
rect 3629 13024 3693 13028
rect 3709 13084 3773 13088
rect 3709 13028 3713 13084
rect 3713 13028 3769 13084
rect 3769 13028 3773 13084
rect 3709 13024 3773 13028
rect 3789 13084 3853 13088
rect 3789 13028 3793 13084
rect 3793 13028 3849 13084
rect 3849 13028 3853 13084
rect 3789 13024 3853 13028
rect 6146 13084 6210 13088
rect 6146 13028 6150 13084
rect 6150 13028 6206 13084
rect 6206 13028 6210 13084
rect 6146 13024 6210 13028
rect 6226 13084 6290 13088
rect 6226 13028 6230 13084
rect 6230 13028 6286 13084
rect 6286 13028 6290 13084
rect 6226 13024 6290 13028
rect 6306 13084 6370 13088
rect 6306 13028 6310 13084
rect 6310 13028 6366 13084
rect 6366 13028 6370 13084
rect 6306 13024 6370 13028
rect 6386 13084 6450 13088
rect 6386 13028 6390 13084
rect 6390 13028 6446 13084
rect 6446 13028 6450 13084
rect 6386 13024 6450 13028
rect 5948 12744 6012 12748
rect 5948 12688 5998 12744
rect 5998 12688 6012 12744
rect 5948 12684 6012 12688
rect 2250 12540 2314 12544
rect 2250 12484 2254 12540
rect 2254 12484 2310 12540
rect 2310 12484 2314 12540
rect 2250 12480 2314 12484
rect 2330 12540 2394 12544
rect 2330 12484 2334 12540
rect 2334 12484 2390 12540
rect 2390 12484 2394 12540
rect 2330 12480 2394 12484
rect 2410 12540 2474 12544
rect 2410 12484 2414 12540
rect 2414 12484 2470 12540
rect 2470 12484 2474 12540
rect 2410 12480 2474 12484
rect 2490 12540 2554 12544
rect 2490 12484 2494 12540
rect 2494 12484 2550 12540
rect 2550 12484 2554 12540
rect 2490 12480 2554 12484
rect 4848 12540 4912 12544
rect 4848 12484 4852 12540
rect 4852 12484 4908 12540
rect 4908 12484 4912 12540
rect 4848 12480 4912 12484
rect 4928 12540 4992 12544
rect 4928 12484 4932 12540
rect 4932 12484 4988 12540
rect 4988 12484 4992 12540
rect 4928 12480 4992 12484
rect 5008 12540 5072 12544
rect 5008 12484 5012 12540
rect 5012 12484 5068 12540
rect 5068 12484 5072 12540
rect 5008 12480 5072 12484
rect 5088 12540 5152 12544
rect 5088 12484 5092 12540
rect 5092 12484 5148 12540
rect 5148 12484 5152 12540
rect 5088 12480 5152 12484
rect 7445 12540 7509 12544
rect 7445 12484 7449 12540
rect 7449 12484 7505 12540
rect 7505 12484 7509 12540
rect 7445 12480 7509 12484
rect 7525 12540 7589 12544
rect 7525 12484 7529 12540
rect 7529 12484 7585 12540
rect 7585 12484 7589 12540
rect 7525 12480 7589 12484
rect 7605 12540 7669 12544
rect 7605 12484 7609 12540
rect 7609 12484 7665 12540
rect 7665 12484 7669 12540
rect 7605 12480 7669 12484
rect 7685 12540 7749 12544
rect 7685 12484 7689 12540
rect 7689 12484 7745 12540
rect 7745 12484 7749 12540
rect 7685 12480 7749 12484
rect 3549 11996 3613 12000
rect 3549 11940 3553 11996
rect 3553 11940 3609 11996
rect 3609 11940 3613 11996
rect 3549 11936 3613 11940
rect 3629 11996 3693 12000
rect 3629 11940 3633 11996
rect 3633 11940 3689 11996
rect 3689 11940 3693 11996
rect 3629 11936 3693 11940
rect 3709 11996 3773 12000
rect 3709 11940 3713 11996
rect 3713 11940 3769 11996
rect 3769 11940 3773 11996
rect 3709 11936 3773 11940
rect 3789 11996 3853 12000
rect 3789 11940 3793 11996
rect 3793 11940 3849 11996
rect 3849 11940 3853 11996
rect 3789 11936 3853 11940
rect 6146 11996 6210 12000
rect 6146 11940 6150 11996
rect 6150 11940 6206 11996
rect 6206 11940 6210 11996
rect 6146 11936 6210 11940
rect 6226 11996 6290 12000
rect 6226 11940 6230 11996
rect 6230 11940 6286 11996
rect 6286 11940 6290 11996
rect 6226 11936 6290 11940
rect 6306 11996 6370 12000
rect 6306 11940 6310 11996
rect 6310 11940 6366 11996
rect 6366 11940 6370 11996
rect 6306 11936 6370 11940
rect 6386 11996 6450 12000
rect 6386 11940 6390 11996
rect 6390 11940 6446 11996
rect 6446 11940 6450 11996
rect 6386 11936 6450 11940
rect 2250 11452 2314 11456
rect 2250 11396 2254 11452
rect 2254 11396 2310 11452
rect 2310 11396 2314 11452
rect 2250 11392 2314 11396
rect 2330 11452 2394 11456
rect 2330 11396 2334 11452
rect 2334 11396 2390 11452
rect 2390 11396 2394 11452
rect 2330 11392 2394 11396
rect 2410 11452 2474 11456
rect 2410 11396 2414 11452
rect 2414 11396 2470 11452
rect 2470 11396 2474 11452
rect 2410 11392 2474 11396
rect 2490 11452 2554 11456
rect 2490 11396 2494 11452
rect 2494 11396 2550 11452
rect 2550 11396 2554 11452
rect 2490 11392 2554 11396
rect 4848 11452 4912 11456
rect 4848 11396 4852 11452
rect 4852 11396 4908 11452
rect 4908 11396 4912 11452
rect 4848 11392 4912 11396
rect 4928 11452 4992 11456
rect 4928 11396 4932 11452
rect 4932 11396 4988 11452
rect 4988 11396 4992 11452
rect 4928 11392 4992 11396
rect 5008 11452 5072 11456
rect 5008 11396 5012 11452
rect 5012 11396 5068 11452
rect 5068 11396 5072 11452
rect 5008 11392 5072 11396
rect 5088 11452 5152 11456
rect 5088 11396 5092 11452
rect 5092 11396 5148 11452
rect 5148 11396 5152 11452
rect 5088 11392 5152 11396
rect 7445 11452 7509 11456
rect 7445 11396 7449 11452
rect 7449 11396 7505 11452
rect 7505 11396 7509 11452
rect 7445 11392 7509 11396
rect 7525 11452 7589 11456
rect 7525 11396 7529 11452
rect 7529 11396 7585 11452
rect 7585 11396 7589 11452
rect 7525 11392 7589 11396
rect 7605 11452 7669 11456
rect 7605 11396 7609 11452
rect 7609 11396 7665 11452
rect 7665 11396 7669 11452
rect 7605 11392 7669 11396
rect 7685 11452 7749 11456
rect 7685 11396 7689 11452
rect 7689 11396 7745 11452
rect 7745 11396 7749 11452
rect 7685 11392 7749 11396
rect 3549 10908 3613 10912
rect 3549 10852 3553 10908
rect 3553 10852 3609 10908
rect 3609 10852 3613 10908
rect 3549 10848 3613 10852
rect 3629 10908 3693 10912
rect 3629 10852 3633 10908
rect 3633 10852 3689 10908
rect 3689 10852 3693 10908
rect 3629 10848 3693 10852
rect 3709 10908 3773 10912
rect 3709 10852 3713 10908
rect 3713 10852 3769 10908
rect 3769 10852 3773 10908
rect 3709 10848 3773 10852
rect 3789 10908 3853 10912
rect 3789 10852 3793 10908
rect 3793 10852 3849 10908
rect 3849 10852 3853 10908
rect 3789 10848 3853 10852
rect 6146 10908 6210 10912
rect 6146 10852 6150 10908
rect 6150 10852 6206 10908
rect 6206 10852 6210 10908
rect 6146 10848 6210 10852
rect 6226 10908 6290 10912
rect 6226 10852 6230 10908
rect 6230 10852 6286 10908
rect 6286 10852 6290 10908
rect 6226 10848 6290 10852
rect 6306 10908 6370 10912
rect 6306 10852 6310 10908
rect 6310 10852 6366 10908
rect 6366 10852 6370 10908
rect 6306 10848 6370 10852
rect 6386 10908 6450 10912
rect 6386 10852 6390 10908
rect 6390 10852 6446 10908
rect 6446 10852 6450 10908
rect 6386 10848 6450 10852
rect 2250 10364 2314 10368
rect 2250 10308 2254 10364
rect 2254 10308 2310 10364
rect 2310 10308 2314 10364
rect 2250 10304 2314 10308
rect 2330 10364 2394 10368
rect 2330 10308 2334 10364
rect 2334 10308 2390 10364
rect 2390 10308 2394 10364
rect 2330 10304 2394 10308
rect 2410 10364 2474 10368
rect 2410 10308 2414 10364
rect 2414 10308 2470 10364
rect 2470 10308 2474 10364
rect 2410 10304 2474 10308
rect 2490 10364 2554 10368
rect 2490 10308 2494 10364
rect 2494 10308 2550 10364
rect 2550 10308 2554 10364
rect 2490 10304 2554 10308
rect 4848 10364 4912 10368
rect 4848 10308 4852 10364
rect 4852 10308 4908 10364
rect 4908 10308 4912 10364
rect 4848 10304 4912 10308
rect 4928 10364 4992 10368
rect 4928 10308 4932 10364
rect 4932 10308 4988 10364
rect 4988 10308 4992 10364
rect 4928 10304 4992 10308
rect 5008 10364 5072 10368
rect 5008 10308 5012 10364
rect 5012 10308 5068 10364
rect 5068 10308 5072 10364
rect 5008 10304 5072 10308
rect 5088 10364 5152 10368
rect 5088 10308 5092 10364
rect 5092 10308 5148 10364
rect 5148 10308 5152 10364
rect 5088 10304 5152 10308
rect 7445 10364 7509 10368
rect 7445 10308 7449 10364
rect 7449 10308 7505 10364
rect 7505 10308 7509 10364
rect 7445 10304 7509 10308
rect 7525 10364 7589 10368
rect 7525 10308 7529 10364
rect 7529 10308 7585 10364
rect 7585 10308 7589 10364
rect 7525 10304 7589 10308
rect 7605 10364 7669 10368
rect 7605 10308 7609 10364
rect 7609 10308 7665 10364
rect 7665 10308 7669 10364
rect 7605 10304 7669 10308
rect 7685 10364 7749 10368
rect 7685 10308 7689 10364
rect 7689 10308 7745 10364
rect 7745 10308 7749 10364
rect 7685 10304 7749 10308
rect 3549 9820 3613 9824
rect 3549 9764 3553 9820
rect 3553 9764 3609 9820
rect 3609 9764 3613 9820
rect 3549 9760 3613 9764
rect 3629 9820 3693 9824
rect 3629 9764 3633 9820
rect 3633 9764 3689 9820
rect 3689 9764 3693 9820
rect 3629 9760 3693 9764
rect 3709 9820 3773 9824
rect 3709 9764 3713 9820
rect 3713 9764 3769 9820
rect 3769 9764 3773 9820
rect 3709 9760 3773 9764
rect 3789 9820 3853 9824
rect 3789 9764 3793 9820
rect 3793 9764 3849 9820
rect 3849 9764 3853 9820
rect 3789 9760 3853 9764
rect 6146 9820 6210 9824
rect 6146 9764 6150 9820
rect 6150 9764 6206 9820
rect 6206 9764 6210 9820
rect 6146 9760 6210 9764
rect 6226 9820 6290 9824
rect 6226 9764 6230 9820
rect 6230 9764 6286 9820
rect 6286 9764 6290 9820
rect 6226 9760 6290 9764
rect 6306 9820 6370 9824
rect 6306 9764 6310 9820
rect 6310 9764 6366 9820
rect 6366 9764 6370 9820
rect 6306 9760 6370 9764
rect 6386 9820 6450 9824
rect 6386 9764 6390 9820
rect 6390 9764 6446 9820
rect 6446 9764 6450 9820
rect 6386 9760 6450 9764
rect 2250 9276 2314 9280
rect 2250 9220 2254 9276
rect 2254 9220 2310 9276
rect 2310 9220 2314 9276
rect 2250 9216 2314 9220
rect 2330 9276 2394 9280
rect 2330 9220 2334 9276
rect 2334 9220 2390 9276
rect 2390 9220 2394 9276
rect 2330 9216 2394 9220
rect 2410 9276 2474 9280
rect 2410 9220 2414 9276
rect 2414 9220 2470 9276
rect 2470 9220 2474 9276
rect 2410 9216 2474 9220
rect 2490 9276 2554 9280
rect 2490 9220 2494 9276
rect 2494 9220 2550 9276
rect 2550 9220 2554 9276
rect 2490 9216 2554 9220
rect 4848 9276 4912 9280
rect 4848 9220 4852 9276
rect 4852 9220 4908 9276
rect 4908 9220 4912 9276
rect 4848 9216 4912 9220
rect 4928 9276 4992 9280
rect 4928 9220 4932 9276
rect 4932 9220 4988 9276
rect 4988 9220 4992 9276
rect 4928 9216 4992 9220
rect 5008 9276 5072 9280
rect 5008 9220 5012 9276
rect 5012 9220 5068 9276
rect 5068 9220 5072 9276
rect 5008 9216 5072 9220
rect 5088 9276 5152 9280
rect 5088 9220 5092 9276
rect 5092 9220 5148 9276
rect 5148 9220 5152 9276
rect 5088 9216 5152 9220
rect 7445 9276 7509 9280
rect 7445 9220 7449 9276
rect 7449 9220 7505 9276
rect 7505 9220 7509 9276
rect 7445 9216 7509 9220
rect 7525 9276 7589 9280
rect 7525 9220 7529 9276
rect 7529 9220 7585 9276
rect 7585 9220 7589 9276
rect 7525 9216 7589 9220
rect 7605 9276 7669 9280
rect 7605 9220 7609 9276
rect 7609 9220 7665 9276
rect 7665 9220 7669 9276
rect 7605 9216 7669 9220
rect 7685 9276 7749 9280
rect 7685 9220 7689 9276
rect 7689 9220 7745 9276
rect 7745 9220 7749 9276
rect 7685 9216 7749 9220
rect 3549 8732 3613 8736
rect 3549 8676 3553 8732
rect 3553 8676 3609 8732
rect 3609 8676 3613 8732
rect 3549 8672 3613 8676
rect 3629 8732 3693 8736
rect 3629 8676 3633 8732
rect 3633 8676 3689 8732
rect 3689 8676 3693 8732
rect 3629 8672 3693 8676
rect 3709 8732 3773 8736
rect 3709 8676 3713 8732
rect 3713 8676 3769 8732
rect 3769 8676 3773 8732
rect 3709 8672 3773 8676
rect 3789 8732 3853 8736
rect 3789 8676 3793 8732
rect 3793 8676 3849 8732
rect 3849 8676 3853 8732
rect 3789 8672 3853 8676
rect 6146 8732 6210 8736
rect 6146 8676 6150 8732
rect 6150 8676 6206 8732
rect 6206 8676 6210 8732
rect 6146 8672 6210 8676
rect 6226 8732 6290 8736
rect 6226 8676 6230 8732
rect 6230 8676 6286 8732
rect 6286 8676 6290 8732
rect 6226 8672 6290 8676
rect 6306 8732 6370 8736
rect 6306 8676 6310 8732
rect 6310 8676 6366 8732
rect 6366 8676 6370 8732
rect 6306 8672 6370 8676
rect 6386 8732 6450 8736
rect 6386 8676 6390 8732
rect 6390 8676 6446 8732
rect 6446 8676 6450 8732
rect 6386 8672 6450 8676
rect 2250 8188 2314 8192
rect 2250 8132 2254 8188
rect 2254 8132 2310 8188
rect 2310 8132 2314 8188
rect 2250 8128 2314 8132
rect 2330 8188 2394 8192
rect 2330 8132 2334 8188
rect 2334 8132 2390 8188
rect 2390 8132 2394 8188
rect 2330 8128 2394 8132
rect 2410 8188 2474 8192
rect 2410 8132 2414 8188
rect 2414 8132 2470 8188
rect 2470 8132 2474 8188
rect 2410 8128 2474 8132
rect 2490 8188 2554 8192
rect 2490 8132 2494 8188
rect 2494 8132 2550 8188
rect 2550 8132 2554 8188
rect 2490 8128 2554 8132
rect 4848 8188 4912 8192
rect 4848 8132 4852 8188
rect 4852 8132 4908 8188
rect 4908 8132 4912 8188
rect 4848 8128 4912 8132
rect 4928 8188 4992 8192
rect 4928 8132 4932 8188
rect 4932 8132 4988 8188
rect 4988 8132 4992 8188
rect 4928 8128 4992 8132
rect 5008 8188 5072 8192
rect 5008 8132 5012 8188
rect 5012 8132 5068 8188
rect 5068 8132 5072 8188
rect 5008 8128 5072 8132
rect 5088 8188 5152 8192
rect 5088 8132 5092 8188
rect 5092 8132 5148 8188
rect 5148 8132 5152 8188
rect 5088 8128 5152 8132
rect 7445 8188 7509 8192
rect 7445 8132 7449 8188
rect 7449 8132 7505 8188
rect 7505 8132 7509 8188
rect 7445 8128 7509 8132
rect 7525 8188 7589 8192
rect 7525 8132 7529 8188
rect 7529 8132 7585 8188
rect 7585 8132 7589 8188
rect 7525 8128 7589 8132
rect 7605 8188 7669 8192
rect 7605 8132 7609 8188
rect 7609 8132 7665 8188
rect 7665 8132 7669 8188
rect 7605 8128 7669 8132
rect 7685 8188 7749 8192
rect 7685 8132 7689 8188
rect 7689 8132 7745 8188
rect 7745 8132 7749 8188
rect 7685 8128 7749 8132
rect 3549 7644 3613 7648
rect 3549 7588 3553 7644
rect 3553 7588 3609 7644
rect 3609 7588 3613 7644
rect 3549 7584 3613 7588
rect 3629 7644 3693 7648
rect 3629 7588 3633 7644
rect 3633 7588 3689 7644
rect 3689 7588 3693 7644
rect 3629 7584 3693 7588
rect 3709 7644 3773 7648
rect 3709 7588 3713 7644
rect 3713 7588 3769 7644
rect 3769 7588 3773 7644
rect 3709 7584 3773 7588
rect 3789 7644 3853 7648
rect 3789 7588 3793 7644
rect 3793 7588 3849 7644
rect 3849 7588 3853 7644
rect 3789 7584 3853 7588
rect 6146 7644 6210 7648
rect 6146 7588 6150 7644
rect 6150 7588 6206 7644
rect 6206 7588 6210 7644
rect 6146 7584 6210 7588
rect 6226 7644 6290 7648
rect 6226 7588 6230 7644
rect 6230 7588 6286 7644
rect 6286 7588 6290 7644
rect 6226 7584 6290 7588
rect 6306 7644 6370 7648
rect 6306 7588 6310 7644
rect 6310 7588 6366 7644
rect 6366 7588 6370 7644
rect 6306 7584 6370 7588
rect 6386 7644 6450 7648
rect 6386 7588 6390 7644
rect 6390 7588 6446 7644
rect 6446 7588 6450 7644
rect 6386 7584 6450 7588
rect 2250 7100 2314 7104
rect 2250 7044 2254 7100
rect 2254 7044 2310 7100
rect 2310 7044 2314 7100
rect 2250 7040 2314 7044
rect 2330 7100 2394 7104
rect 2330 7044 2334 7100
rect 2334 7044 2390 7100
rect 2390 7044 2394 7100
rect 2330 7040 2394 7044
rect 2410 7100 2474 7104
rect 2410 7044 2414 7100
rect 2414 7044 2470 7100
rect 2470 7044 2474 7100
rect 2410 7040 2474 7044
rect 2490 7100 2554 7104
rect 2490 7044 2494 7100
rect 2494 7044 2550 7100
rect 2550 7044 2554 7100
rect 2490 7040 2554 7044
rect 4848 7100 4912 7104
rect 4848 7044 4852 7100
rect 4852 7044 4908 7100
rect 4908 7044 4912 7100
rect 4848 7040 4912 7044
rect 4928 7100 4992 7104
rect 4928 7044 4932 7100
rect 4932 7044 4988 7100
rect 4988 7044 4992 7100
rect 4928 7040 4992 7044
rect 5008 7100 5072 7104
rect 5008 7044 5012 7100
rect 5012 7044 5068 7100
rect 5068 7044 5072 7100
rect 5008 7040 5072 7044
rect 5088 7100 5152 7104
rect 5088 7044 5092 7100
rect 5092 7044 5148 7100
rect 5148 7044 5152 7100
rect 5088 7040 5152 7044
rect 7445 7100 7509 7104
rect 7445 7044 7449 7100
rect 7449 7044 7505 7100
rect 7505 7044 7509 7100
rect 7445 7040 7509 7044
rect 7525 7100 7589 7104
rect 7525 7044 7529 7100
rect 7529 7044 7585 7100
rect 7585 7044 7589 7100
rect 7525 7040 7589 7044
rect 7605 7100 7669 7104
rect 7605 7044 7609 7100
rect 7609 7044 7665 7100
rect 7665 7044 7669 7100
rect 7605 7040 7669 7044
rect 7685 7100 7749 7104
rect 7685 7044 7689 7100
rect 7689 7044 7745 7100
rect 7745 7044 7749 7100
rect 7685 7040 7749 7044
rect 3549 6556 3613 6560
rect 3549 6500 3553 6556
rect 3553 6500 3609 6556
rect 3609 6500 3613 6556
rect 3549 6496 3613 6500
rect 3629 6556 3693 6560
rect 3629 6500 3633 6556
rect 3633 6500 3689 6556
rect 3689 6500 3693 6556
rect 3629 6496 3693 6500
rect 3709 6556 3773 6560
rect 3709 6500 3713 6556
rect 3713 6500 3769 6556
rect 3769 6500 3773 6556
rect 3709 6496 3773 6500
rect 3789 6556 3853 6560
rect 3789 6500 3793 6556
rect 3793 6500 3849 6556
rect 3849 6500 3853 6556
rect 3789 6496 3853 6500
rect 6146 6556 6210 6560
rect 6146 6500 6150 6556
rect 6150 6500 6206 6556
rect 6206 6500 6210 6556
rect 6146 6496 6210 6500
rect 6226 6556 6290 6560
rect 6226 6500 6230 6556
rect 6230 6500 6286 6556
rect 6286 6500 6290 6556
rect 6226 6496 6290 6500
rect 6306 6556 6370 6560
rect 6306 6500 6310 6556
rect 6310 6500 6366 6556
rect 6366 6500 6370 6556
rect 6306 6496 6370 6500
rect 6386 6556 6450 6560
rect 6386 6500 6390 6556
rect 6390 6500 6446 6556
rect 6446 6500 6450 6556
rect 6386 6496 6450 6500
rect 2250 6012 2314 6016
rect 2250 5956 2254 6012
rect 2254 5956 2310 6012
rect 2310 5956 2314 6012
rect 2250 5952 2314 5956
rect 2330 6012 2394 6016
rect 2330 5956 2334 6012
rect 2334 5956 2390 6012
rect 2390 5956 2394 6012
rect 2330 5952 2394 5956
rect 2410 6012 2474 6016
rect 2410 5956 2414 6012
rect 2414 5956 2470 6012
rect 2470 5956 2474 6012
rect 2410 5952 2474 5956
rect 2490 6012 2554 6016
rect 2490 5956 2494 6012
rect 2494 5956 2550 6012
rect 2550 5956 2554 6012
rect 2490 5952 2554 5956
rect 4848 6012 4912 6016
rect 4848 5956 4852 6012
rect 4852 5956 4908 6012
rect 4908 5956 4912 6012
rect 4848 5952 4912 5956
rect 4928 6012 4992 6016
rect 4928 5956 4932 6012
rect 4932 5956 4988 6012
rect 4988 5956 4992 6012
rect 4928 5952 4992 5956
rect 5008 6012 5072 6016
rect 5008 5956 5012 6012
rect 5012 5956 5068 6012
rect 5068 5956 5072 6012
rect 5008 5952 5072 5956
rect 5088 6012 5152 6016
rect 5088 5956 5092 6012
rect 5092 5956 5148 6012
rect 5148 5956 5152 6012
rect 5088 5952 5152 5956
rect 7445 6012 7509 6016
rect 7445 5956 7449 6012
rect 7449 5956 7505 6012
rect 7505 5956 7509 6012
rect 7445 5952 7509 5956
rect 7525 6012 7589 6016
rect 7525 5956 7529 6012
rect 7529 5956 7585 6012
rect 7585 5956 7589 6012
rect 7525 5952 7589 5956
rect 7605 6012 7669 6016
rect 7605 5956 7609 6012
rect 7609 5956 7665 6012
rect 7665 5956 7669 6012
rect 7605 5952 7669 5956
rect 7685 6012 7749 6016
rect 7685 5956 7689 6012
rect 7689 5956 7745 6012
rect 7745 5956 7749 6012
rect 7685 5952 7749 5956
rect 3549 5468 3613 5472
rect 3549 5412 3553 5468
rect 3553 5412 3609 5468
rect 3609 5412 3613 5468
rect 3549 5408 3613 5412
rect 3629 5468 3693 5472
rect 3629 5412 3633 5468
rect 3633 5412 3689 5468
rect 3689 5412 3693 5468
rect 3629 5408 3693 5412
rect 3709 5468 3773 5472
rect 3709 5412 3713 5468
rect 3713 5412 3769 5468
rect 3769 5412 3773 5468
rect 3709 5408 3773 5412
rect 3789 5468 3853 5472
rect 3789 5412 3793 5468
rect 3793 5412 3849 5468
rect 3849 5412 3853 5468
rect 3789 5408 3853 5412
rect 6146 5468 6210 5472
rect 6146 5412 6150 5468
rect 6150 5412 6206 5468
rect 6206 5412 6210 5468
rect 6146 5408 6210 5412
rect 6226 5468 6290 5472
rect 6226 5412 6230 5468
rect 6230 5412 6286 5468
rect 6286 5412 6290 5468
rect 6226 5408 6290 5412
rect 6306 5468 6370 5472
rect 6306 5412 6310 5468
rect 6310 5412 6366 5468
rect 6366 5412 6370 5468
rect 6306 5408 6370 5412
rect 6386 5468 6450 5472
rect 6386 5412 6390 5468
rect 6390 5412 6446 5468
rect 6446 5412 6450 5468
rect 6386 5408 6450 5412
rect 2250 4924 2314 4928
rect 2250 4868 2254 4924
rect 2254 4868 2310 4924
rect 2310 4868 2314 4924
rect 2250 4864 2314 4868
rect 2330 4924 2394 4928
rect 2330 4868 2334 4924
rect 2334 4868 2390 4924
rect 2390 4868 2394 4924
rect 2330 4864 2394 4868
rect 2410 4924 2474 4928
rect 2410 4868 2414 4924
rect 2414 4868 2470 4924
rect 2470 4868 2474 4924
rect 2410 4864 2474 4868
rect 2490 4924 2554 4928
rect 2490 4868 2494 4924
rect 2494 4868 2550 4924
rect 2550 4868 2554 4924
rect 2490 4864 2554 4868
rect 4848 4924 4912 4928
rect 4848 4868 4852 4924
rect 4852 4868 4908 4924
rect 4908 4868 4912 4924
rect 4848 4864 4912 4868
rect 4928 4924 4992 4928
rect 4928 4868 4932 4924
rect 4932 4868 4988 4924
rect 4988 4868 4992 4924
rect 4928 4864 4992 4868
rect 5008 4924 5072 4928
rect 5008 4868 5012 4924
rect 5012 4868 5068 4924
rect 5068 4868 5072 4924
rect 5008 4864 5072 4868
rect 5088 4924 5152 4928
rect 5088 4868 5092 4924
rect 5092 4868 5148 4924
rect 5148 4868 5152 4924
rect 5088 4864 5152 4868
rect 7445 4924 7509 4928
rect 7445 4868 7449 4924
rect 7449 4868 7505 4924
rect 7505 4868 7509 4924
rect 7445 4864 7509 4868
rect 7525 4924 7589 4928
rect 7525 4868 7529 4924
rect 7529 4868 7585 4924
rect 7585 4868 7589 4924
rect 7525 4864 7589 4868
rect 7605 4924 7669 4928
rect 7605 4868 7609 4924
rect 7609 4868 7665 4924
rect 7665 4868 7669 4924
rect 7605 4864 7669 4868
rect 7685 4924 7749 4928
rect 7685 4868 7689 4924
rect 7689 4868 7745 4924
rect 7745 4868 7749 4924
rect 7685 4864 7749 4868
rect 3549 4380 3613 4384
rect 3549 4324 3553 4380
rect 3553 4324 3609 4380
rect 3609 4324 3613 4380
rect 3549 4320 3613 4324
rect 3629 4380 3693 4384
rect 3629 4324 3633 4380
rect 3633 4324 3689 4380
rect 3689 4324 3693 4380
rect 3629 4320 3693 4324
rect 3709 4380 3773 4384
rect 3709 4324 3713 4380
rect 3713 4324 3769 4380
rect 3769 4324 3773 4380
rect 3709 4320 3773 4324
rect 3789 4380 3853 4384
rect 3789 4324 3793 4380
rect 3793 4324 3849 4380
rect 3849 4324 3853 4380
rect 3789 4320 3853 4324
rect 6146 4380 6210 4384
rect 6146 4324 6150 4380
rect 6150 4324 6206 4380
rect 6206 4324 6210 4380
rect 6146 4320 6210 4324
rect 6226 4380 6290 4384
rect 6226 4324 6230 4380
rect 6230 4324 6286 4380
rect 6286 4324 6290 4380
rect 6226 4320 6290 4324
rect 6306 4380 6370 4384
rect 6306 4324 6310 4380
rect 6310 4324 6366 4380
rect 6366 4324 6370 4380
rect 6306 4320 6370 4324
rect 6386 4380 6450 4384
rect 6386 4324 6390 4380
rect 6390 4324 6446 4380
rect 6446 4324 6450 4380
rect 6386 4320 6450 4324
rect 2250 3836 2314 3840
rect 2250 3780 2254 3836
rect 2254 3780 2310 3836
rect 2310 3780 2314 3836
rect 2250 3776 2314 3780
rect 2330 3836 2394 3840
rect 2330 3780 2334 3836
rect 2334 3780 2390 3836
rect 2390 3780 2394 3836
rect 2330 3776 2394 3780
rect 2410 3836 2474 3840
rect 2410 3780 2414 3836
rect 2414 3780 2470 3836
rect 2470 3780 2474 3836
rect 2410 3776 2474 3780
rect 2490 3836 2554 3840
rect 2490 3780 2494 3836
rect 2494 3780 2550 3836
rect 2550 3780 2554 3836
rect 2490 3776 2554 3780
rect 4848 3836 4912 3840
rect 4848 3780 4852 3836
rect 4852 3780 4908 3836
rect 4908 3780 4912 3836
rect 4848 3776 4912 3780
rect 4928 3836 4992 3840
rect 4928 3780 4932 3836
rect 4932 3780 4988 3836
rect 4988 3780 4992 3836
rect 4928 3776 4992 3780
rect 5008 3836 5072 3840
rect 5008 3780 5012 3836
rect 5012 3780 5068 3836
rect 5068 3780 5072 3836
rect 5008 3776 5072 3780
rect 5088 3836 5152 3840
rect 5088 3780 5092 3836
rect 5092 3780 5148 3836
rect 5148 3780 5152 3836
rect 5088 3776 5152 3780
rect 7445 3836 7509 3840
rect 7445 3780 7449 3836
rect 7449 3780 7505 3836
rect 7505 3780 7509 3836
rect 7445 3776 7509 3780
rect 7525 3836 7589 3840
rect 7525 3780 7529 3836
rect 7529 3780 7585 3836
rect 7585 3780 7589 3836
rect 7525 3776 7589 3780
rect 7605 3836 7669 3840
rect 7605 3780 7609 3836
rect 7609 3780 7665 3836
rect 7665 3780 7669 3836
rect 7605 3776 7669 3780
rect 7685 3836 7749 3840
rect 7685 3780 7689 3836
rect 7689 3780 7745 3836
rect 7745 3780 7749 3836
rect 7685 3776 7749 3780
rect 3549 3292 3613 3296
rect 3549 3236 3553 3292
rect 3553 3236 3609 3292
rect 3609 3236 3613 3292
rect 3549 3232 3613 3236
rect 3629 3292 3693 3296
rect 3629 3236 3633 3292
rect 3633 3236 3689 3292
rect 3689 3236 3693 3292
rect 3629 3232 3693 3236
rect 3709 3292 3773 3296
rect 3709 3236 3713 3292
rect 3713 3236 3769 3292
rect 3769 3236 3773 3292
rect 3709 3232 3773 3236
rect 3789 3292 3853 3296
rect 3789 3236 3793 3292
rect 3793 3236 3849 3292
rect 3849 3236 3853 3292
rect 3789 3232 3853 3236
rect 6146 3292 6210 3296
rect 6146 3236 6150 3292
rect 6150 3236 6206 3292
rect 6206 3236 6210 3292
rect 6146 3232 6210 3236
rect 6226 3292 6290 3296
rect 6226 3236 6230 3292
rect 6230 3236 6286 3292
rect 6286 3236 6290 3292
rect 6226 3232 6290 3236
rect 6306 3292 6370 3296
rect 6306 3236 6310 3292
rect 6310 3236 6366 3292
rect 6366 3236 6370 3292
rect 6306 3232 6370 3236
rect 6386 3292 6450 3296
rect 6386 3236 6390 3292
rect 6390 3236 6446 3292
rect 6446 3236 6450 3292
rect 6386 3232 6450 3236
rect 2250 2748 2314 2752
rect 2250 2692 2254 2748
rect 2254 2692 2310 2748
rect 2310 2692 2314 2748
rect 2250 2688 2314 2692
rect 2330 2748 2394 2752
rect 2330 2692 2334 2748
rect 2334 2692 2390 2748
rect 2390 2692 2394 2748
rect 2330 2688 2394 2692
rect 2410 2748 2474 2752
rect 2410 2692 2414 2748
rect 2414 2692 2470 2748
rect 2470 2692 2474 2748
rect 2410 2688 2474 2692
rect 2490 2748 2554 2752
rect 2490 2692 2494 2748
rect 2494 2692 2550 2748
rect 2550 2692 2554 2748
rect 2490 2688 2554 2692
rect 4848 2748 4912 2752
rect 4848 2692 4852 2748
rect 4852 2692 4908 2748
rect 4908 2692 4912 2748
rect 4848 2688 4912 2692
rect 4928 2748 4992 2752
rect 4928 2692 4932 2748
rect 4932 2692 4988 2748
rect 4988 2692 4992 2748
rect 4928 2688 4992 2692
rect 5008 2748 5072 2752
rect 5008 2692 5012 2748
rect 5012 2692 5068 2748
rect 5068 2692 5072 2748
rect 5008 2688 5072 2692
rect 5088 2748 5152 2752
rect 5088 2692 5092 2748
rect 5092 2692 5148 2748
rect 5148 2692 5152 2748
rect 5088 2688 5152 2692
rect 7445 2748 7509 2752
rect 7445 2692 7449 2748
rect 7449 2692 7505 2748
rect 7505 2692 7509 2748
rect 7445 2688 7509 2692
rect 7525 2748 7589 2752
rect 7525 2692 7529 2748
rect 7529 2692 7585 2748
rect 7585 2692 7589 2748
rect 7525 2688 7589 2692
rect 7605 2748 7669 2752
rect 7605 2692 7609 2748
rect 7609 2692 7665 2748
rect 7665 2692 7669 2748
rect 7605 2688 7669 2692
rect 7685 2748 7749 2752
rect 7685 2692 7689 2748
rect 7689 2692 7745 2748
rect 7745 2692 7749 2748
rect 7685 2688 7749 2692
rect 3549 2204 3613 2208
rect 3549 2148 3553 2204
rect 3553 2148 3609 2204
rect 3609 2148 3613 2204
rect 3549 2144 3613 2148
rect 3629 2204 3693 2208
rect 3629 2148 3633 2204
rect 3633 2148 3689 2204
rect 3689 2148 3693 2204
rect 3629 2144 3693 2148
rect 3709 2204 3773 2208
rect 3709 2148 3713 2204
rect 3713 2148 3769 2204
rect 3769 2148 3773 2204
rect 3709 2144 3773 2148
rect 3789 2204 3853 2208
rect 3789 2148 3793 2204
rect 3793 2148 3849 2204
rect 3849 2148 3853 2204
rect 3789 2144 3853 2148
rect 6146 2204 6210 2208
rect 6146 2148 6150 2204
rect 6150 2148 6206 2204
rect 6206 2148 6210 2204
rect 6146 2144 6210 2148
rect 6226 2204 6290 2208
rect 6226 2148 6230 2204
rect 6230 2148 6286 2204
rect 6286 2148 6290 2204
rect 6226 2144 6290 2148
rect 6306 2204 6370 2208
rect 6306 2148 6310 2204
rect 6310 2148 6366 2204
rect 6366 2148 6370 2204
rect 6306 2144 6370 2148
rect 6386 2204 6450 2208
rect 6386 2148 6390 2204
rect 6390 2148 6446 2204
rect 6446 2148 6450 2204
rect 6386 2144 6450 2148
<< metal4 >>
rect 2242 27776 2563 27792
rect 2242 27712 2250 27776
rect 2314 27712 2330 27776
rect 2394 27712 2410 27776
rect 2474 27712 2490 27776
rect 2554 27712 2563 27776
rect 2242 26688 2563 27712
rect 2242 26624 2250 26688
rect 2314 26624 2330 26688
rect 2394 26624 2410 26688
rect 2474 26624 2490 26688
rect 2554 26624 2563 26688
rect 2242 25600 2563 26624
rect 2242 25536 2250 25600
rect 2314 25536 2330 25600
rect 2394 25536 2410 25600
rect 2474 25536 2490 25600
rect 2554 25536 2563 25600
rect 2242 24512 2563 25536
rect 2242 24448 2250 24512
rect 2314 24448 2330 24512
rect 2394 24448 2410 24512
rect 2474 24448 2490 24512
rect 2554 24448 2563 24512
rect 2242 23424 2563 24448
rect 2242 23360 2250 23424
rect 2314 23360 2330 23424
rect 2394 23360 2410 23424
rect 2474 23360 2490 23424
rect 2554 23360 2563 23424
rect 2242 22336 2563 23360
rect 2242 22272 2250 22336
rect 2314 22272 2330 22336
rect 2394 22272 2410 22336
rect 2474 22272 2490 22336
rect 2554 22272 2563 22336
rect 2242 21248 2563 22272
rect 2242 21184 2250 21248
rect 2314 21184 2330 21248
rect 2394 21184 2410 21248
rect 2474 21184 2490 21248
rect 2554 21184 2563 21248
rect 2242 20160 2563 21184
rect 2242 20096 2250 20160
rect 2314 20096 2330 20160
rect 2394 20096 2410 20160
rect 2474 20096 2490 20160
rect 2554 20096 2563 20160
rect 2242 19072 2563 20096
rect 2242 19008 2250 19072
rect 2314 19008 2330 19072
rect 2394 19008 2410 19072
rect 2474 19008 2490 19072
rect 2554 19008 2563 19072
rect 2242 17984 2563 19008
rect 2242 17920 2250 17984
rect 2314 17920 2330 17984
rect 2394 17920 2410 17984
rect 2474 17920 2490 17984
rect 2554 17920 2563 17984
rect 2242 16896 2563 17920
rect 2242 16832 2250 16896
rect 2314 16832 2330 16896
rect 2394 16832 2410 16896
rect 2474 16832 2490 16896
rect 2554 16832 2563 16896
rect 2242 15808 2563 16832
rect 2242 15744 2250 15808
rect 2314 15744 2330 15808
rect 2394 15744 2410 15808
rect 2474 15744 2490 15808
rect 2554 15744 2563 15808
rect 2242 14720 2563 15744
rect 2242 14656 2250 14720
rect 2314 14656 2330 14720
rect 2394 14656 2410 14720
rect 2474 14656 2490 14720
rect 2554 14656 2563 14720
rect 2242 13632 2563 14656
rect 2242 13568 2250 13632
rect 2314 13568 2330 13632
rect 2394 13568 2410 13632
rect 2474 13568 2490 13632
rect 2554 13568 2563 13632
rect 2242 12544 2563 13568
rect 2242 12480 2250 12544
rect 2314 12480 2330 12544
rect 2394 12480 2410 12544
rect 2474 12480 2490 12544
rect 2554 12480 2563 12544
rect 2242 11456 2563 12480
rect 2242 11392 2250 11456
rect 2314 11392 2330 11456
rect 2394 11392 2410 11456
rect 2474 11392 2490 11456
rect 2554 11392 2563 11456
rect 2242 10368 2563 11392
rect 2242 10304 2250 10368
rect 2314 10304 2330 10368
rect 2394 10304 2410 10368
rect 2474 10304 2490 10368
rect 2554 10304 2563 10368
rect 2242 9280 2563 10304
rect 2242 9216 2250 9280
rect 2314 9216 2330 9280
rect 2394 9216 2410 9280
rect 2474 9216 2490 9280
rect 2554 9216 2563 9280
rect 2242 8192 2563 9216
rect 2242 8128 2250 8192
rect 2314 8128 2330 8192
rect 2394 8128 2410 8192
rect 2474 8128 2490 8192
rect 2554 8128 2563 8192
rect 2242 7104 2563 8128
rect 2242 7040 2250 7104
rect 2314 7040 2330 7104
rect 2394 7040 2410 7104
rect 2474 7040 2490 7104
rect 2554 7040 2563 7104
rect 2242 6016 2563 7040
rect 2242 5952 2250 6016
rect 2314 5952 2330 6016
rect 2394 5952 2410 6016
rect 2474 5952 2490 6016
rect 2554 5952 2563 6016
rect 2242 4928 2563 5952
rect 2242 4864 2250 4928
rect 2314 4864 2330 4928
rect 2394 4864 2410 4928
rect 2474 4864 2490 4928
rect 2554 4864 2563 4928
rect 2242 3840 2563 4864
rect 2242 3776 2250 3840
rect 2314 3776 2330 3840
rect 2394 3776 2410 3840
rect 2474 3776 2490 3840
rect 2554 3776 2563 3840
rect 2242 2752 2563 3776
rect 2242 2688 2250 2752
rect 2314 2688 2330 2752
rect 2394 2688 2410 2752
rect 2474 2688 2490 2752
rect 2554 2688 2563 2752
rect 2242 2128 2563 2688
rect 3541 27232 3861 27792
rect 3541 27168 3549 27232
rect 3613 27168 3629 27232
rect 3693 27168 3709 27232
rect 3773 27168 3789 27232
rect 3853 27168 3861 27232
rect 3541 26144 3861 27168
rect 3541 26080 3549 26144
rect 3613 26080 3629 26144
rect 3693 26080 3709 26144
rect 3773 26080 3789 26144
rect 3853 26080 3861 26144
rect 3541 25056 3861 26080
rect 3541 24992 3549 25056
rect 3613 24992 3629 25056
rect 3693 24992 3709 25056
rect 3773 24992 3789 25056
rect 3853 24992 3861 25056
rect 3541 23968 3861 24992
rect 3541 23904 3549 23968
rect 3613 23904 3629 23968
rect 3693 23904 3709 23968
rect 3773 23904 3789 23968
rect 3853 23904 3861 23968
rect 3541 22880 3861 23904
rect 3541 22816 3549 22880
rect 3613 22816 3629 22880
rect 3693 22816 3709 22880
rect 3773 22816 3789 22880
rect 3853 22816 3861 22880
rect 3541 21792 3861 22816
rect 3541 21728 3549 21792
rect 3613 21728 3629 21792
rect 3693 21728 3709 21792
rect 3773 21728 3789 21792
rect 3853 21728 3861 21792
rect 3541 20704 3861 21728
rect 3541 20640 3549 20704
rect 3613 20640 3629 20704
rect 3693 20640 3709 20704
rect 3773 20640 3789 20704
rect 3853 20640 3861 20704
rect 3541 19616 3861 20640
rect 3541 19552 3549 19616
rect 3613 19552 3629 19616
rect 3693 19552 3709 19616
rect 3773 19552 3789 19616
rect 3853 19552 3861 19616
rect 3541 18528 3861 19552
rect 3541 18464 3549 18528
rect 3613 18464 3629 18528
rect 3693 18464 3709 18528
rect 3773 18464 3789 18528
rect 3853 18464 3861 18528
rect 3541 17440 3861 18464
rect 3541 17376 3549 17440
rect 3613 17376 3629 17440
rect 3693 17376 3709 17440
rect 3773 17376 3789 17440
rect 3853 17376 3861 17440
rect 3541 16352 3861 17376
rect 3541 16288 3549 16352
rect 3613 16288 3629 16352
rect 3693 16288 3709 16352
rect 3773 16288 3789 16352
rect 3853 16288 3861 16352
rect 3541 15264 3861 16288
rect 3541 15200 3549 15264
rect 3613 15200 3629 15264
rect 3693 15200 3709 15264
rect 3773 15200 3789 15264
rect 3853 15200 3861 15264
rect 3541 14176 3861 15200
rect 3541 14112 3549 14176
rect 3613 14112 3629 14176
rect 3693 14112 3709 14176
rect 3773 14112 3789 14176
rect 3853 14112 3861 14176
rect 3541 13088 3861 14112
rect 3541 13024 3549 13088
rect 3613 13024 3629 13088
rect 3693 13024 3709 13088
rect 3773 13024 3789 13088
rect 3853 13024 3861 13088
rect 3541 12000 3861 13024
rect 3541 11936 3549 12000
rect 3613 11936 3629 12000
rect 3693 11936 3709 12000
rect 3773 11936 3789 12000
rect 3853 11936 3861 12000
rect 3541 10912 3861 11936
rect 3541 10848 3549 10912
rect 3613 10848 3629 10912
rect 3693 10848 3709 10912
rect 3773 10848 3789 10912
rect 3853 10848 3861 10912
rect 3541 9824 3861 10848
rect 3541 9760 3549 9824
rect 3613 9760 3629 9824
rect 3693 9760 3709 9824
rect 3773 9760 3789 9824
rect 3853 9760 3861 9824
rect 3541 8736 3861 9760
rect 3541 8672 3549 8736
rect 3613 8672 3629 8736
rect 3693 8672 3709 8736
rect 3773 8672 3789 8736
rect 3853 8672 3861 8736
rect 3541 7648 3861 8672
rect 3541 7584 3549 7648
rect 3613 7584 3629 7648
rect 3693 7584 3709 7648
rect 3773 7584 3789 7648
rect 3853 7584 3861 7648
rect 3541 6560 3861 7584
rect 3541 6496 3549 6560
rect 3613 6496 3629 6560
rect 3693 6496 3709 6560
rect 3773 6496 3789 6560
rect 3853 6496 3861 6560
rect 3541 5472 3861 6496
rect 3541 5408 3549 5472
rect 3613 5408 3629 5472
rect 3693 5408 3709 5472
rect 3773 5408 3789 5472
rect 3853 5408 3861 5472
rect 3541 4384 3861 5408
rect 3541 4320 3549 4384
rect 3613 4320 3629 4384
rect 3693 4320 3709 4384
rect 3773 4320 3789 4384
rect 3853 4320 3861 4384
rect 3541 3296 3861 4320
rect 3541 3232 3549 3296
rect 3613 3232 3629 3296
rect 3693 3232 3709 3296
rect 3773 3232 3789 3296
rect 3853 3232 3861 3296
rect 3541 2208 3861 3232
rect 3541 2144 3549 2208
rect 3613 2144 3629 2208
rect 3693 2144 3709 2208
rect 3773 2144 3789 2208
rect 3853 2144 3861 2208
rect 3541 2128 3861 2144
rect 4840 27776 5160 27792
rect 4840 27712 4848 27776
rect 4912 27712 4928 27776
rect 4992 27712 5008 27776
rect 5072 27712 5088 27776
rect 5152 27712 5160 27776
rect 4840 26688 5160 27712
rect 4840 26624 4848 26688
rect 4912 26624 4928 26688
rect 4992 26624 5008 26688
rect 5072 26624 5088 26688
rect 5152 26624 5160 26688
rect 4840 25600 5160 26624
rect 4840 25536 4848 25600
rect 4912 25536 4928 25600
rect 4992 25536 5008 25600
rect 5072 25536 5088 25600
rect 5152 25536 5160 25600
rect 4840 24512 5160 25536
rect 4840 24448 4848 24512
rect 4912 24448 4928 24512
rect 4992 24448 5008 24512
rect 5072 24448 5088 24512
rect 5152 24448 5160 24512
rect 4840 23424 5160 24448
rect 4840 23360 4848 23424
rect 4912 23360 4928 23424
rect 4992 23360 5008 23424
rect 5072 23360 5088 23424
rect 5152 23360 5160 23424
rect 4840 22336 5160 23360
rect 4840 22272 4848 22336
rect 4912 22272 4928 22336
rect 4992 22272 5008 22336
rect 5072 22272 5088 22336
rect 5152 22272 5160 22336
rect 4840 21248 5160 22272
rect 4840 21184 4848 21248
rect 4912 21184 4928 21248
rect 4992 21184 5008 21248
rect 5072 21184 5088 21248
rect 5152 21184 5160 21248
rect 4840 20160 5160 21184
rect 4840 20096 4848 20160
rect 4912 20096 4928 20160
rect 4992 20096 5008 20160
rect 5072 20096 5088 20160
rect 5152 20096 5160 20160
rect 4840 19072 5160 20096
rect 4840 19008 4848 19072
rect 4912 19008 4928 19072
rect 4992 19008 5008 19072
rect 5072 19008 5088 19072
rect 5152 19008 5160 19072
rect 4840 17984 5160 19008
rect 4840 17920 4848 17984
rect 4912 17920 4928 17984
rect 4992 17920 5008 17984
rect 5072 17920 5088 17984
rect 5152 17920 5160 17984
rect 4840 16896 5160 17920
rect 6138 27232 6458 27792
rect 6138 27168 6146 27232
rect 6210 27168 6226 27232
rect 6290 27168 6306 27232
rect 6370 27168 6386 27232
rect 6450 27168 6458 27232
rect 6138 26144 6458 27168
rect 6138 26080 6146 26144
rect 6210 26080 6226 26144
rect 6290 26080 6306 26144
rect 6370 26080 6386 26144
rect 6450 26080 6458 26144
rect 6138 25056 6458 26080
rect 6138 24992 6146 25056
rect 6210 24992 6226 25056
rect 6290 24992 6306 25056
rect 6370 24992 6386 25056
rect 6450 24992 6458 25056
rect 6138 23968 6458 24992
rect 6138 23904 6146 23968
rect 6210 23904 6226 23968
rect 6290 23904 6306 23968
rect 6370 23904 6386 23968
rect 6450 23904 6458 23968
rect 6138 22880 6458 23904
rect 6138 22816 6146 22880
rect 6210 22816 6226 22880
rect 6290 22816 6306 22880
rect 6370 22816 6386 22880
rect 6450 22816 6458 22880
rect 6138 21792 6458 22816
rect 6138 21728 6146 21792
rect 6210 21728 6226 21792
rect 6290 21728 6306 21792
rect 6370 21728 6386 21792
rect 6450 21728 6458 21792
rect 6138 20704 6458 21728
rect 6138 20640 6146 20704
rect 6210 20640 6226 20704
rect 6290 20640 6306 20704
rect 6370 20640 6386 20704
rect 6450 20640 6458 20704
rect 6138 19616 6458 20640
rect 6138 19552 6146 19616
rect 6210 19552 6226 19616
rect 6290 19552 6306 19616
rect 6370 19552 6386 19616
rect 6450 19552 6458 19616
rect 6138 18528 6458 19552
rect 6138 18464 6146 18528
rect 6210 18464 6226 18528
rect 6290 18464 6306 18528
rect 6370 18464 6386 18528
rect 6450 18464 6458 18528
rect 5947 17916 6013 17917
rect 5947 17852 5948 17916
rect 6012 17852 6013 17916
rect 5947 17851 6013 17852
rect 4840 16832 4848 16896
rect 4912 16832 4928 16896
rect 4992 16832 5008 16896
rect 5072 16832 5088 16896
rect 5152 16832 5160 16896
rect 4840 15808 5160 16832
rect 4840 15744 4848 15808
rect 4912 15744 4928 15808
rect 4992 15744 5008 15808
rect 5072 15744 5088 15808
rect 5152 15744 5160 15808
rect 4840 14720 5160 15744
rect 4840 14656 4848 14720
rect 4912 14656 4928 14720
rect 4992 14656 5008 14720
rect 5072 14656 5088 14720
rect 5152 14656 5160 14720
rect 4840 13632 5160 14656
rect 4840 13568 4848 13632
rect 4912 13568 4928 13632
rect 4992 13568 5008 13632
rect 5072 13568 5088 13632
rect 5152 13568 5160 13632
rect 4840 12544 5160 13568
rect 5950 12749 6010 17851
rect 6138 17440 6458 18464
rect 6138 17376 6146 17440
rect 6210 17376 6226 17440
rect 6290 17376 6306 17440
rect 6370 17376 6386 17440
rect 6450 17376 6458 17440
rect 6138 16352 6458 17376
rect 6138 16288 6146 16352
rect 6210 16288 6226 16352
rect 6290 16288 6306 16352
rect 6370 16288 6386 16352
rect 6450 16288 6458 16352
rect 6138 15264 6458 16288
rect 6138 15200 6146 15264
rect 6210 15200 6226 15264
rect 6290 15200 6306 15264
rect 6370 15200 6386 15264
rect 6450 15200 6458 15264
rect 6138 14176 6458 15200
rect 6138 14112 6146 14176
rect 6210 14112 6226 14176
rect 6290 14112 6306 14176
rect 6370 14112 6386 14176
rect 6450 14112 6458 14176
rect 6138 13088 6458 14112
rect 6138 13024 6146 13088
rect 6210 13024 6226 13088
rect 6290 13024 6306 13088
rect 6370 13024 6386 13088
rect 6450 13024 6458 13088
rect 5947 12748 6013 12749
rect 5947 12684 5948 12748
rect 6012 12684 6013 12748
rect 5947 12683 6013 12684
rect 4840 12480 4848 12544
rect 4912 12480 4928 12544
rect 4992 12480 5008 12544
rect 5072 12480 5088 12544
rect 5152 12480 5160 12544
rect 4840 11456 5160 12480
rect 4840 11392 4848 11456
rect 4912 11392 4928 11456
rect 4992 11392 5008 11456
rect 5072 11392 5088 11456
rect 5152 11392 5160 11456
rect 4840 10368 5160 11392
rect 4840 10304 4848 10368
rect 4912 10304 4928 10368
rect 4992 10304 5008 10368
rect 5072 10304 5088 10368
rect 5152 10304 5160 10368
rect 4840 9280 5160 10304
rect 4840 9216 4848 9280
rect 4912 9216 4928 9280
rect 4992 9216 5008 9280
rect 5072 9216 5088 9280
rect 5152 9216 5160 9280
rect 4840 8192 5160 9216
rect 4840 8128 4848 8192
rect 4912 8128 4928 8192
rect 4992 8128 5008 8192
rect 5072 8128 5088 8192
rect 5152 8128 5160 8192
rect 4840 7104 5160 8128
rect 4840 7040 4848 7104
rect 4912 7040 4928 7104
rect 4992 7040 5008 7104
rect 5072 7040 5088 7104
rect 5152 7040 5160 7104
rect 4840 6016 5160 7040
rect 4840 5952 4848 6016
rect 4912 5952 4928 6016
rect 4992 5952 5008 6016
rect 5072 5952 5088 6016
rect 5152 5952 5160 6016
rect 4840 4928 5160 5952
rect 4840 4864 4848 4928
rect 4912 4864 4928 4928
rect 4992 4864 5008 4928
rect 5072 4864 5088 4928
rect 5152 4864 5160 4928
rect 4840 3840 5160 4864
rect 4840 3776 4848 3840
rect 4912 3776 4928 3840
rect 4992 3776 5008 3840
rect 5072 3776 5088 3840
rect 5152 3776 5160 3840
rect 4840 2752 5160 3776
rect 4840 2688 4848 2752
rect 4912 2688 4928 2752
rect 4992 2688 5008 2752
rect 5072 2688 5088 2752
rect 5152 2688 5160 2752
rect 4840 2128 5160 2688
rect 6138 12000 6458 13024
rect 6138 11936 6146 12000
rect 6210 11936 6226 12000
rect 6290 11936 6306 12000
rect 6370 11936 6386 12000
rect 6450 11936 6458 12000
rect 6138 10912 6458 11936
rect 6138 10848 6146 10912
rect 6210 10848 6226 10912
rect 6290 10848 6306 10912
rect 6370 10848 6386 10912
rect 6450 10848 6458 10912
rect 6138 9824 6458 10848
rect 6138 9760 6146 9824
rect 6210 9760 6226 9824
rect 6290 9760 6306 9824
rect 6370 9760 6386 9824
rect 6450 9760 6458 9824
rect 6138 8736 6458 9760
rect 6138 8672 6146 8736
rect 6210 8672 6226 8736
rect 6290 8672 6306 8736
rect 6370 8672 6386 8736
rect 6450 8672 6458 8736
rect 6138 7648 6458 8672
rect 6138 7584 6146 7648
rect 6210 7584 6226 7648
rect 6290 7584 6306 7648
rect 6370 7584 6386 7648
rect 6450 7584 6458 7648
rect 6138 6560 6458 7584
rect 6138 6496 6146 6560
rect 6210 6496 6226 6560
rect 6290 6496 6306 6560
rect 6370 6496 6386 6560
rect 6450 6496 6458 6560
rect 6138 5472 6458 6496
rect 6138 5408 6146 5472
rect 6210 5408 6226 5472
rect 6290 5408 6306 5472
rect 6370 5408 6386 5472
rect 6450 5408 6458 5472
rect 6138 4384 6458 5408
rect 6138 4320 6146 4384
rect 6210 4320 6226 4384
rect 6290 4320 6306 4384
rect 6370 4320 6386 4384
rect 6450 4320 6458 4384
rect 6138 3296 6458 4320
rect 6138 3232 6146 3296
rect 6210 3232 6226 3296
rect 6290 3232 6306 3296
rect 6370 3232 6386 3296
rect 6450 3232 6458 3296
rect 6138 2208 6458 3232
rect 6138 2144 6146 2208
rect 6210 2144 6226 2208
rect 6290 2144 6306 2208
rect 6370 2144 6386 2208
rect 6450 2144 6458 2208
rect 6138 2128 6458 2144
rect 7437 27776 7757 27792
rect 7437 27712 7445 27776
rect 7509 27712 7525 27776
rect 7589 27712 7605 27776
rect 7669 27712 7685 27776
rect 7749 27712 7757 27776
rect 7437 26688 7757 27712
rect 7437 26624 7445 26688
rect 7509 26624 7525 26688
rect 7589 26624 7605 26688
rect 7669 26624 7685 26688
rect 7749 26624 7757 26688
rect 7437 25600 7757 26624
rect 7437 25536 7445 25600
rect 7509 25536 7525 25600
rect 7589 25536 7605 25600
rect 7669 25536 7685 25600
rect 7749 25536 7757 25600
rect 7437 24512 7757 25536
rect 7437 24448 7445 24512
rect 7509 24448 7525 24512
rect 7589 24448 7605 24512
rect 7669 24448 7685 24512
rect 7749 24448 7757 24512
rect 7437 23424 7757 24448
rect 7437 23360 7445 23424
rect 7509 23360 7525 23424
rect 7589 23360 7605 23424
rect 7669 23360 7685 23424
rect 7749 23360 7757 23424
rect 7437 22336 7757 23360
rect 7437 22272 7445 22336
rect 7509 22272 7525 22336
rect 7589 22272 7605 22336
rect 7669 22272 7685 22336
rect 7749 22272 7757 22336
rect 7437 21248 7757 22272
rect 7437 21184 7445 21248
rect 7509 21184 7525 21248
rect 7589 21184 7605 21248
rect 7669 21184 7685 21248
rect 7749 21184 7757 21248
rect 7437 20160 7757 21184
rect 7437 20096 7445 20160
rect 7509 20096 7525 20160
rect 7589 20096 7605 20160
rect 7669 20096 7685 20160
rect 7749 20096 7757 20160
rect 7437 19072 7757 20096
rect 7437 19008 7445 19072
rect 7509 19008 7525 19072
rect 7589 19008 7605 19072
rect 7669 19008 7685 19072
rect 7749 19008 7757 19072
rect 7437 17984 7757 19008
rect 7437 17920 7445 17984
rect 7509 17920 7525 17984
rect 7589 17920 7605 17984
rect 7669 17920 7685 17984
rect 7749 17920 7757 17984
rect 7437 16896 7757 17920
rect 7437 16832 7445 16896
rect 7509 16832 7525 16896
rect 7589 16832 7605 16896
rect 7669 16832 7685 16896
rect 7749 16832 7757 16896
rect 7437 15808 7757 16832
rect 7437 15744 7445 15808
rect 7509 15744 7525 15808
rect 7589 15744 7605 15808
rect 7669 15744 7685 15808
rect 7749 15744 7757 15808
rect 7437 14720 7757 15744
rect 7437 14656 7445 14720
rect 7509 14656 7525 14720
rect 7589 14656 7605 14720
rect 7669 14656 7685 14720
rect 7749 14656 7757 14720
rect 7437 13632 7757 14656
rect 7437 13568 7445 13632
rect 7509 13568 7525 13632
rect 7589 13568 7605 13632
rect 7669 13568 7685 13632
rect 7749 13568 7757 13632
rect 7437 12544 7757 13568
rect 7437 12480 7445 12544
rect 7509 12480 7525 12544
rect 7589 12480 7605 12544
rect 7669 12480 7685 12544
rect 7749 12480 7757 12544
rect 7437 11456 7757 12480
rect 7437 11392 7445 11456
rect 7509 11392 7525 11456
rect 7589 11392 7605 11456
rect 7669 11392 7685 11456
rect 7749 11392 7757 11456
rect 7437 10368 7757 11392
rect 7437 10304 7445 10368
rect 7509 10304 7525 10368
rect 7589 10304 7605 10368
rect 7669 10304 7685 10368
rect 7749 10304 7757 10368
rect 7437 9280 7757 10304
rect 7437 9216 7445 9280
rect 7509 9216 7525 9280
rect 7589 9216 7605 9280
rect 7669 9216 7685 9280
rect 7749 9216 7757 9280
rect 7437 8192 7757 9216
rect 7437 8128 7445 8192
rect 7509 8128 7525 8192
rect 7589 8128 7605 8192
rect 7669 8128 7685 8192
rect 7749 8128 7757 8192
rect 7437 7104 7757 8128
rect 7437 7040 7445 7104
rect 7509 7040 7525 7104
rect 7589 7040 7605 7104
rect 7669 7040 7685 7104
rect 7749 7040 7757 7104
rect 7437 6016 7757 7040
rect 7437 5952 7445 6016
rect 7509 5952 7525 6016
rect 7589 5952 7605 6016
rect 7669 5952 7685 6016
rect 7749 5952 7757 6016
rect 7437 4928 7757 5952
rect 7437 4864 7445 4928
rect 7509 4864 7525 4928
rect 7589 4864 7605 4928
rect 7669 4864 7685 4928
rect 7749 4864 7757 4928
rect 7437 3840 7757 4864
rect 7437 3776 7445 3840
rect 7509 3776 7525 3840
rect 7589 3776 7605 3840
rect 7669 3776 7685 3840
rect 7749 3776 7757 3840
rect 7437 2752 7757 3776
rect 7437 2688 7445 2752
rect 7509 2688 7525 2752
rect 7589 2688 7605 2752
rect 7669 2688 7685 2752
rect 7749 2688 7757 2752
rect 7437 2128 7757 2688
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.dstage\[1\].id.delayenb0_TE_B $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635306529
transform -1 0 2760 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635306529
transform 1 0 2484 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635306529
transform 1 0 3036 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635306529
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_15
timestamp 1635306529
transform 1 0 2484 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_18 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635306529
transform 1 0 2760 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1635306529
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635306529
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1635306529
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635306529
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_30
timestamp 1635306529
transform 1 0 3864 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_24
timestamp 1635306529
transform 1 0 3312 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635306529
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24
timestamp 1635306529
transform 1 0 3312 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.dstage\[1\].id.delayen0_TE
timestamp 1635306529
transform 1 0 3128 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__26__RESET_B
timestamp 1635306529
transform -1 0 3312 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__21__C
timestamp 1635306529
transform 1 0 3956 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__12__A
timestamp 1635306529
transform 1 0 3680 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__nor3_2  _21_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635306529
transform 1 0 4508 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _12_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635306529
transform 1 0 4232 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_41
timestamp 1635306529
transform 1 0 4876 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_37
timestamp 1635306529
transform 1 0 4508 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33
timestamp 1635306529
transform 1 0 4140 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _23_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635306529
transform 1 0 4968 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _16_
timestamp 1635306529
transform 1 0 5612 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 1635306529
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52
timestamp 1635306529
transform 1 0 5888 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45
timestamp 1635306529
transform 1 0 5244 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_2  ring.dstage\[1\].id.delayen0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635306529
transform -1 0 7728 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _17_
timestamp 1635306529
transform -1 0 6624 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1635306529
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1635306529
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_57
timestamp 1635306529
transform 1 0 6348 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1635306529
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64
timestamp 1635306529
transform 1 0 6992 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_60
timestamp 1635306529
transform 1 0 6624 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__einvn_8  ring.dstage\[1\].id.delayenb0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635306529
transform 1 0 6532 0 -1 3264
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_8  FILLER_0_72 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635306529
transform 1 0 7728 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80
timestamp 1635306529
transform 1 0 8464 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_77
timestamp 1635306529
transform 1 0 8188 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1635306529
transform -1 0 8832 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1635306529
transform -1 0 8832 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__18__C
timestamp 1635306529
transform -1 0 2760 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_15
timestamp 1635306529
transform 1 0 2484 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_18
timestamp 1635306529
transform 1 0 2760 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1635306529
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1635306529
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__18__A
timestamp 1635306529
transform 1 0 3772 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__18__B
timestamp 1635306529
transform 1 0 3128 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_24
timestamp 1635306529
transform 1 0 3312 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_31
timestamp 1635306529
transform 1 0 3956 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_43
timestamp 1635306529
transform 1 0 5060 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1635306529
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__nor3_2  _18_
timestamp 1635306529
transform 1 0 4324 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_2  _26_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635306529
transform 1 0 5428 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_4  FILLER_2_68
timestamp 1635306529
transform 1 0 7360 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_72
timestamp 1635306529
transform 1 0 7728 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_77
timestamp 1635306529
transform 1 0 8188 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1635306529
transform -1 0 8832 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ring.dstage\[2\].id.delaybuf0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635306529
transform -1 0 8188 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__20__A
timestamp 1635306529
transform 1 0 2208 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.dstage\[2\].id.delayenb0_TE_B
timestamp 1635306529
transform -1 0 1840 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_14
timestamp 1635306529
transform 1 0 2392 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_3_3
timestamp 1635306529
transform 1 0 1380 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_8
timestamp 1635306529
transform 1 0 1840 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1635306529
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_2  _20_
timestamp 1635306529
transform 1 0 2760 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_26
timestamp 1635306529
transform 1 0 3496 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_39
timestamp 1635306529
transform 1 0 4692 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _22_
timestamp 1635306529
transform 1 0 5060 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _24_
timestamp 1635306529
transform -1 0 4692 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_3_52
timestamp 1635306529
transform 1 0 5888 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_57
timestamp 1635306529
transform 1 0 6348 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1635306529
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__einvn_8  ring.dstage\[2\].id.delayenb0
timestamp 1635306529
transform -1 0 8188 0 -1 4352
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_4  FILLER_3_77
timestamp 1635306529
transform 1 0 8188 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1635306529
transform -1 0 8832 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__20__C
timestamp 1635306529
transform -1 0 2760 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_15
timestamp 1635306529
transform 1 0 2484 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_18
timestamp 1635306529
transform 1 0 2760 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1635306529
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1635306529
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__19__B
timestamp 1635306529
transform 1 0 3128 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_24
timestamp 1635306529
transform 1 0 3312 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_29
timestamp 1635306529
transform 1 0 3772 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_41
timestamp 1635306529
transform 1 0 4876 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1635306529
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__nor3_2  _19_
timestamp 1635306529
transform -1 0 4876 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_2  _27_
timestamp 1635306529
transform -1 0 7176 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_4  FILLER_4_66
timestamp 1635306529
transform 1 0 7176 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_77
timestamp 1635306529
transform 1 0 8188 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1635306529
transform -1 0 8832 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ring.dstage\[2\].id.delayen0
timestamp 1635306529
transform -1 0 8188 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.dstage\[2\].id.delayen0_TE
timestamp 1635306529
transform -1 0 3220 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.dstage\[2\].id.delayenb1_TE_B
timestamp 1635306529
transform -1 0 2668 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_17
timestamp 1635306529
transform 1 0 2668 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1635306529
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1635306529
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__13__A
timestamp 1635306529
transform 1 0 3588 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_23
timestamp 1635306529
transform 1 0 3220 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_29
timestamp 1635306529
transform 1 0 3772 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_36
timestamp 1635306529
transform 1 0 4416 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _13_
timestamp 1635306529
transform -1 0 4416 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _25_
timestamp 1635306529
transform -1 0 5612 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_5_49
timestamp 1635306529
transform 1 0 5612 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1635306529
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_57
timestamp 1635306529
transform 1 0 6348 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_62
timestamp 1635306529
transform 1 0 6808 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1635306529
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  ring.dstage\[3\].id.delaybuf0
timestamp 1635306529
transform -1 0 6808 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_77
timestamp 1635306529
transform 1 0 8188 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1635306529
transform -1 0 8832 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__einvn_4  ring.dstage\[2\].id.delayenb1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635306529
transform -1 0 8188 0 -1 5440
box -38 -48 1050 592
use sky130_fd_sc_hd__decap_6  FILLER_6_15
timestamp 1635306529
transform 1 0 2484 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_21
timestamp 1635306529
transform 1 0 3036 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1635306529
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1635306529
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1635306529
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1635306529
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1635306529
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_24
timestamp 1635306529
transform 1 0 3312 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.dstage\[2\].id.delayen1_TE
timestamp 1635306529
transform 1 0 3128 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1635306529
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_31
timestamp 1635306529
transform 1 0 3956 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_27
timestamp 1635306529
transform 1 0 3588 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_29
timestamp 1635306529
transform 1 0 3772 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.dstage\[1\].id.delayenb1_TE_B
timestamp 1635306529
transform -1 0 3956 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__19__C
timestamp 1635306529
transform -1 0 4140 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_33
timestamp 1635306529
transform 1 0 4140 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.dstage\[1\].id.delayen1_TE
timestamp 1635306529
transform 1 0 4324 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__clkinv_1  ring.dstage\[2\].id.delayint0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635306529
transform -1 0 5152 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ring.dstage\[2\].id.delaybuf1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635306529
transform -1 0 4784 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_37
timestamp 1635306529
transform 1 0 4508 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_40
timestamp 1635306529
transform 1 0 4784 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_2  ring.dstage\[2\].id.delayen1
timestamp 1635306529
transform -1 0 6440 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_1  ring.dstage\[1\].id.delayint0
timestamp 1635306529
transform -1 0 5428 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ring.dstage\[1\].id.delaybuf0
timestamp 1635306529
transform 1 0 5520 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_52
timestamp 1635306529
transform 1 0 5888 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_44
timestamp 1635306529
transform 1 0 5152 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_47
timestamp 1635306529
transform 1 0 5428 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_2  ring.dstage\[1\].id.delayen1
timestamp 1635306529
transform 1 0 6900 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1635306529
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_59
timestamp 1635306529
transform 1 0 6532 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_58
timestamp 1635306529
transform 1 0 6440 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__27__RESET_B
timestamp 1635306529
transform 1 0 6348 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__einvn_4  ring.dstage\[1\].id.delayenb1
timestamp 1635306529
transform -1 0 7820 0 1 5440
box -38 -48 1050 592
use sky130_fd_sc_hd__decap_8  FILLER_6_73
timestamp 1635306529
transform 1 0 7820 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_70
timestamp 1635306529
transform 1 0 7544 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_77
timestamp 1635306529
transform 1 0 8188 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1635306529
transform -1 0 8832 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1635306529
transform -1 0 8832 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ring.dstage\[1\].id.delaybuf1
timestamp 1635306529
transform 1 0 7912 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1635306529
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1635306529
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1635306529
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1635306529
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_29
timestamp 1635306529
transform 1 0 3772 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_35
timestamp 1635306529
transform 1 0 4324 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_39
timestamp 1635306529
transform 1 0 4692 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1635306529
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _15_
timestamp 1635306529
transform 1 0 4416 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _28_
timestamp 1635306529
transform 1 0 5060 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_4  FILLER_8_64
timestamp 1635306529
transform 1 0 6992 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_75
timestamp 1635306529
transform 1 0 8004 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1635306529
transform -1 0 8832 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ring.dstage\[0\].id.delayen0
timestamp 1635306529
transform -1 0 8004 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1635306529
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1635306529
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1635306529
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__28__RESET_B
timestamp 1635306529
transform 1 0 4968 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.dstage\[0\].id.delayen0_TE
timestamp 1635306529
transform 1 0 4416 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.dstage\[0\].id.delayenb0_TE_B
timestamp 1635306529
transform -1 0 4048 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_27
timestamp 1635306529
transform 1 0 3588 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_32
timestamp 1635306529
transform 1 0 4048 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_38
timestamp 1635306529
transform 1 0 4600 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_44
timestamp 1635306529
transform 1 0 5152 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_52
timestamp 1635306529
transform 1 0 5888 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1635306529
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__einvn_8  ring.dstage\[0\].id.delayenb0
timestamp 1635306529
transform 1 0 6348 0 -1 7616
box -38 -48 1694 592
use sky130_fd_sc_hd__clkinv_2  ring.ibufp00 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635306529
transform 1 0 5520 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_75
timestamp 1635306529
transform 1 0 8004 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1635306529
transform -1 0 8832 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_10_15
timestamp 1635306529
transform 1 0 2484 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_21
timestamp 1635306529
transform 1 0 3036 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1635306529
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1635306529
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__14__A
timestamp 1635306529
transform -1 0 4416 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.dstage\[3\].id.delayenb1_TE_B
timestamp 1635306529
transform -1 0 3312 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_24
timestamp 1635306529
transform 1 0 3312 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_29
timestamp 1635306529
transform 1 0 3772 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_33
timestamp 1635306529
transform 1 0 4140 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_36
timestamp 1635306529
transform 1 0 4416 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_43
timestamp 1635306529
transform 1 0 5060 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1635306529
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _14_
timestamp 1635306529
transform 1 0 4784 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_10_60
timestamp 1635306529
transform 1 0 6624 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkinv_8  ring.ibufp01 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635306529
transform 1 0 5428 0 1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_10_77
timestamp 1635306529
transform 1 0 8188 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1635306529
transform -1 0 8832 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__einvn_4  ring.dstage\[3\].id.delayenb1
timestamp 1635306529
transform -1 0 8188 0 1 7616
box -38 -48 1050 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1635306529
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1635306529
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1635306529
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.dstage\[3\].id.delayen0_TE
timestamp 1635306529
transform -1 0 4232 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_27
timestamp 1635306529
transform 1 0 3588 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_31
timestamp 1635306529
transform 1 0 3956 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_34
timestamp 1635306529
transform 1 0 4232 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_41
timestamp 1635306529
transform 1 0 4876 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ring.dstage\[3\].id.delaybuf1
timestamp 1635306529
transform -1 0 4876 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_52
timestamp 1635306529
transform 1 0 5888 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_57
timestamp 1635306529
transform 1 0 6348 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1635306529
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__einvp_2  ring.dstage\[3\].id.delayen0
timestamp 1635306529
transform 1 0 5244 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ring.dstage\[3\].id.delayenb0
timestamp 1635306529
transform -1 0 8188 0 -1 8704
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_4  FILLER_11_77
timestamp 1635306529
transform 1 0 8188 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1635306529
transform -1 0 8832 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1635306529
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1635306529
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1635306529
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.dstage\[3\].id.delayenb0_TE_B
timestamp 1635306529
transform -1 0 5060 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1635306529
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_29
timestamp 1635306529
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_43
timestamp 1635306529
transform 1 0 5060 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1635306529
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.dstage\[0\].id.delayen1_TE
timestamp 1635306529
transform -1 0 5612 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_49
timestamp 1635306529
transform 1 0 5612 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_56
timestamp 1635306529
transform 1 0 6256 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_2  ring.dstage\[0\].id.delayen1
timestamp 1635306529
transform 1 0 6624 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_1  ring.dstage\[0\].id.delayint0
timestamp 1635306529
transform -1 0 6256 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_67
timestamp 1635306529
transform 1 0 7268 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_75
timestamp 1635306529
transform 1 0 8004 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1635306529
transform -1 0 8832 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ring.dstage\[0\].id.delaybuf0
timestamp 1635306529
transform 1 0 7636 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1635306529
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1635306529
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1635306529
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1635306529
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1635306529
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1635306529
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1635306529
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_39
timestamp 1635306529
transform 1 0 4692 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1635306529
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_29
timestamp 1635306529
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_41
timestamp 1635306529
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1635306529
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_53
timestamp 1635306529
transform 1 0 5980 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_52
timestamp 1635306529
transform 1 0 5888 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_13_47
timestamp 1635306529
transform 1 0 5428 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.dstage\[0\].id.delayenb1_TE_B
timestamp 1635306529
transform 1 0 5704 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__clkinv_1  ring.dstage\[3\].id.delayint0
timestamp 1635306529
transform -1 0 7176 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1635306529
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_59
timestamp 1635306529
transform 1 0 6532 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_57
timestamp 1635306529
transform 1 0 6348 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.dstage\[3\].id.delayen1_TE
timestamp 1635306529
transform 1 0 6348 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__einvn_4  ring.dstage\[0\].id.delayenb1
timestamp 1635306529
transform 1 0 6440 0 -1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__decap_4  FILLER_13_69
timestamp 1635306529
transform 1 0 7452 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_76
timestamp 1635306529
transform 1 0 8096 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_80
timestamp 1635306529
transform 1 0 8464 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_66
timestamp 1635306529
transform 1 0 7176 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_77
timestamp 1635306529
transform 1 0 8188 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1635306529
transform -1 0 8832 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1635306529
transform -1 0 8832 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ring.dstage\[0\].id.delaybuf1
timestamp 1635306529
transform 1 0 7820 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ring.dstage\[3\].id.delayen1
timestamp 1635306529
transform -1 0 8188 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1635306529
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1635306529
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1635306529
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_27
timestamp 1635306529
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_39
timestamp 1635306529
transform 1 0 4692 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.dstage\[4\].id.delayenb1_TE_B
timestamp 1635306529
transform -1 0 5888 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_47
timestamp 1635306529
transform 1 0 5428 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_52
timestamp 1635306529
transform 1 0 5888 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_61
timestamp 1635306529
transform 1 0 6716 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1635306529
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  ring.dstage\[4\].id.delaybuf0
timestamp 1635306529
transform 1 0 6348 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__einvn_4  ring.dstage\[4\].id.delayenb1
timestamp 1635306529
transform -1 0 8096 0 -1 10880
box -38 -48 1050 592
use sky130_fd_sc_hd__decap_4  FILLER_15_76
timestamp 1635306529
transform 1 0 8096 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_80
timestamp 1635306529
transform 1 0 8464 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1635306529
transform -1 0 8832 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1635306529
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1635306529
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1635306529
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1635306529
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_29
timestamp 1635306529
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_41
timestamp 1635306529
transform 1 0 4876 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1635306529
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.dstage\[4\].id.delayenb0_TE_B
timestamp 1635306529
transform -1 0 5520 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_45
timestamp 1635306529
transform 1 0 5244 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_48
timestamp 1635306529
transform 1 0 5520 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_55
timestamp 1635306529
transform 1 0 6164 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__einvn_8  ring.dstage\[4\].id.delayenb0
timestamp 1635306529
transform -1 0 8188 0 1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__clkinv_1  ring.dstage\[4\].id.delayint0
timestamp 1635306529
transform -1 0 6164 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_77
timestamp 1635306529
transform 1 0 8188 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1635306529
transform -1 0 8832 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1635306529
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1635306529
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1635306529
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_27
timestamp 1635306529
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_39
timestamp 1635306529
transform 1 0 4692 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.dstage\[4\].id.delayen0_TE
timestamp 1635306529
transform 1 0 5704 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_47
timestamp 1635306529
transform 1 0 5428 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_52
timestamp 1635306529
transform 1 0 5888 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_57
timestamp 1635306529
transform 1 0 6348 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_65
timestamp 1635306529
transform 1 0 7084 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1635306529
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  ring.dstage\[5\].id.delaybuf0
timestamp 1635306529
transform 1 0 6716 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_76
timestamp 1635306529
transform 1 0 8096 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_80
timestamp 1635306529
transform 1 0 8464 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1635306529
transform -1 0 8832 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ring.dstage\[4\].id.delayen0
timestamp 1635306529
transform -1 0 8096 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1635306529
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1635306529
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1635306529
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1635306529
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_29
timestamp 1635306529
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_41
timestamp 1635306529
transform 1 0 4876 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1635306529
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.dstage\[4\].id.delayen1_TE
timestamp 1635306529
transform 1 0 5796 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_49
timestamp 1635306529
transform 1 0 5612 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_53
timestamp 1635306529
transform 1 0 5980 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_62
timestamp 1635306529
transform 1 0 6808 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_1  ring.iss.reseten0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635306529
transform 1 0 6348 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__decap_8  FILLER_18_73
timestamp 1635306529
transform 1 0 7820 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1635306529
transform -1 0 8832 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ring.dstage\[4\].id.delayen1
timestamp 1635306529
transform 1 0 7176 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1635306529
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1635306529
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1635306529
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1635306529
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1635306529
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1635306529
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_27
timestamp 1635306529
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_39
timestamp 1635306529
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1635306529
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_29
timestamp 1635306529
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_41
timestamp 1635306529
transform 1 0 4876 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1635306529
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_52
timestamp 1635306529
transform 1 0 5888 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_49
timestamp 1635306529
transform 1 0 5612 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1635306529
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.iss.delayen0_TE
timestamp 1635306529
transform -1 0 5888 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1635306529
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_56
timestamp 1635306529
transform 1 0 6256 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_57
timestamp 1635306529
transform 1 0 6348 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1635306529
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.dstage\[5\].id.delayen0_TE
timestamp 1635306529
transform 1 0 6348 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  ring.iss.const1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635306529
transform -1 0 6808 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ring.dstage\[5\].id.delaybuf1
timestamp 1635306529
transform -1 0 7176 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_59
timestamp 1635306529
transform 1 0 6532 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_62
timestamp 1635306529
transform 1 0 6808 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_1  ring.dstage\[5\].id.delayint0
timestamp 1635306529
transform -1 0 7452 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ring.dstage\[5\].id.delayen0
timestamp 1635306529
transform -1 0 8188 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  ring.dstage\[4\].id.delaybuf1
timestamp 1635306529
transform 1 0 7820 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_66
timestamp 1635306529
transform 1 0 7176 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_69
timestamp 1635306529
transform 1 0 7452 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1635306529
transform -1 0 8832 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1635306529
transform -1 0 8832 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_77
timestamp 1635306529
transform 1 0 8188 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_80
timestamp 1635306529
transform 1 0 8464 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_76
timestamp 1635306529
transform 1 0 8096 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1635306529
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1635306529
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1635306529
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_27
timestamp 1635306529
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_39
timestamp 1635306529
transform 1 0 4692 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.dstage\[5\].id.delayenb0_TE_B
timestamp 1635306529
transform -1 0 5888 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_47
timestamp 1635306529
transform 1 0 5428 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_52
timestamp 1635306529
transform 1 0 5888 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_57
timestamp 1635306529
transform 1 0 6348 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1635306529
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__einvn_8  ring.dstage\[5\].id.delayenb0
timestamp 1635306529
transform 1 0 6532 0 -1 14144
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_4  FILLER_21_77
timestamp 1635306529
transform 1 0 8188 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1635306529
transform -1 0 8832 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1635306529
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1635306529
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1635306529
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1635306529
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_29
timestamp 1635306529
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_41
timestamp 1635306529
transform 1 0 4876 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1635306529
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__einvp_2  ring.iss.delayen0
timestamp 1635306529
transform 1 0 5060 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_22_50
timestamp 1635306529
transform 1 0 5704 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__einvn_8  ring.iss.delayenb0
timestamp 1635306529
transform 1 0 6072 0 1 14144
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_8  FILLER_22_72
timestamp 1635306529
transform 1 0 7728 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_80
timestamp 1635306529
transform 1 0 8464 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1635306529
transform -1 0 8832 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1635306529
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1635306529
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1635306529
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.dstage\[5\].id.delayenb1_TE_B
timestamp 1635306529
transform -1 0 5152 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.iss.ctrlen0_B
timestamp 1635306529
transform -1 0 4600 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_27
timestamp 1635306529
transform 1 0 3588 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_35
timestamp 1635306529
transform 1 0 4324 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_38
timestamp 1635306529
transform 1 0 4600 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_44
timestamp 1635306529
transform 1 0 5152 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_52
timestamp 1635306529
transform 1 0 5888 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_62
timestamp 1635306529
transform 1 0 6808 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1635306529
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  ring.dstage\[6\].id.delaybuf0
timestamp 1635306529
transform 1 0 5520 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__or2_2  ring.iss.ctrlen0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635306529
transform -1 0 6808 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_23_77
timestamp 1635306529
transform 1 0 8188 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1635306529
transform -1 0 8832 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__einvn_4  ring.dstage\[5\].id.delayenb1
timestamp 1635306529
transform -1 0 8188 0 -1 15232
box -38 -48 1050 592
use sky130_fd_sc_hd__decap_12  FILLER_24_15
timestamp 1635306529
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1635306529
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1635306529
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.iss.delayen1_TE
timestamp 1635306529
transform -1 0 4876 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1635306529
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_29
timestamp 1635306529
transform 1 0 3772 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_37
timestamp 1635306529
transform 1 0 4508 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_41
timestamp 1635306529
transform 1 0 4876 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1635306529
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.dstage\[5\].id.delayen1_TE
timestamp 1635306529
transform 1 0 5244 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_47
timestamp 1635306529
transform 1 0 5428 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_54
timestamp 1635306529
transform 1 0 6072 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_65
timestamp 1635306529
transform 1 0 7084 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_2  ring.iss.delayen1
timestamp 1635306529
transform -1 0 7084 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_1  ring.iss.delayint0
timestamp 1635306529
transform -1 0 6072 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_76
timestamp 1635306529
transform 1 0 8096 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_80
timestamp 1635306529
transform 1 0 8464 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1635306529
transform -1 0 8832 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ring.dstage\[5\].id.delayen1
timestamp 1635306529
transform -1 0 8096 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_25_15
timestamp 1635306529
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1635306529
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1635306529
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.iss.delayenb1_TE_B
timestamp 1635306529
transform 1 0 5060 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_27
timestamp 1635306529
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_39
timestamp 1635306529
transform 1 0 4692 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_45
timestamp 1635306529
transform 1 0 5244 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_52
timestamp 1635306529
transform 1 0 5888 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_57
timestamp 1635306529
transform 1 0 6348 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1635306529
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  ring.iss.delaybuf0
timestamp 1635306529
transform -1 0 5888 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__einvn_4  ring.iss.delayenb1
timestamp 1635306529
transform -1 0 7544 0 -1 16320
box -38 -48 1050 592
use sky130_fd_sc_hd__decap_4  FILLER_25_70
timestamp 1635306529
transform 1 0 7544 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_77
timestamp 1635306529
transform 1 0 8188 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1635306529
transform -1 0 8832 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  ring.dstage\[6\].id.delayint0
timestamp 1635306529
transform 1 0 7912 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1635306529
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1635306529
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_15
timestamp 1635306529
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_3
timestamp 1635306529
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1635306529
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1635306529
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.dstage\[6\].id.delayenb1_TE_B
timestamp 1635306529
transform -1 0 5244 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1635306529
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_29
timestamp 1635306529
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_41
timestamp 1635306529
transform 1 0 4876 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_27
timestamp 1635306529
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_39
timestamp 1635306529
transform 1 0 4692 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1635306529
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_52
timestamp 1635306529
transform 1 0 5888 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_27_47
timestamp 1635306529
transform 1 0 5428 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_51
timestamp 1635306529
transform 1 0 5796 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_45
timestamp 1635306529
transform 1 0 5244 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.dstage\[6\].id.delayenb0_TE_B
timestamp 1635306529
transform 1 0 5704 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.dstage\[6\].id.delayen0_TE
timestamp 1635306529
transform -1 0 5796 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_2  ring.dstage\[6\].id.delayen0
timestamp 1635306529
transform 1 0 6164 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1635306529
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_57
timestamp 1635306529
transform 1 0 6348 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_62
timestamp 1635306529
transform 1 0 6808 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__einvn_8  ring.dstage\[6\].id.delayenb0
timestamp 1635306529
transform -1 0 8188 0 -1 17408
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_4  FILLER_26_77
timestamp 1635306529
transform 1 0 8188 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_77
timestamp 1635306529
transform 1 0 8188 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1635306529
transform -1 0 8832 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1635306529
transform -1 0 8832 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__einvn_4  ring.dstage\[6\].id.delayenb1
timestamp 1635306529
transform -1 0 8188 0 1 16320
box -38 -48 1050 592
use sky130_fd_sc_hd__decap_12  FILLER_28_15
timestamp 1635306529
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_3
timestamp 1635306529
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1635306529
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1635306529
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_29
timestamp 1635306529
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_41
timestamp 1635306529
transform 1 0 4876 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1635306529
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.dstage\[6\].id.delayen1_TE
timestamp 1635306529
transform 1 0 5244 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_47
timestamp 1635306529
transform 1 0 5428 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_58
timestamp 1635306529
transform 1 0 6440 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_2  ring.dstage\[11\].id.delayen0
timestamp 1635306529
transform 1 0 6808 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ring.dstage\[6\].id.delayen1
timestamp 1635306529
transform 1 0 5796 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_28_69
timestamp 1635306529
transform 1 0 7452 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_73
timestamp 1635306529
transform 1 0 7820 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_77
timestamp 1635306529
transform 1 0 8188 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1635306529
transform -1 0 8832 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ring.dstage\[6\].id.delaybuf1
timestamp 1635306529
transform 1 0 7912 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_15
timestamp 1635306529
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_3
timestamp 1635306529
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1635306529
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_27
timestamp 1635306529
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_39
timestamp 1635306529
transform 1 0 4692 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.dstage\[11\].id.delayenb0_TE_B
timestamp 1635306529
transform -1 0 5888 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_47
timestamp 1635306529
transform 1 0 5428 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_52
timestamp 1635306529
transform 1 0 5888 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1635306529
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__einvn_8  ring.dstage\[11\].id.delayenb0
timestamp 1635306529
transform 1 0 6348 0 -1 18496
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_6  FILLER_29_75
timestamp 1635306529
transform 1 0 8004 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1635306529
transform -1 0 8832 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_15
timestamp 1635306529
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_3
timestamp 1635306529
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1635306529
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1635306529
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_29
timestamp 1635306529
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_41
timestamp 1635306529
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1635306529
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.dstage\[11\].id.delayen1_TE
timestamp 1635306529
transform -1 0 6808 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_53
timestamp 1635306529
transform 1 0 5980 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_59
timestamp 1635306529
transform 1 0 6532 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_62
timestamp 1635306529
transform 1 0 6808 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.dstage\[11\].id.delayen0_TE
timestamp 1635306529
transform -1 0 8004 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_69
timestamp 1635306529
transform 1 0 7452 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_75
timestamp 1635306529
transform 1 0 8004 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1635306529
transform -1 0 8832 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  ring.dstage\[11\].id.delayint0
timestamp 1635306529
transform 1 0 7176 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_15
timestamp 1635306529
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_3
timestamp 1635306529
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1635306529
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_27
timestamp 1635306529
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_39
timestamp 1635306529
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1635306529
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1635306529
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_57
timestamp 1635306529
transform 1 0 6348 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1635306529
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__einvp_2  ring.dstage\[11\].id.delayen1
timestamp 1635306529
transform 1 0 6716 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_31_68
timestamp 1635306529
transform 1 0 7360 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_72
timestamp 1635306529
transform 1 0 7728 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_77
timestamp 1635306529
transform 1 0 8188 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1635306529
transform -1 0 8832 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ring.dstage\[7\].id.delaybuf0
timestamp 1635306529
transform 1 0 7820 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_15
timestamp 1635306529
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1635306529
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1635306529
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1635306529
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_29
timestamp 1635306529
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_41
timestamp 1635306529
transform 1 0 4876 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1635306529
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.dstage\[11\].id.delayenb1_TE_B
timestamp 1635306529
transform -1 0 6164 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.dstage\[7\].id.delayenb0_TE_B
timestamp 1635306529
transform 1 0 5428 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_49
timestamp 1635306529
transform 1 0 5612 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_55
timestamp 1635306529
transform 1 0 6164 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__einvn_4  ring.dstage\[11\].id.delayenb1
timestamp 1635306529
transform 1 0 6532 0 1 19584
box -38 -48 1050 592
use sky130_fd_sc_hd__decap_4  FILLER_32_70
timestamp 1635306529
transform 1 0 7544 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_77
timestamp 1635306529
transform 1 0 8188 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1635306529
transform -1 0 8832 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ring.dstage\[11\].id.delaybuf1
timestamp 1635306529
transform 1 0 7912 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_15
timestamp 1635306529
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_3
timestamp 1635306529
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_15
timestamp 1635306529
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3
timestamp 1635306529
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1635306529
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1635306529
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.dstage\[7\].id.delayen0_TE
timestamp 1635306529
transform -1 0 4784 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.dstage\[7\].id.delayen1_TE
timestamp 1635306529
transform -1 0 5244 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_27
timestamp 1635306529
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_39
timestamp 1635306529
transform 1 0 4692 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1635306529
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_29
timestamp 1635306529
transform 1 0 3772 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_37
timestamp 1635306529
transform 1 0 4508 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_40
timestamp 1635306529
transform 1 0 4784 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1635306529
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__einvp_2  ring.dstage\[7\].id.delayen1
timestamp 1635306529
transform 1 0 5152 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  ring.dstage\[7\].id.delaybuf1
timestamp 1635306529
transform 1 0 5612 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_51
timestamp 1635306529
transform 1 0 5796 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_52
timestamp 1635306529
transform 1 0 5888 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_45
timestamp 1635306529
transform 1 0 5244 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_2  ring.dstage\[7\].id.delayen0
timestamp 1635306529
transform -1 0 6808 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1635306529
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_62
timestamp 1635306529
transform 1 0 6808 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_57
timestamp 1635306529
transform 1 0 6348 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__einvn_8  ring.dstage\[7\].id.delayenb0
timestamp 1635306529
transform -1 0 8188 0 -1 20672
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_4  FILLER_33_77
timestamp 1635306529
transform 1 0 8188 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_77
timestamp 1635306529
transform 1 0 8188 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1635306529
transform -1 0 8832 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1635306529
transform -1 0 8832 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__einvn_4  ring.dstage\[7\].id.delayenb1
timestamp 1635306529
transform -1 0 8188 0 1 20672
box -38 -48 1050 592
use sky130_fd_sc_hd__decap_12  FILLER_35_15
timestamp 1635306529
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_3
timestamp 1635306529
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1635306529
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.dstage\[7\].id.delayenb1_TE_B
timestamp 1635306529
transform -1 0 5244 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_35_27
timestamp 1635306529
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_39
timestamp 1635306529
transform 1 0 4692 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_45
timestamp 1635306529
transform 1 0 5244 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_52
timestamp 1635306529
transform 1 0 5888 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_57
timestamp 1635306529
transform 1 0 6348 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_61
timestamp 1635306529
transform 1 0 6716 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1635306529
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__einvp_2  ring.dstage\[10\].id.delayen0
timestamp 1635306529
transform -1 0 7452 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_1  ring.dstage\[7\].id.delayint0
timestamp 1635306529
transform 1 0 5612 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_69
timestamp 1635306529
transform 1 0 7452 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_77
timestamp 1635306529
transform 1 0 8188 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1635306529
transform -1 0 8832 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ring.dstage\[11\].id.delaybuf0
timestamp 1635306529
transform 1 0 7820 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_15
timestamp 1635306529
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_3
timestamp 1635306529
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1635306529
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1635306529
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_29
timestamp 1635306529
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_41
timestamp 1635306529
transform 1 0 4876 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1635306529
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.dstage\[10\].id.delayen0_TE
timestamp 1635306529
transform -1 0 5980 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.dstage\[10\].id.delayenb0_TE_B
timestamp 1635306529
transform -1 0 5428 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_47
timestamp 1635306529
transform 1 0 5428 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_53
timestamp 1635306529
transform 1 0 5980 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__einvn_8  ring.dstage\[10\].id.delayenb0
timestamp 1635306529
transform 1 0 6348 0 1 21760
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_6  FILLER_36_75
timestamp 1635306529
transform 1 0 8004 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1635306529
transform -1 0 8832 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_15
timestamp 1635306529
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_3
timestamp 1635306529
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1635306529
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.dstage\[10\].id.delayen1_TE
timestamp 1635306529
transform -1 0 5244 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_27
timestamp 1635306529
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_39
timestamp 1635306529
transform 1 0 4692 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_45
timestamp 1635306529
transform 1 0 5244 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_52
timestamp 1635306529
transform 1 0 5888 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_57
timestamp 1635306529
transform 1 0 6348 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_61
timestamp 1635306529
transform 1 0 6716 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1635306529
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__einvp_2  ring.dstage\[10\].id.delayen1
timestamp 1635306529
transform -1 0 7452 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_1  ring.dstage\[10\].id.delayint0
timestamp 1635306529
transform -1 0 5888 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_69
timestamp 1635306529
transform 1 0 7452 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_77
timestamp 1635306529
transform 1 0 8188 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1635306529
transform -1 0 8832 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ring.dstage\[10\].id.delaybuf0
timestamp 1635306529
transform -1 0 8188 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_15
timestamp 1635306529
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_3
timestamp 1635306529
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1635306529
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1635306529
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_29
timestamp 1635306529
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_41
timestamp 1635306529
transform 1 0 4876 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1635306529
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.dstage\[10\].id.delayenb1_TE_B
timestamp 1635306529
transform 1 0 5520 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_47
timestamp 1635306529
transform 1 0 5428 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_50
timestamp 1635306529
transform 1 0 5704 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_57
timestamp 1635306529
transform 1 0 6348 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ring.dstage\[10\].id.delaybuf1
timestamp 1635306529
transform -1 0 6348 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__einvn_4  ring.dstage\[10\].id.delayenb1
timestamp 1635306529
transform -1 0 7728 0 1 22848
box -38 -48 1050 592
use sky130_fd_sc_hd__decap_8  FILLER_38_72
timestamp 1635306529
transform 1 0 7728 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_80
timestamp 1635306529
transform 1 0 8464 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1635306529
transform -1 0 8832 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_39_15
timestamp 1635306529
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_3
timestamp 1635306529
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_15
timestamp 1635306529
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_3
timestamp 1635306529
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1635306529
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1635306529
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_39_27
timestamp 1635306529
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_39
timestamp 1635306529
transform 1 0 4692 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1635306529
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_29
timestamp 1635306529
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_41
timestamp 1635306529
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1635306529
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_39_47
timestamp 1635306529
transform 1 0 5428 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_52
timestamp 1635306529
transform 1 0 5888 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.dstage\[8\].id.delayenb1_TE_B
timestamp 1635306529
transform 1 0 5980 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.dstage\[8\].id.delayen1_TE
timestamp 1635306529
transform -1 0 5888 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1635306529
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_55
timestamp 1635306529
transform 1 0 6164 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_57
timestamp 1635306529
transform 1 0 6348 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ring.dstage\[8\].id.delaybuf1
timestamp 1635306529
transform -1 0 6808 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ring.dstage\[8\].id.delaybuf0
timestamp 1635306529
transform -1 0 7176 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_62
timestamp 1635306529
transform 1 0 6808 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_61
timestamp 1635306529
transform 1 0 6716 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_66
timestamp 1635306529
transform 1 0 7176 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_77
timestamp 1635306529
transform 1 0 8188 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_77
timestamp 1635306529
transform 1 0 8188 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1635306529
transform -1 0 8832 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1635306529
transform -1 0 8832 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ring.dstage\[8\].id.delayen1
timestamp 1635306529
transform -1 0 8188 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_4  ring.dstage\[8\].id.delayenb1
timestamp 1635306529
transform -1 0 8188 0 1 23936
box -38 -48 1050 592
use sky130_fd_sc_hd__decap_12  FILLER_41_15
timestamp 1635306529
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_3
timestamp 1635306529
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1635306529
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_27
timestamp 1635306529
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_39
timestamp 1635306529
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.dstage\[8\].id.delayen0_TE
timestamp 1635306529
transform 1 0 6348 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1635306529
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1635306529
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_59
timestamp 1635306529
transform 1 0 6532 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1635306529
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_1  ring.dstage\[8\].id.delayint0
timestamp 1635306529
transform -1 0 7176 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_66
timestamp 1635306529
transform 1 0 7176 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_77
timestamp 1635306529
transform 1 0 8188 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1635306529
transform -1 0 8832 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ring.dstage\[8\].id.delayen0
timestamp 1635306529
transform -1 0 8188 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_42_15
timestamp 1635306529
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_3
timestamp 1635306529
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1635306529
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1635306529
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_29
timestamp 1635306529
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_41
timestamp 1635306529
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1635306529
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.dstage\[8\].id.delayenb0_TE_B
timestamp 1635306529
transform -1 0 6164 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_55
timestamp 1635306529
transform 1 0 6164 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__einvn_8  ring.dstage\[8\].id.delayenb0
timestamp 1635306529
transform -1 0 8188 0 1 25024
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_4  FILLER_42_77
timestamp 1635306529
transform 1 0 8188 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1635306529
transform -1 0 8832 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_43_15
timestamp 1635306529
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_3
timestamp 1635306529
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1635306529
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_43_27
timestamp 1635306529
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_39
timestamp 1635306529
transform 1 0 4692 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.dstage\[9\].id.delayenb1_TE_B
timestamp 1635306529
transform -1 0 5888 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_43_47
timestamp 1635306529
transform 1 0 5428 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_52
timestamp 1635306529
transform 1 0 5888 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_57
timestamp 1635306529
transform 1 0 6348 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_61
timestamp 1635306529
transform 1 0 6716 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1635306529
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__einvn_4  ring.dstage\[9\].id.delayenb1
timestamp 1635306529
transform -1 0 7820 0 -1 26112
box -38 -48 1050 592
use sky130_fd_sc_hd__decap_8  FILLER_43_73
timestamp 1635306529
transform 1 0 7820 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1635306529
transform -1 0 8832 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_44_15
timestamp 1635306529
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_3
timestamp 1635306529
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1635306529
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1635306529
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_29
timestamp 1635306529
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_44_41
timestamp 1635306529
transform 1 0 4876 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1635306529
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_47
timestamp 1635306529
transform 1 0 5428 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_55
timestamp 1635306529
transform 1 0 6164 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  ring.dstage\[9\].id.delaybuf0
timestamp 1635306529
transform 1 0 5796 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__einvn_8  ring.dstage\[9\].id.delayenb0
timestamp 1635306529
transform -1 0 8188 0 1 26112
box -38 -48 1694 592
use sky130_fd_sc_hd__clkinv_1  ring.dstage\[9\].id.delayint0
timestamp 1635306529
transform -1 0 5428 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_77
timestamp 1635306529
transform 1 0 8188 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1635306529
transform -1 0 8832 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_45_15
timestamp 1635306529
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_3
timestamp 1635306529
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1635306529
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_45_27
timestamp 1635306529
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_39
timestamp 1635306529
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1635306529
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1635306529
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_60
timestamp 1635306529
transform 1 0 6624 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1635306529
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  ring.dstage\[9\].id.delaybuf1
timestamp 1635306529
transform -1 0 6624 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ring.dstage\[9\].id.delayen0
timestamp 1635306529
transform -1 0 7636 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.dstage\[9\].id.delayen0_TE
timestamp 1635306529
transform 1 0 8004 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_71
timestamp 1635306529
transform 1 0 7636 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_77
timestamp 1635306529
transform 1 0 8188 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1635306529
transform -1 0 8832 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_46_15
timestamp 1635306529
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_3
timestamp 1635306529
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1635306529
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1635306529
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_29
timestamp 1635306529
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_41
timestamp 1635306529
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1635306529
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.dstage\[9\].id.delayenb0_TE_B
timestamp 1635306529
transform -1 0 6624 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_46_53
timestamp 1635306529
transform 1 0 5980 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_46_57
timestamp 1635306529
transform 1 0 6348 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_60
timestamp 1635306529
transform 1 0 6624 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1635306529
transform 1 0 6256 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__einvp_2  ring.dstage\[9\].id.delayen1
timestamp 1635306529
transform -1 0 7636 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.dstage\[9\].id.delayen1_TE
timestamp 1635306529
transform -1 0 8188 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_71
timestamp 1635306529
transform 1 0 7636 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_77
timestamp 1635306529
transform 1 0 8188 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1635306529
transform -1 0 8832 0 1 27200
box -38 -48 314 592
<< labels >>
rlabel metal2 s 6918 0 6974 800 6 clk_out
port 0 nsew signal tristate
rlabel metal2 s 938 0 994 800 6 clkmux[0]
port 1 nsew signal input
rlabel metal2 s 2870 0 2926 800 6 clkmux[1]
port 2 nsew signal input
rlabel metal2 s 4894 0 4950 800 6 clkmux[2]
port 3 nsew signal input
rlabel metal2 s 8942 0 8998 800 6 start
port 4 nsew signal input
rlabel metal3 s 9200 552 10000 672 6 trim_a[0]
port 5 nsew signal input
rlabel metal3 s 9200 12112 10000 12232 6 trim_a[10]
port 6 nsew signal input
rlabel metal3 s 9200 13200 10000 13320 6 trim_a[11]
port 7 nsew signal input
rlabel metal3 s 9200 14424 10000 14544 6 trim_a[12]
port 8 nsew signal input
rlabel metal3 s 9200 15512 10000 15632 6 trim_a[13]
port 9 nsew signal input
rlabel metal3 s 9200 16736 10000 16856 6 trim_a[14]
port 10 nsew signal input
rlabel metal3 s 9200 17824 10000 17944 6 trim_a[15]
port 11 nsew signal input
rlabel metal3 s 9200 19048 10000 19168 6 trim_a[16]
port 12 nsew signal input
rlabel metal3 s 9200 20136 10000 20256 6 trim_a[17]
port 13 nsew signal input
rlabel metal3 s 9200 21360 10000 21480 6 trim_a[18]
port 14 nsew signal input
rlabel metal3 s 9200 22448 10000 22568 6 trim_a[19]
port 15 nsew signal input
rlabel metal3 s 9200 1640 10000 1760 6 trim_a[1]
port 16 nsew signal input
rlabel metal3 s 9200 23672 10000 23792 6 trim_a[20]
port 17 nsew signal input
rlabel metal3 s 9200 24760 10000 24880 6 trim_a[21]
port 18 nsew signal input
rlabel metal3 s 9200 25984 10000 26104 6 trim_a[22]
port 19 nsew signal input
rlabel metal3 s 9200 27072 10000 27192 6 trim_a[23]
port 20 nsew signal input
rlabel metal3 s 9200 28296 10000 28416 6 trim_a[24]
port 21 nsew signal input
rlabel metal3 s 9200 29384 10000 29504 6 trim_a[25]
port 22 nsew signal input
rlabel metal3 s 9200 2864 10000 2984 6 trim_a[2]
port 23 nsew signal input
rlabel metal3 s 9200 3952 10000 4072 6 trim_a[3]
port 24 nsew signal input
rlabel metal3 s 9200 5176 10000 5296 6 trim_a[4]
port 25 nsew signal input
rlabel metal3 s 9200 6264 10000 6384 6 trim_a[5]
port 26 nsew signal input
rlabel metal3 s 9200 7488 10000 7608 6 trim_a[6]
port 27 nsew signal input
rlabel metal3 s 9200 8576 10000 8696 6 trim_a[7]
port 28 nsew signal input
rlabel metal3 s 9200 9800 10000 9920 6 trim_a[8]
port 29 nsew signal input
rlabel metal3 s 9200 10888 10000 11008 6 trim_a[9]
port 30 nsew signal input
rlabel metal4 s 2243 2128 2563 27792 6 vccd1
port 31 nsew power input
rlabel metal4 s 4840 2128 5160 27792 6 vccd1
port 31 nsew power input
rlabel metal4 s 7437 2128 7757 27792 6 vccd1
port 31 nsew power input
rlabel metal4 s 3541 2128 3861 27792 6 vssd1
port 32 nsew ground input
rlabel metal4 s 6138 2128 6458 27792 6 vssd1
port 32 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 10000 30000
<< end >>
