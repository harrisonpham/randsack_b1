magic
tech sky130A
magscale 1 2
timestamp 1635110680
<< locali >>
rect 5181 8279 5215 8585
rect 3801 6715 3835 6953
<< viali >>
rect 3249 27557 3283 27591
rect 2145 27489 2179 27523
rect 4997 27489 5031 27523
rect 3801 27421 3835 27455
rect 7297 27421 7331 27455
rect 7849 27421 7883 27455
rect 4445 27353 4479 27387
rect 4537 27353 4571 27387
rect 5733 27353 5767 27387
rect 6745 27353 6779 27387
rect 7389 27353 7423 27387
rect 2697 27285 2731 27319
rect 3985 27285 4019 27319
rect 5641 27285 5675 27319
rect 6653 27285 6687 27319
rect 2053 27081 2087 27115
rect 3893 27081 3927 27115
rect 6653 27013 6687 27047
rect 3249 26945 3283 26979
rect 4353 26945 4387 26979
rect 4537 26945 4571 26979
rect 5273 26945 5307 26979
rect 7113 26945 7147 26979
rect 3801 26877 3835 26911
rect 6561 26877 6595 26911
rect 7573 26877 7607 26911
rect 8125 26877 8159 26911
rect 7665 26809 7699 26843
rect 2605 26741 2639 26775
rect 3157 26741 3191 26775
rect 5825 26741 5859 26775
rect 2605 26537 2639 26571
rect 2053 26469 2087 26503
rect 4077 26469 4111 26503
rect 6469 26469 6503 26503
rect 3985 26401 4019 26435
rect 3065 26333 3099 26367
rect 4537 26333 4571 26367
rect 5181 26333 5215 26367
rect 5917 26333 5951 26367
rect 6469 26333 6503 26367
rect 7941 26333 7975 26367
rect 4997 26265 5031 26299
rect 3249 26197 3283 26231
rect 1777 25993 1811 26027
rect 6469 25993 6503 26027
rect 2329 25925 2363 25959
rect 3801 25925 3835 25959
rect 7021 25925 7055 25959
rect 7297 25925 7331 25959
rect 2881 25857 2915 25891
rect 3065 25857 3099 25891
rect 3617 25857 3651 25891
rect 4261 25857 4295 25891
rect 5273 25857 5307 25891
rect 6561 25857 6595 25891
rect 7941 25857 7975 25891
rect 5549 25721 5583 25755
rect 2053 25449 2087 25483
rect 5273 25381 5307 25415
rect 6837 25381 6871 25415
rect 5181 25313 5215 25347
rect 5733 25313 5767 25347
rect 2605 25245 2639 25279
rect 3249 25245 3283 25279
rect 4721 25245 4755 25279
rect 7205 25245 7239 25279
rect 8125 25245 8159 25279
rect 3157 25177 3191 25211
rect 4169 25177 4203 25211
rect 4261 25177 4295 25211
rect 3433 24769 3467 24803
rect 4169 24769 4203 24803
rect 5641 24769 5675 24803
rect 6377 24769 6411 24803
rect 6561 24769 6595 24803
rect 7297 24769 7331 24803
rect 8033 24769 8067 24803
rect 1869 24701 1903 24735
rect 2421 24701 2455 24735
rect 3617 24633 3651 24667
rect 4169 24633 4203 24667
rect 7849 24633 7883 24667
rect 2973 24565 3007 24599
rect 4629 24293 4663 24327
rect 7665 24293 7699 24327
rect 5549 24225 5583 24259
rect 8125 24225 8159 24259
rect 4077 24157 4111 24191
rect 5089 24157 5123 24191
rect 5641 24157 5675 24191
rect 7113 24157 7147 24191
rect 2697 24089 2731 24123
rect 4537 24089 4571 24123
rect 7573 24089 7607 24123
rect 2145 24021 2179 24055
rect 3249 24021 3283 24055
rect 3985 24021 4019 24055
rect 4169 23817 4203 23851
rect 4813 23817 4847 23851
rect 5273 23749 5307 23783
rect 5365 23749 5399 23783
rect 6469 23749 6503 23783
rect 7205 23749 7239 23783
rect 7389 23749 7423 23783
rect 3985 23681 4019 23715
rect 4629 23681 4663 23715
rect 6653 23681 6687 23715
rect 8125 23681 8159 23715
rect 5825 23613 5859 23647
rect 3525 23545 3559 23579
rect 2973 23477 3007 23511
rect 3893 23273 3927 23307
rect 7205 23205 7239 23239
rect 4445 23137 4479 23171
rect 7113 23137 7147 23171
rect 2697 23069 2731 23103
rect 5549 23069 5583 23103
rect 6653 23069 6687 23103
rect 7665 23069 7699 23103
rect 4997 23001 5031 23035
rect 5089 23001 5123 23035
rect 6101 23001 6135 23035
rect 6193 23001 6227 23035
rect 3249 22933 3283 22967
rect 4537 22933 4571 22967
rect 3065 22729 3099 22763
rect 3709 22729 3743 22763
rect 4261 22661 4295 22695
rect 3525 22593 3559 22627
rect 7205 22593 7239 22627
rect 8125 22593 8159 22627
rect 4905 22525 4939 22559
rect 5457 22525 5491 22559
rect 4445 22457 4479 22491
rect 4997 22457 5031 22491
rect 6653 22457 6687 22491
rect 2513 22389 2547 22423
rect 3249 22185 3283 22219
rect 2697 22117 2731 22151
rect 4721 22117 4755 22151
rect 3893 22049 3927 22083
rect 4905 21981 4939 22015
rect 6009 21981 6043 22015
rect 7021 21981 7055 22015
rect 7757 21981 7791 22015
rect 6837 21913 6871 21947
rect 3985 21845 4019 21879
rect 2605 21641 2639 21675
rect 4445 21641 4479 21675
rect 4905 21573 4939 21607
rect 5089 21573 5123 21607
rect 4261 21505 4295 21539
rect 5825 21505 5859 21539
rect 6469 21505 6503 21539
rect 7573 21437 7607 21471
rect 8125 21437 8159 21471
rect 6653 21369 6687 21403
rect 7665 21369 7699 21403
rect 3157 21301 3191 21335
rect 3801 21301 3835 21335
rect 3249 21097 3283 21131
rect 4353 21029 4387 21063
rect 7849 21029 7883 21063
rect 5549 20961 5583 20995
rect 6101 20961 6135 20995
rect 4169 20893 4203 20927
rect 4997 20893 5031 20927
rect 6561 20893 6595 20927
rect 7481 20893 7515 20927
rect 5641 20825 5675 20859
rect 2605 20757 2639 20791
rect 4905 20757 4939 20791
rect 3157 20553 3191 20587
rect 4445 20485 4479 20519
rect 5181 20485 5215 20519
rect 2973 20417 3007 20451
rect 3801 20417 3835 20451
rect 4905 20417 4939 20451
rect 5825 20417 5859 20451
rect 6653 20417 6687 20451
rect 7941 20417 7975 20451
rect 6469 20281 6503 20315
rect 2513 20213 2547 20247
rect 3709 20213 3743 20247
rect 4353 20213 4387 20247
rect 2697 20009 2731 20043
rect 4261 20009 4295 20043
rect 6469 19873 6503 19907
rect 3249 19805 3283 19839
rect 4905 19805 4939 19839
rect 5825 19805 5859 19839
rect 7205 19805 7239 19839
rect 7389 19805 7423 19839
rect 8125 19805 8159 19839
rect 4353 19737 4387 19771
rect 1593 19669 1627 19703
rect 2053 19669 2087 19703
rect 2973 19465 3007 19499
rect 4077 19465 4111 19499
rect 6469 19397 6503 19431
rect 7573 19397 7607 19431
rect 4169 19329 4203 19363
rect 4813 19329 4847 19363
rect 5273 19329 5307 19363
rect 8125 19329 8159 19363
rect 2421 19261 2455 19295
rect 4721 19261 4755 19295
rect 6377 19261 6411 19295
rect 6929 19261 6963 19295
rect 7665 19261 7699 19295
rect 1869 19193 1903 19227
rect 3525 19193 3559 19227
rect 5825 19125 5859 19159
rect 2697 18921 2731 18955
rect 3249 18853 3283 18887
rect 4445 18853 4479 18887
rect 6561 18853 6595 18887
rect 6469 18785 6503 18819
rect 8125 18785 8159 18819
rect 4445 18717 4479 18751
rect 5733 18717 5767 18751
rect 7021 18717 7055 18751
rect 7665 18717 7699 18751
rect 1593 18649 1627 18683
rect 7573 18649 7607 18683
rect 2145 18581 2179 18615
rect 3801 18377 3835 18411
rect 3893 18309 3927 18343
rect 4537 18309 4571 18343
rect 7573 18309 7607 18343
rect 3249 18241 3283 18275
rect 4353 18241 4387 18275
rect 5273 18241 5307 18275
rect 6929 18241 6963 18275
rect 8125 18241 8159 18275
rect 6377 18173 6411 18207
rect 7665 18173 7699 18207
rect 6469 18105 6503 18139
rect 1501 18037 1535 18071
rect 2053 18037 2087 18071
rect 2605 18037 2639 18071
rect 3157 18037 3191 18071
rect 5825 18037 5859 18071
rect 2605 17833 2639 17867
rect 3249 17833 3283 17867
rect 2145 17765 2179 17799
rect 6837 17765 6871 17799
rect 4629 17697 4663 17731
rect 4169 17629 4203 17663
rect 4721 17629 4755 17663
rect 5365 17629 5399 17663
rect 6101 17629 6135 17663
rect 7205 17629 7239 17663
rect 8125 17629 8159 17663
rect 5181 17561 5215 17595
rect 1593 17493 1627 17527
rect 1685 17289 1719 17323
rect 4813 17289 4847 17323
rect 5365 17221 5399 17255
rect 6561 17221 6595 17255
rect 2881 17153 2915 17187
rect 3341 17153 3375 17187
rect 3985 17153 4019 17187
rect 4629 17153 4663 17187
rect 6377 17153 6411 17187
rect 7297 17153 7331 17187
rect 7941 17153 7975 17187
rect 2789 17085 2823 17119
rect 5273 17085 5307 17119
rect 5825 17085 5859 17119
rect 2237 17017 2271 17051
rect 3525 17017 3559 17051
rect 7757 17017 7791 17051
rect 4169 16949 4203 16983
rect 2605 16745 2639 16779
rect 1501 16677 1535 16711
rect 3065 16541 3099 16575
rect 4261 16541 4295 16575
rect 4445 16541 4479 16575
rect 4997 16541 5031 16575
rect 5457 16541 5491 16575
rect 6193 16541 6227 16575
rect 7113 16541 7147 16575
rect 4905 16473 4939 16507
rect 7757 16473 7791 16507
rect 2053 16405 2087 16439
rect 3249 16405 3283 16439
rect 2605 16201 2639 16235
rect 3249 16201 3283 16235
rect 3893 16201 3927 16235
rect 6377 16133 6411 16167
rect 7205 16133 7239 16167
rect 7389 16133 7423 16167
rect 3709 16065 3743 16099
rect 4537 16065 4571 16099
rect 5089 16065 5123 16099
rect 6561 16065 6595 16099
rect 8125 16065 8159 16099
rect 4445 15997 4479 16031
rect 4997 15997 5031 16031
rect 5549 15997 5583 16031
rect 1593 15861 1627 15895
rect 2145 15861 2179 15895
rect 2697 15657 2731 15691
rect 3249 15657 3283 15691
rect 7481 15589 7515 15623
rect 7389 15521 7423 15555
rect 7941 15521 7975 15555
rect 4721 15453 4755 15487
rect 5917 15453 5951 15487
rect 6929 15453 6963 15487
rect 4353 15385 4387 15419
rect 6377 15385 6411 15419
rect 6469 15385 6503 15419
rect 1593 15317 1627 15351
rect 2145 15317 2179 15351
rect 3893 15317 3927 15351
rect 3065 15113 3099 15147
rect 4905 15045 4939 15079
rect 4077 14977 4111 15011
rect 4721 14977 4755 15011
rect 5641 14977 5675 15011
rect 6469 14977 6503 15011
rect 7941 14977 7975 15011
rect 6377 14909 6411 14943
rect 1869 14773 1903 14807
rect 2513 14773 2547 14807
rect 3617 14773 3651 14807
rect 4261 14773 4295 14807
rect 3249 14501 3283 14535
rect 5089 14433 5123 14467
rect 5181 14433 5215 14467
rect 3893 14365 3927 14399
rect 4537 14365 4571 14399
rect 5641 14365 5675 14399
rect 6101 14365 6135 14399
rect 6285 14365 6319 14399
rect 7021 14365 7055 14399
rect 8125 14365 8159 14399
rect 2145 14297 2179 14331
rect 7573 14297 7607 14331
rect 7665 14297 7699 14331
rect 1593 14229 1627 14263
rect 2697 14229 2731 14263
rect 4445 14229 4479 14263
rect 3709 14025 3743 14059
rect 4353 14025 4387 14059
rect 4261 13957 4295 13991
rect 5733 13957 5767 13991
rect 6561 13957 6595 13991
rect 1501 13889 1535 13923
rect 3065 13889 3099 13923
rect 4813 13889 4847 13923
rect 4997 13889 5031 13923
rect 7021 13889 7055 13923
rect 8125 13889 8159 13923
rect 5549 13821 5583 13855
rect 1961 13685 1995 13719
rect 2605 13685 2639 13719
rect 2145 13481 2179 13515
rect 3249 13413 3283 13447
rect 3801 13277 3835 13311
rect 4997 13277 5031 13311
rect 5457 13277 5491 13311
rect 6377 13277 6411 13311
rect 7205 13277 7239 13311
rect 8125 13277 8159 13311
rect 4445 13209 4479 13243
rect 4537 13209 4571 13243
rect 5733 13209 5767 13243
rect 7389 13209 7423 13243
rect 1593 13141 1627 13175
rect 2697 13141 2731 13175
rect 3985 13141 4019 13175
rect 1777 12937 1811 12971
rect 2421 12937 2455 12971
rect 5733 12937 5767 12971
rect 3065 12869 3099 12903
rect 4445 12869 4479 12903
rect 5825 12869 5859 12903
rect 7665 12869 7699 12903
rect 2237 12801 2271 12835
rect 3709 12801 3743 12835
rect 4261 12801 4295 12835
rect 5181 12801 5215 12835
rect 7573 12801 7607 12835
rect 8125 12801 8159 12835
rect 3525 12733 3559 12767
rect 6561 12733 6595 12767
rect 7113 12733 7147 12767
rect 2973 12665 3007 12699
rect 6653 12665 6687 12699
rect 3249 12393 3283 12427
rect 4721 12325 4755 12359
rect 6469 12257 6503 12291
rect 2421 12189 2455 12223
rect 3065 12189 3099 12223
rect 5089 12189 5123 12223
rect 6009 12189 6043 12223
rect 6561 12189 6595 12223
rect 8033 12189 8067 12223
rect 1961 12053 1995 12087
rect 2605 12053 2639 12087
rect 3893 12053 3927 12087
rect 3985 12053 4019 12087
rect 6377 11849 6411 11883
rect 3433 11781 3467 11815
rect 6929 11781 6963 11815
rect 7113 11781 7147 11815
rect 4261 11713 4295 11747
rect 5457 11713 5491 11747
rect 7849 11713 7883 11747
rect 2789 11645 2823 11679
rect 4169 11577 4203 11611
rect 1685 11509 1719 11543
rect 2145 11509 2179 11543
rect 3341 11509 3375 11543
rect 3249 11305 3283 11339
rect 7941 11305 7975 11339
rect 4445 11237 4479 11271
rect 6929 11237 6963 11271
rect 3893 11169 3927 11203
rect 4353 11169 4387 11203
rect 5457 11169 5491 11203
rect 6837 11169 6871 11203
rect 1593 11101 1627 11135
rect 4905 11101 4939 11135
rect 6009 11101 6043 11135
rect 7389 11101 7423 11135
rect 2697 11033 2731 11067
rect 5549 11033 5583 11067
rect 8033 11033 8067 11067
rect 2145 10965 2179 10999
rect 2329 10761 2363 10795
rect 4629 10761 4663 10795
rect 4077 10693 4111 10727
rect 6469 10693 6503 10727
rect 4721 10625 4755 10659
rect 6377 10625 6411 10659
rect 6929 10625 6963 10659
rect 5273 10557 5307 10591
rect 5825 10557 5859 10591
rect 7573 10557 7607 10591
rect 8125 10557 8159 10591
rect 3341 10489 3375 10523
rect 5365 10489 5399 10523
rect 7665 10489 7699 10523
rect 1777 10421 1811 10455
rect 2881 10421 2915 10455
rect 3985 10421 4019 10455
rect 5365 10217 5399 10251
rect 3157 10149 3191 10183
rect 7297 10081 7331 10115
rect 2605 10013 2639 10047
rect 4077 10013 4111 10047
rect 4905 10013 4939 10047
rect 5181 10013 5215 10047
rect 6101 10013 6135 10047
rect 6837 10013 6871 10047
rect 7849 10013 7883 10047
rect 2053 9945 2087 9979
rect 4261 9945 4295 9979
rect 5917 9945 5951 9979
rect 7389 9945 7423 9979
rect 1501 9877 1535 9911
rect 3249 9877 3283 9911
rect 4353 9673 4387 9707
rect 3249 9605 3283 9639
rect 6377 9605 6411 9639
rect 2421 9537 2455 9571
rect 4997 9537 5031 9571
rect 5549 9537 5583 9571
rect 6469 9537 6503 9571
rect 7941 9537 7975 9571
rect 4261 9469 4295 9503
rect 4445 9469 4479 9503
rect 5365 9469 5399 9503
rect 2605 9401 2639 9435
rect 3065 9401 3099 9435
rect 1961 9333 1995 9367
rect 3893 9333 3927 9367
rect 2053 9129 2087 9163
rect 4169 9129 4203 9163
rect 3249 9061 3283 9095
rect 5641 9061 5675 9095
rect 7849 9061 7883 9095
rect 5549 8993 5583 9027
rect 6101 8993 6135 9027
rect 3065 8925 3099 8959
rect 4261 8925 4295 8959
rect 4997 8925 5031 8959
rect 6561 8925 6595 8959
rect 7481 8925 7515 8959
rect 1501 8789 1535 8823
rect 2513 8789 2547 8823
rect 4905 8789 4939 8823
rect 1501 8585 1535 8619
rect 3157 8585 3191 8619
rect 5181 8585 5215 8619
rect 3801 8517 3835 8551
rect 3249 8449 3283 8483
rect 2053 8381 2087 8415
rect 4537 8381 4571 8415
rect 2605 8313 2639 8347
rect 6377 8517 6411 8551
rect 7205 8517 7239 8551
rect 7389 8517 7423 8551
rect 5273 8449 5307 8483
rect 6561 8449 6595 8483
rect 8125 8449 8159 8483
rect 5825 8381 5859 8415
rect 5365 8313 5399 8347
rect 5181 8245 5215 8279
rect 1961 8041 1995 8075
rect 5641 7905 5675 7939
rect 2421 7837 2455 7871
rect 3065 7837 3099 7871
rect 4905 7837 4939 7871
rect 5733 7837 5767 7871
rect 6193 7837 6227 7871
rect 7665 7837 7699 7871
rect 4353 7769 4387 7803
rect 4445 7769 4479 7803
rect 6745 7769 6779 7803
rect 6929 7769 6963 7803
rect 2605 7701 2639 7735
rect 3249 7701 3283 7735
rect 3893 7701 3927 7735
rect 2053 7497 2087 7531
rect 3249 7429 3283 7463
rect 3341 7429 3375 7463
rect 4261 7429 4295 7463
rect 4445 7429 4479 7463
rect 5641 7429 5675 7463
rect 6377 7429 6411 7463
rect 2697 7361 2731 7395
rect 5181 7361 5215 7395
rect 6745 7361 6779 7395
rect 7941 7361 7975 7395
rect 1961 7293 1995 7327
rect 3801 7293 3835 7327
rect 2513 7225 2547 7259
rect 5733 7157 5767 7191
rect 1501 6953 1535 6987
rect 3801 6953 3835 6987
rect 3157 6885 3191 6919
rect 3249 6817 3283 6851
rect 1593 6749 1627 6783
rect 2053 6749 2087 6783
rect 2697 6749 2731 6783
rect 4261 6885 4295 6919
rect 6101 6885 6135 6919
rect 4261 6749 4295 6783
rect 5549 6749 5583 6783
rect 6193 6749 6227 6783
rect 7573 6749 7607 6783
rect 3801 6681 3835 6715
rect 2237 6613 2271 6647
rect 8033 6613 8067 6647
rect 2237 6409 2271 6443
rect 4997 6341 5031 6375
rect 1409 6273 1443 6307
rect 4270 6273 4304 6307
rect 6653 6273 6687 6307
rect 8125 6273 8159 6307
rect 2789 6205 2823 6239
rect 4537 6205 4571 6239
rect 5089 6205 5123 6239
rect 5549 6205 5583 6239
rect 6653 6137 6687 6171
rect 1593 6069 1627 6103
rect 2145 6069 2179 6103
rect 3157 6069 3191 6103
rect 2513 5865 2547 5899
rect 1869 5797 1903 5831
rect 4261 5729 4295 5763
rect 4813 5729 4847 5763
rect 1685 5661 1719 5695
rect 2329 5661 2363 5695
rect 3157 5661 3191 5695
rect 5457 5661 5491 5695
rect 6193 5661 6227 5695
rect 7205 5661 7239 5695
rect 8119 5661 8153 5695
rect 4353 5593 4387 5627
rect 5273 5593 5307 5627
rect 7389 5593 7423 5627
rect 3065 5525 3099 5559
rect 6745 5525 6779 5559
rect 5089 5321 5123 5355
rect 7389 5253 7423 5287
rect 1676 5185 1710 5219
rect 3976 5185 4010 5219
rect 7941 5185 7975 5219
rect 1409 5117 1443 5151
rect 3157 5117 3191 5151
rect 3709 5117 3743 5151
rect 5457 5117 5491 5151
rect 6377 5117 6411 5151
rect 6929 5117 6963 5151
rect 6469 5049 6503 5083
rect 7481 5049 7515 5083
rect 2789 4981 2823 5015
rect 1685 4777 1719 4811
rect 2237 4641 2271 4675
rect 7389 4641 7423 4675
rect 1777 4573 1811 4607
rect 2421 4573 2455 4607
rect 4353 4573 4387 4607
rect 5365 4573 5399 4607
rect 6101 4573 6135 4607
rect 6837 4573 6871 4607
rect 7849 4573 7883 4607
rect 3157 4505 3191 4539
rect 3801 4505 3835 4539
rect 3893 4505 3927 4539
rect 4813 4505 4847 4539
rect 4905 4505 4939 4539
rect 5917 4505 5951 4539
rect 7297 4505 7331 4539
rect 3065 4437 3099 4471
rect 1685 4233 1719 4267
rect 1593 4165 1627 4199
rect 2412 4097 2446 4131
rect 4445 4097 4479 4131
rect 4629 4097 4663 4131
rect 5365 4097 5399 4131
rect 6469 4097 6503 4131
rect 7941 4097 7975 4131
rect 2145 4029 2179 4063
rect 3893 4029 3927 4063
rect 6469 3961 6503 3995
rect 3525 3893 3559 3927
rect 1869 3689 1903 3723
rect 4353 3621 4387 3655
rect 1501 3553 1535 3587
rect 3249 3553 3283 3587
rect 2982 3485 3016 3519
rect 4445 3485 4479 3519
rect 5825 3485 5859 3519
rect 6653 3485 6687 3519
rect 8125 3485 8159 3519
rect 6561 3417 6595 3451
rect 6377 3145 6411 3179
rect 1869 3077 1903 3111
rect 2053 3077 2087 3111
rect 6929 3077 6963 3111
rect 7205 3077 7239 3111
rect 2605 3009 2639 3043
rect 2872 3009 2906 3043
rect 4905 3009 4939 3043
rect 7849 3009 7883 3043
rect 4353 2941 4387 2975
rect 5733 2941 5767 2975
rect 3985 2805 4019 2839
rect 2513 2601 2547 2635
rect 5273 2601 5307 2635
rect 6653 2533 6687 2567
rect 7665 2533 7699 2567
rect 1777 2465 1811 2499
rect 6561 2465 6595 2499
rect 7113 2465 7147 2499
rect 8125 2465 8159 2499
rect 2329 2397 2363 2431
rect 4353 2397 4387 2431
rect 4721 2397 4755 2431
rect 3065 2329 3099 2363
rect 3985 2329 4019 2363
rect 4261 2329 4295 2363
rect 5089 2329 5123 2363
rect 7573 2329 7607 2363
rect 1869 2261 1903 2295
rect 3157 2261 3191 2295
<< metal1 >>
rect 1104 27770 8832 27792
rect 1104 27718 2248 27770
rect 2300 27718 2312 27770
rect 2364 27718 2376 27770
rect 2428 27718 2440 27770
rect 2492 27718 2504 27770
rect 2556 27718 4846 27770
rect 4898 27718 4910 27770
rect 4962 27718 4974 27770
rect 5026 27718 5038 27770
rect 5090 27718 5102 27770
rect 5154 27718 7443 27770
rect 7495 27718 7507 27770
rect 7559 27718 7571 27770
rect 7623 27718 7635 27770
rect 7687 27718 7699 27770
rect 7751 27718 8832 27770
rect 1104 27696 8832 27718
rect 2590 27548 2596 27600
rect 2648 27588 2654 27600
rect 3237 27591 3295 27597
rect 3237 27588 3249 27591
rect 2648 27560 3249 27588
rect 2648 27548 2654 27560
rect 3237 27557 3249 27560
rect 3283 27588 3295 27591
rect 5810 27588 5816 27600
rect 3283 27560 5816 27588
rect 3283 27557 3295 27560
rect 3237 27551 3295 27557
rect 5810 27548 5816 27560
rect 5868 27548 5874 27600
rect 2038 27480 2044 27532
rect 2096 27520 2102 27532
rect 2133 27523 2191 27529
rect 2133 27520 2145 27523
rect 2096 27492 2145 27520
rect 2096 27480 2102 27492
rect 2133 27489 2145 27492
rect 2179 27520 2191 27523
rect 4985 27523 5043 27529
rect 4985 27520 4997 27523
rect 2179 27492 4997 27520
rect 2179 27489 2191 27492
rect 2133 27483 2191 27489
rect 4985 27489 4997 27492
rect 5031 27520 5043 27523
rect 5534 27520 5540 27532
rect 5031 27492 5540 27520
rect 5031 27489 5043 27492
rect 4985 27483 5043 27489
rect 5534 27480 5540 27492
rect 5592 27480 5598 27532
rect 3789 27455 3847 27461
rect 3789 27421 3801 27455
rect 3835 27452 3847 27455
rect 4062 27452 4068 27464
rect 3835 27424 4068 27452
rect 3835 27421 3847 27424
rect 3789 27415 3847 27421
rect 4062 27412 4068 27424
rect 4120 27412 4126 27464
rect 4154 27412 4160 27464
rect 4212 27452 4218 27464
rect 7285 27455 7343 27461
rect 7285 27452 7297 27455
rect 4212 27424 7297 27452
rect 4212 27412 4218 27424
rect 7285 27421 7297 27424
rect 7331 27421 7343 27455
rect 7834 27452 7840 27464
rect 7795 27424 7840 27452
rect 7285 27415 7343 27421
rect 7834 27412 7840 27424
rect 7892 27412 7898 27464
rect 3878 27344 3884 27396
rect 3936 27384 3942 27396
rect 4433 27387 4491 27393
rect 4433 27384 4445 27387
rect 3936 27356 4445 27384
rect 3936 27344 3942 27356
rect 4433 27353 4445 27356
rect 4479 27353 4491 27387
rect 4433 27347 4491 27353
rect 4522 27344 4528 27396
rect 4580 27384 4586 27396
rect 4580 27356 4625 27384
rect 4580 27344 4586 27356
rect 5442 27344 5448 27396
rect 5500 27384 5506 27396
rect 5721 27387 5779 27393
rect 5721 27384 5733 27387
rect 5500 27356 5733 27384
rect 5500 27344 5506 27356
rect 5721 27353 5733 27356
rect 5767 27353 5779 27387
rect 5721 27347 5779 27353
rect 6733 27387 6791 27393
rect 6733 27353 6745 27387
rect 6779 27384 6791 27387
rect 6822 27384 6828 27396
rect 6779 27356 6828 27384
rect 6779 27353 6791 27356
rect 6733 27347 6791 27353
rect 6822 27344 6828 27356
rect 6880 27344 6886 27396
rect 7374 27384 7380 27396
rect 7335 27356 7380 27384
rect 7374 27344 7380 27356
rect 7432 27344 7438 27396
rect 2682 27316 2688 27328
rect 2643 27288 2688 27316
rect 2682 27276 2688 27288
rect 2740 27276 2746 27328
rect 3970 27316 3976 27328
rect 3931 27288 3976 27316
rect 3970 27276 3976 27288
rect 4028 27276 4034 27328
rect 5626 27316 5632 27328
rect 5587 27288 5632 27316
rect 5626 27276 5632 27288
rect 5684 27276 5690 27328
rect 6641 27319 6699 27325
rect 6641 27285 6653 27319
rect 6687 27316 6699 27319
rect 6914 27316 6920 27328
rect 6687 27288 6920 27316
rect 6687 27285 6699 27288
rect 6641 27279 6699 27285
rect 6914 27276 6920 27288
rect 6972 27276 6978 27328
rect 1104 27226 8832 27248
rect 1104 27174 3547 27226
rect 3599 27174 3611 27226
rect 3663 27174 3675 27226
rect 3727 27174 3739 27226
rect 3791 27174 3803 27226
rect 3855 27174 6144 27226
rect 6196 27174 6208 27226
rect 6260 27174 6272 27226
rect 6324 27174 6336 27226
rect 6388 27174 6400 27226
rect 6452 27174 8832 27226
rect 1104 27152 8832 27174
rect 2038 27112 2044 27124
rect 1999 27084 2044 27112
rect 2038 27072 2044 27084
rect 2096 27072 2102 27124
rect 3881 27115 3939 27121
rect 3881 27081 3893 27115
rect 3927 27112 3939 27115
rect 7374 27112 7380 27124
rect 3927 27084 7380 27112
rect 3927 27081 3939 27084
rect 3881 27075 3939 27081
rect 7374 27072 7380 27084
rect 7432 27072 7438 27124
rect 5442 27004 5448 27056
rect 5500 27044 5506 27056
rect 6454 27044 6460 27056
rect 5500 27016 6460 27044
rect 5500 27004 5506 27016
rect 6454 27004 6460 27016
rect 6512 27044 6518 27056
rect 6641 27047 6699 27053
rect 6641 27044 6653 27047
rect 6512 27016 6653 27044
rect 6512 27004 6518 27016
rect 6641 27013 6653 27016
rect 6687 27013 6699 27047
rect 6641 27007 6699 27013
rect 3234 26976 3240 26988
rect 3195 26948 3240 26976
rect 3234 26936 3240 26948
rect 3292 26936 3298 26988
rect 3418 26936 3424 26988
rect 3476 26976 3482 26988
rect 4341 26979 4399 26985
rect 4341 26976 4353 26979
rect 3476 26948 4353 26976
rect 3476 26936 3482 26948
rect 4341 26945 4353 26948
rect 4387 26945 4399 26979
rect 4522 26976 4528 26988
rect 4483 26948 4528 26976
rect 4341 26939 4399 26945
rect 4522 26936 4528 26948
rect 4580 26936 4586 26988
rect 5261 26979 5319 26985
rect 5261 26945 5273 26979
rect 5307 26976 5319 26979
rect 5534 26976 5540 26988
rect 5307 26948 5540 26976
rect 5307 26945 5319 26948
rect 5261 26939 5319 26945
rect 5534 26936 5540 26948
rect 5592 26936 5598 26988
rect 5810 26936 5816 26988
rect 5868 26976 5874 26988
rect 7101 26979 7159 26985
rect 7101 26976 7113 26979
rect 5868 26948 7113 26976
rect 5868 26936 5874 26948
rect 7101 26945 7113 26948
rect 7147 26976 7159 26979
rect 7926 26976 7932 26988
rect 7147 26948 7932 26976
rect 7147 26945 7159 26948
rect 7101 26939 7159 26945
rect 7926 26936 7932 26948
rect 7984 26936 7990 26988
rect 3789 26911 3847 26917
rect 3789 26877 3801 26911
rect 3835 26908 3847 26911
rect 6549 26911 6607 26917
rect 6549 26908 6561 26911
rect 3835 26880 6561 26908
rect 3835 26877 3847 26880
rect 3789 26871 3847 26877
rect 6549 26877 6561 26880
rect 6595 26877 6607 26911
rect 6549 26871 6607 26877
rect 7190 26868 7196 26920
rect 7248 26908 7254 26920
rect 7561 26911 7619 26917
rect 7561 26908 7573 26911
rect 7248 26880 7573 26908
rect 7248 26868 7254 26880
rect 7561 26877 7573 26880
rect 7607 26877 7619 26911
rect 7561 26871 7619 26877
rect 8113 26911 8171 26917
rect 8113 26877 8125 26911
rect 8159 26908 8171 26911
rect 8202 26908 8208 26920
rect 8159 26880 8208 26908
rect 8159 26877 8171 26880
rect 8113 26871 8171 26877
rect 5902 26840 5908 26852
rect 2746 26812 5908 26840
rect 2746 26784 2774 26812
rect 5902 26800 5908 26812
rect 5960 26800 5966 26852
rect 6822 26800 6828 26852
rect 6880 26840 6886 26852
rect 7653 26843 7711 26849
rect 7653 26840 7665 26843
rect 6880 26812 7665 26840
rect 6880 26800 6886 26812
rect 7653 26809 7665 26812
rect 7699 26809 7711 26843
rect 7653 26803 7711 26809
rect 2593 26775 2651 26781
rect 2593 26741 2605 26775
rect 2639 26772 2651 26775
rect 2746 26772 2780 26784
rect 2639 26744 2780 26772
rect 2639 26741 2651 26744
rect 2593 26735 2651 26741
rect 2774 26732 2780 26744
rect 2832 26732 2838 26784
rect 3145 26775 3203 26781
rect 3145 26741 3157 26775
rect 3191 26772 3203 26775
rect 5166 26772 5172 26784
rect 3191 26744 5172 26772
rect 3191 26741 3203 26744
rect 3145 26735 3203 26741
rect 5166 26732 5172 26744
rect 5224 26732 5230 26784
rect 5813 26775 5871 26781
rect 5813 26741 5825 26775
rect 5859 26772 5871 26775
rect 8128 26772 8156 26871
rect 8202 26868 8208 26880
rect 8260 26868 8266 26920
rect 5859 26744 8156 26772
rect 5859 26741 5871 26744
rect 5813 26735 5871 26741
rect 1104 26682 8832 26704
rect 1104 26630 2248 26682
rect 2300 26630 2312 26682
rect 2364 26630 2376 26682
rect 2428 26630 2440 26682
rect 2492 26630 2504 26682
rect 2556 26630 4846 26682
rect 4898 26630 4910 26682
rect 4962 26630 4974 26682
rect 5026 26630 5038 26682
rect 5090 26630 5102 26682
rect 5154 26630 7443 26682
rect 7495 26630 7507 26682
rect 7559 26630 7571 26682
rect 7623 26630 7635 26682
rect 7687 26630 7699 26682
rect 7751 26630 8832 26682
rect 1104 26608 8832 26630
rect 2590 26568 2596 26580
rect 2551 26540 2596 26568
rect 2590 26528 2596 26540
rect 2648 26528 2654 26580
rect 2774 26568 2780 26580
rect 2700 26540 2780 26568
rect 2041 26503 2099 26509
rect 2041 26469 2053 26503
rect 2087 26500 2099 26503
rect 2700 26500 2728 26540
rect 2774 26528 2780 26540
rect 2832 26528 2838 26580
rect 3068 26540 6040 26568
rect 2087 26472 2728 26500
rect 2087 26469 2099 26472
rect 2041 26463 2099 26469
rect 3068 26373 3096 26540
rect 3234 26460 3240 26512
rect 3292 26500 3298 26512
rect 4065 26503 4123 26509
rect 4065 26500 4077 26503
rect 3292 26472 4077 26500
rect 3292 26460 3298 26472
rect 4065 26469 4077 26472
rect 4111 26469 4123 26503
rect 4065 26463 4123 26469
rect 3970 26432 3976 26444
rect 3931 26404 3976 26432
rect 3970 26392 3976 26404
rect 4028 26392 4034 26444
rect 4080 26432 4108 26463
rect 4080 26404 5212 26432
rect 3053 26367 3111 26373
rect 3053 26333 3065 26367
rect 3099 26333 3111 26367
rect 4154 26364 4160 26376
rect 3053 26327 3111 26333
rect 3988 26336 4160 26364
rect 3988 26296 4016 26336
rect 4154 26324 4160 26336
rect 4212 26324 4218 26376
rect 5184 26373 5212 26404
rect 4525 26367 4583 26373
rect 4525 26333 4537 26367
rect 4571 26364 4583 26367
rect 5169 26367 5227 26373
rect 4571 26336 5120 26364
rect 4571 26333 4583 26336
rect 4525 26327 4583 26333
rect 3252 26268 4016 26296
rect 3252 26237 3280 26268
rect 4062 26256 4068 26308
rect 4120 26296 4126 26308
rect 4985 26299 5043 26305
rect 4985 26296 4997 26299
rect 4120 26268 4997 26296
rect 4120 26256 4126 26268
rect 4985 26265 4997 26268
rect 5031 26265 5043 26299
rect 5092 26296 5120 26336
rect 5169 26333 5181 26367
rect 5215 26333 5227 26367
rect 5902 26364 5908 26376
rect 5863 26336 5908 26364
rect 5169 26327 5227 26333
rect 5902 26324 5908 26336
rect 5960 26324 5966 26376
rect 6012 26364 6040 26540
rect 6454 26500 6460 26512
rect 6415 26472 6460 26500
rect 6454 26460 6460 26472
rect 6512 26460 6518 26512
rect 6457 26367 6515 26373
rect 6457 26364 6469 26367
rect 6012 26336 6469 26364
rect 6457 26333 6469 26336
rect 6503 26364 6515 26367
rect 6914 26364 6920 26376
rect 6503 26336 6920 26364
rect 6503 26333 6515 26336
rect 6457 26327 6515 26333
rect 6914 26324 6920 26336
rect 6972 26324 6978 26376
rect 7926 26364 7932 26376
rect 7887 26336 7932 26364
rect 7926 26324 7932 26336
rect 7984 26324 7990 26376
rect 5920 26296 5948 26324
rect 5092 26268 5948 26296
rect 4985 26259 5043 26265
rect 3237 26231 3295 26237
rect 3237 26197 3249 26231
rect 3283 26197 3295 26231
rect 5000 26228 5028 26259
rect 5258 26228 5264 26240
rect 5000 26200 5264 26228
rect 3237 26191 3295 26197
rect 5258 26188 5264 26200
rect 5316 26188 5322 26240
rect 5902 26188 5908 26240
rect 5960 26228 5966 26240
rect 6638 26228 6644 26240
rect 5960 26200 6644 26228
rect 5960 26188 5966 26200
rect 6638 26188 6644 26200
rect 6696 26188 6702 26240
rect 1104 26138 8832 26160
rect 1104 26086 3547 26138
rect 3599 26086 3611 26138
rect 3663 26086 3675 26138
rect 3727 26086 3739 26138
rect 3791 26086 3803 26138
rect 3855 26086 6144 26138
rect 6196 26086 6208 26138
rect 6260 26086 6272 26138
rect 6324 26086 6336 26138
rect 6388 26086 6400 26138
rect 6452 26086 8832 26138
rect 1104 26064 8832 26086
rect 1765 26027 1823 26033
rect 1765 25993 1777 26027
rect 1811 26024 1823 26027
rect 2038 26024 2044 26036
rect 1811 25996 2044 26024
rect 1811 25993 1823 25996
rect 1765 25987 1823 25993
rect 2038 25984 2044 25996
rect 2096 26024 2102 26036
rect 6457 26027 6515 26033
rect 2096 25996 4292 26024
rect 2096 25984 2102 25996
rect 2317 25959 2375 25965
rect 2317 25925 2329 25959
rect 2363 25956 2375 25959
rect 2682 25956 2688 25968
rect 2363 25928 2688 25956
rect 2363 25925 2375 25928
rect 2317 25919 2375 25925
rect 2682 25916 2688 25928
rect 2740 25956 2746 25968
rect 3789 25959 3847 25965
rect 2740 25916 2774 25956
rect 3789 25925 3801 25959
rect 3835 25956 3847 25959
rect 4062 25956 4068 25968
rect 3835 25928 4068 25956
rect 3835 25925 3847 25928
rect 3789 25919 3847 25925
rect 4062 25916 4068 25928
rect 4120 25916 4126 25968
rect 2746 25684 2774 25916
rect 2869 25891 2927 25897
rect 2869 25857 2881 25891
rect 2915 25857 2927 25891
rect 2869 25851 2927 25857
rect 3053 25891 3111 25897
rect 3053 25857 3065 25891
rect 3099 25888 3111 25891
rect 3418 25888 3424 25900
rect 3099 25860 3424 25888
rect 3099 25857 3111 25860
rect 3053 25851 3111 25857
rect 2884 25820 2912 25851
rect 3418 25848 3424 25860
rect 3476 25848 3482 25900
rect 3605 25891 3663 25897
rect 3605 25857 3617 25891
rect 3651 25888 3663 25891
rect 4154 25888 4160 25900
rect 3651 25860 4160 25888
rect 3651 25857 3663 25860
rect 3605 25851 3663 25857
rect 4154 25848 4160 25860
rect 4212 25848 4218 25900
rect 4264 25897 4292 25996
rect 6457 25993 6469 26027
rect 6503 26024 6515 26027
rect 7190 26024 7196 26036
rect 6503 25996 7196 26024
rect 6503 25993 6515 25996
rect 6457 25987 6515 25993
rect 7190 25984 7196 25996
rect 7248 25984 7254 26036
rect 7006 25956 7012 25968
rect 6967 25928 7012 25956
rect 7006 25916 7012 25928
rect 7064 25916 7070 25968
rect 7282 25956 7288 25968
rect 7243 25928 7288 25956
rect 7282 25916 7288 25928
rect 7340 25916 7346 25968
rect 4249 25891 4307 25897
rect 4249 25857 4261 25891
rect 4295 25888 4307 25891
rect 4540 25888 4660 25894
rect 4295 25866 5120 25888
rect 4295 25860 4568 25866
rect 4632 25860 5120 25866
rect 4295 25857 4307 25860
rect 4249 25851 4307 25857
rect 5092 25820 5120 25860
rect 5258 25848 5264 25900
rect 5316 25888 5322 25900
rect 6549 25891 6607 25897
rect 5316 25860 5361 25888
rect 5316 25848 5322 25860
rect 6549 25857 6561 25891
rect 6595 25888 6607 25891
rect 6914 25888 6920 25900
rect 6595 25860 6920 25888
rect 6595 25857 6607 25860
rect 6549 25851 6607 25857
rect 6914 25848 6920 25860
rect 6972 25848 6978 25900
rect 7834 25848 7840 25900
rect 7892 25888 7898 25900
rect 7929 25891 7987 25897
rect 7929 25888 7941 25891
rect 7892 25860 7941 25888
rect 7892 25848 7898 25860
rect 7929 25857 7941 25860
rect 7975 25857 7987 25891
rect 7929 25851 7987 25857
rect 5718 25820 5724 25832
rect 2884 25792 3464 25820
rect 5092 25792 5724 25820
rect 3436 25752 3464 25792
rect 5718 25780 5724 25792
rect 5776 25780 5782 25832
rect 5258 25752 5264 25764
rect 3436 25724 5264 25752
rect 5258 25712 5264 25724
rect 5316 25752 5322 25764
rect 5537 25755 5595 25761
rect 5537 25752 5549 25755
rect 5316 25724 5549 25752
rect 5316 25712 5322 25724
rect 5537 25721 5549 25724
rect 5583 25721 5595 25755
rect 5537 25715 5595 25721
rect 7944 25684 7972 25851
rect 2746 25656 7972 25684
rect 1104 25594 8832 25616
rect 1104 25542 2248 25594
rect 2300 25542 2312 25594
rect 2364 25542 2376 25594
rect 2428 25542 2440 25594
rect 2492 25542 2504 25594
rect 2556 25542 4846 25594
rect 4898 25542 4910 25594
rect 4962 25542 4974 25594
rect 5026 25542 5038 25594
rect 5090 25542 5102 25594
rect 5154 25542 7443 25594
rect 7495 25542 7507 25594
rect 7559 25542 7571 25594
rect 7623 25542 7635 25594
rect 7687 25542 7699 25594
rect 7751 25542 8832 25594
rect 1104 25520 8832 25542
rect 2038 25480 2044 25492
rect 1999 25452 2044 25480
rect 2038 25440 2044 25452
rect 2096 25440 2102 25492
rect 5258 25412 5264 25424
rect 5219 25384 5264 25412
rect 5258 25372 5264 25384
rect 5316 25372 5322 25424
rect 6822 25412 6828 25424
rect 6783 25384 6828 25412
rect 6822 25372 6828 25384
rect 6880 25372 6886 25424
rect 5166 25344 5172 25356
rect 5127 25316 5172 25344
rect 5166 25304 5172 25316
rect 5224 25304 5230 25356
rect 5718 25344 5724 25356
rect 5679 25316 5724 25344
rect 5718 25304 5724 25316
rect 5776 25304 5782 25356
rect 2593 25279 2651 25285
rect 2593 25245 2605 25279
rect 2639 25276 2651 25279
rect 3237 25279 3295 25285
rect 2639 25248 2774 25276
rect 2639 25245 2651 25248
rect 2593 25239 2651 25245
rect 2746 25140 2774 25248
rect 3237 25245 3249 25279
rect 3283 25276 3295 25279
rect 4522 25276 4528 25288
rect 3283 25248 4528 25276
rect 3283 25245 3295 25248
rect 3237 25239 3295 25245
rect 4522 25236 4528 25248
rect 4580 25236 4586 25288
rect 4709 25279 4767 25285
rect 4709 25245 4721 25279
rect 4755 25276 4767 25279
rect 5994 25276 6000 25288
rect 4755 25248 6000 25276
rect 4755 25245 4767 25248
rect 4709 25239 4767 25245
rect 5994 25236 6000 25248
rect 6052 25236 6058 25288
rect 7190 25276 7196 25288
rect 7151 25248 7196 25276
rect 7190 25236 7196 25248
rect 7248 25236 7254 25288
rect 8113 25279 8171 25285
rect 8113 25245 8125 25279
rect 8159 25276 8171 25279
rect 8202 25276 8208 25288
rect 8159 25248 8208 25276
rect 8159 25245 8171 25248
rect 8113 25239 8171 25245
rect 3145 25211 3203 25217
rect 3145 25177 3157 25211
rect 3191 25208 3203 25211
rect 4157 25211 4215 25217
rect 4157 25208 4169 25211
rect 3191 25180 4169 25208
rect 3191 25177 3203 25180
rect 3145 25171 3203 25177
rect 4157 25177 4169 25180
rect 4203 25177 4215 25211
rect 4157 25171 4215 25177
rect 4246 25168 4252 25220
rect 4304 25208 4310 25220
rect 4304 25180 4349 25208
rect 4304 25168 4310 25180
rect 8128 25140 8156 25239
rect 8202 25236 8208 25248
rect 8260 25236 8266 25288
rect 2746 25112 8156 25140
rect 1104 25050 8832 25072
rect 1104 24998 3547 25050
rect 3599 24998 3611 25050
rect 3663 24998 3675 25050
rect 3727 24998 3739 25050
rect 3791 24998 3803 25050
rect 3855 24998 6144 25050
rect 6196 24998 6208 25050
rect 6260 24998 6272 25050
rect 6324 24998 6336 25050
rect 6388 24998 6400 25050
rect 6452 24998 8832 25050
rect 1104 24976 8832 24998
rect 6546 24896 6552 24948
rect 6604 24896 6610 24948
rect 5994 24868 6000 24880
rect 5644 24840 6000 24868
rect 3418 24800 3424 24812
rect 3379 24772 3424 24800
rect 3418 24760 3424 24772
rect 3476 24800 3482 24812
rect 5644 24809 5672 24840
rect 5994 24828 6000 24840
rect 6052 24828 6058 24880
rect 6086 24828 6092 24880
rect 6144 24868 6150 24880
rect 6564 24868 6592 24896
rect 6144 24840 6592 24868
rect 6144 24828 6150 24840
rect 4157 24803 4215 24809
rect 4157 24800 4169 24803
rect 3476 24772 4169 24800
rect 3476 24760 3482 24772
rect 4157 24769 4169 24772
rect 4203 24769 4215 24803
rect 4157 24763 4215 24769
rect 5629 24803 5687 24809
rect 5629 24769 5641 24803
rect 5675 24769 5687 24803
rect 5629 24763 5687 24769
rect 1857 24735 1915 24741
rect 1857 24701 1869 24735
rect 1903 24732 1915 24735
rect 2409 24735 2467 24741
rect 2409 24732 2421 24735
rect 1903 24704 2421 24732
rect 1903 24701 1915 24704
rect 1857 24695 1915 24701
rect 2409 24701 2421 24704
rect 2455 24732 2467 24735
rect 5644 24732 5672 24763
rect 5718 24760 5724 24812
rect 5776 24800 5782 24812
rect 6365 24803 6423 24809
rect 6365 24800 6377 24803
rect 5776 24772 6377 24800
rect 5776 24760 5782 24772
rect 6365 24769 6377 24772
rect 6411 24769 6423 24803
rect 6546 24800 6552 24812
rect 6507 24772 6552 24800
rect 6365 24763 6423 24769
rect 6546 24760 6552 24772
rect 6604 24760 6610 24812
rect 6730 24760 6736 24812
rect 6788 24800 6794 24812
rect 7285 24803 7343 24809
rect 7285 24800 7297 24803
rect 6788 24772 7297 24800
rect 6788 24760 6794 24772
rect 7285 24769 7297 24772
rect 7331 24769 7343 24803
rect 7285 24763 7343 24769
rect 7834 24760 7840 24812
rect 7892 24800 7898 24812
rect 8021 24803 8079 24809
rect 8021 24800 8033 24803
rect 7892 24772 8033 24800
rect 7892 24760 7898 24772
rect 8021 24769 8033 24772
rect 8067 24769 8079 24803
rect 8021 24763 8079 24769
rect 2455 24704 5672 24732
rect 2455 24701 2467 24704
rect 2409 24695 2467 24701
rect 3605 24667 3663 24673
rect 3605 24633 3617 24667
rect 3651 24664 3663 24667
rect 3878 24664 3884 24676
rect 3651 24636 3884 24664
rect 3651 24633 3663 24636
rect 3605 24627 3663 24633
rect 3878 24624 3884 24636
rect 3936 24624 3942 24676
rect 4157 24667 4215 24673
rect 4157 24633 4169 24667
rect 4203 24664 4215 24667
rect 4246 24664 4252 24676
rect 4203 24636 4252 24664
rect 4203 24633 4215 24636
rect 4157 24627 4215 24633
rect 4246 24624 4252 24636
rect 4304 24624 4310 24676
rect 7282 24624 7288 24676
rect 7340 24664 7346 24676
rect 7837 24667 7895 24673
rect 7837 24664 7849 24667
rect 7340 24636 7849 24664
rect 7340 24624 7346 24636
rect 7837 24633 7849 24636
rect 7883 24633 7895 24667
rect 7837 24627 7895 24633
rect 2958 24596 2964 24608
rect 2919 24568 2964 24596
rect 2958 24556 2964 24568
rect 3016 24556 3022 24608
rect 1104 24506 8832 24528
rect 1104 24454 2248 24506
rect 2300 24454 2312 24506
rect 2364 24454 2376 24506
rect 2428 24454 2440 24506
rect 2492 24454 2504 24506
rect 2556 24454 4846 24506
rect 4898 24454 4910 24506
rect 4962 24454 4974 24506
rect 5026 24454 5038 24506
rect 5090 24454 5102 24506
rect 5154 24454 7443 24506
rect 7495 24454 7507 24506
rect 7559 24454 7571 24506
rect 7623 24454 7635 24506
rect 7687 24454 7699 24506
rect 7751 24454 8832 24506
rect 1104 24432 8832 24454
rect 4617 24327 4675 24333
rect 4617 24324 4629 24327
rect 4080 24296 4629 24324
rect 4080 24197 4108 24296
rect 4617 24293 4629 24296
rect 4663 24324 4675 24327
rect 6546 24324 6552 24336
rect 4663 24296 6552 24324
rect 4663 24293 4675 24296
rect 4617 24287 4675 24293
rect 6546 24284 6552 24296
rect 6604 24284 6610 24336
rect 6914 24284 6920 24336
rect 6972 24324 6978 24336
rect 7374 24324 7380 24336
rect 6972 24296 7380 24324
rect 6972 24284 6978 24296
rect 7374 24284 7380 24296
rect 7432 24324 7438 24336
rect 7653 24327 7711 24333
rect 7653 24324 7665 24327
rect 7432 24296 7665 24324
rect 7432 24284 7438 24296
rect 7653 24293 7665 24296
rect 7699 24293 7711 24327
rect 7653 24287 7711 24293
rect 4154 24216 4160 24268
rect 4212 24256 4218 24268
rect 5350 24256 5356 24268
rect 4212 24228 5356 24256
rect 4212 24216 4218 24228
rect 5350 24216 5356 24228
rect 5408 24256 5414 24268
rect 5537 24259 5595 24265
rect 5537 24256 5549 24259
rect 5408 24228 5549 24256
rect 5408 24216 5414 24228
rect 5537 24225 5549 24228
rect 5583 24225 5595 24259
rect 8110 24256 8116 24268
rect 8071 24228 8116 24256
rect 5537 24219 5595 24225
rect 8110 24216 8116 24228
rect 8168 24216 8174 24268
rect 4065 24191 4123 24197
rect 4065 24157 4077 24191
rect 4111 24157 4123 24191
rect 4065 24151 4123 24157
rect 5077 24191 5135 24197
rect 5077 24157 5089 24191
rect 5123 24157 5135 24191
rect 5626 24188 5632 24200
rect 5587 24160 5632 24188
rect 5077 24151 5135 24157
rect 2685 24123 2743 24129
rect 2685 24089 2697 24123
rect 2731 24120 2743 24123
rect 2958 24120 2964 24132
rect 2731 24092 2964 24120
rect 2731 24089 2743 24092
rect 2685 24083 2743 24089
rect 2958 24080 2964 24092
rect 3016 24120 3022 24132
rect 3016 24092 4108 24120
rect 3016 24080 3022 24092
rect 2130 24052 2136 24064
rect 2091 24024 2136 24052
rect 2130 24012 2136 24024
rect 2188 24012 2194 24064
rect 3234 24052 3240 24064
rect 3195 24024 3240 24052
rect 3234 24012 3240 24024
rect 3292 24012 3298 24064
rect 3970 24052 3976 24064
rect 3931 24024 3976 24052
rect 3970 24012 3976 24024
rect 4028 24012 4034 24064
rect 4080 24052 4108 24092
rect 4154 24080 4160 24132
rect 4212 24120 4218 24132
rect 4525 24123 4583 24129
rect 4525 24120 4537 24123
rect 4212 24092 4537 24120
rect 4212 24080 4218 24092
rect 4525 24089 4537 24092
rect 4571 24089 4583 24123
rect 4525 24083 4583 24089
rect 5092 24120 5120 24151
rect 5626 24148 5632 24160
rect 5684 24148 5690 24200
rect 6638 24148 6644 24200
rect 6696 24188 6702 24200
rect 7101 24191 7159 24197
rect 7101 24188 7113 24191
rect 6696 24160 7113 24188
rect 6696 24148 6702 24160
rect 7101 24157 7113 24160
rect 7147 24157 7159 24191
rect 7101 24151 7159 24157
rect 6730 24120 6736 24132
rect 5092 24092 6736 24120
rect 5092 24052 5120 24092
rect 6730 24080 6736 24092
rect 6788 24080 6794 24132
rect 7558 24120 7564 24132
rect 7519 24092 7564 24120
rect 7558 24080 7564 24092
rect 7616 24080 7622 24132
rect 4080 24024 5120 24052
rect 1104 23962 8832 23984
rect 1104 23910 3547 23962
rect 3599 23910 3611 23962
rect 3663 23910 3675 23962
rect 3727 23910 3739 23962
rect 3791 23910 3803 23962
rect 3855 23910 6144 23962
rect 6196 23910 6208 23962
rect 6260 23910 6272 23962
rect 6324 23910 6336 23962
rect 6388 23910 6400 23962
rect 6452 23910 8832 23962
rect 1104 23888 8832 23910
rect 3970 23808 3976 23860
rect 4028 23808 4034 23860
rect 4154 23848 4160 23860
rect 4115 23820 4160 23848
rect 4154 23808 4160 23820
rect 4212 23808 4218 23860
rect 4801 23851 4859 23857
rect 4801 23817 4813 23851
rect 4847 23848 4859 23851
rect 7558 23848 7564 23860
rect 4847 23820 7564 23848
rect 4847 23817 4859 23820
rect 4801 23811 4859 23817
rect 7558 23808 7564 23820
rect 7616 23808 7622 23860
rect 3988 23780 4016 23808
rect 5261 23783 5319 23789
rect 5261 23780 5273 23783
rect 3988 23752 5273 23780
rect 5261 23749 5273 23752
rect 5307 23749 5319 23783
rect 5261 23743 5319 23749
rect 5350 23740 5356 23792
rect 5408 23780 5414 23792
rect 6457 23783 6515 23789
rect 5408 23752 5453 23780
rect 5408 23740 5414 23752
rect 6457 23749 6469 23783
rect 6503 23780 6515 23783
rect 7190 23780 7196 23792
rect 6503 23752 7196 23780
rect 6503 23749 6515 23752
rect 6457 23743 6515 23749
rect 3973 23715 4031 23721
rect 3973 23681 3985 23715
rect 4019 23681 4031 23715
rect 3973 23675 4031 23681
rect 4617 23715 4675 23721
rect 4617 23681 4629 23715
rect 4663 23712 4675 23715
rect 6472 23712 6500 23743
rect 7190 23740 7196 23752
rect 7248 23740 7254 23792
rect 7374 23780 7380 23792
rect 7335 23752 7380 23780
rect 7374 23740 7380 23752
rect 7432 23740 7438 23792
rect 6638 23712 6644 23724
rect 4663 23684 6500 23712
rect 6599 23684 6644 23712
rect 4663 23681 4675 23684
rect 4617 23675 4675 23681
rect 3988 23644 4016 23675
rect 6638 23672 6644 23684
rect 6696 23672 6702 23724
rect 8110 23712 8116 23724
rect 8071 23684 8116 23712
rect 8110 23672 8116 23684
rect 8168 23672 8174 23724
rect 5626 23644 5632 23656
rect 3988 23616 5632 23644
rect 5626 23604 5632 23616
rect 5684 23604 5690 23656
rect 5810 23604 5816 23656
rect 5868 23644 5874 23656
rect 6546 23644 6552 23656
rect 5868 23616 6552 23644
rect 5868 23604 5874 23616
rect 6546 23604 6552 23616
rect 6604 23604 6610 23656
rect 2130 23536 2136 23588
rect 2188 23576 2194 23588
rect 2188 23548 2774 23576
rect 2188 23536 2194 23548
rect 2746 23508 2774 23548
rect 3234 23536 3240 23588
rect 3292 23576 3298 23588
rect 3513 23579 3571 23585
rect 3513 23576 3525 23579
rect 3292 23548 3525 23576
rect 3292 23536 3298 23548
rect 3513 23545 3525 23548
rect 3559 23576 3571 23579
rect 8128 23576 8156 23672
rect 3559 23548 8156 23576
rect 3559 23545 3571 23548
rect 3513 23539 3571 23545
rect 2961 23511 3019 23517
rect 2961 23508 2973 23511
rect 2746 23480 2973 23508
rect 2961 23477 2973 23480
rect 3007 23508 3019 23511
rect 5810 23508 5816 23520
rect 3007 23480 5816 23508
rect 3007 23477 3019 23480
rect 2961 23471 3019 23477
rect 5810 23468 5816 23480
rect 5868 23468 5874 23520
rect 1104 23418 8832 23440
rect 1104 23366 2248 23418
rect 2300 23366 2312 23418
rect 2364 23366 2376 23418
rect 2428 23366 2440 23418
rect 2492 23366 2504 23418
rect 2556 23366 4846 23418
rect 4898 23366 4910 23418
rect 4962 23366 4974 23418
rect 5026 23366 5038 23418
rect 5090 23366 5102 23418
rect 5154 23366 7443 23418
rect 7495 23366 7507 23418
rect 7559 23366 7571 23418
rect 7623 23366 7635 23418
rect 7687 23366 7699 23418
rect 7751 23366 8832 23418
rect 1104 23344 8832 23366
rect 3050 23264 3056 23316
rect 3108 23304 3114 23316
rect 3881 23307 3939 23313
rect 3881 23304 3893 23307
rect 3108 23276 3893 23304
rect 3108 23264 3114 23276
rect 3881 23273 3893 23276
rect 3927 23304 3939 23307
rect 3927 23276 7696 23304
rect 3927 23273 3939 23276
rect 3881 23267 3939 23273
rect 6638 23196 6644 23248
rect 6696 23236 6702 23248
rect 7193 23239 7251 23245
rect 7193 23236 7205 23239
rect 6696 23208 7205 23236
rect 6696 23196 6702 23208
rect 7193 23205 7205 23208
rect 7239 23205 7251 23239
rect 7193 23199 7251 23205
rect 4433 23171 4491 23177
rect 4433 23137 4445 23171
rect 4479 23168 4491 23171
rect 7101 23171 7159 23177
rect 7101 23168 7113 23171
rect 4479 23140 7113 23168
rect 4479 23137 4491 23140
rect 4433 23131 4491 23137
rect 7101 23137 7113 23140
rect 7147 23137 7159 23171
rect 7101 23131 7159 23137
rect 2590 23060 2596 23112
rect 2648 23100 2654 23112
rect 2685 23103 2743 23109
rect 2685 23100 2697 23103
rect 2648 23072 2697 23100
rect 2648 23060 2654 23072
rect 2685 23069 2697 23072
rect 2731 23100 2743 23103
rect 5537 23103 5595 23109
rect 5537 23100 5549 23103
rect 2731 23072 5549 23100
rect 2731 23069 2743 23072
rect 2685 23063 2743 23069
rect 5537 23069 5549 23072
rect 5583 23100 5595 23103
rect 5902 23100 5908 23112
rect 5583 23072 5908 23100
rect 5583 23069 5595 23072
rect 5537 23063 5595 23069
rect 5902 23060 5908 23072
rect 5960 23060 5966 23112
rect 6641 23103 6699 23109
rect 6641 23069 6653 23103
rect 6687 23100 6699 23103
rect 6730 23100 6736 23112
rect 6687 23072 6736 23100
rect 6687 23069 6699 23072
rect 6641 23063 6699 23069
rect 6730 23060 6736 23072
rect 6788 23060 6794 23112
rect 7668 23109 7696 23276
rect 7653 23103 7711 23109
rect 7653 23069 7665 23103
rect 7699 23100 7711 23103
rect 8110 23100 8116 23112
rect 7699 23072 8116 23100
rect 7699 23069 7711 23072
rect 7653 23063 7711 23069
rect 8110 23060 8116 23072
rect 8168 23060 8174 23112
rect 4614 22992 4620 23044
rect 4672 23032 4678 23044
rect 4985 23035 5043 23041
rect 4985 23032 4997 23035
rect 4672 23004 4997 23032
rect 4672 22992 4678 23004
rect 4985 23001 4997 23004
rect 5031 23001 5043 23035
rect 4985 22995 5043 23001
rect 5077 23035 5135 23041
rect 5077 23001 5089 23035
rect 5123 23032 5135 23035
rect 5166 23032 5172 23044
rect 5123 23004 5172 23032
rect 5123 23001 5135 23004
rect 5077 22995 5135 23001
rect 5166 22992 5172 23004
rect 5224 22992 5230 23044
rect 5258 22992 5264 23044
rect 5316 23032 5322 23044
rect 6089 23035 6147 23041
rect 6089 23032 6101 23035
rect 5316 23004 6101 23032
rect 5316 22992 5322 23004
rect 6089 23001 6101 23004
rect 6135 23001 6147 23035
rect 6089 22995 6147 23001
rect 6181 23035 6239 23041
rect 6181 23001 6193 23035
rect 6227 23032 6239 23035
rect 7006 23032 7012 23044
rect 6227 23004 7012 23032
rect 6227 23001 6239 23004
rect 6181 22995 6239 23001
rect 3234 22964 3240 22976
rect 3195 22936 3240 22964
rect 3234 22924 3240 22936
rect 3292 22924 3298 22976
rect 4525 22967 4583 22973
rect 4525 22933 4537 22967
rect 4571 22964 4583 22967
rect 6196 22964 6224 22995
rect 7006 22992 7012 23004
rect 7064 22992 7070 23044
rect 4571 22936 6224 22964
rect 4571 22933 4583 22936
rect 4525 22927 4583 22933
rect 1104 22874 8832 22896
rect 1104 22822 3547 22874
rect 3599 22822 3611 22874
rect 3663 22822 3675 22874
rect 3727 22822 3739 22874
rect 3791 22822 3803 22874
rect 3855 22822 6144 22874
rect 6196 22822 6208 22874
rect 6260 22822 6272 22874
rect 6324 22822 6336 22874
rect 6388 22822 6400 22874
rect 6452 22822 8832 22874
rect 1104 22800 8832 22822
rect 3050 22760 3056 22772
rect 3011 22732 3056 22760
rect 3050 22720 3056 22732
rect 3108 22720 3114 22772
rect 3697 22763 3755 22769
rect 3697 22729 3709 22763
rect 3743 22760 3755 22763
rect 5258 22760 5264 22772
rect 3743 22732 5264 22760
rect 3743 22729 3755 22732
rect 3697 22723 3755 22729
rect 5258 22720 5264 22732
rect 5316 22720 5322 22772
rect 4246 22692 4252 22704
rect 4207 22664 4252 22692
rect 4246 22652 4252 22664
rect 4304 22652 4310 22704
rect 3513 22627 3571 22633
rect 3513 22593 3525 22627
rect 3559 22624 3571 22627
rect 6914 22624 6920 22636
rect 3559 22596 6920 22624
rect 3559 22593 3571 22596
rect 3513 22587 3571 22593
rect 6914 22584 6920 22596
rect 6972 22624 6978 22636
rect 7193 22627 7251 22633
rect 7193 22624 7205 22627
rect 6972 22596 7205 22624
rect 6972 22584 6978 22596
rect 7193 22593 7205 22596
rect 7239 22624 7251 22627
rect 7282 22624 7288 22636
rect 7239 22596 7288 22624
rect 7239 22593 7251 22596
rect 7193 22587 7251 22593
rect 7282 22584 7288 22596
rect 7340 22584 7346 22636
rect 8110 22624 8116 22636
rect 8071 22596 8116 22624
rect 8110 22584 8116 22596
rect 8168 22584 8174 22636
rect 4154 22516 4160 22568
rect 4212 22556 4218 22568
rect 4893 22559 4951 22565
rect 4893 22556 4905 22559
rect 4212 22528 4905 22556
rect 4212 22516 4218 22528
rect 4893 22525 4905 22528
rect 4939 22525 4951 22559
rect 4893 22519 4951 22525
rect 5445 22559 5503 22565
rect 5445 22525 5457 22559
rect 5491 22556 5503 22559
rect 5994 22556 6000 22568
rect 5491 22528 6000 22556
rect 5491 22525 5503 22528
rect 5445 22519 5503 22525
rect 4433 22491 4491 22497
rect 4433 22457 4445 22491
rect 4479 22488 4491 22491
rect 4522 22488 4528 22500
rect 4479 22460 4528 22488
rect 4479 22457 4491 22460
rect 4433 22451 4491 22457
rect 4522 22448 4528 22460
rect 4580 22448 4586 22500
rect 4706 22448 4712 22500
rect 4764 22488 4770 22500
rect 4985 22491 5043 22497
rect 4985 22488 4997 22491
rect 4764 22460 4997 22488
rect 4764 22448 4770 22460
rect 4985 22457 4997 22460
rect 5031 22457 5043 22491
rect 4985 22451 5043 22457
rect 2501 22423 2559 22429
rect 2501 22389 2513 22423
rect 2547 22420 2559 22423
rect 2682 22420 2688 22432
rect 2547 22392 2688 22420
rect 2547 22389 2559 22392
rect 2501 22383 2559 22389
rect 2682 22380 2688 22392
rect 2740 22380 2746 22432
rect 4062 22380 4068 22432
rect 4120 22420 4126 22432
rect 5460 22420 5488 22519
rect 5994 22516 6000 22528
rect 6052 22516 6058 22568
rect 6638 22488 6644 22500
rect 6599 22460 6644 22488
rect 6638 22448 6644 22460
rect 6696 22448 6702 22500
rect 4120 22392 5488 22420
rect 4120 22380 4126 22392
rect 1104 22330 8832 22352
rect 1104 22278 2248 22330
rect 2300 22278 2312 22330
rect 2364 22278 2376 22330
rect 2428 22278 2440 22330
rect 2492 22278 2504 22330
rect 2556 22278 4846 22330
rect 4898 22278 4910 22330
rect 4962 22278 4974 22330
rect 5026 22278 5038 22330
rect 5090 22278 5102 22330
rect 5154 22278 7443 22330
rect 7495 22278 7507 22330
rect 7559 22278 7571 22330
rect 7623 22278 7635 22330
rect 7687 22278 7699 22330
rect 7751 22278 8832 22330
rect 1104 22256 8832 22278
rect 3234 22216 3240 22228
rect 3147 22188 3240 22216
rect 3234 22176 3240 22188
rect 3292 22216 3298 22228
rect 6730 22216 6736 22228
rect 3292 22188 6736 22216
rect 3292 22176 3298 22188
rect 6730 22176 6736 22188
rect 6788 22176 6794 22228
rect 2682 22148 2688 22160
rect 2595 22120 2688 22148
rect 2682 22108 2688 22120
rect 2740 22148 2746 22160
rect 4062 22148 4068 22160
rect 2740 22120 4068 22148
rect 2740 22108 2746 22120
rect 4062 22108 4068 22120
rect 4120 22108 4126 22160
rect 4246 22108 4252 22160
rect 4304 22148 4310 22160
rect 4706 22148 4712 22160
rect 4304 22120 4712 22148
rect 4304 22108 4310 22120
rect 4706 22108 4712 22120
rect 4764 22108 4770 22160
rect 3881 22083 3939 22089
rect 3881 22049 3893 22083
rect 3927 22080 3939 22083
rect 4154 22080 4160 22092
rect 3927 22052 4160 22080
rect 3927 22049 3939 22052
rect 3881 22043 3939 22049
rect 4154 22040 4160 22052
rect 4212 22040 4218 22092
rect 6638 22040 6644 22092
rect 6696 22080 6702 22092
rect 6696 22052 7788 22080
rect 6696 22040 6702 22052
rect 4522 21972 4528 22024
rect 4580 22012 4586 22024
rect 4890 22012 4896 22024
rect 4580 21984 4896 22012
rect 4580 21972 4586 21984
rect 4890 21972 4896 21984
rect 4948 21972 4954 22024
rect 5994 22012 6000 22024
rect 5955 21984 6000 22012
rect 5994 21972 6000 21984
rect 6052 21972 6058 22024
rect 7006 22012 7012 22024
rect 6967 21984 7012 22012
rect 7006 21972 7012 21984
rect 7064 21972 7070 22024
rect 7760 22021 7788 22052
rect 7745 22015 7803 22021
rect 7745 21981 7757 22015
rect 7791 21981 7803 22015
rect 7745 21975 7803 21981
rect 6825 21947 6883 21953
rect 6825 21913 6837 21947
rect 6871 21944 6883 21947
rect 6914 21944 6920 21956
rect 6871 21916 6920 21944
rect 6871 21913 6883 21916
rect 6825 21907 6883 21913
rect 6914 21904 6920 21916
rect 6972 21904 6978 21956
rect 3973 21879 4031 21885
rect 3973 21845 3985 21879
rect 4019 21876 4031 21879
rect 5074 21876 5080 21888
rect 4019 21848 5080 21876
rect 4019 21845 4031 21848
rect 3973 21839 4031 21845
rect 5074 21836 5080 21848
rect 5132 21836 5138 21888
rect 1104 21786 8832 21808
rect 1104 21734 3547 21786
rect 3599 21734 3611 21786
rect 3663 21734 3675 21786
rect 3727 21734 3739 21786
rect 3791 21734 3803 21786
rect 3855 21734 6144 21786
rect 6196 21734 6208 21786
rect 6260 21734 6272 21786
rect 6324 21734 6336 21786
rect 6388 21734 6400 21786
rect 6452 21734 8832 21786
rect 1104 21712 8832 21734
rect 2590 21672 2596 21684
rect 2551 21644 2596 21672
rect 2590 21632 2596 21644
rect 2648 21632 2654 21684
rect 4433 21675 4491 21681
rect 4433 21641 4445 21675
rect 4479 21672 4491 21675
rect 4614 21672 4620 21684
rect 4479 21644 4620 21672
rect 4479 21641 4491 21644
rect 4433 21635 4491 21641
rect 4614 21632 4620 21644
rect 4672 21632 4678 21684
rect 4890 21604 4896 21616
rect 4851 21576 4896 21604
rect 4890 21564 4896 21576
rect 4948 21564 4954 21616
rect 5074 21604 5080 21616
rect 5035 21576 5080 21604
rect 5074 21564 5080 21576
rect 5132 21564 5138 21616
rect 4249 21539 4307 21545
rect 4249 21505 4261 21539
rect 4295 21536 4307 21539
rect 4908 21536 4936 21564
rect 4295 21508 4936 21536
rect 5813 21539 5871 21545
rect 4295 21505 4307 21508
rect 4249 21499 4307 21505
rect 5813 21505 5825 21539
rect 5859 21536 5871 21539
rect 5902 21536 5908 21548
rect 5859 21508 5908 21536
rect 5859 21505 5871 21508
rect 5813 21499 5871 21505
rect 5902 21496 5908 21508
rect 5960 21496 5966 21548
rect 6457 21539 6515 21545
rect 6457 21505 6469 21539
rect 6503 21536 6515 21539
rect 6546 21536 6552 21548
rect 6503 21508 6552 21536
rect 6503 21505 6515 21508
rect 6457 21499 6515 21505
rect 6546 21496 6552 21508
rect 6604 21496 6610 21548
rect 4338 21428 4344 21480
rect 4396 21468 4402 21480
rect 7561 21471 7619 21477
rect 7561 21468 7573 21471
rect 4396 21440 7573 21468
rect 4396 21428 4402 21440
rect 7561 21437 7573 21440
rect 7607 21437 7619 21471
rect 7561 21431 7619 21437
rect 8113 21471 8171 21477
rect 8113 21437 8125 21471
rect 8159 21437 8171 21471
rect 8113 21431 8171 21437
rect 6638 21400 6644 21412
rect 3160 21372 6500 21400
rect 6599 21372 6644 21400
rect 3160 21344 3188 21372
rect 3142 21332 3148 21344
rect 3103 21304 3148 21332
rect 3142 21292 3148 21304
rect 3200 21292 3206 21344
rect 3234 21292 3240 21344
rect 3292 21332 3298 21344
rect 3789 21335 3847 21341
rect 3789 21332 3801 21335
rect 3292 21304 3801 21332
rect 3292 21292 3298 21304
rect 3789 21301 3801 21304
rect 3835 21332 3847 21335
rect 5810 21332 5816 21344
rect 3835 21304 5816 21332
rect 3835 21301 3847 21304
rect 3789 21295 3847 21301
rect 5810 21292 5816 21304
rect 5868 21292 5874 21344
rect 6472 21332 6500 21372
rect 6638 21360 6644 21372
rect 6696 21360 6702 21412
rect 7282 21360 7288 21412
rect 7340 21400 7346 21412
rect 7653 21403 7711 21409
rect 7653 21400 7665 21403
rect 7340 21372 7665 21400
rect 7340 21360 7346 21372
rect 7653 21369 7665 21372
rect 7699 21369 7711 21403
rect 7653 21363 7711 21369
rect 8128 21344 8156 21431
rect 8110 21332 8116 21344
rect 6472 21304 8116 21332
rect 8110 21292 8116 21304
rect 8168 21292 8174 21344
rect 1104 21242 8832 21264
rect 1104 21190 2248 21242
rect 2300 21190 2312 21242
rect 2364 21190 2376 21242
rect 2428 21190 2440 21242
rect 2492 21190 2504 21242
rect 2556 21190 4846 21242
rect 4898 21190 4910 21242
rect 4962 21190 4974 21242
rect 5026 21190 5038 21242
rect 5090 21190 5102 21242
rect 5154 21190 7443 21242
rect 7495 21190 7507 21242
rect 7559 21190 7571 21242
rect 7623 21190 7635 21242
rect 7687 21190 7699 21242
rect 7751 21190 8832 21242
rect 1104 21168 8832 21190
rect 3234 21128 3240 21140
rect 3195 21100 3240 21128
rect 3234 21088 3240 21100
rect 3292 21088 3298 21140
rect 6730 21128 6736 21140
rect 4264 21100 6736 21128
rect 2590 21020 2596 21072
rect 2648 21060 2654 21072
rect 4264 21060 4292 21100
rect 6730 21088 6736 21100
rect 6788 21088 6794 21140
rect 2648 21032 4292 21060
rect 4341 21063 4399 21069
rect 2648 21020 2654 21032
rect 4341 21029 4353 21063
rect 4387 21060 4399 21063
rect 7834 21060 7840 21072
rect 4387 21032 5580 21060
rect 7795 21032 7840 21060
rect 4387 21029 4399 21032
rect 4341 21023 4399 21029
rect 5552 21001 5580 21032
rect 7834 21020 7840 21032
rect 7892 21020 7898 21072
rect 5537 20995 5595 21001
rect 5537 20961 5549 20995
rect 5583 20961 5595 20995
rect 5537 20955 5595 20961
rect 5810 20952 5816 21004
rect 5868 20992 5874 21004
rect 6089 20995 6147 21001
rect 6089 20992 6101 20995
rect 5868 20964 6101 20992
rect 5868 20952 5874 20964
rect 6089 20961 6101 20964
rect 6135 20961 6147 20995
rect 6089 20955 6147 20961
rect 4154 20924 4160 20936
rect 4115 20896 4160 20924
rect 4154 20884 4160 20896
rect 4212 20884 4218 20936
rect 4985 20927 5043 20933
rect 4985 20893 4997 20927
rect 5031 20924 5043 20927
rect 6549 20927 6607 20933
rect 5031 20896 6040 20924
rect 5031 20893 5043 20896
rect 4985 20887 5043 20893
rect 5626 20856 5632 20868
rect 5587 20828 5632 20856
rect 5626 20816 5632 20828
rect 5684 20816 5690 20868
rect 6012 20856 6040 20896
rect 6549 20893 6561 20927
rect 6595 20924 6607 20927
rect 6730 20924 6736 20936
rect 6595 20896 6736 20924
rect 6595 20893 6607 20896
rect 6549 20887 6607 20893
rect 6730 20884 6736 20896
rect 6788 20884 6794 20936
rect 6822 20884 6828 20936
rect 6880 20924 6886 20936
rect 7469 20927 7527 20933
rect 7469 20924 7481 20927
rect 6880 20896 7481 20924
rect 6880 20884 6886 20896
rect 7469 20893 7481 20896
rect 7515 20893 7527 20927
rect 7469 20887 7527 20893
rect 7006 20856 7012 20868
rect 6012 20828 7012 20856
rect 7006 20816 7012 20828
rect 7064 20816 7070 20868
rect 2590 20788 2596 20800
rect 2551 20760 2596 20788
rect 2590 20748 2596 20760
rect 2648 20748 2654 20800
rect 4062 20748 4068 20800
rect 4120 20788 4126 20800
rect 4893 20791 4951 20797
rect 4893 20788 4905 20791
rect 4120 20760 4905 20788
rect 4120 20748 4126 20760
rect 4893 20757 4905 20760
rect 4939 20788 4951 20791
rect 6822 20788 6828 20800
rect 4939 20760 6828 20788
rect 4939 20757 4951 20760
rect 4893 20751 4951 20757
rect 6822 20748 6828 20760
rect 6880 20748 6886 20800
rect 1104 20698 8832 20720
rect 1104 20646 3547 20698
rect 3599 20646 3611 20698
rect 3663 20646 3675 20698
rect 3727 20646 3739 20698
rect 3791 20646 3803 20698
rect 3855 20646 6144 20698
rect 6196 20646 6208 20698
rect 6260 20646 6272 20698
rect 6324 20646 6336 20698
rect 6388 20646 6400 20698
rect 6452 20646 8832 20698
rect 1104 20624 8832 20646
rect 3145 20587 3203 20593
rect 3145 20553 3157 20587
rect 3191 20584 3203 20587
rect 4338 20584 4344 20596
rect 3191 20556 4344 20584
rect 3191 20553 3203 20556
rect 3145 20547 3203 20553
rect 4338 20544 4344 20556
rect 4396 20544 4402 20596
rect 4062 20516 4068 20528
rect 2976 20488 4068 20516
rect 2976 20457 3004 20488
rect 4062 20476 4068 20488
rect 4120 20476 4126 20528
rect 4433 20519 4491 20525
rect 4433 20485 4445 20519
rect 4479 20516 4491 20519
rect 5169 20519 5227 20525
rect 5169 20516 5181 20519
rect 4479 20488 5181 20516
rect 4479 20485 4491 20488
rect 4433 20479 4491 20485
rect 5169 20485 5181 20488
rect 5215 20516 5227 20519
rect 5626 20516 5632 20528
rect 5215 20488 5632 20516
rect 5215 20485 5227 20488
rect 5169 20479 5227 20485
rect 5626 20476 5632 20488
rect 5684 20476 5690 20528
rect 2961 20451 3019 20457
rect 2961 20417 2973 20451
rect 3007 20417 3019 20451
rect 2961 20411 3019 20417
rect 3789 20451 3847 20457
rect 3789 20417 3801 20451
rect 3835 20417 3847 20451
rect 3789 20411 3847 20417
rect 3804 20312 3832 20411
rect 4154 20408 4160 20460
rect 4212 20448 4218 20460
rect 4893 20451 4951 20457
rect 4893 20448 4905 20451
rect 4212 20420 4905 20448
rect 4212 20408 4218 20420
rect 4893 20417 4905 20420
rect 4939 20417 4951 20451
rect 5810 20448 5816 20460
rect 5771 20420 5816 20448
rect 4893 20411 4951 20417
rect 4908 20380 4936 20411
rect 5810 20408 5816 20420
rect 5868 20408 5874 20460
rect 6638 20448 6644 20460
rect 6599 20420 6644 20448
rect 6638 20408 6644 20420
rect 6696 20408 6702 20460
rect 7190 20408 7196 20460
rect 7248 20448 7254 20460
rect 7929 20451 7987 20457
rect 7929 20448 7941 20451
rect 7248 20420 7941 20448
rect 7248 20408 7254 20420
rect 7929 20417 7941 20420
rect 7975 20417 7987 20451
rect 7929 20411 7987 20417
rect 6656 20380 6684 20408
rect 4908 20352 6684 20380
rect 6454 20312 6460 20324
rect 3804 20284 6316 20312
rect 6415 20284 6460 20312
rect 2501 20247 2559 20253
rect 2501 20213 2513 20247
rect 2547 20244 2559 20247
rect 2682 20244 2688 20256
rect 2547 20216 2688 20244
rect 2547 20213 2559 20216
rect 2501 20207 2559 20213
rect 2682 20204 2688 20216
rect 2740 20204 2746 20256
rect 3697 20247 3755 20253
rect 3697 20213 3709 20247
rect 3743 20244 3755 20247
rect 4246 20244 4252 20256
rect 3743 20216 4252 20244
rect 3743 20213 3755 20216
rect 3697 20207 3755 20213
rect 4246 20204 4252 20216
rect 4304 20204 4310 20256
rect 4341 20247 4399 20253
rect 4341 20213 4353 20247
rect 4387 20244 4399 20247
rect 5994 20244 6000 20256
rect 4387 20216 6000 20244
rect 4387 20213 4399 20216
rect 4341 20207 4399 20213
rect 5994 20204 6000 20216
rect 6052 20204 6058 20256
rect 6288 20244 6316 20284
rect 6454 20272 6460 20284
rect 6512 20272 6518 20324
rect 7282 20244 7288 20256
rect 6288 20216 7288 20244
rect 7282 20204 7288 20216
rect 7340 20204 7346 20256
rect 1104 20154 8832 20176
rect 1104 20102 2248 20154
rect 2300 20102 2312 20154
rect 2364 20102 2376 20154
rect 2428 20102 2440 20154
rect 2492 20102 2504 20154
rect 2556 20102 4846 20154
rect 4898 20102 4910 20154
rect 4962 20102 4974 20154
rect 5026 20102 5038 20154
rect 5090 20102 5102 20154
rect 5154 20102 7443 20154
rect 7495 20102 7507 20154
rect 7559 20102 7571 20154
rect 7623 20102 7635 20154
rect 7687 20102 7699 20154
rect 7751 20102 8832 20154
rect 1104 20080 8832 20102
rect 2685 20043 2743 20049
rect 2685 20009 2697 20043
rect 2731 20040 2743 20043
rect 3142 20040 3148 20052
rect 2731 20012 3148 20040
rect 2731 20009 2743 20012
rect 2685 20003 2743 20009
rect 3142 20000 3148 20012
rect 3200 20000 3206 20052
rect 4249 20043 4307 20049
rect 4249 20009 4261 20043
rect 4295 20040 4307 20043
rect 4338 20040 4344 20052
rect 4295 20012 4344 20040
rect 4295 20009 4307 20012
rect 4249 20003 4307 20009
rect 4338 20000 4344 20012
rect 4396 20000 4402 20052
rect 4062 19864 4068 19916
rect 4120 19904 4126 19916
rect 6457 19907 6515 19913
rect 4120 19876 5856 19904
rect 4120 19864 4126 19876
rect 2958 19796 2964 19848
rect 3016 19836 3022 19848
rect 3237 19839 3295 19845
rect 3237 19836 3249 19839
rect 3016 19808 3249 19836
rect 3016 19796 3022 19808
rect 3237 19805 3249 19808
rect 3283 19836 3295 19839
rect 4893 19839 4951 19845
rect 4893 19836 4905 19839
rect 3283 19808 4905 19836
rect 3283 19805 3295 19808
rect 3237 19799 3295 19805
rect 4893 19805 4905 19808
rect 4939 19836 4951 19839
rect 5534 19836 5540 19848
rect 4939 19808 5540 19836
rect 4939 19805 4951 19808
rect 4893 19799 4951 19805
rect 5534 19796 5540 19808
rect 5592 19796 5598 19848
rect 5828 19845 5856 19876
rect 6457 19873 6469 19907
rect 6503 19904 6515 19907
rect 6546 19904 6552 19916
rect 6503 19876 6552 19904
rect 6503 19873 6515 19876
rect 6457 19867 6515 19873
rect 6546 19864 6552 19876
rect 6604 19864 6610 19916
rect 5813 19839 5871 19845
rect 5813 19805 5825 19839
rect 5859 19805 5871 19839
rect 5813 19799 5871 19805
rect 6822 19796 6828 19848
rect 6880 19836 6886 19848
rect 7193 19839 7251 19845
rect 7193 19836 7205 19839
rect 6880 19808 7205 19836
rect 6880 19796 6886 19808
rect 7193 19805 7205 19808
rect 7239 19805 7251 19839
rect 7193 19799 7251 19805
rect 7282 19796 7288 19848
rect 7340 19836 7346 19848
rect 7377 19839 7435 19845
rect 7377 19836 7389 19839
rect 7340 19808 7389 19836
rect 7340 19796 7346 19808
rect 7377 19805 7389 19808
rect 7423 19805 7435 19839
rect 8110 19836 8116 19848
rect 8071 19808 8116 19836
rect 7377 19799 7435 19805
rect 8110 19796 8116 19808
rect 8168 19796 8174 19848
rect 4341 19771 4399 19777
rect 4341 19737 4353 19771
rect 4387 19768 4399 19771
rect 6454 19768 6460 19780
rect 4387 19740 6460 19768
rect 4387 19737 4399 19740
rect 4341 19731 4399 19737
rect 6454 19728 6460 19740
rect 6512 19768 6518 19780
rect 6638 19768 6644 19780
rect 6512 19740 6644 19768
rect 6512 19728 6518 19740
rect 6638 19728 6644 19740
rect 6696 19728 6702 19780
rect 1578 19700 1584 19712
rect 1539 19672 1584 19700
rect 1578 19660 1584 19672
rect 1636 19660 1642 19712
rect 2038 19700 2044 19712
rect 1999 19672 2044 19700
rect 2038 19660 2044 19672
rect 2096 19660 2102 19712
rect 1104 19610 8832 19632
rect 1104 19558 3547 19610
rect 3599 19558 3611 19610
rect 3663 19558 3675 19610
rect 3727 19558 3739 19610
rect 3791 19558 3803 19610
rect 3855 19558 6144 19610
rect 6196 19558 6208 19610
rect 6260 19558 6272 19610
rect 6324 19558 6336 19610
rect 6388 19558 6400 19610
rect 6452 19558 8832 19610
rect 1104 19536 8832 19558
rect 2958 19496 2964 19508
rect 2919 19468 2964 19496
rect 2958 19456 2964 19468
rect 3016 19456 3022 19508
rect 4062 19496 4068 19508
rect 4023 19468 4068 19496
rect 4062 19456 4068 19468
rect 4120 19456 4126 19508
rect 4246 19456 4252 19508
rect 4304 19496 4310 19508
rect 4304 19468 7604 19496
rect 4304 19456 4310 19468
rect 6457 19431 6515 19437
rect 6457 19397 6469 19431
rect 6503 19428 6515 19431
rect 6546 19428 6552 19440
rect 6503 19400 6552 19428
rect 6503 19397 6515 19400
rect 6457 19391 6515 19397
rect 6546 19388 6552 19400
rect 6604 19388 6610 19440
rect 7576 19437 7604 19468
rect 7561 19431 7619 19437
rect 7561 19397 7573 19431
rect 7607 19397 7619 19431
rect 7561 19391 7619 19397
rect 4157 19363 4215 19369
rect 4157 19329 4169 19363
rect 4203 19360 4215 19363
rect 4430 19360 4436 19372
rect 4203 19332 4436 19360
rect 4203 19329 4215 19332
rect 4157 19323 4215 19329
rect 4430 19320 4436 19332
rect 4488 19360 4494 19372
rect 4801 19363 4859 19369
rect 4801 19360 4813 19363
rect 4488 19332 4813 19360
rect 4488 19320 4494 19332
rect 4801 19329 4813 19332
rect 4847 19329 4859 19363
rect 4801 19323 4859 19329
rect 5261 19363 5319 19369
rect 5261 19329 5273 19363
rect 5307 19329 5319 19363
rect 5261 19323 5319 19329
rect 2409 19295 2467 19301
rect 2409 19261 2421 19295
rect 2455 19292 2467 19295
rect 2590 19292 2596 19304
rect 2455 19264 2596 19292
rect 2455 19261 2467 19264
rect 2409 19255 2467 19261
rect 2590 19252 2596 19264
rect 2648 19252 2654 19304
rect 4706 19292 4712 19304
rect 4667 19264 4712 19292
rect 4706 19252 4712 19264
rect 4764 19252 4770 19304
rect 1578 19184 1584 19236
rect 1636 19224 1642 19236
rect 1857 19227 1915 19233
rect 1857 19224 1869 19227
rect 1636 19196 1869 19224
rect 1636 19184 1642 19196
rect 1857 19193 1869 19196
rect 1903 19224 1915 19227
rect 1903 19196 2774 19224
rect 1903 19193 1915 19196
rect 1857 19187 1915 19193
rect 2746 19156 2774 19196
rect 3234 19184 3240 19236
rect 3292 19224 3298 19236
rect 3513 19227 3571 19233
rect 3513 19224 3525 19227
rect 3292 19196 3525 19224
rect 3292 19184 3298 19196
rect 3513 19193 3525 19196
rect 3559 19224 3571 19227
rect 5276 19224 5304 19323
rect 5534 19320 5540 19372
rect 5592 19360 5598 19372
rect 5592 19332 6500 19360
rect 5592 19320 5598 19332
rect 5626 19252 5632 19304
rect 5684 19292 5690 19304
rect 6365 19295 6423 19301
rect 6365 19292 6377 19295
rect 5684 19264 6377 19292
rect 5684 19252 5690 19264
rect 6365 19261 6377 19264
rect 6411 19261 6423 19295
rect 6472 19292 6500 19332
rect 6730 19320 6736 19372
rect 6788 19360 6794 19372
rect 8113 19363 8171 19369
rect 8113 19360 8125 19363
rect 6788 19332 8125 19360
rect 6788 19320 6794 19332
rect 8113 19329 8125 19332
rect 8159 19329 8171 19363
rect 8113 19323 8171 19329
rect 6917 19295 6975 19301
rect 6917 19292 6929 19295
rect 6472 19264 6929 19292
rect 6365 19255 6423 19261
rect 5718 19224 5724 19236
rect 3559 19196 5724 19224
rect 3559 19193 3571 19196
rect 3513 19187 3571 19193
rect 5718 19184 5724 19196
rect 5776 19184 5782 19236
rect 6840 19168 6868 19264
rect 6917 19261 6929 19264
rect 6963 19261 6975 19295
rect 6917 19255 6975 19261
rect 7653 19295 7711 19301
rect 7653 19261 7665 19295
rect 7699 19292 7711 19295
rect 7834 19292 7840 19304
rect 7699 19264 7840 19292
rect 7699 19261 7711 19264
rect 7653 19255 7711 19261
rect 7834 19252 7840 19264
rect 7892 19252 7898 19304
rect 5534 19156 5540 19168
rect 2746 19128 5540 19156
rect 5534 19116 5540 19128
rect 5592 19116 5598 19168
rect 5810 19156 5816 19168
rect 5771 19128 5816 19156
rect 5810 19116 5816 19128
rect 5868 19116 5874 19168
rect 6822 19116 6828 19168
rect 6880 19116 6886 19168
rect 1104 19066 8832 19088
rect 1104 19014 2248 19066
rect 2300 19014 2312 19066
rect 2364 19014 2376 19066
rect 2428 19014 2440 19066
rect 2492 19014 2504 19066
rect 2556 19014 4846 19066
rect 4898 19014 4910 19066
rect 4962 19014 4974 19066
rect 5026 19014 5038 19066
rect 5090 19014 5102 19066
rect 5154 19014 7443 19066
rect 7495 19014 7507 19066
rect 7559 19014 7571 19066
rect 7623 19014 7635 19066
rect 7687 19014 7699 19066
rect 7751 19014 8832 19066
rect 1104 18992 8832 19014
rect 2682 18952 2688 18964
rect 2595 18924 2688 18952
rect 2682 18912 2688 18924
rect 2740 18952 2746 18964
rect 7190 18952 7196 18964
rect 2740 18924 7196 18952
rect 2740 18912 2746 18924
rect 7190 18912 7196 18924
rect 7248 18912 7254 18964
rect 3234 18884 3240 18896
rect 3195 18856 3240 18884
rect 3234 18844 3240 18856
rect 3292 18844 3298 18896
rect 4430 18884 4436 18896
rect 4391 18856 4436 18884
rect 4430 18844 4436 18856
rect 4488 18844 4494 18896
rect 6549 18887 6607 18893
rect 6549 18853 6561 18887
rect 6595 18884 6607 18887
rect 6638 18884 6644 18896
rect 6595 18856 6644 18884
rect 6595 18853 6607 18856
rect 6549 18847 6607 18853
rect 6638 18844 6644 18856
rect 6696 18844 6702 18896
rect 5994 18776 6000 18828
rect 6052 18816 6058 18828
rect 6457 18819 6515 18825
rect 6457 18816 6469 18819
rect 6052 18788 6469 18816
rect 6052 18776 6058 18788
rect 6457 18785 6469 18788
rect 6503 18785 6515 18819
rect 6457 18779 6515 18785
rect 8018 18776 8024 18828
rect 8076 18816 8082 18828
rect 8113 18819 8171 18825
rect 8113 18816 8125 18819
rect 8076 18788 8125 18816
rect 8076 18776 8082 18788
rect 8113 18785 8125 18788
rect 8159 18785 8171 18819
rect 8113 18779 8171 18785
rect 4430 18748 4436 18760
rect 4391 18720 4436 18748
rect 4430 18708 4436 18720
rect 4488 18708 4494 18760
rect 5718 18748 5724 18760
rect 5631 18720 5724 18748
rect 5718 18708 5724 18720
rect 5776 18748 5782 18760
rect 6546 18748 6552 18760
rect 5776 18720 6552 18748
rect 5776 18708 5782 18720
rect 6546 18708 6552 18720
rect 6604 18708 6610 18760
rect 7009 18751 7067 18757
rect 7009 18717 7021 18751
rect 7055 18748 7067 18751
rect 7190 18748 7196 18760
rect 7055 18720 7196 18748
rect 7055 18717 7067 18720
rect 7009 18711 7067 18717
rect 7190 18708 7196 18720
rect 7248 18708 7254 18760
rect 7282 18708 7288 18760
rect 7340 18748 7346 18760
rect 7653 18751 7711 18757
rect 7653 18748 7665 18751
rect 7340 18720 7665 18748
rect 7340 18708 7346 18720
rect 7653 18717 7665 18720
rect 7699 18717 7711 18751
rect 7653 18711 7711 18717
rect 1581 18683 1639 18689
rect 1581 18649 1593 18683
rect 1627 18680 1639 18683
rect 2038 18680 2044 18692
rect 1627 18652 2044 18680
rect 1627 18649 1639 18652
rect 1581 18643 1639 18649
rect 2038 18640 2044 18652
rect 2096 18680 2102 18692
rect 2774 18680 2780 18692
rect 2096 18652 2780 18680
rect 2096 18640 2102 18652
rect 2774 18640 2780 18652
rect 2832 18640 2838 18692
rect 7098 18640 7104 18692
rect 7156 18680 7162 18692
rect 7561 18683 7619 18689
rect 7561 18680 7573 18683
rect 7156 18652 7573 18680
rect 7156 18640 7162 18652
rect 7561 18649 7573 18652
rect 7607 18649 7619 18683
rect 7561 18643 7619 18649
rect 2130 18612 2136 18624
rect 2091 18584 2136 18612
rect 2130 18572 2136 18584
rect 2188 18572 2194 18624
rect 1104 18522 8832 18544
rect 1104 18470 3547 18522
rect 3599 18470 3611 18522
rect 3663 18470 3675 18522
rect 3727 18470 3739 18522
rect 3791 18470 3803 18522
rect 3855 18470 6144 18522
rect 6196 18470 6208 18522
rect 6260 18470 6272 18522
rect 6324 18470 6336 18522
rect 6388 18470 6400 18522
rect 6452 18470 8832 18522
rect 1104 18448 8832 18470
rect 3789 18411 3847 18417
rect 3789 18377 3801 18411
rect 3835 18408 3847 18411
rect 4706 18408 4712 18420
rect 3835 18380 4712 18408
rect 3835 18377 3847 18380
rect 3789 18371 3847 18377
rect 4706 18368 4712 18380
rect 4764 18368 4770 18420
rect 5810 18408 5816 18420
rect 5092 18380 5816 18408
rect 3881 18343 3939 18349
rect 3881 18309 3893 18343
rect 3927 18340 3939 18343
rect 4525 18343 4583 18349
rect 4525 18340 4537 18343
rect 3927 18312 4537 18340
rect 3927 18309 3939 18312
rect 3881 18303 3939 18309
rect 4525 18309 4537 18312
rect 4571 18340 4583 18343
rect 4614 18340 4620 18352
rect 4571 18312 4620 18340
rect 4571 18309 4583 18312
rect 4525 18303 4583 18309
rect 4614 18300 4620 18312
rect 4672 18300 4678 18352
rect 3237 18275 3295 18281
rect 3237 18241 3249 18275
rect 3283 18241 3295 18275
rect 3237 18235 3295 18241
rect 4341 18275 4399 18281
rect 4341 18241 4353 18275
rect 4387 18272 4399 18275
rect 4430 18272 4436 18284
rect 4387 18244 4436 18272
rect 4387 18241 4399 18244
rect 4341 18235 4399 18241
rect 3252 18136 3280 18235
rect 4356 18204 4384 18235
rect 4430 18232 4436 18244
rect 4488 18232 4494 18284
rect 5092 18272 5120 18380
rect 5810 18368 5816 18380
rect 5868 18368 5874 18420
rect 5166 18300 5172 18352
rect 5224 18340 5230 18352
rect 7561 18343 7619 18349
rect 7561 18340 7573 18343
rect 5224 18312 7573 18340
rect 5224 18300 5230 18312
rect 7561 18309 7573 18312
rect 7607 18309 7619 18343
rect 7561 18303 7619 18309
rect 5261 18275 5319 18281
rect 5261 18272 5273 18275
rect 5092 18244 5273 18272
rect 5261 18241 5273 18244
rect 5307 18241 5319 18275
rect 5718 18272 5724 18284
rect 5261 18235 5319 18241
rect 5368 18244 5724 18272
rect 5368 18204 5396 18244
rect 5718 18232 5724 18244
rect 5776 18232 5782 18284
rect 6914 18272 6920 18284
rect 6827 18244 6920 18272
rect 6914 18232 6920 18244
rect 6972 18272 6978 18284
rect 7834 18272 7840 18284
rect 6972 18244 7840 18272
rect 6972 18232 6978 18244
rect 7834 18232 7840 18244
rect 7892 18232 7898 18284
rect 8113 18275 8171 18281
rect 8113 18241 8125 18275
rect 8159 18272 8171 18275
rect 8202 18272 8208 18284
rect 8159 18244 8208 18272
rect 8159 18241 8171 18244
rect 8113 18235 8171 18241
rect 8202 18232 8208 18244
rect 8260 18232 8266 18284
rect 4356 18176 5396 18204
rect 5534 18164 5540 18216
rect 5592 18204 5598 18216
rect 6365 18207 6423 18213
rect 6365 18204 6377 18207
rect 5592 18176 6377 18204
rect 5592 18164 5598 18176
rect 6365 18173 6377 18176
rect 6411 18173 6423 18207
rect 6365 18167 6423 18173
rect 7006 18164 7012 18216
rect 7064 18204 7070 18216
rect 7653 18207 7711 18213
rect 7653 18204 7665 18207
rect 7064 18176 7665 18204
rect 7064 18164 7070 18176
rect 7653 18173 7665 18176
rect 7699 18173 7711 18207
rect 7653 18167 7711 18173
rect 5350 18136 5356 18148
rect 3252 18108 5356 18136
rect 5350 18096 5356 18108
rect 5408 18136 5414 18148
rect 6457 18139 6515 18145
rect 6457 18136 6469 18139
rect 5408 18108 6469 18136
rect 5408 18096 5414 18108
rect 6457 18105 6469 18108
rect 6503 18105 6515 18139
rect 6457 18099 6515 18105
rect 1489 18071 1547 18077
rect 1489 18037 1501 18071
rect 1535 18068 1547 18071
rect 1670 18068 1676 18080
rect 1535 18040 1676 18068
rect 1535 18037 1547 18040
rect 1489 18031 1547 18037
rect 1670 18028 1676 18040
rect 1728 18028 1734 18080
rect 2038 18068 2044 18080
rect 1999 18040 2044 18068
rect 2038 18028 2044 18040
rect 2096 18028 2102 18080
rect 2590 18068 2596 18080
rect 2551 18040 2596 18068
rect 2590 18028 2596 18040
rect 2648 18028 2654 18080
rect 3145 18071 3203 18077
rect 3145 18037 3157 18071
rect 3191 18068 3203 18071
rect 5626 18068 5632 18080
rect 3191 18040 5632 18068
rect 3191 18037 3203 18040
rect 3145 18031 3203 18037
rect 5626 18028 5632 18040
rect 5684 18028 5690 18080
rect 5813 18071 5871 18077
rect 5813 18037 5825 18071
rect 5859 18068 5871 18071
rect 5902 18068 5908 18080
rect 5859 18040 5908 18068
rect 5859 18037 5871 18040
rect 5813 18031 5871 18037
rect 5902 18028 5908 18040
rect 5960 18028 5966 18080
rect 1104 17978 8832 18000
rect 1104 17926 2248 17978
rect 2300 17926 2312 17978
rect 2364 17926 2376 17978
rect 2428 17926 2440 17978
rect 2492 17926 2504 17978
rect 2556 17926 4846 17978
rect 4898 17926 4910 17978
rect 4962 17926 4974 17978
rect 5026 17926 5038 17978
rect 5090 17926 5102 17978
rect 5154 17926 7443 17978
rect 7495 17926 7507 17978
rect 7559 17926 7571 17978
rect 7623 17926 7635 17978
rect 7687 17926 7699 17978
rect 7751 17926 8832 17978
rect 1104 17904 8832 17926
rect 2590 17864 2596 17876
rect 2551 17836 2596 17864
rect 2590 17824 2596 17836
rect 2648 17824 2654 17876
rect 3237 17867 3295 17873
rect 3237 17833 3249 17867
rect 3283 17864 3295 17867
rect 3970 17864 3976 17876
rect 3283 17836 3976 17864
rect 3283 17833 3295 17836
rect 3237 17827 3295 17833
rect 3970 17824 3976 17836
rect 4028 17864 4034 17876
rect 5810 17864 5816 17876
rect 4028 17836 5816 17864
rect 4028 17824 4034 17836
rect 5810 17824 5816 17836
rect 5868 17824 5874 17876
rect 2038 17756 2044 17808
rect 2096 17796 2102 17808
rect 2133 17799 2191 17805
rect 2133 17796 2145 17799
rect 2096 17768 2145 17796
rect 2096 17756 2102 17768
rect 2133 17765 2145 17768
rect 2179 17796 2191 17799
rect 6825 17799 6883 17805
rect 2179 17768 6776 17796
rect 2179 17765 2191 17768
rect 2133 17759 2191 17765
rect 2590 17688 2596 17740
rect 2648 17728 2654 17740
rect 4522 17728 4528 17740
rect 2648 17700 4528 17728
rect 2648 17688 2654 17700
rect 4522 17688 4528 17700
rect 4580 17688 4586 17740
rect 4614 17688 4620 17740
rect 4672 17728 4678 17740
rect 4672 17700 4717 17728
rect 4672 17688 4678 17700
rect 4798 17688 4804 17740
rect 4856 17728 4862 17740
rect 6748 17728 6776 17768
rect 6825 17765 6837 17799
rect 6871 17796 6883 17799
rect 7006 17796 7012 17808
rect 6871 17768 7012 17796
rect 6871 17765 6883 17768
rect 6825 17759 6883 17765
rect 7006 17756 7012 17768
rect 7064 17756 7070 17808
rect 4856 17700 6132 17728
rect 6748 17700 8156 17728
rect 4856 17688 4862 17700
rect 3970 17620 3976 17672
rect 4028 17660 4034 17672
rect 4157 17663 4215 17669
rect 4157 17660 4169 17663
rect 4028 17632 4169 17660
rect 4028 17620 4034 17632
rect 4157 17629 4169 17632
rect 4203 17629 4215 17663
rect 4157 17623 4215 17629
rect 4709 17663 4767 17669
rect 4709 17629 4721 17663
rect 4755 17660 4767 17663
rect 5350 17660 5356 17672
rect 4755 17632 4844 17660
rect 5311 17632 5356 17660
rect 4755 17629 4767 17632
rect 4709 17623 4767 17629
rect 1670 17552 1676 17604
rect 1728 17592 1734 17604
rect 4430 17592 4436 17604
rect 1728 17564 4436 17592
rect 1728 17552 1734 17564
rect 4430 17552 4436 17564
rect 4488 17552 4494 17604
rect 4816 17536 4844 17632
rect 5350 17620 5356 17632
rect 5408 17620 5414 17672
rect 6104 17669 6132 17700
rect 6089 17663 6147 17669
rect 6089 17629 6101 17663
rect 6135 17660 6147 17663
rect 6914 17660 6920 17672
rect 6135 17632 6920 17660
rect 6135 17629 6147 17632
rect 6089 17623 6147 17629
rect 6914 17620 6920 17632
rect 6972 17620 6978 17672
rect 7190 17660 7196 17672
rect 7151 17632 7196 17660
rect 7190 17620 7196 17632
rect 7248 17620 7254 17672
rect 8128 17669 8156 17700
rect 8113 17663 8171 17669
rect 8113 17629 8125 17663
rect 8159 17660 8171 17663
rect 8202 17660 8208 17672
rect 8159 17632 8208 17660
rect 8159 17629 8171 17632
rect 8113 17623 8171 17629
rect 8202 17620 8208 17632
rect 8260 17620 8266 17672
rect 5074 17552 5080 17604
rect 5132 17592 5138 17604
rect 5169 17595 5227 17601
rect 5169 17592 5181 17595
rect 5132 17564 5181 17592
rect 5132 17552 5138 17564
rect 5169 17561 5181 17564
rect 5215 17561 5227 17595
rect 5169 17555 5227 17561
rect 5258 17552 5264 17604
rect 5316 17592 5322 17604
rect 7926 17592 7932 17604
rect 5316 17564 7932 17592
rect 5316 17552 5322 17564
rect 7926 17552 7932 17564
rect 7984 17552 7990 17604
rect 1578 17524 1584 17536
rect 1539 17496 1584 17524
rect 1578 17484 1584 17496
rect 1636 17484 1642 17536
rect 4798 17484 4804 17536
rect 4856 17484 4862 17536
rect 1104 17434 8832 17456
rect 1104 17382 3547 17434
rect 3599 17382 3611 17434
rect 3663 17382 3675 17434
rect 3727 17382 3739 17434
rect 3791 17382 3803 17434
rect 3855 17382 6144 17434
rect 6196 17382 6208 17434
rect 6260 17382 6272 17434
rect 6324 17382 6336 17434
rect 6388 17382 6400 17434
rect 6452 17382 8832 17434
rect 1104 17360 8832 17382
rect 1670 17320 1676 17332
rect 1631 17292 1676 17320
rect 1670 17280 1676 17292
rect 1728 17280 1734 17332
rect 4798 17320 4804 17332
rect 4759 17292 4804 17320
rect 4798 17280 4804 17292
rect 4856 17280 4862 17332
rect 4338 17252 4344 17264
rect 3344 17224 4344 17252
rect 2866 17184 2872 17196
rect 2827 17156 2872 17184
rect 2866 17144 2872 17156
rect 2924 17144 2930 17196
rect 3344 17193 3372 17224
rect 4338 17212 4344 17224
rect 4396 17212 4402 17264
rect 4430 17212 4436 17264
rect 4488 17252 4494 17264
rect 5353 17255 5411 17261
rect 5353 17252 5365 17255
rect 4488 17224 5365 17252
rect 4488 17212 4494 17224
rect 5353 17221 5365 17224
rect 5399 17252 5411 17255
rect 6549 17255 6607 17261
rect 6549 17252 6561 17255
rect 5399 17224 6561 17252
rect 5399 17221 5411 17224
rect 5353 17215 5411 17221
rect 6549 17221 6561 17224
rect 6595 17221 6607 17255
rect 6549 17215 6607 17221
rect 3329 17187 3387 17193
rect 3329 17153 3341 17187
rect 3375 17153 3387 17187
rect 3329 17147 3387 17153
rect 3973 17187 4031 17193
rect 3973 17153 3985 17187
rect 4019 17184 4031 17187
rect 4062 17184 4068 17196
rect 4019 17156 4068 17184
rect 4019 17153 4031 17156
rect 3973 17147 4031 17153
rect 4062 17144 4068 17156
rect 4120 17144 4126 17196
rect 4617 17187 4675 17193
rect 4617 17153 4629 17187
rect 4663 17184 4675 17187
rect 5626 17184 5632 17196
rect 4663 17156 5632 17184
rect 4663 17153 4675 17156
rect 4617 17147 4675 17153
rect 5626 17144 5632 17156
rect 5684 17144 5690 17196
rect 6362 17184 6368 17196
rect 6323 17156 6368 17184
rect 6362 17144 6368 17156
rect 6420 17144 6426 17196
rect 6730 17144 6736 17196
rect 6788 17184 6794 17196
rect 7285 17187 7343 17193
rect 7285 17184 7297 17187
rect 6788 17156 7297 17184
rect 6788 17144 6794 17156
rect 7285 17153 7297 17156
rect 7331 17153 7343 17187
rect 7285 17147 7343 17153
rect 7834 17144 7840 17196
rect 7892 17184 7898 17196
rect 7929 17187 7987 17193
rect 7929 17184 7941 17187
rect 7892 17156 7941 17184
rect 7892 17144 7898 17156
rect 7929 17153 7941 17156
rect 7975 17153 7987 17187
rect 7929 17147 7987 17153
rect 2777 17119 2835 17125
rect 2777 17085 2789 17119
rect 2823 17116 2835 17119
rect 5166 17116 5172 17128
rect 2823 17088 5172 17116
rect 2823 17085 2835 17088
rect 2777 17079 2835 17085
rect 5166 17076 5172 17088
rect 5224 17076 5230 17128
rect 5261 17119 5319 17125
rect 5261 17085 5273 17119
rect 5307 17085 5319 17119
rect 5261 17079 5319 17085
rect 2225 17051 2283 17057
rect 2225 17017 2237 17051
rect 2271 17048 2283 17051
rect 2590 17048 2596 17060
rect 2271 17020 2596 17048
rect 2271 17017 2283 17020
rect 2225 17011 2283 17017
rect 2590 17008 2596 17020
rect 2648 17008 2654 17060
rect 3513 17051 3571 17057
rect 3513 17017 3525 17051
rect 3559 17048 3571 17051
rect 5276 17048 5304 17079
rect 5350 17076 5356 17128
rect 5408 17116 5414 17128
rect 5813 17119 5871 17125
rect 5813 17116 5825 17119
rect 5408 17088 5825 17116
rect 5408 17076 5414 17088
rect 5813 17085 5825 17088
rect 5859 17116 5871 17119
rect 6748 17116 6776 17144
rect 5859 17088 6776 17116
rect 5859 17085 5871 17088
rect 5813 17079 5871 17085
rect 3559 17020 5304 17048
rect 3559 17017 3571 17020
rect 3513 17011 3571 17017
rect 7190 17008 7196 17060
rect 7248 17048 7254 17060
rect 7745 17051 7803 17057
rect 7745 17048 7757 17051
rect 7248 17020 7757 17048
rect 7248 17008 7254 17020
rect 7745 17017 7757 17020
rect 7791 17017 7803 17051
rect 7745 17011 7803 17017
rect 4157 16983 4215 16989
rect 4157 16949 4169 16983
rect 4203 16980 4215 16983
rect 5534 16980 5540 16992
rect 4203 16952 5540 16980
rect 4203 16949 4215 16952
rect 4157 16943 4215 16949
rect 5534 16940 5540 16952
rect 5592 16940 5598 16992
rect 1104 16890 8832 16912
rect 1104 16838 2248 16890
rect 2300 16838 2312 16890
rect 2364 16838 2376 16890
rect 2428 16838 2440 16890
rect 2492 16838 2504 16890
rect 2556 16838 4846 16890
rect 4898 16838 4910 16890
rect 4962 16838 4974 16890
rect 5026 16838 5038 16890
rect 5090 16838 5102 16890
rect 5154 16838 7443 16890
rect 7495 16838 7507 16890
rect 7559 16838 7571 16890
rect 7623 16838 7635 16890
rect 7687 16838 7699 16890
rect 7751 16838 8832 16890
rect 1104 16816 8832 16838
rect 2590 16776 2596 16788
rect 2551 16748 2596 16776
rect 2590 16736 2596 16748
rect 2648 16736 2654 16788
rect 2866 16736 2872 16788
rect 2924 16776 2930 16788
rect 7282 16776 7288 16788
rect 2924 16748 7288 16776
rect 2924 16736 2930 16748
rect 7282 16736 7288 16748
rect 7340 16736 7346 16788
rect 1489 16711 1547 16717
rect 1489 16677 1501 16711
rect 1535 16708 1547 16711
rect 1578 16708 1584 16720
rect 1535 16680 1584 16708
rect 1535 16677 1547 16680
rect 1489 16671 1547 16677
rect 1578 16668 1584 16680
rect 1636 16708 1642 16720
rect 6730 16708 6736 16720
rect 1636 16680 6736 16708
rect 1636 16668 1642 16680
rect 6730 16668 6736 16680
rect 6788 16668 6794 16720
rect 4062 16600 4068 16652
rect 4120 16640 4126 16652
rect 4120 16612 4292 16640
rect 4120 16600 4126 16612
rect 3053 16575 3111 16581
rect 3053 16541 3065 16575
rect 3099 16572 3111 16575
rect 3970 16572 3976 16584
rect 3099 16544 3976 16572
rect 3099 16541 3111 16544
rect 3053 16535 3111 16541
rect 3970 16532 3976 16544
rect 4028 16532 4034 16584
rect 4264 16581 4292 16612
rect 4338 16600 4344 16652
rect 4396 16640 4402 16652
rect 4396 16612 6408 16640
rect 4396 16600 4402 16612
rect 6380 16584 6408 16612
rect 4249 16575 4307 16581
rect 4249 16541 4261 16575
rect 4295 16541 4307 16575
rect 4430 16572 4436 16584
rect 4391 16544 4436 16572
rect 4249 16535 4307 16541
rect 4430 16532 4436 16544
rect 4488 16532 4494 16584
rect 4522 16532 4528 16584
rect 4580 16572 4586 16584
rect 4985 16575 5043 16581
rect 4985 16572 4997 16575
rect 4580 16544 4997 16572
rect 4580 16532 4586 16544
rect 4985 16541 4997 16544
rect 5031 16541 5043 16575
rect 4985 16535 5043 16541
rect 5445 16575 5503 16581
rect 5445 16541 5457 16575
rect 5491 16572 5503 16575
rect 5718 16572 5724 16584
rect 5491 16544 5724 16572
rect 5491 16541 5503 16544
rect 5445 16535 5503 16541
rect 5718 16532 5724 16544
rect 5776 16532 5782 16584
rect 5994 16532 6000 16584
rect 6052 16572 6058 16584
rect 6181 16575 6239 16581
rect 6181 16572 6193 16575
rect 6052 16544 6193 16572
rect 6052 16532 6058 16544
rect 6181 16541 6193 16544
rect 6227 16541 6239 16575
rect 6181 16535 6239 16541
rect 6362 16532 6368 16584
rect 6420 16572 6426 16584
rect 7101 16575 7159 16581
rect 7101 16572 7113 16575
rect 6420 16544 7113 16572
rect 6420 16532 6426 16544
rect 7101 16541 7113 16544
rect 7147 16541 7159 16575
rect 7101 16535 7159 16541
rect 3878 16464 3884 16516
rect 3936 16504 3942 16516
rect 4893 16507 4951 16513
rect 4893 16504 4905 16507
rect 3936 16476 4905 16504
rect 3936 16464 3942 16476
rect 4893 16473 4905 16476
rect 4939 16473 4951 16507
rect 4893 16467 4951 16473
rect 5534 16464 5540 16516
rect 5592 16504 5598 16516
rect 5902 16504 5908 16516
rect 5592 16476 5908 16504
rect 5592 16464 5598 16476
rect 5902 16464 5908 16476
rect 5960 16464 5966 16516
rect 7745 16507 7803 16513
rect 7745 16473 7757 16507
rect 7791 16504 7803 16507
rect 7834 16504 7840 16516
rect 7791 16476 7840 16504
rect 7791 16473 7803 16476
rect 7745 16467 7803 16473
rect 7834 16464 7840 16476
rect 7892 16464 7898 16516
rect 2041 16439 2099 16445
rect 2041 16405 2053 16439
rect 2087 16436 2099 16439
rect 2590 16436 2596 16448
rect 2087 16408 2596 16436
rect 2087 16405 2099 16408
rect 2041 16399 2099 16405
rect 2590 16396 2596 16408
rect 2648 16396 2654 16448
rect 3237 16439 3295 16445
rect 3237 16405 3249 16439
rect 3283 16436 3295 16439
rect 7098 16436 7104 16448
rect 3283 16408 7104 16436
rect 3283 16405 3295 16408
rect 3237 16399 3295 16405
rect 7098 16396 7104 16408
rect 7156 16396 7162 16448
rect 1104 16346 8832 16368
rect 1104 16294 3547 16346
rect 3599 16294 3611 16346
rect 3663 16294 3675 16346
rect 3727 16294 3739 16346
rect 3791 16294 3803 16346
rect 3855 16294 6144 16346
rect 6196 16294 6208 16346
rect 6260 16294 6272 16346
rect 6324 16294 6336 16346
rect 6388 16294 6400 16346
rect 6452 16294 8832 16346
rect 1104 16272 8832 16294
rect 2590 16232 2596 16244
rect 2551 16204 2596 16232
rect 2590 16192 2596 16204
rect 2648 16192 2654 16244
rect 3237 16235 3295 16241
rect 3237 16201 3249 16235
rect 3283 16232 3295 16235
rect 3878 16232 3884 16244
rect 3283 16204 3648 16232
rect 3839 16204 3884 16232
rect 3283 16201 3295 16204
rect 3237 16195 3295 16201
rect 2608 16164 2636 16192
rect 3510 16164 3516 16176
rect 2608 16136 3516 16164
rect 3510 16124 3516 16136
rect 3568 16124 3574 16176
rect 3620 16028 3648 16204
rect 3878 16192 3884 16204
rect 3936 16192 3942 16244
rect 3970 16192 3976 16244
rect 4028 16232 4034 16244
rect 4028 16204 6500 16232
rect 4028 16192 4034 16204
rect 4706 16164 4712 16176
rect 3712 16136 4712 16164
rect 3712 16105 3740 16136
rect 4706 16124 4712 16136
rect 4764 16124 4770 16176
rect 5626 16124 5632 16176
rect 5684 16164 5690 16176
rect 6365 16167 6423 16173
rect 6365 16164 6377 16167
rect 5684 16136 6377 16164
rect 5684 16124 5690 16136
rect 6365 16133 6377 16136
rect 6411 16133 6423 16167
rect 6472 16164 6500 16204
rect 7190 16164 7196 16176
rect 6472 16136 7196 16164
rect 6365 16127 6423 16133
rect 7190 16124 7196 16136
rect 7248 16124 7254 16176
rect 7282 16124 7288 16176
rect 7340 16164 7346 16176
rect 7377 16167 7435 16173
rect 7377 16164 7389 16167
rect 7340 16136 7389 16164
rect 7340 16124 7346 16136
rect 7377 16133 7389 16136
rect 7423 16133 7435 16167
rect 7377 16127 7435 16133
rect 3697 16099 3755 16105
rect 3697 16065 3709 16099
rect 3743 16065 3755 16099
rect 4522 16096 4528 16108
rect 4483 16068 4528 16096
rect 3697 16059 3755 16065
rect 4522 16056 4528 16068
rect 4580 16056 4586 16108
rect 4614 16056 4620 16108
rect 4672 16096 4678 16108
rect 5077 16099 5135 16105
rect 5077 16096 5089 16099
rect 4672 16068 5089 16096
rect 4672 16056 4678 16068
rect 5077 16065 5089 16068
rect 5123 16096 5135 16099
rect 6549 16099 6607 16105
rect 6549 16096 6561 16099
rect 5123 16068 6561 16096
rect 5123 16065 5135 16068
rect 5077 16059 5135 16065
rect 6549 16065 6561 16068
rect 6595 16065 6607 16099
rect 6549 16059 6607 16065
rect 7006 16056 7012 16108
rect 7064 16096 7070 16108
rect 8018 16096 8024 16108
rect 7064 16068 8024 16096
rect 7064 16056 7070 16068
rect 8018 16056 8024 16068
rect 8076 16096 8082 16108
rect 8113 16099 8171 16105
rect 8113 16096 8125 16099
rect 8076 16068 8125 16096
rect 8076 16056 8082 16068
rect 8113 16065 8125 16068
rect 8159 16065 8171 16099
rect 8113 16059 8171 16065
rect 4433 16031 4491 16037
rect 2746 16000 4384 16028
rect 2746 15972 2774 16000
rect 2682 15920 2688 15972
rect 2740 15932 2774 15972
rect 4356 15960 4384 16000
rect 4433 15997 4445 16031
rect 4479 16028 4491 16031
rect 4985 16031 5043 16037
rect 4985 16028 4997 16031
rect 4479 16000 4997 16028
rect 4479 15997 4491 16000
rect 4433 15991 4491 15997
rect 4985 15997 4997 16000
rect 5031 15997 5043 16031
rect 5534 16028 5540 16040
rect 5495 16000 5540 16028
rect 4985 15991 5043 15997
rect 5534 15988 5540 16000
rect 5592 15988 5598 16040
rect 5552 15960 5580 15988
rect 4356 15932 5580 15960
rect 2740 15920 2746 15932
rect 1581 15895 1639 15901
rect 1581 15861 1593 15895
rect 1627 15892 1639 15895
rect 1946 15892 1952 15904
rect 1627 15864 1952 15892
rect 1627 15861 1639 15864
rect 1581 15855 1639 15861
rect 1946 15852 1952 15864
rect 2004 15852 2010 15904
rect 2130 15892 2136 15904
rect 2043 15864 2136 15892
rect 2130 15852 2136 15864
rect 2188 15892 2194 15904
rect 3142 15892 3148 15904
rect 2188 15864 3148 15892
rect 2188 15852 2194 15864
rect 3142 15852 3148 15864
rect 3200 15852 3206 15904
rect 3510 15852 3516 15904
rect 3568 15892 3574 15904
rect 5994 15892 6000 15904
rect 3568 15864 6000 15892
rect 3568 15852 3574 15864
rect 5994 15852 6000 15864
rect 6052 15852 6058 15904
rect 1104 15802 8832 15824
rect 1104 15750 2248 15802
rect 2300 15750 2312 15802
rect 2364 15750 2376 15802
rect 2428 15750 2440 15802
rect 2492 15750 2504 15802
rect 2556 15750 4846 15802
rect 4898 15750 4910 15802
rect 4962 15750 4974 15802
rect 5026 15750 5038 15802
rect 5090 15750 5102 15802
rect 5154 15750 7443 15802
rect 7495 15750 7507 15802
rect 7559 15750 7571 15802
rect 7623 15750 7635 15802
rect 7687 15750 7699 15802
rect 7751 15750 8832 15802
rect 1104 15728 8832 15750
rect 2682 15688 2688 15700
rect 2643 15660 2688 15688
rect 2682 15648 2688 15660
rect 2740 15648 2746 15700
rect 3237 15691 3295 15697
rect 3237 15657 3249 15691
rect 3283 15688 3295 15691
rect 5718 15688 5724 15700
rect 3283 15660 5724 15688
rect 3283 15657 3295 15660
rect 3237 15651 3295 15657
rect 5718 15648 5724 15660
rect 5776 15648 5782 15700
rect 5994 15648 6000 15700
rect 6052 15688 6058 15700
rect 6052 15660 7972 15688
rect 6052 15648 6058 15660
rect 3142 15580 3148 15632
rect 3200 15620 3206 15632
rect 7006 15620 7012 15632
rect 3200 15592 7012 15620
rect 3200 15580 3206 15592
rect 7006 15580 7012 15592
rect 7064 15580 7070 15632
rect 7469 15623 7527 15629
rect 7469 15589 7481 15623
rect 7515 15620 7527 15623
rect 7834 15620 7840 15632
rect 7515 15592 7840 15620
rect 7515 15589 7527 15592
rect 7469 15583 7527 15589
rect 7834 15580 7840 15592
rect 7892 15580 7898 15632
rect 4062 15512 4068 15564
rect 4120 15552 4126 15564
rect 7944 15561 7972 15660
rect 7377 15555 7435 15561
rect 7377 15552 7389 15555
rect 4120 15524 7389 15552
rect 4120 15512 4126 15524
rect 7377 15521 7389 15524
rect 7423 15521 7435 15555
rect 7377 15515 7435 15521
rect 7929 15555 7987 15561
rect 7929 15521 7941 15555
rect 7975 15521 7987 15555
rect 7929 15515 7987 15521
rect 4706 15484 4712 15496
rect 4667 15456 4712 15484
rect 4706 15444 4712 15456
rect 4764 15444 4770 15496
rect 5534 15444 5540 15496
rect 5592 15484 5598 15496
rect 5905 15487 5963 15493
rect 5905 15484 5917 15487
rect 5592 15456 5917 15484
rect 5592 15444 5598 15456
rect 5905 15453 5917 15456
rect 5951 15484 5963 15487
rect 6638 15484 6644 15496
rect 5951 15456 6644 15484
rect 5951 15453 5963 15456
rect 5905 15447 5963 15453
rect 6638 15444 6644 15456
rect 6696 15444 6702 15496
rect 6917 15487 6975 15493
rect 6917 15453 6929 15487
rect 6963 15453 6975 15487
rect 6917 15447 6975 15453
rect 4341 15419 4399 15425
rect 4341 15385 4353 15419
rect 4387 15416 4399 15419
rect 4614 15416 4620 15428
rect 4387 15388 4620 15416
rect 4387 15385 4399 15388
rect 4341 15379 4399 15385
rect 4614 15376 4620 15388
rect 4672 15376 4678 15428
rect 5626 15376 5632 15428
rect 5684 15416 5690 15428
rect 6365 15419 6423 15425
rect 6365 15416 6377 15419
rect 5684 15388 6377 15416
rect 5684 15376 5690 15388
rect 6365 15385 6377 15388
rect 6411 15385 6423 15419
rect 6365 15379 6423 15385
rect 6457 15419 6515 15425
rect 6457 15385 6469 15419
rect 6503 15416 6515 15419
rect 6546 15416 6552 15428
rect 6503 15388 6552 15416
rect 6503 15385 6515 15388
rect 6457 15379 6515 15385
rect 6546 15376 6552 15388
rect 6604 15376 6610 15428
rect 6932 15416 6960 15447
rect 8110 15416 8116 15428
rect 6932 15388 8116 15416
rect 1581 15351 1639 15357
rect 1581 15317 1593 15351
rect 1627 15348 1639 15351
rect 1854 15348 1860 15360
rect 1627 15320 1860 15348
rect 1627 15317 1639 15320
rect 1581 15311 1639 15317
rect 1854 15308 1860 15320
rect 1912 15308 1918 15360
rect 1946 15308 1952 15360
rect 2004 15348 2010 15360
rect 2133 15351 2191 15357
rect 2133 15348 2145 15351
rect 2004 15320 2145 15348
rect 2004 15308 2010 15320
rect 2133 15317 2145 15320
rect 2179 15348 2191 15351
rect 2866 15348 2872 15360
rect 2179 15320 2872 15348
rect 2179 15317 2191 15320
rect 2133 15311 2191 15317
rect 2866 15308 2872 15320
rect 2924 15308 2930 15360
rect 3050 15308 3056 15360
rect 3108 15348 3114 15360
rect 3881 15351 3939 15357
rect 3881 15348 3893 15351
rect 3108 15320 3893 15348
rect 3108 15308 3114 15320
rect 3881 15317 3893 15320
rect 3927 15348 3939 15351
rect 6932 15348 6960 15388
rect 8110 15376 8116 15388
rect 8168 15376 8174 15428
rect 3927 15320 6960 15348
rect 3927 15317 3939 15320
rect 3881 15311 3939 15317
rect 1104 15258 8832 15280
rect 1104 15206 3547 15258
rect 3599 15206 3611 15258
rect 3663 15206 3675 15258
rect 3727 15206 3739 15258
rect 3791 15206 3803 15258
rect 3855 15206 6144 15258
rect 6196 15206 6208 15258
rect 6260 15206 6272 15258
rect 6324 15206 6336 15258
rect 6388 15206 6400 15258
rect 6452 15206 8832 15258
rect 1104 15184 8832 15206
rect 3050 15144 3056 15156
rect 3011 15116 3056 15144
rect 3050 15104 3056 15116
rect 3108 15104 3114 15156
rect 6730 15104 6736 15156
rect 6788 15144 6794 15156
rect 6788 15116 6868 15144
rect 6788 15104 6794 15116
rect 4522 15036 4528 15088
rect 4580 15076 4586 15088
rect 4893 15079 4951 15085
rect 4893 15076 4905 15079
rect 4580 15048 4905 15076
rect 4580 15036 4586 15048
rect 4893 15045 4905 15048
rect 4939 15045 4951 15079
rect 4893 15039 4951 15045
rect 4065 15011 4123 15017
rect 4065 14977 4077 15011
rect 4111 15008 4123 15011
rect 4111 14980 4660 15008
rect 4111 14977 4123 14980
rect 4065 14971 4123 14977
rect 4632 14872 4660 14980
rect 4706 14968 4712 15020
rect 4764 15008 4770 15020
rect 5629 15011 5687 15017
rect 4764 14980 4809 15008
rect 4764 14968 4770 14980
rect 5629 14977 5641 15011
rect 5675 15008 5687 15011
rect 5718 15008 5724 15020
rect 5675 14980 5724 15008
rect 5675 14977 5687 14980
rect 5629 14971 5687 14977
rect 5718 14968 5724 14980
rect 5776 14968 5782 15020
rect 6086 14968 6092 15020
rect 6144 15008 6150 15020
rect 6457 15011 6515 15017
rect 6457 15008 6469 15011
rect 6144 14980 6469 15008
rect 6144 14968 6150 14980
rect 6457 14977 6469 14980
rect 6503 14977 6515 15011
rect 6457 14971 6515 14977
rect 6840 14952 6868 15116
rect 7929 15011 7987 15017
rect 7929 14977 7941 15011
rect 7975 15008 7987 15011
rect 8110 15008 8116 15020
rect 7975 14980 8116 15008
rect 7975 14977 7987 14980
rect 7929 14971 7987 14977
rect 8110 14968 8116 14980
rect 8168 14968 8174 15020
rect 5534 14900 5540 14952
rect 5592 14940 5598 14952
rect 6365 14943 6423 14949
rect 6365 14940 6377 14943
rect 5592 14912 6377 14940
rect 5592 14900 5598 14912
rect 6365 14909 6377 14912
rect 6411 14940 6423 14943
rect 6546 14940 6552 14952
rect 6411 14912 6552 14940
rect 6411 14909 6423 14912
rect 6365 14903 6423 14909
rect 6546 14900 6552 14912
rect 6604 14900 6610 14952
rect 6822 14900 6828 14952
rect 6880 14900 6886 14952
rect 6086 14872 6092 14884
rect 4632 14844 6092 14872
rect 6086 14832 6092 14844
rect 6144 14832 6150 14884
rect 1854 14804 1860 14816
rect 1815 14776 1860 14804
rect 1854 14764 1860 14776
rect 1912 14764 1918 14816
rect 2501 14807 2559 14813
rect 2501 14773 2513 14807
rect 2547 14804 2559 14807
rect 2590 14804 2596 14816
rect 2547 14776 2596 14804
rect 2547 14773 2559 14776
rect 2501 14767 2559 14773
rect 2590 14764 2596 14776
rect 2648 14764 2654 14816
rect 3602 14804 3608 14816
rect 3563 14776 3608 14804
rect 3602 14764 3608 14776
rect 3660 14764 3666 14816
rect 4246 14804 4252 14816
rect 4207 14776 4252 14804
rect 4246 14764 4252 14776
rect 4304 14764 4310 14816
rect 4338 14764 4344 14816
rect 4396 14804 4402 14816
rect 8202 14804 8208 14816
rect 4396 14776 8208 14804
rect 4396 14764 4402 14776
rect 8202 14764 8208 14776
rect 8260 14764 8266 14816
rect 1104 14714 8832 14736
rect 1104 14662 2248 14714
rect 2300 14662 2312 14714
rect 2364 14662 2376 14714
rect 2428 14662 2440 14714
rect 2492 14662 2504 14714
rect 2556 14662 4846 14714
rect 4898 14662 4910 14714
rect 4962 14662 4974 14714
rect 5026 14662 5038 14714
rect 5090 14662 5102 14714
rect 5154 14662 7443 14714
rect 7495 14662 7507 14714
rect 7559 14662 7571 14714
rect 7623 14662 7635 14714
rect 7687 14662 7699 14714
rect 7751 14662 8832 14714
rect 1104 14640 8832 14662
rect 3237 14535 3295 14541
rect 3237 14501 3249 14535
rect 3283 14532 3295 14535
rect 3602 14532 3608 14544
rect 3283 14504 3608 14532
rect 3283 14501 3295 14504
rect 3237 14495 3295 14501
rect 3602 14492 3608 14504
rect 3660 14532 3666 14544
rect 5718 14532 5724 14544
rect 3660 14504 5724 14532
rect 3660 14492 3666 14504
rect 5718 14492 5724 14504
rect 5776 14492 5782 14544
rect 4246 14424 4252 14476
rect 4304 14464 4310 14476
rect 5077 14467 5135 14473
rect 5077 14464 5089 14467
rect 4304 14436 5089 14464
rect 4304 14424 4310 14436
rect 5077 14433 5089 14436
rect 5123 14433 5135 14467
rect 5077 14427 5135 14433
rect 5166 14424 5172 14476
rect 5224 14464 5230 14476
rect 5224 14436 6316 14464
rect 5224 14424 5230 14436
rect 3878 14396 3884 14408
rect 3791 14368 3884 14396
rect 3878 14356 3884 14368
rect 3936 14396 3942 14408
rect 4338 14396 4344 14408
rect 3936 14368 4344 14396
rect 3936 14356 3942 14368
rect 4338 14356 4344 14368
rect 4396 14356 4402 14408
rect 4525 14399 4583 14405
rect 4525 14365 4537 14399
rect 4571 14396 4583 14399
rect 5534 14396 5540 14408
rect 4571 14368 5540 14396
rect 4571 14365 4583 14368
rect 4525 14359 4583 14365
rect 5534 14356 5540 14368
rect 5592 14356 5598 14408
rect 5629 14399 5687 14405
rect 5629 14365 5641 14399
rect 5675 14396 5687 14399
rect 5718 14396 5724 14408
rect 5675 14368 5724 14396
rect 5675 14365 5687 14368
rect 5629 14359 5687 14365
rect 5718 14356 5724 14368
rect 5776 14356 5782 14408
rect 6086 14396 6092 14408
rect 6047 14368 6092 14396
rect 6086 14356 6092 14368
rect 6144 14356 6150 14408
rect 6288 14405 6316 14436
rect 6273 14399 6331 14405
rect 6273 14365 6285 14399
rect 6319 14365 6331 14399
rect 6273 14359 6331 14365
rect 6822 14356 6828 14408
rect 6880 14396 6886 14408
rect 7009 14399 7067 14405
rect 7009 14396 7021 14399
rect 6880 14368 7021 14396
rect 6880 14356 6886 14368
rect 7009 14365 7021 14368
rect 7055 14365 7067 14399
rect 7009 14359 7067 14365
rect 8113 14399 8171 14405
rect 8113 14365 8125 14399
rect 8159 14396 8171 14399
rect 8202 14396 8208 14408
rect 8159 14368 8208 14396
rect 8159 14365 8171 14368
rect 8113 14359 8171 14365
rect 8202 14356 8208 14368
rect 8260 14356 8266 14408
rect 2133 14331 2191 14337
rect 2133 14297 2145 14331
rect 2179 14328 2191 14331
rect 2590 14328 2596 14340
rect 2179 14300 2596 14328
rect 2179 14297 2191 14300
rect 2133 14291 2191 14297
rect 2590 14288 2596 14300
rect 2648 14288 2654 14340
rect 4798 14288 4804 14340
rect 4856 14328 4862 14340
rect 6104 14328 6132 14356
rect 4856 14300 6132 14328
rect 4856 14288 4862 14300
rect 6914 14288 6920 14340
rect 6972 14328 6978 14340
rect 7561 14331 7619 14337
rect 7561 14328 7573 14331
rect 6972 14300 7573 14328
rect 6972 14288 6978 14300
rect 7561 14297 7573 14300
rect 7607 14297 7619 14331
rect 7561 14291 7619 14297
rect 7650 14288 7656 14340
rect 7708 14328 7714 14340
rect 7708 14300 7753 14328
rect 7708 14288 7714 14300
rect 1578 14260 1584 14272
rect 1539 14232 1584 14260
rect 1578 14220 1584 14232
rect 1636 14220 1642 14272
rect 2682 14260 2688 14272
rect 2643 14232 2688 14260
rect 2682 14220 2688 14232
rect 2740 14220 2746 14272
rect 4433 14263 4491 14269
rect 4433 14229 4445 14263
rect 4479 14260 4491 14263
rect 5442 14260 5448 14272
rect 4479 14232 5448 14260
rect 4479 14229 4491 14232
rect 4433 14223 4491 14229
rect 5442 14220 5448 14232
rect 5500 14220 5506 14272
rect 5718 14220 5724 14272
rect 5776 14260 5782 14272
rect 6822 14260 6828 14272
rect 5776 14232 6828 14260
rect 5776 14220 5782 14232
rect 6822 14220 6828 14232
rect 6880 14220 6886 14272
rect 1104 14170 8832 14192
rect 1104 14118 3547 14170
rect 3599 14118 3611 14170
rect 3663 14118 3675 14170
rect 3727 14118 3739 14170
rect 3791 14118 3803 14170
rect 3855 14118 6144 14170
rect 6196 14118 6208 14170
rect 6260 14118 6272 14170
rect 6324 14118 6336 14170
rect 6388 14118 6400 14170
rect 6452 14118 8832 14170
rect 1104 14096 8832 14118
rect 3697 14059 3755 14065
rect 3697 14025 3709 14059
rect 3743 14056 3755 14059
rect 3878 14056 3884 14068
rect 3743 14028 3884 14056
rect 3743 14025 3755 14028
rect 3697 14019 3755 14025
rect 3878 14016 3884 14028
rect 3936 14016 3942 14068
rect 4341 14059 4399 14065
rect 4341 14025 4353 14059
rect 4387 14056 4399 14059
rect 5166 14056 5172 14068
rect 4387 14028 5172 14056
rect 4387 14025 4399 14028
rect 4341 14019 4399 14025
rect 5166 14016 5172 14028
rect 5224 14016 5230 14068
rect 4249 13991 4307 13997
rect 4249 13957 4261 13991
rect 4295 13988 4307 13991
rect 5626 13988 5632 14000
rect 4295 13960 5632 13988
rect 4295 13957 4307 13960
rect 4249 13951 4307 13957
rect 5626 13948 5632 13960
rect 5684 13948 5690 14000
rect 5721 13991 5779 13997
rect 5721 13957 5733 13991
rect 5767 13988 5779 13991
rect 6549 13991 6607 13997
rect 6549 13988 6561 13991
rect 5767 13960 6561 13988
rect 5767 13957 5779 13960
rect 5721 13951 5779 13957
rect 6549 13957 6561 13960
rect 6595 13988 6607 13991
rect 7650 13988 7656 14000
rect 6595 13960 7656 13988
rect 6595 13957 6607 13960
rect 6549 13951 6607 13957
rect 7650 13948 7656 13960
rect 7708 13948 7714 14000
rect 1489 13923 1547 13929
rect 1489 13889 1501 13923
rect 1535 13920 1547 13923
rect 1578 13920 1584 13932
rect 1535 13892 1584 13920
rect 1535 13889 1547 13892
rect 1489 13883 1547 13889
rect 1578 13880 1584 13892
rect 1636 13920 1642 13932
rect 1636 13892 2774 13920
rect 1636 13880 1642 13892
rect 2746 13852 2774 13892
rect 2958 13880 2964 13932
rect 3016 13920 3022 13932
rect 3053 13923 3111 13929
rect 3053 13920 3065 13923
rect 3016 13892 3065 13920
rect 3016 13880 3022 13892
rect 3053 13889 3065 13892
rect 3099 13889 3111 13923
rect 4798 13920 4804 13932
rect 4759 13892 4804 13920
rect 3053 13883 3111 13889
rect 4798 13880 4804 13892
rect 4856 13880 4862 13932
rect 4985 13923 5043 13929
rect 4985 13889 4997 13923
rect 5031 13920 5043 13923
rect 5350 13920 5356 13932
rect 5031 13892 5356 13920
rect 5031 13889 5043 13892
rect 4985 13883 5043 13889
rect 5350 13880 5356 13892
rect 5408 13880 5414 13932
rect 7006 13920 7012 13932
rect 6967 13892 7012 13920
rect 7006 13880 7012 13892
rect 7064 13880 7070 13932
rect 8113 13923 8171 13929
rect 8113 13889 8125 13923
rect 8159 13920 8171 13923
rect 8202 13920 8208 13932
rect 8159 13892 8208 13920
rect 8159 13889 8171 13892
rect 8113 13883 8171 13889
rect 8202 13880 8208 13892
rect 8260 13880 8266 13932
rect 5534 13852 5540 13864
rect 2746 13824 4476 13852
rect 5495 13824 5540 13852
rect 1578 13676 1584 13728
rect 1636 13716 1642 13728
rect 1949 13719 2007 13725
rect 1949 13716 1961 13719
rect 1636 13688 1961 13716
rect 1636 13676 1642 13688
rect 1949 13685 1961 13688
rect 1995 13685 2007 13719
rect 1949 13679 2007 13685
rect 2593 13719 2651 13725
rect 2593 13685 2605 13719
rect 2639 13716 2651 13719
rect 2682 13716 2688 13728
rect 2639 13688 2688 13716
rect 2639 13685 2651 13688
rect 2593 13679 2651 13685
rect 2682 13676 2688 13688
rect 2740 13676 2746 13728
rect 4448 13716 4476 13824
rect 5534 13812 5540 13824
rect 5592 13812 5598 13864
rect 4706 13716 4712 13728
rect 4448 13688 4712 13716
rect 4706 13676 4712 13688
rect 4764 13676 4770 13728
rect 1104 13626 8832 13648
rect 1104 13574 2248 13626
rect 2300 13574 2312 13626
rect 2364 13574 2376 13626
rect 2428 13574 2440 13626
rect 2492 13574 2504 13626
rect 2556 13574 4846 13626
rect 4898 13574 4910 13626
rect 4962 13574 4974 13626
rect 5026 13574 5038 13626
rect 5090 13574 5102 13626
rect 5154 13574 7443 13626
rect 7495 13574 7507 13626
rect 7559 13574 7571 13626
rect 7623 13574 7635 13626
rect 7687 13574 7699 13626
rect 7751 13574 8832 13626
rect 1104 13552 8832 13574
rect 1762 13472 1768 13524
rect 1820 13512 1826 13524
rect 2133 13515 2191 13521
rect 2133 13512 2145 13515
rect 1820 13484 2145 13512
rect 1820 13472 1826 13484
rect 2133 13481 2145 13484
rect 2179 13512 2191 13515
rect 5810 13512 5816 13524
rect 2179 13484 5816 13512
rect 2179 13481 2191 13484
rect 2133 13475 2191 13481
rect 5810 13472 5816 13484
rect 5868 13472 5874 13524
rect 6086 13472 6092 13524
rect 6144 13512 6150 13524
rect 8386 13512 8392 13524
rect 6144 13484 8392 13512
rect 6144 13472 6150 13484
rect 8386 13472 8392 13484
rect 8444 13472 8450 13524
rect 3237 13447 3295 13453
rect 3237 13413 3249 13447
rect 3283 13444 3295 13447
rect 5994 13444 6000 13456
rect 3283 13416 6000 13444
rect 3283 13413 3295 13416
rect 3237 13407 3295 13413
rect 5994 13404 6000 13416
rect 6052 13444 6058 13456
rect 6052 13416 8156 13444
rect 6052 13404 6058 13416
rect 7006 13376 7012 13388
rect 3804 13348 7012 13376
rect 3804 13317 3832 13348
rect 7006 13336 7012 13348
rect 7064 13376 7070 13388
rect 7064 13348 7236 13376
rect 7064 13336 7070 13348
rect 3789 13311 3847 13317
rect 3789 13277 3801 13311
rect 3835 13277 3847 13311
rect 3789 13271 3847 13277
rect 4985 13311 5043 13317
rect 4985 13277 4997 13311
rect 5031 13277 5043 13311
rect 5442 13308 5448 13320
rect 5403 13280 5448 13308
rect 4985 13271 5043 13277
rect 2406 13200 2412 13252
rect 2464 13240 2470 13252
rect 4433 13243 4491 13249
rect 4433 13240 4445 13243
rect 2464 13212 4445 13240
rect 2464 13200 2470 13212
rect 4433 13209 4445 13212
rect 4479 13209 4491 13243
rect 4433 13203 4491 13209
rect 4522 13200 4528 13252
rect 4580 13240 4586 13252
rect 5000 13240 5028 13271
rect 5442 13268 5448 13280
rect 5500 13268 5506 13320
rect 5810 13308 5816 13320
rect 5552 13280 5816 13308
rect 5552 13240 5580 13280
rect 5810 13268 5816 13280
rect 5868 13268 5874 13320
rect 6365 13311 6423 13317
rect 6365 13277 6377 13311
rect 6411 13308 6423 13311
rect 7098 13308 7104 13320
rect 6411 13280 7104 13308
rect 6411 13277 6423 13280
rect 6365 13271 6423 13277
rect 7098 13268 7104 13280
rect 7156 13268 7162 13320
rect 7208 13317 7236 13348
rect 8128 13320 8156 13416
rect 7193 13311 7251 13317
rect 7193 13277 7205 13311
rect 7239 13308 7251 13311
rect 7926 13308 7932 13320
rect 7239 13280 7932 13308
rect 7239 13277 7251 13280
rect 7193 13271 7251 13277
rect 7926 13268 7932 13280
rect 7984 13268 7990 13320
rect 8110 13268 8116 13320
rect 8168 13308 8174 13320
rect 8168 13280 8261 13308
rect 8168 13268 8174 13280
rect 4580 13212 4625 13240
rect 5000 13212 5580 13240
rect 5721 13243 5779 13249
rect 4580 13200 4586 13212
rect 5721 13209 5733 13243
rect 5767 13240 5779 13243
rect 7006 13240 7012 13252
rect 5767 13212 7012 13240
rect 5767 13209 5779 13212
rect 5721 13203 5779 13209
rect 7006 13200 7012 13212
rect 7064 13200 7070 13252
rect 7374 13240 7380 13252
rect 7335 13212 7380 13240
rect 7374 13200 7380 13212
rect 7432 13200 7438 13252
rect 1578 13172 1584 13184
rect 1539 13144 1584 13172
rect 1578 13132 1584 13144
rect 1636 13132 1642 13184
rect 2685 13175 2743 13181
rect 2685 13141 2697 13175
rect 2731 13172 2743 13175
rect 3050 13172 3056 13184
rect 2731 13144 3056 13172
rect 2731 13141 2743 13144
rect 2685 13135 2743 13141
rect 3050 13132 3056 13144
rect 3108 13132 3114 13184
rect 3973 13175 4031 13181
rect 3973 13141 3985 13175
rect 4019 13172 4031 13175
rect 7558 13172 7564 13184
rect 4019 13144 7564 13172
rect 4019 13141 4031 13144
rect 3973 13135 4031 13141
rect 7558 13132 7564 13144
rect 7616 13132 7622 13184
rect 1104 13082 8832 13104
rect 1104 13030 3547 13082
rect 3599 13030 3611 13082
rect 3663 13030 3675 13082
rect 3727 13030 3739 13082
rect 3791 13030 3803 13082
rect 3855 13030 6144 13082
rect 6196 13030 6208 13082
rect 6260 13030 6272 13082
rect 6324 13030 6336 13082
rect 6388 13030 6400 13082
rect 6452 13030 8832 13082
rect 1104 13008 8832 13030
rect 1762 12968 1768 12980
rect 1723 12940 1768 12968
rect 1762 12928 1768 12940
rect 1820 12928 1826 12980
rect 2406 12968 2412 12980
rect 2367 12940 2412 12968
rect 2406 12928 2412 12940
rect 2464 12928 2470 12980
rect 2866 12928 2872 12980
rect 2924 12968 2930 12980
rect 5626 12968 5632 12980
rect 2924 12940 5632 12968
rect 2924 12928 2930 12940
rect 5626 12928 5632 12940
rect 5684 12928 5690 12980
rect 5721 12971 5779 12977
rect 5721 12937 5733 12971
rect 5767 12968 5779 12971
rect 6914 12968 6920 12980
rect 5767 12940 6920 12968
rect 5767 12937 5779 12940
rect 5721 12931 5779 12937
rect 6914 12928 6920 12940
rect 6972 12928 6978 12980
rect 3053 12903 3111 12909
rect 3053 12869 3065 12903
rect 3099 12900 3111 12903
rect 4433 12903 4491 12909
rect 4433 12900 4445 12903
rect 3099 12872 4445 12900
rect 3099 12869 3111 12872
rect 3053 12863 3111 12869
rect 4433 12869 4445 12872
rect 4479 12900 4491 12903
rect 4522 12900 4528 12912
rect 4479 12872 4528 12900
rect 4479 12869 4491 12872
rect 4433 12863 4491 12869
rect 4522 12860 4528 12872
rect 4580 12860 4586 12912
rect 5813 12903 5871 12909
rect 5813 12869 5825 12903
rect 5859 12900 5871 12903
rect 7374 12900 7380 12912
rect 5859 12872 7380 12900
rect 5859 12869 5871 12872
rect 5813 12863 5871 12869
rect 7374 12860 7380 12872
rect 7432 12900 7438 12912
rect 7653 12903 7711 12909
rect 7653 12900 7665 12903
rect 7432 12872 7665 12900
rect 7432 12860 7438 12872
rect 7653 12869 7665 12872
rect 7699 12869 7711 12903
rect 7653 12863 7711 12869
rect 2225 12835 2283 12841
rect 2225 12801 2237 12835
rect 2271 12832 2283 12835
rect 3694 12832 3700 12844
rect 2271 12804 3556 12832
rect 3655 12804 3700 12832
rect 2271 12801 2283 12804
rect 2225 12795 2283 12801
rect 3528 12773 3556 12804
rect 3694 12792 3700 12804
rect 3752 12792 3758 12844
rect 4246 12832 4252 12844
rect 4207 12804 4252 12832
rect 4246 12792 4252 12804
rect 4304 12792 4310 12844
rect 5169 12835 5227 12841
rect 5169 12801 5181 12835
rect 5215 12832 5227 12835
rect 7558 12832 7564 12844
rect 5215 12804 5856 12832
rect 7519 12804 7564 12832
rect 5215 12801 5227 12804
rect 5169 12795 5227 12801
rect 3513 12767 3571 12773
rect 3513 12733 3525 12767
rect 3559 12764 3571 12767
rect 4264 12764 4292 12792
rect 5828 12776 5856 12804
rect 7558 12792 7564 12804
rect 7616 12792 7622 12844
rect 8110 12832 8116 12844
rect 8071 12804 8116 12832
rect 8110 12792 8116 12804
rect 8168 12792 8174 12844
rect 3559 12736 4292 12764
rect 3559 12733 3571 12736
rect 3513 12727 3571 12733
rect 5810 12724 5816 12776
rect 5868 12724 5874 12776
rect 6549 12767 6607 12773
rect 6549 12733 6561 12767
rect 6595 12733 6607 12767
rect 6549 12727 6607 12733
rect 2961 12699 3019 12705
rect 2961 12665 2973 12699
rect 3007 12696 3019 12699
rect 4338 12696 4344 12708
rect 3007 12668 4344 12696
rect 3007 12665 3019 12668
rect 2961 12659 3019 12665
rect 4338 12656 4344 12668
rect 4396 12656 4402 12708
rect 4154 12588 4160 12640
rect 4212 12628 4218 12640
rect 6564 12628 6592 12727
rect 7006 12724 7012 12776
rect 7064 12764 7070 12776
rect 7101 12767 7159 12773
rect 7101 12764 7113 12767
rect 7064 12736 7113 12764
rect 7064 12724 7070 12736
rect 7101 12733 7113 12736
rect 7147 12733 7159 12767
rect 7101 12727 7159 12733
rect 6641 12699 6699 12705
rect 6641 12665 6653 12699
rect 6687 12696 6699 12699
rect 7282 12696 7288 12708
rect 6687 12668 7288 12696
rect 6687 12665 6699 12668
rect 6641 12659 6699 12665
rect 7282 12656 7288 12668
rect 7340 12656 7346 12708
rect 4212 12600 6592 12628
rect 4212 12588 4218 12600
rect 1104 12538 8832 12560
rect 1104 12486 2248 12538
rect 2300 12486 2312 12538
rect 2364 12486 2376 12538
rect 2428 12486 2440 12538
rect 2492 12486 2504 12538
rect 2556 12486 4846 12538
rect 4898 12486 4910 12538
rect 4962 12486 4974 12538
rect 5026 12486 5038 12538
rect 5090 12486 5102 12538
rect 5154 12486 7443 12538
rect 7495 12486 7507 12538
rect 7559 12486 7571 12538
rect 7623 12486 7635 12538
rect 7687 12486 7699 12538
rect 7751 12486 8832 12538
rect 1104 12464 8832 12486
rect 3237 12427 3295 12433
rect 3237 12393 3249 12427
rect 3283 12424 3295 12427
rect 4154 12424 4160 12436
rect 3283 12396 4160 12424
rect 3283 12393 3295 12396
rect 3237 12387 3295 12393
rect 4154 12384 4160 12396
rect 4212 12384 4218 12436
rect 5442 12424 5448 12436
rect 4816 12396 5448 12424
rect 3694 12316 3700 12368
rect 3752 12356 3758 12368
rect 4706 12356 4712 12368
rect 3752 12328 4712 12356
rect 3752 12316 3758 12328
rect 4706 12316 4712 12328
rect 4764 12316 4770 12368
rect 4816 12288 4844 12396
rect 5442 12384 5448 12396
rect 5500 12384 5506 12436
rect 5534 12356 5540 12368
rect 2424 12260 4844 12288
rect 5000 12328 5540 12356
rect 2424 12229 2452 12260
rect 2409 12223 2467 12229
rect 2409 12189 2421 12223
rect 2455 12189 2467 12223
rect 2409 12183 2467 12189
rect 3053 12223 3111 12229
rect 3053 12189 3065 12223
rect 3099 12220 3111 12223
rect 5000 12220 5028 12328
rect 5534 12316 5540 12328
rect 5592 12356 5598 12368
rect 5592 12328 6592 12356
rect 5592 12316 5598 12328
rect 5350 12248 5356 12300
rect 5408 12288 5414 12300
rect 6457 12291 6515 12297
rect 6457 12288 6469 12291
rect 5408 12260 6469 12288
rect 5408 12248 5414 12260
rect 6457 12257 6469 12260
rect 6503 12257 6515 12291
rect 6457 12251 6515 12257
rect 6564 12232 6592 12328
rect 3099 12192 5028 12220
rect 5077 12223 5135 12229
rect 3099 12189 3111 12192
rect 3053 12183 3111 12189
rect 5077 12189 5089 12223
rect 5123 12220 5135 12223
rect 5442 12220 5448 12232
rect 5123 12192 5448 12220
rect 5123 12189 5135 12192
rect 5077 12183 5135 12189
rect 5442 12180 5448 12192
rect 5500 12180 5506 12232
rect 5810 12180 5816 12232
rect 5868 12220 5874 12232
rect 5997 12223 6055 12229
rect 5997 12220 6009 12223
rect 5868 12192 6009 12220
rect 5868 12180 5874 12192
rect 5997 12189 6009 12192
rect 6043 12189 6055 12223
rect 6546 12220 6552 12232
rect 6459 12192 6552 12220
rect 5997 12183 6055 12189
rect 5902 12152 5908 12164
rect 2608 12124 5908 12152
rect 1946 12084 1952 12096
rect 1907 12056 1952 12084
rect 1946 12044 1952 12056
rect 2004 12044 2010 12096
rect 2608 12093 2636 12124
rect 5902 12112 5908 12124
rect 5960 12112 5966 12164
rect 6012 12152 6040 12183
rect 6546 12180 6552 12192
rect 6604 12180 6610 12232
rect 6730 12180 6736 12232
rect 6788 12220 6794 12232
rect 8021 12223 8079 12229
rect 8021 12220 8033 12223
rect 6788 12192 8033 12220
rect 6788 12180 6794 12192
rect 8021 12189 8033 12192
rect 8067 12189 8079 12223
rect 8021 12183 8079 12189
rect 6638 12152 6644 12164
rect 6012 12124 6644 12152
rect 6638 12112 6644 12124
rect 6696 12112 6702 12164
rect 2593 12087 2651 12093
rect 2593 12053 2605 12087
rect 2639 12053 2651 12087
rect 3878 12084 3884 12096
rect 3839 12056 3884 12084
rect 2593 12047 2651 12053
rect 3878 12044 3884 12056
rect 3936 12044 3942 12096
rect 3973 12087 4031 12093
rect 3973 12053 3985 12087
rect 4019 12084 4031 12087
rect 7098 12084 7104 12096
rect 4019 12056 7104 12084
rect 4019 12053 4031 12056
rect 3973 12047 4031 12053
rect 7098 12044 7104 12056
rect 7156 12084 7162 12096
rect 7282 12084 7288 12096
rect 7156 12056 7288 12084
rect 7156 12044 7162 12056
rect 7282 12044 7288 12056
rect 7340 12044 7346 12096
rect 1104 11994 8832 12016
rect 1104 11942 3547 11994
rect 3599 11942 3611 11994
rect 3663 11942 3675 11994
rect 3727 11942 3739 11994
rect 3791 11942 3803 11994
rect 3855 11942 6144 11994
rect 6196 11942 6208 11994
rect 6260 11942 6272 11994
rect 6324 11942 6336 11994
rect 6388 11942 6400 11994
rect 6452 11942 8832 11994
rect 1104 11920 8832 11942
rect 3142 11840 3148 11892
rect 3200 11880 3206 11892
rect 3970 11880 3976 11892
rect 3200 11852 3976 11880
rect 3200 11840 3206 11852
rect 3970 11840 3976 11852
rect 4028 11880 4034 11892
rect 4028 11852 5856 11880
rect 4028 11840 4034 11852
rect 3421 11815 3479 11821
rect 3421 11781 3433 11815
rect 3467 11812 3479 11815
rect 5534 11812 5540 11824
rect 3467 11784 5540 11812
rect 3467 11781 3479 11784
rect 3421 11775 3479 11781
rect 5534 11772 5540 11784
rect 5592 11772 5598 11824
rect 4246 11744 4252 11756
rect 4207 11716 4252 11744
rect 4246 11704 4252 11716
rect 4304 11704 4310 11756
rect 5258 11704 5264 11756
rect 5316 11744 5322 11756
rect 5445 11747 5503 11753
rect 5445 11744 5457 11747
rect 5316 11716 5457 11744
rect 5316 11704 5322 11716
rect 5445 11713 5457 11716
rect 5491 11713 5503 11747
rect 5828 11744 5856 11852
rect 5994 11840 6000 11892
rect 6052 11880 6058 11892
rect 6365 11883 6423 11889
rect 6365 11880 6377 11883
rect 6052 11852 6377 11880
rect 6052 11840 6058 11852
rect 6365 11849 6377 11852
rect 6411 11849 6423 11883
rect 6365 11843 6423 11849
rect 6546 11772 6552 11824
rect 6604 11812 6610 11824
rect 6917 11815 6975 11821
rect 6917 11812 6929 11815
rect 6604 11784 6929 11812
rect 6604 11772 6610 11784
rect 6917 11781 6929 11784
rect 6963 11781 6975 11815
rect 7098 11812 7104 11824
rect 7059 11784 7104 11812
rect 6917 11775 6975 11781
rect 7098 11772 7104 11784
rect 7156 11772 7162 11824
rect 7006 11744 7012 11756
rect 5828 11716 7012 11744
rect 5445 11707 5503 11713
rect 7006 11704 7012 11716
rect 7064 11744 7070 11756
rect 7834 11744 7840 11756
rect 7064 11716 7840 11744
rect 7064 11704 7070 11716
rect 7834 11704 7840 11716
rect 7892 11704 7898 11756
rect 2777 11679 2835 11685
rect 2777 11645 2789 11679
rect 2823 11676 2835 11679
rect 3234 11676 3240 11688
rect 2823 11648 3240 11676
rect 2823 11645 2835 11648
rect 2777 11639 2835 11645
rect 3234 11636 3240 11648
rect 3292 11676 3298 11688
rect 6730 11676 6736 11688
rect 3292 11648 6736 11676
rect 3292 11636 3298 11648
rect 6730 11636 6736 11648
rect 6788 11636 6794 11688
rect 4154 11608 4160 11620
rect 4115 11580 4160 11608
rect 4154 11568 4160 11580
rect 4212 11568 4218 11620
rect 1670 11540 1676 11552
rect 1631 11512 1676 11540
rect 1670 11500 1676 11512
rect 1728 11500 1734 11552
rect 1854 11500 1860 11552
rect 1912 11540 1918 11552
rect 2133 11543 2191 11549
rect 2133 11540 2145 11543
rect 1912 11512 2145 11540
rect 1912 11500 1918 11512
rect 2133 11509 2145 11512
rect 2179 11509 2191 11543
rect 2133 11503 2191 11509
rect 3329 11543 3387 11549
rect 3329 11509 3341 11543
rect 3375 11540 3387 11543
rect 5442 11540 5448 11552
rect 3375 11512 5448 11540
rect 3375 11509 3387 11512
rect 3329 11503 3387 11509
rect 5442 11500 5448 11512
rect 5500 11500 5506 11552
rect 1104 11450 8832 11472
rect 1104 11398 2248 11450
rect 2300 11398 2312 11450
rect 2364 11398 2376 11450
rect 2428 11398 2440 11450
rect 2492 11398 2504 11450
rect 2556 11398 4846 11450
rect 4898 11398 4910 11450
rect 4962 11398 4974 11450
rect 5026 11398 5038 11450
rect 5090 11398 5102 11450
rect 5154 11398 7443 11450
rect 7495 11398 7507 11450
rect 7559 11398 7571 11450
rect 7623 11398 7635 11450
rect 7687 11398 7699 11450
rect 7751 11398 8832 11450
rect 1104 11376 8832 11398
rect 3234 11336 3240 11348
rect 3195 11308 3240 11336
rect 3234 11296 3240 11308
rect 3292 11296 3298 11348
rect 3878 11296 3884 11348
rect 3936 11336 3942 11348
rect 7926 11336 7932 11348
rect 3936 11308 7052 11336
rect 7887 11308 7932 11336
rect 3936 11296 3942 11308
rect 4154 11228 4160 11280
rect 4212 11268 4218 11280
rect 4433 11271 4491 11277
rect 4433 11268 4445 11271
rect 4212 11240 4445 11268
rect 4212 11228 4218 11240
rect 4433 11237 4445 11240
rect 4479 11237 4491 11271
rect 4433 11231 4491 11237
rect 5350 11228 5356 11280
rect 5408 11268 5414 11280
rect 6917 11271 6975 11277
rect 6917 11268 6929 11271
rect 5408 11240 6929 11268
rect 5408 11228 5414 11240
rect 6917 11237 6929 11240
rect 6963 11237 6975 11271
rect 6917 11231 6975 11237
rect 3881 11203 3939 11209
rect 3881 11169 3893 11203
rect 3927 11200 3939 11203
rect 3970 11200 3976 11212
rect 3927 11172 3976 11200
rect 3927 11169 3939 11172
rect 3881 11163 3939 11169
rect 3970 11160 3976 11172
rect 4028 11160 4034 11212
rect 4338 11200 4344 11212
rect 4299 11172 4344 11200
rect 4338 11160 4344 11172
rect 4396 11160 4402 11212
rect 5442 11200 5448 11212
rect 5403 11172 5448 11200
rect 5442 11160 5448 11172
rect 5500 11160 5506 11212
rect 6825 11203 6883 11209
rect 6825 11169 6837 11203
rect 6871 11200 6883 11203
rect 7024 11200 7052 11308
rect 7926 11296 7932 11308
rect 7984 11296 7990 11348
rect 6871 11172 7052 11200
rect 6871 11169 6883 11172
rect 6825 11163 6883 11169
rect 1581 11135 1639 11141
rect 1581 11101 1593 11135
rect 1627 11132 1639 11135
rect 1670 11132 1676 11144
rect 1627 11104 1676 11132
rect 1627 11101 1639 11104
rect 1581 11095 1639 11101
rect 1670 11092 1676 11104
rect 1728 11132 1734 11144
rect 4893 11135 4951 11141
rect 4893 11132 4905 11135
rect 1728 11104 4905 11132
rect 1728 11092 1734 11104
rect 4893 11101 4905 11104
rect 4939 11132 4951 11135
rect 5258 11132 5264 11144
rect 4939 11104 5264 11132
rect 4939 11101 4951 11104
rect 4893 11095 4951 11101
rect 5258 11092 5264 11104
rect 5316 11092 5322 11144
rect 5997 11135 6055 11141
rect 5997 11101 6009 11135
rect 6043 11101 6055 11135
rect 5997 11095 6055 11101
rect 1946 11024 1952 11076
rect 2004 11064 2010 11076
rect 2685 11067 2743 11073
rect 2685 11064 2697 11067
rect 2004 11036 2697 11064
rect 2004 11024 2010 11036
rect 2685 11033 2697 11036
rect 2731 11064 2743 11067
rect 2731 11036 4660 11064
rect 2731 11033 2743 11036
rect 2685 11027 2743 11033
rect 2130 10996 2136 11008
rect 2091 10968 2136 10996
rect 2130 10956 2136 10968
rect 2188 10956 2194 11008
rect 4632 10996 4660 11036
rect 4706 11024 4712 11076
rect 4764 11064 4770 11076
rect 5537 11067 5595 11073
rect 5537 11064 5549 11067
rect 4764 11036 5549 11064
rect 4764 11024 4770 11036
rect 5537 11033 5549 11036
rect 5583 11033 5595 11067
rect 5537 11027 5595 11033
rect 5810 11024 5816 11076
rect 5868 11024 5874 11076
rect 5828 10996 5856 11024
rect 6012 10996 6040 11095
rect 6730 11092 6736 11144
rect 6788 11132 6794 11144
rect 7374 11132 7380 11144
rect 6788 11104 7380 11132
rect 6788 11092 6794 11104
rect 7374 11092 7380 11104
rect 7432 11092 7438 11144
rect 7834 11024 7840 11076
rect 7892 11064 7898 11076
rect 8021 11067 8079 11073
rect 8021 11064 8033 11067
rect 7892 11036 8033 11064
rect 7892 11024 7898 11036
rect 8021 11033 8033 11036
rect 8067 11033 8079 11067
rect 8021 11027 8079 11033
rect 4632 10968 6040 10996
rect 8202 10956 8208 11008
rect 8260 10996 8266 11008
rect 8386 10996 8392 11008
rect 8260 10968 8392 10996
rect 8260 10956 8266 10968
rect 8386 10956 8392 10968
rect 8444 10956 8450 11008
rect 1104 10906 8832 10928
rect 1104 10854 3547 10906
rect 3599 10854 3611 10906
rect 3663 10854 3675 10906
rect 3727 10854 3739 10906
rect 3791 10854 3803 10906
rect 3855 10854 6144 10906
rect 6196 10854 6208 10906
rect 6260 10854 6272 10906
rect 6324 10854 6336 10906
rect 6388 10854 6400 10906
rect 6452 10854 8832 10906
rect 1104 10832 8832 10854
rect 2317 10795 2375 10801
rect 2317 10761 2329 10795
rect 2363 10792 2375 10795
rect 3050 10792 3056 10804
rect 2363 10764 3056 10792
rect 2363 10761 2375 10764
rect 2317 10755 2375 10761
rect 3050 10752 3056 10764
rect 3108 10752 3114 10804
rect 4614 10792 4620 10804
rect 4575 10764 4620 10792
rect 4614 10752 4620 10764
rect 4672 10752 4678 10804
rect 5534 10752 5540 10804
rect 5592 10792 5598 10804
rect 6914 10792 6920 10804
rect 5592 10764 6920 10792
rect 5592 10752 5598 10764
rect 4065 10727 4123 10733
rect 4065 10693 4077 10727
rect 4111 10724 4123 10727
rect 6086 10724 6092 10736
rect 4111 10696 6092 10724
rect 4111 10693 4123 10696
rect 4065 10687 4123 10693
rect 6086 10684 6092 10696
rect 6144 10684 6150 10736
rect 6472 10733 6500 10764
rect 6914 10752 6920 10764
rect 6972 10752 6978 10804
rect 6457 10727 6515 10733
rect 6457 10693 6469 10727
rect 6503 10693 6515 10727
rect 6457 10687 6515 10693
rect 4706 10656 4712 10668
rect 4667 10628 4712 10656
rect 4706 10616 4712 10628
rect 4764 10616 4770 10668
rect 5902 10616 5908 10668
rect 5960 10656 5966 10668
rect 6365 10659 6423 10665
rect 6365 10656 6377 10659
rect 5960 10628 6377 10656
rect 5960 10616 5966 10628
rect 6365 10625 6377 10628
rect 6411 10625 6423 10659
rect 6365 10619 6423 10625
rect 6917 10659 6975 10665
rect 6917 10625 6929 10659
rect 6963 10656 6975 10659
rect 7190 10656 7196 10668
rect 6963 10628 7196 10656
rect 6963 10625 6975 10628
rect 6917 10619 6975 10625
rect 7190 10616 7196 10628
rect 7248 10616 7254 10668
rect 4338 10548 4344 10600
rect 4396 10588 4402 10600
rect 5261 10591 5319 10597
rect 5261 10588 5273 10591
rect 4396 10560 5273 10588
rect 4396 10548 4402 10560
rect 5261 10557 5273 10560
rect 5307 10557 5319 10591
rect 5810 10588 5816 10600
rect 5771 10560 5816 10588
rect 5261 10551 5319 10557
rect 5810 10548 5816 10560
rect 5868 10548 5874 10600
rect 6546 10548 6552 10600
rect 6604 10588 6610 10600
rect 7561 10591 7619 10597
rect 7561 10588 7573 10591
rect 6604 10560 7573 10588
rect 6604 10548 6610 10560
rect 7561 10557 7573 10560
rect 7607 10557 7619 10591
rect 7561 10551 7619 10557
rect 8113 10591 8171 10597
rect 8113 10557 8125 10591
rect 8159 10588 8171 10591
rect 8202 10588 8208 10600
rect 8159 10560 8208 10588
rect 8159 10557 8171 10560
rect 8113 10551 8171 10557
rect 8202 10548 8208 10560
rect 8260 10548 8266 10600
rect 2038 10480 2044 10532
rect 2096 10520 2102 10532
rect 3329 10523 3387 10529
rect 3329 10520 3341 10523
rect 2096 10492 3341 10520
rect 2096 10480 2102 10492
rect 3329 10489 3341 10492
rect 3375 10489 3387 10523
rect 4614 10520 4620 10532
rect 3329 10483 3387 10489
rect 3896 10492 4620 10520
rect 1765 10455 1823 10461
rect 1765 10421 1777 10455
rect 1811 10452 1823 10455
rect 1854 10452 1860 10464
rect 1811 10424 1860 10452
rect 1811 10421 1823 10424
rect 1765 10415 1823 10421
rect 1854 10412 1860 10424
rect 1912 10452 1918 10464
rect 2774 10452 2780 10464
rect 1912 10424 2780 10452
rect 1912 10412 1918 10424
rect 2774 10412 2780 10424
rect 2832 10412 2838 10464
rect 2869 10455 2927 10461
rect 2869 10421 2881 10455
rect 2915 10452 2927 10455
rect 3896 10452 3924 10492
rect 4614 10480 4620 10492
rect 4672 10480 4678 10532
rect 5353 10523 5411 10529
rect 5353 10489 5365 10523
rect 5399 10520 5411 10523
rect 5442 10520 5448 10532
rect 5399 10492 5448 10520
rect 5399 10489 5411 10492
rect 5353 10483 5411 10489
rect 5442 10480 5448 10492
rect 5500 10480 5506 10532
rect 7653 10523 7711 10529
rect 7653 10489 7665 10523
rect 7699 10520 7711 10523
rect 7834 10520 7840 10532
rect 7699 10492 7840 10520
rect 7699 10489 7711 10492
rect 7653 10483 7711 10489
rect 7834 10480 7840 10492
rect 7892 10480 7898 10532
rect 2915 10424 3924 10452
rect 3973 10455 4031 10461
rect 2915 10421 2927 10424
rect 2869 10415 2927 10421
rect 3973 10421 3985 10455
rect 4019 10452 4031 10455
rect 7282 10452 7288 10464
rect 4019 10424 7288 10452
rect 4019 10421 4031 10424
rect 3973 10415 4031 10421
rect 7282 10412 7288 10424
rect 7340 10412 7346 10464
rect 1104 10362 8832 10384
rect 1104 10310 2248 10362
rect 2300 10310 2312 10362
rect 2364 10310 2376 10362
rect 2428 10310 2440 10362
rect 2492 10310 2504 10362
rect 2556 10310 4846 10362
rect 4898 10310 4910 10362
rect 4962 10310 4974 10362
rect 5026 10310 5038 10362
rect 5090 10310 5102 10362
rect 5154 10310 7443 10362
rect 7495 10310 7507 10362
rect 7559 10310 7571 10362
rect 7623 10310 7635 10362
rect 7687 10310 7699 10362
rect 7751 10310 8832 10362
rect 1104 10288 8832 10310
rect 2774 10208 2780 10260
rect 2832 10248 2838 10260
rect 4430 10248 4436 10260
rect 2832 10220 4436 10248
rect 2832 10208 2838 10220
rect 4430 10208 4436 10220
rect 4488 10208 4494 10260
rect 4706 10208 4712 10260
rect 4764 10248 4770 10260
rect 5353 10251 5411 10257
rect 5353 10248 5365 10251
rect 4764 10220 5365 10248
rect 4764 10208 4770 10220
rect 5353 10217 5365 10220
rect 5399 10217 5411 10251
rect 5353 10211 5411 10217
rect 3145 10183 3203 10189
rect 3145 10149 3157 10183
rect 3191 10180 3203 10183
rect 6546 10180 6552 10192
rect 3191 10152 6552 10180
rect 3191 10149 3203 10152
rect 3145 10143 3203 10149
rect 6546 10140 6552 10152
rect 6604 10140 6610 10192
rect 7282 10112 7288 10124
rect 4172 10084 5212 10112
rect 7243 10084 7288 10112
rect 4172 10056 4200 10084
rect 2593 10047 2651 10053
rect 2593 10013 2605 10047
rect 2639 10044 2651 10047
rect 2866 10044 2872 10056
rect 2639 10016 2872 10044
rect 2639 10013 2651 10016
rect 2593 10007 2651 10013
rect 2866 10004 2872 10016
rect 2924 10004 2930 10056
rect 4065 10047 4123 10053
rect 4065 10013 4077 10047
rect 4111 10044 4123 10047
rect 4154 10044 4160 10056
rect 4111 10016 4160 10044
rect 4111 10013 4123 10016
rect 4065 10007 4123 10013
rect 4154 10004 4160 10016
rect 4212 10004 4218 10056
rect 5184 10053 5212 10084
rect 7282 10072 7288 10084
rect 7340 10072 7346 10124
rect 4893 10047 4951 10053
rect 4893 10013 4905 10047
rect 4939 10013 4951 10047
rect 4893 10007 4951 10013
rect 5169 10047 5227 10053
rect 5169 10013 5181 10047
rect 5215 10013 5227 10047
rect 6086 10044 6092 10056
rect 6047 10016 6092 10044
rect 5169 10007 5227 10013
rect 2041 9979 2099 9985
rect 2041 9945 2053 9979
rect 2087 9976 2099 9979
rect 3050 9976 3056 9988
rect 2087 9948 3056 9976
rect 2087 9945 2099 9948
rect 2041 9939 2099 9945
rect 3050 9936 3056 9948
rect 3108 9936 3114 9988
rect 4246 9976 4252 9988
rect 4207 9948 4252 9976
rect 4246 9936 4252 9948
rect 4304 9936 4310 9988
rect 4908 9976 4936 10007
rect 6086 10004 6092 10016
rect 6144 10004 6150 10056
rect 6638 10004 6644 10056
rect 6696 10044 6702 10056
rect 6822 10044 6828 10056
rect 6696 10016 6828 10044
rect 6696 10004 6702 10016
rect 6822 10004 6828 10016
rect 6880 10004 6886 10056
rect 7837 10047 7895 10053
rect 7837 10013 7849 10047
rect 7883 10044 7895 10047
rect 7926 10044 7932 10056
rect 7883 10016 7932 10044
rect 7883 10013 7895 10016
rect 7837 10007 7895 10013
rect 7926 10004 7932 10016
rect 7984 10004 7990 10056
rect 5534 9976 5540 9988
rect 4908 9948 5540 9976
rect 5534 9936 5540 9948
rect 5592 9936 5598 9988
rect 5902 9976 5908 9988
rect 5863 9948 5908 9976
rect 5902 9936 5908 9948
rect 5960 9936 5966 9988
rect 7374 9976 7380 9988
rect 7335 9948 7380 9976
rect 7374 9936 7380 9948
rect 7432 9936 7438 9988
rect 1489 9911 1547 9917
rect 1489 9877 1501 9911
rect 1535 9908 1547 9911
rect 2130 9908 2136 9920
rect 1535 9880 2136 9908
rect 1535 9877 1547 9880
rect 1489 9871 1547 9877
rect 2130 9868 2136 9880
rect 2188 9908 2194 9920
rect 2590 9908 2596 9920
rect 2188 9880 2596 9908
rect 2188 9868 2194 9880
rect 2590 9868 2596 9880
rect 2648 9868 2654 9920
rect 3237 9911 3295 9917
rect 3237 9877 3249 9911
rect 3283 9908 3295 9911
rect 5442 9908 5448 9920
rect 3283 9880 5448 9908
rect 3283 9877 3295 9880
rect 3237 9871 3295 9877
rect 5442 9868 5448 9880
rect 5500 9868 5506 9920
rect 1104 9818 8832 9840
rect 1104 9766 3547 9818
rect 3599 9766 3611 9818
rect 3663 9766 3675 9818
rect 3727 9766 3739 9818
rect 3791 9766 3803 9818
rect 3855 9766 6144 9818
rect 6196 9766 6208 9818
rect 6260 9766 6272 9818
rect 6324 9766 6336 9818
rect 6388 9766 6400 9818
rect 6452 9766 8832 9818
rect 1104 9744 8832 9766
rect 4246 9664 4252 9716
rect 4304 9704 4310 9716
rect 4341 9707 4399 9713
rect 4341 9704 4353 9707
rect 4304 9676 4353 9704
rect 4304 9664 4310 9676
rect 4341 9673 4353 9676
rect 4387 9673 4399 9707
rect 4341 9667 4399 9673
rect 4430 9664 4436 9716
rect 4488 9704 4494 9716
rect 6546 9704 6552 9716
rect 4488 9676 6552 9704
rect 4488 9664 4494 9676
rect 6546 9664 6552 9676
rect 6604 9664 6610 9716
rect 3237 9639 3295 9645
rect 3237 9605 3249 9639
rect 3283 9636 3295 9639
rect 6365 9639 6423 9645
rect 6365 9636 6377 9639
rect 3283 9608 6377 9636
rect 3283 9605 3295 9608
rect 3237 9599 3295 9605
rect 6365 9605 6377 9608
rect 6411 9636 6423 9639
rect 7374 9636 7380 9648
rect 6411 9608 7380 9636
rect 6411 9605 6423 9608
rect 6365 9599 6423 9605
rect 7374 9596 7380 9608
rect 7432 9596 7438 9648
rect 2409 9571 2467 9577
rect 2409 9537 2421 9571
rect 2455 9537 2467 9571
rect 4338 9568 4344 9580
rect 2409 9531 2467 9537
rect 2746 9540 4344 9568
rect 1946 9364 1952 9376
rect 1907 9336 1952 9364
rect 1946 9324 1952 9336
rect 2004 9324 2010 9376
rect 2424 9364 2452 9531
rect 2593 9435 2651 9441
rect 2593 9401 2605 9435
rect 2639 9432 2651 9435
rect 2746 9432 2774 9540
rect 4338 9528 4344 9540
rect 4396 9528 4402 9580
rect 4522 9528 4528 9580
rect 4580 9568 4586 9580
rect 4985 9571 5043 9577
rect 4985 9568 4997 9571
rect 4580 9540 4997 9568
rect 4580 9528 4586 9540
rect 4985 9537 4997 9540
rect 5031 9537 5043 9571
rect 5534 9568 5540 9580
rect 5495 9540 5540 9568
rect 4985 9531 5043 9537
rect 5534 9528 5540 9540
rect 5592 9528 5598 9580
rect 5902 9528 5908 9580
rect 5960 9568 5966 9580
rect 6457 9571 6515 9577
rect 6457 9568 6469 9571
rect 5960 9540 6469 9568
rect 5960 9528 5966 9540
rect 6457 9537 6469 9540
rect 6503 9537 6515 9571
rect 7926 9568 7932 9580
rect 7887 9540 7932 9568
rect 6457 9531 6515 9537
rect 7926 9528 7932 9540
rect 7984 9528 7990 9580
rect 4154 9460 4160 9512
rect 4212 9500 4218 9512
rect 4249 9503 4307 9509
rect 4249 9500 4261 9503
rect 4212 9472 4261 9500
rect 4212 9460 4218 9472
rect 4249 9469 4261 9472
rect 4295 9469 4307 9503
rect 4249 9463 4307 9469
rect 4433 9503 4491 9509
rect 4433 9469 4445 9503
rect 4479 9500 4491 9503
rect 4614 9500 4620 9512
rect 4479 9472 4620 9500
rect 4479 9469 4491 9472
rect 4433 9463 4491 9469
rect 4614 9460 4620 9472
rect 4672 9460 4678 9512
rect 5350 9500 5356 9512
rect 5311 9472 5356 9500
rect 5350 9460 5356 9472
rect 5408 9460 5414 9512
rect 2639 9404 2774 9432
rect 3053 9435 3111 9441
rect 2639 9401 2651 9404
rect 2593 9395 2651 9401
rect 3053 9401 3065 9435
rect 3099 9432 3111 9435
rect 7190 9432 7196 9444
rect 3099 9404 7196 9432
rect 3099 9401 3111 9404
rect 3053 9395 3111 9401
rect 3068 9364 3096 9395
rect 7190 9392 7196 9404
rect 7248 9392 7254 9444
rect 3878 9364 3884 9376
rect 2424 9336 3096 9364
rect 3839 9336 3884 9364
rect 3878 9324 3884 9336
rect 3936 9324 3942 9376
rect 5810 9324 5816 9376
rect 5868 9364 5874 9376
rect 8110 9364 8116 9376
rect 5868 9336 8116 9364
rect 5868 9324 5874 9336
rect 8110 9324 8116 9336
rect 8168 9324 8174 9376
rect 1104 9274 8832 9296
rect 1104 9222 2248 9274
rect 2300 9222 2312 9274
rect 2364 9222 2376 9274
rect 2428 9222 2440 9274
rect 2492 9222 2504 9274
rect 2556 9222 4846 9274
rect 4898 9222 4910 9274
rect 4962 9222 4974 9274
rect 5026 9222 5038 9274
rect 5090 9222 5102 9274
rect 5154 9222 7443 9274
rect 7495 9222 7507 9274
rect 7559 9222 7571 9274
rect 7623 9222 7635 9274
rect 7687 9222 7699 9274
rect 7751 9222 8832 9274
rect 1104 9200 8832 9222
rect 2038 9160 2044 9172
rect 1999 9132 2044 9160
rect 2038 9120 2044 9132
rect 2096 9120 2102 9172
rect 4154 9160 4160 9172
rect 4115 9132 4160 9160
rect 4154 9120 4160 9132
rect 4212 9120 4218 9172
rect 3237 9095 3295 9101
rect 3237 9061 3249 9095
rect 3283 9092 3295 9095
rect 5629 9095 5687 9101
rect 3283 9064 5580 9092
rect 3283 9061 3295 9064
rect 3237 9055 3295 9061
rect 5552 9033 5580 9064
rect 5629 9061 5641 9095
rect 5675 9092 5687 9095
rect 5994 9092 6000 9104
rect 5675 9064 6000 9092
rect 5675 9061 5687 9064
rect 5629 9055 5687 9061
rect 5994 9052 6000 9064
rect 6052 9052 6058 9104
rect 7834 9092 7840 9104
rect 7795 9064 7840 9092
rect 7834 9052 7840 9064
rect 7892 9052 7898 9104
rect 5537 9027 5595 9033
rect 5537 8993 5549 9027
rect 5583 8993 5595 9027
rect 5537 8987 5595 8993
rect 6089 9027 6147 9033
rect 6089 8993 6101 9027
rect 6135 9024 6147 9027
rect 6638 9024 6644 9036
rect 6135 8996 6644 9024
rect 6135 8993 6147 8996
rect 6089 8987 6147 8993
rect 6638 8984 6644 8996
rect 6696 8984 6702 9036
rect 3053 8959 3111 8965
rect 3053 8925 3065 8959
rect 3099 8925 3111 8959
rect 3053 8919 3111 8925
rect 4249 8959 4307 8965
rect 4249 8925 4261 8959
rect 4295 8956 4307 8959
rect 4522 8956 4528 8968
rect 4295 8928 4528 8956
rect 4295 8925 4307 8928
rect 4249 8919 4307 8925
rect 3068 8888 3096 8919
rect 4522 8916 4528 8928
rect 4580 8916 4586 8968
rect 4985 8959 5043 8965
rect 4985 8925 4997 8959
rect 5031 8956 5043 8959
rect 5350 8956 5356 8968
rect 5031 8928 5356 8956
rect 5031 8925 5043 8928
rect 4985 8919 5043 8925
rect 5350 8916 5356 8928
rect 5408 8916 5414 8968
rect 6549 8959 6607 8965
rect 6549 8925 6561 8959
rect 6595 8956 6607 8959
rect 6822 8956 6828 8968
rect 6595 8928 6828 8956
rect 6595 8925 6607 8928
rect 6549 8919 6607 8925
rect 6822 8916 6828 8928
rect 6880 8916 6886 8968
rect 7190 8916 7196 8968
rect 7248 8956 7254 8968
rect 7469 8959 7527 8965
rect 7469 8956 7481 8959
rect 7248 8928 7481 8956
rect 7248 8916 7254 8928
rect 7469 8925 7481 8928
rect 7515 8925 7527 8959
rect 7469 8919 7527 8925
rect 3142 8888 3148 8900
rect 3055 8860 3148 8888
rect 3142 8848 3148 8860
rect 3200 8888 3206 8900
rect 5902 8888 5908 8900
rect 3200 8860 5908 8888
rect 3200 8848 3206 8860
rect 5902 8848 5908 8860
rect 5960 8848 5966 8900
rect 6178 8848 6184 8900
rect 6236 8888 6242 8900
rect 8294 8888 8300 8900
rect 6236 8860 8300 8888
rect 6236 8848 6242 8860
rect 8294 8848 8300 8860
rect 8352 8848 8358 8900
rect 1486 8820 1492 8832
rect 1447 8792 1492 8820
rect 1486 8780 1492 8792
rect 1544 8780 1550 8832
rect 2038 8780 2044 8832
rect 2096 8820 2102 8832
rect 2501 8823 2559 8829
rect 2501 8820 2513 8823
rect 2096 8792 2513 8820
rect 2096 8780 2102 8792
rect 2501 8789 2513 8792
rect 2547 8789 2559 8823
rect 2501 8783 2559 8789
rect 4246 8780 4252 8832
rect 4304 8820 4310 8832
rect 4893 8823 4951 8829
rect 4893 8820 4905 8823
rect 4304 8792 4905 8820
rect 4304 8780 4310 8792
rect 4893 8789 4905 8792
rect 4939 8789 4951 8823
rect 4893 8783 4951 8789
rect 1104 8730 8832 8752
rect 1104 8678 3547 8730
rect 3599 8678 3611 8730
rect 3663 8678 3675 8730
rect 3727 8678 3739 8730
rect 3791 8678 3803 8730
rect 3855 8678 6144 8730
rect 6196 8678 6208 8730
rect 6260 8678 6272 8730
rect 6324 8678 6336 8730
rect 6388 8678 6400 8730
rect 6452 8678 8832 8730
rect 1104 8656 8832 8678
rect 1486 8616 1492 8628
rect 1447 8588 1492 8616
rect 1486 8576 1492 8588
rect 1544 8616 1550 8628
rect 3142 8616 3148 8628
rect 1544 8588 2774 8616
rect 3103 8588 3148 8616
rect 1544 8576 1550 8588
rect 2746 8548 2774 8588
rect 3142 8576 3148 8588
rect 3200 8576 3206 8628
rect 5169 8619 5227 8625
rect 5169 8616 5181 8619
rect 3252 8588 5181 8616
rect 3252 8548 3280 8588
rect 5169 8585 5181 8588
rect 5215 8585 5227 8619
rect 5169 8579 5227 8585
rect 5442 8576 5448 8628
rect 5500 8616 5506 8628
rect 5500 8588 7420 8616
rect 5500 8576 5506 8588
rect 2746 8520 3280 8548
rect 3789 8551 3847 8557
rect 3789 8517 3801 8551
rect 3835 8548 3847 8551
rect 3878 8548 3884 8560
rect 3835 8520 3884 8548
rect 3835 8517 3847 8520
rect 3789 8511 3847 8517
rect 3878 8508 3884 8520
rect 3936 8508 3942 8560
rect 4706 8508 4712 8560
rect 4764 8548 4770 8560
rect 6365 8551 6423 8557
rect 6365 8548 6377 8551
rect 4764 8520 6377 8548
rect 4764 8508 4770 8520
rect 6365 8517 6377 8520
rect 6411 8517 6423 8551
rect 7190 8548 7196 8560
rect 7151 8520 7196 8548
rect 6365 8511 6423 8517
rect 7190 8508 7196 8520
rect 7248 8508 7254 8560
rect 7392 8557 7420 8588
rect 7377 8551 7435 8557
rect 7377 8517 7389 8551
rect 7423 8517 7435 8551
rect 7377 8511 7435 8517
rect 3237 8483 3295 8489
rect 3237 8449 3249 8483
rect 3283 8480 3295 8483
rect 3283 8452 4108 8480
rect 3283 8449 3295 8452
rect 3237 8443 3295 8449
rect 2041 8415 2099 8421
rect 2041 8381 2053 8415
rect 2087 8412 2099 8415
rect 3878 8412 3884 8424
rect 2087 8384 3884 8412
rect 2087 8381 2099 8384
rect 2041 8375 2099 8381
rect 3878 8372 3884 8384
rect 3936 8372 3942 8424
rect 2593 8347 2651 8353
rect 2593 8313 2605 8347
rect 2639 8344 2651 8347
rect 4080 8344 4108 8452
rect 4154 8440 4160 8492
rect 4212 8480 4218 8492
rect 5261 8483 5319 8489
rect 5261 8480 5273 8483
rect 4212 8452 5273 8480
rect 4212 8440 4218 8452
rect 5261 8449 5273 8452
rect 5307 8449 5319 8483
rect 5261 8443 5319 8449
rect 5442 8440 5448 8492
rect 5500 8480 5506 8492
rect 6549 8483 6607 8489
rect 6549 8480 6561 8483
rect 5500 8452 6561 8480
rect 5500 8440 5506 8452
rect 6549 8449 6561 8452
rect 6595 8449 6607 8483
rect 8110 8480 8116 8492
rect 8071 8452 8116 8480
rect 6549 8443 6607 8449
rect 8110 8440 8116 8452
rect 8168 8440 8174 8492
rect 4522 8412 4528 8424
rect 4483 8384 4528 8412
rect 4522 8372 4528 8384
rect 4580 8372 4586 8424
rect 5718 8372 5724 8424
rect 5776 8412 5782 8424
rect 5813 8415 5871 8421
rect 5813 8412 5825 8415
rect 5776 8384 5825 8412
rect 5776 8372 5782 8384
rect 5813 8381 5825 8384
rect 5859 8381 5871 8415
rect 5813 8375 5871 8381
rect 5350 8344 5356 8356
rect 2639 8316 2774 8344
rect 4080 8316 5356 8344
rect 2639 8313 2651 8316
rect 2593 8307 2651 8313
rect 2746 8276 2774 8316
rect 5350 8304 5356 8316
rect 5408 8304 5414 8356
rect 5828 8344 5856 8375
rect 5828 8316 6960 8344
rect 3970 8276 3976 8288
rect 2746 8248 3976 8276
rect 3970 8236 3976 8248
rect 4028 8236 4034 8288
rect 5169 8279 5227 8285
rect 5169 8245 5181 8279
rect 5215 8276 5227 8279
rect 6178 8276 6184 8288
rect 5215 8248 6184 8276
rect 5215 8245 5227 8248
rect 5169 8239 5227 8245
rect 6178 8236 6184 8248
rect 6236 8236 6242 8288
rect 6932 8276 6960 8316
rect 7282 8276 7288 8288
rect 6932 8248 7288 8276
rect 7282 8236 7288 8248
rect 7340 8236 7346 8288
rect 1104 8186 8832 8208
rect 1104 8134 2248 8186
rect 2300 8134 2312 8186
rect 2364 8134 2376 8186
rect 2428 8134 2440 8186
rect 2492 8134 2504 8186
rect 2556 8134 4846 8186
rect 4898 8134 4910 8186
rect 4962 8134 4974 8186
rect 5026 8134 5038 8186
rect 5090 8134 5102 8186
rect 5154 8134 7443 8186
rect 7495 8134 7507 8186
rect 7559 8134 7571 8186
rect 7623 8134 7635 8186
rect 7687 8134 7699 8186
rect 7751 8134 8832 8186
rect 1104 8112 8832 8134
rect 1854 8032 1860 8084
rect 1912 8072 1918 8084
rect 1949 8075 2007 8081
rect 1949 8072 1961 8075
rect 1912 8044 1961 8072
rect 1912 8032 1918 8044
rect 1949 8041 1961 8044
rect 1995 8072 2007 8075
rect 2038 8072 2044 8084
rect 1995 8044 2044 8072
rect 1995 8041 2007 8044
rect 1949 8035 2007 8041
rect 2038 8032 2044 8044
rect 2096 8032 2102 8084
rect 3418 7964 3424 8016
rect 3476 8004 3482 8016
rect 4522 8004 4528 8016
rect 3476 7976 4528 8004
rect 3476 7964 3482 7976
rect 4522 7964 4528 7976
rect 4580 7964 4586 8016
rect 5166 7964 5172 8016
rect 5224 8004 5230 8016
rect 5902 8004 5908 8016
rect 5224 7976 5908 8004
rect 5224 7964 5230 7976
rect 5902 7964 5908 7976
rect 5960 7964 5966 8016
rect 1486 7896 1492 7948
rect 1544 7936 1550 7948
rect 5629 7939 5687 7945
rect 5629 7936 5641 7939
rect 1544 7908 5641 7936
rect 1544 7896 1550 7908
rect 5629 7905 5641 7908
rect 5675 7905 5687 7939
rect 5629 7899 5687 7905
rect 2406 7868 2412 7880
rect 2367 7840 2412 7868
rect 2406 7828 2412 7840
rect 2464 7828 2470 7880
rect 3053 7871 3111 7877
rect 3053 7837 3065 7871
rect 3099 7868 3111 7871
rect 4522 7868 4528 7880
rect 3099 7840 4528 7868
rect 3099 7837 3111 7840
rect 3053 7831 3111 7837
rect 4522 7828 4528 7840
rect 4580 7828 4586 7880
rect 4893 7871 4951 7877
rect 4893 7837 4905 7871
rect 4939 7837 4951 7871
rect 4893 7831 4951 7837
rect 4338 7800 4344 7812
rect 4299 7772 4344 7800
rect 4338 7760 4344 7772
rect 4396 7760 4402 7812
rect 4430 7760 4436 7812
rect 4488 7800 4494 7812
rect 4488 7772 4533 7800
rect 4488 7760 4494 7772
rect 2590 7732 2596 7744
rect 2551 7704 2596 7732
rect 2590 7692 2596 7704
rect 2648 7692 2654 7744
rect 3234 7732 3240 7744
rect 3195 7704 3240 7732
rect 3234 7692 3240 7704
rect 3292 7692 3298 7744
rect 3881 7735 3939 7741
rect 3881 7701 3893 7735
rect 3927 7732 3939 7735
rect 3970 7732 3976 7744
rect 3927 7704 3976 7732
rect 3927 7701 3939 7704
rect 3881 7695 3939 7701
rect 3970 7692 3976 7704
rect 4028 7732 4034 7744
rect 4908 7732 4936 7831
rect 5258 7828 5264 7880
rect 5316 7868 5322 7880
rect 5721 7871 5779 7877
rect 5721 7868 5733 7871
rect 5316 7840 5733 7868
rect 5316 7828 5322 7840
rect 5721 7837 5733 7840
rect 5767 7837 5779 7871
rect 6178 7868 6184 7880
rect 6091 7840 6184 7868
rect 5721 7831 5779 7837
rect 6178 7828 6184 7840
rect 6236 7868 6242 7880
rect 7006 7868 7012 7880
rect 6236 7840 7012 7868
rect 6236 7828 6242 7840
rect 7006 7828 7012 7840
rect 7064 7828 7070 7880
rect 7653 7871 7711 7877
rect 7653 7837 7665 7871
rect 7699 7868 7711 7871
rect 7834 7868 7840 7880
rect 7699 7840 7840 7868
rect 7699 7837 7711 7840
rect 7653 7831 7711 7837
rect 7834 7828 7840 7840
rect 7892 7828 7898 7880
rect 6730 7800 6736 7812
rect 6691 7772 6736 7800
rect 6730 7760 6736 7772
rect 6788 7760 6794 7812
rect 6914 7800 6920 7812
rect 6875 7772 6920 7800
rect 6914 7760 6920 7772
rect 6972 7760 6978 7812
rect 4028 7704 4936 7732
rect 4028 7692 4034 7704
rect 1104 7642 8832 7664
rect 1104 7590 3547 7642
rect 3599 7590 3611 7642
rect 3663 7590 3675 7642
rect 3727 7590 3739 7642
rect 3791 7590 3803 7642
rect 3855 7590 6144 7642
rect 6196 7590 6208 7642
rect 6260 7590 6272 7642
rect 6324 7590 6336 7642
rect 6388 7590 6400 7642
rect 6452 7590 8832 7642
rect 1104 7568 8832 7590
rect 2041 7531 2099 7537
rect 2041 7497 2053 7531
rect 2087 7528 2099 7531
rect 6914 7528 6920 7540
rect 2087 7500 6920 7528
rect 2087 7497 2099 7500
rect 2041 7491 2099 7497
rect 2590 7420 2596 7472
rect 2648 7460 2654 7472
rect 3344 7469 3372 7500
rect 6914 7488 6920 7500
rect 6972 7488 6978 7540
rect 3237 7463 3295 7469
rect 3237 7460 3249 7463
rect 2648 7432 3249 7460
rect 2648 7420 2654 7432
rect 3237 7429 3249 7432
rect 3283 7429 3295 7463
rect 3237 7423 3295 7429
rect 3329 7463 3387 7469
rect 3329 7429 3341 7463
rect 3375 7429 3387 7463
rect 4062 7460 4068 7472
rect 3329 7423 3387 7429
rect 3620 7432 4068 7460
rect 2685 7395 2743 7401
rect 2685 7361 2697 7395
rect 2731 7392 2743 7395
rect 3620 7392 3648 7432
rect 4062 7420 4068 7432
rect 4120 7420 4126 7472
rect 4246 7460 4252 7472
rect 4207 7432 4252 7460
rect 4246 7420 4252 7432
rect 4304 7420 4310 7472
rect 4430 7460 4436 7472
rect 4391 7432 4436 7460
rect 4430 7420 4436 7432
rect 4488 7460 4494 7472
rect 5629 7463 5687 7469
rect 5629 7460 5641 7463
rect 4488 7432 5641 7460
rect 4488 7420 4494 7432
rect 5629 7429 5641 7432
rect 5675 7429 5687 7463
rect 5629 7423 5687 7429
rect 6365 7463 6423 7469
rect 6365 7429 6377 7463
rect 6411 7429 6423 7463
rect 6365 7423 6423 7429
rect 4154 7392 4160 7404
rect 2731 7364 3648 7392
rect 3712 7364 4160 7392
rect 2731 7361 2743 7364
rect 2685 7355 2743 7361
rect 1949 7327 2007 7333
rect 1949 7293 1961 7327
rect 1995 7324 2007 7327
rect 3712 7324 3740 7364
rect 4154 7352 4160 7364
rect 4212 7352 4218 7404
rect 5169 7395 5227 7401
rect 5169 7392 5181 7395
rect 4264 7364 5181 7392
rect 1995 7296 3740 7324
rect 1995 7293 2007 7296
rect 1949 7287 2007 7293
rect 3786 7284 3792 7336
rect 3844 7324 3850 7336
rect 3844 7296 3889 7324
rect 3844 7284 3850 7296
rect 3970 7284 3976 7336
rect 4028 7324 4034 7336
rect 4264 7324 4292 7364
rect 5169 7361 5181 7364
rect 5215 7361 5227 7395
rect 5169 7355 5227 7361
rect 5350 7352 5356 7404
rect 5408 7392 5414 7404
rect 6380 7392 6408 7423
rect 6730 7392 6736 7404
rect 5408 7364 6408 7392
rect 6691 7364 6736 7392
rect 5408 7352 5414 7364
rect 6730 7352 6736 7364
rect 6788 7352 6794 7404
rect 7282 7352 7288 7404
rect 7340 7392 7346 7404
rect 7926 7392 7932 7404
rect 7340 7364 7932 7392
rect 7340 7352 7346 7364
rect 7926 7352 7932 7364
rect 7984 7352 7990 7404
rect 6748 7324 6776 7352
rect 4028 7296 4292 7324
rect 4540 7296 6776 7324
rect 4028 7284 4034 7296
rect 2406 7216 2412 7268
rect 2464 7256 2470 7268
rect 2501 7259 2559 7265
rect 2501 7256 2513 7259
rect 2464 7228 2513 7256
rect 2464 7216 2470 7228
rect 2501 7225 2513 7228
rect 2547 7256 2559 7259
rect 4540 7256 4568 7296
rect 2547 7228 4568 7256
rect 2547 7225 2559 7228
rect 2501 7219 2559 7225
rect 2038 7148 2044 7200
rect 2096 7188 2102 7200
rect 4246 7188 4252 7200
rect 2096 7160 4252 7188
rect 2096 7148 2102 7160
rect 4246 7148 4252 7160
rect 4304 7148 4310 7200
rect 5166 7148 5172 7200
rect 5224 7188 5230 7200
rect 5721 7191 5779 7197
rect 5721 7188 5733 7191
rect 5224 7160 5733 7188
rect 5224 7148 5230 7160
rect 5721 7157 5733 7160
rect 5767 7157 5779 7191
rect 5721 7151 5779 7157
rect 1104 7098 8832 7120
rect 1104 7046 2248 7098
rect 2300 7046 2312 7098
rect 2364 7046 2376 7098
rect 2428 7046 2440 7098
rect 2492 7046 2504 7098
rect 2556 7046 4846 7098
rect 4898 7046 4910 7098
rect 4962 7046 4974 7098
rect 5026 7046 5038 7098
rect 5090 7046 5102 7098
rect 5154 7046 7443 7098
rect 7495 7046 7507 7098
rect 7559 7046 7571 7098
rect 7623 7046 7635 7098
rect 7687 7046 7699 7098
rect 7751 7046 8832 7098
rect 1104 7024 8832 7046
rect 1486 6984 1492 6996
rect 1447 6956 1492 6984
rect 1486 6944 1492 6956
rect 1544 6944 1550 6996
rect 3789 6987 3847 6993
rect 3789 6984 3801 6987
rect 3160 6956 3801 6984
rect 3160 6925 3188 6956
rect 3789 6953 3801 6956
rect 3835 6953 3847 6987
rect 3789 6947 3847 6953
rect 4430 6944 4436 6996
rect 4488 6984 4494 6996
rect 4706 6984 4712 6996
rect 4488 6956 4712 6984
rect 4488 6944 4494 6956
rect 4706 6944 4712 6956
rect 4764 6944 4770 6996
rect 3145 6919 3203 6925
rect 3145 6916 3157 6919
rect 1596 6888 3157 6916
rect 1596 6789 1624 6888
rect 3145 6885 3157 6888
rect 3191 6885 3203 6919
rect 3145 6879 3203 6885
rect 4249 6919 4307 6925
rect 4249 6885 4261 6919
rect 4295 6916 4307 6919
rect 5442 6916 5448 6928
rect 4295 6888 5448 6916
rect 4295 6885 4307 6888
rect 4249 6879 4307 6885
rect 5442 6876 5448 6888
rect 5500 6876 5506 6928
rect 6089 6919 6147 6925
rect 6089 6916 6101 6919
rect 5552 6888 6101 6916
rect 3234 6848 3240 6860
rect 3195 6820 3240 6848
rect 3234 6808 3240 6820
rect 3292 6808 3298 6860
rect 3326 6808 3332 6860
rect 3384 6848 3390 6860
rect 3384 6820 4660 6848
rect 3384 6808 3390 6820
rect 1581 6783 1639 6789
rect 1581 6749 1593 6783
rect 1627 6749 1639 6783
rect 2038 6780 2044 6792
rect 1999 6752 2044 6780
rect 1581 6743 1639 6749
rect 2038 6740 2044 6752
rect 2096 6740 2102 6792
rect 2590 6740 2596 6792
rect 2648 6780 2654 6792
rect 2685 6783 2743 6789
rect 2685 6780 2697 6783
rect 2648 6752 2697 6780
rect 2648 6740 2654 6752
rect 2685 6749 2697 6752
rect 2731 6749 2743 6783
rect 4246 6780 4252 6792
rect 4207 6752 4252 6780
rect 2685 6743 2743 6749
rect 4246 6740 4252 6752
rect 4304 6740 4310 6792
rect 4632 6780 4660 6820
rect 4706 6808 4712 6860
rect 4764 6848 4770 6860
rect 5258 6848 5264 6860
rect 4764 6820 5264 6848
rect 4764 6808 4770 6820
rect 5258 6808 5264 6820
rect 5316 6848 5322 6860
rect 5552 6848 5580 6888
rect 6089 6885 6101 6888
rect 6135 6885 6147 6919
rect 6089 6879 6147 6885
rect 7098 6848 7104 6860
rect 5316 6820 5580 6848
rect 6104 6820 7104 6848
rect 5316 6808 5322 6820
rect 5537 6783 5595 6789
rect 4632 6752 5488 6780
rect 3789 6715 3847 6721
rect 3789 6681 3801 6715
rect 3835 6712 3847 6715
rect 5350 6712 5356 6724
rect 3835 6684 5356 6712
rect 3835 6681 3847 6684
rect 3789 6675 3847 6681
rect 5350 6672 5356 6684
rect 5408 6672 5414 6724
rect 5460 6712 5488 6752
rect 5537 6749 5549 6783
rect 5583 6780 5595 6783
rect 5718 6780 5724 6792
rect 5583 6752 5724 6780
rect 5583 6749 5595 6752
rect 5537 6743 5595 6749
rect 5718 6740 5724 6752
rect 5776 6740 5782 6792
rect 6104 6712 6132 6820
rect 7098 6808 7104 6820
rect 7156 6808 7162 6860
rect 6181 6783 6239 6789
rect 6181 6749 6193 6783
rect 6227 6749 6239 6783
rect 6181 6743 6239 6749
rect 5460 6684 6132 6712
rect 2225 6647 2283 6653
rect 2225 6613 2237 6647
rect 2271 6644 2283 6647
rect 4338 6644 4344 6656
rect 2271 6616 4344 6644
rect 2271 6613 2283 6616
rect 2225 6607 2283 6613
rect 4338 6604 4344 6616
rect 4396 6604 4402 6656
rect 4522 6604 4528 6656
rect 4580 6644 4586 6656
rect 5258 6644 5264 6656
rect 4580 6616 5264 6644
rect 4580 6604 4586 6616
rect 5258 6604 5264 6616
rect 5316 6644 5322 6656
rect 6196 6644 6224 6743
rect 7006 6740 7012 6792
rect 7064 6780 7070 6792
rect 7561 6783 7619 6789
rect 7561 6780 7573 6783
rect 7064 6752 7573 6780
rect 7064 6740 7070 6752
rect 7561 6749 7573 6752
rect 7607 6780 7619 6783
rect 8018 6780 8024 6792
rect 7607 6752 8024 6780
rect 7607 6749 7619 6752
rect 7561 6743 7619 6749
rect 8018 6740 8024 6752
rect 8076 6740 8082 6792
rect 5316 6616 6224 6644
rect 5316 6604 5322 6616
rect 6730 6604 6736 6656
rect 6788 6644 6794 6656
rect 8021 6647 8079 6653
rect 8021 6644 8033 6647
rect 6788 6616 8033 6644
rect 6788 6604 6794 6616
rect 8021 6613 8033 6616
rect 8067 6613 8079 6647
rect 8021 6607 8079 6613
rect 1104 6554 8832 6576
rect 1104 6502 3547 6554
rect 3599 6502 3611 6554
rect 3663 6502 3675 6554
rect 3727 6502 3739 6554
rect 3791 6502 3803 6554
rect 3855 6502 6144 6554
rect 6196 6502 6208 6554
rect 6260 6502 6272 6554
rect 6324 6502 6336 6554
rect 6388 6502 6400 6554
rect 6452 6502 8832 6554
rect 1104 6480 8832 6502
rect 2225 6443 2283 6449
rect 2225 6409 2237 6443
rect 2271 6440 2283 6443
rect 3234 6440 3240 6452
rect 2271 6412 3240 6440
rect 2271 6409 2283 6412
rect 2225 6403 2283 6409
rect 3234 6400 3240 6412
rect 3292 6400 3298 6452
rect 4985 6375 5043 6381
rect 3344 6344 4384 6372
rect 1397 6307 1455 6313
rect 1397 6273 1409 6307
rect 1443 6304 1455 6307
rect 1670 6304 1676 6316
rect 1443 6276 1676 6304
rect 1443 6273 1455 6276
rect 1397 6267 1455 6273
rect 1670 6264 1676 6276
rect 1728 6304 1734 6316
rect 3344 6304 3372 6344
rect 4258 6307 4316 6313
rect 4258 6304 4270 6307
rect 1728 6276 3372 6304
rect 3528 6276 4270 6304
rect 1728 6264 1734 6276
rect 2777 6239 2835 6245
rect 2777 6205 2789 6239
rect 2823 6236 2835 6239
rect 3528 6236 3556 6276
rect 4258 6273 4270 6276
rect 4304 6273 4316 6307
rect 4356 6304 4384 6344
rect 4985 6341 4997 6375
rect 5031 6372 5043 6375
rect 5166 6372 5172 6384
rect 5031 6344 5172 6372
rect 5031 6341 5043 6344
rect 4985 6335 5043 6341
rect 5166 6332 5172 6344
rect 5224 6332 5230 6384
rect 6641 6307 6699 6313
rect 6641 6304 6653 6307
rect 4356 6276 6653 6304
rect 4258 6267 4316 6273
rect 6641 6273 6653 6276
rect 6687 6304 6699 6307
rect 7190 6304 7196 6316
rect 6687 6276 7196 6304
rect 6687 6273 6699 6276
rect 6641 6267 6699 6273
rect 7190 6264 7196 6276
rect 7248 6264 7254 6316
rect 8113 6307 8171 6313
rect 8113 6273 8125 6307
rect 8159 6304 8171 6307
rect 8202 6304 8208 6316
rect 8159 6276 8208 6304
rect 8159 6273 8171 6276
rect 8113 6267 8171 6273
rect 8202 6264 8208 6276
rect 8260 6264 8266 6316
rect 4522 6236 4528 6248
rect 2823 6208 3556 6236
rect 4483 6208 4528 6236
rect 2823 6205 2835 6208
rect 2777 6199 2835 6205
rect 4522 6196 4528 6208
rect 4580 6196 4586 6248
rect 5077 6239 5135 6245
rect 5077 6205 5089 6239
rect 5123 6236 5135 6239
rect 5442 6236 5448 6248
rect 5123 6208 5448 6236
rect 5123 6205 5135 6208
rect 5077 6199 5135 6205
rect 5442 6196 5448 6208
rect 5500 6196 5506 6248
rect 5537 6239 5595 6245
rect 5537 6205 5549 6239
rect 5583 6236 5595 6239
rect 5718 6236 5724 6248
rect 5583 6208 5724 6236
rect 5583 6205 5595 6208
rect 5537 6199 5595 6205
rect 5718 6196 5724 6208
rect 5776 6236 5782 6248
rect 6730 6236 6736 6248
rect 5776 6208 6736 6236
rect 5776 6196 5782 6208
rect 6730 6196 6736 6208
rect 6788 6196 6794 6248
rect 6641 6171 6699 6177
rect 6641 6137 6653 6171
rect 6687 6137 6699 6171
rect 6641 6131 6699 6137
rect 1578 6100 1584 6112
rect 1539 6072 1584 6100
rect 1578 6060 1584 6072
rect 1636 6060 1642 6112
rect 2130 6100 2136 6112
rect 2091 6072 2136 6100
rect 2130 6060 2136 6072
rect 2188 6060 2194 6112
rect 3145 6103 3203 6109
rect 3145 6069 3157 6103
rect 3191 6100 3203 6103
rect 4246 6100 4252 6112
rect 3191 6072 4252 6100
rect 3191 6069 3203 6072
rect 3145 6063 3203 6069
rect 4246 6060 4252 6072
rect 4304 6060 4310 6112
rect 4338 6060 4344 6112
rect 4396 6100 4402 6112
rect 6656 6100 6684 6131
rect 4396 6072 6684 6100
rect 4396 6060 4402 6072
rect 1104 6010 8832 6032
rect 1104 5958 2248 6010
rect 2300 5958 2312 6010
rect 2364 5958 2376 6010
rect 2428 5958 2440 6010
rect 2492 5958 2504 6010
rect 2556 5958 4846 6010
rect 4898 5958 4910 6010
rect 4962 5958 4974 6010
rect 5026 5958 5038 6010
rect 5090 5958 5102 6010
rect 5154 5958 7443 6010
rect 7495 5958 7507 6010
rect 7559 5958 7571 6010
rect 7623 5958 7635 6010
rect 7687 5958 7699 6010
rect 7751 5958 8832 6010
rect 1104 5936 8832 5958
rect 2501 5899 2559 5905
rect 2501 5865 2513 5899
rect 2547 5896 2559 5899
rect 7282 5896 7288 5908
rect 2547 5868 7288 5896
rect 2547 5865 2559 5868
rect 2501 5859 2559 5865
rect 7282 5856 7288 5868
rect 7340 5856 7346 5908
rect 1857 5831 1915 5837
rect 1857 5797 1869 5831
rect 1903 5828 1915 5831
rect 7374 5828 7380 5840
rect 1903 5800 7380 5828
rect 1903 5797 1915 5800
rect 1857 5791 1915 5797
rect 7374 5788 7380 5800
rect 7432 5788 7438 5840
rect 2130 5720 2136 5772
rect 2188 5760 2194 5772
rect 4249 5763 4307 5769
rect 4249 5760 4261 5763
rect 2188 5732 4261 5760
rect 2188 5720 2194 5732
rect 4249 5729 4261 5732
rect 4295 5729 4307 5763
rect 4249 5723 4307 5729
rect 4801 5763 4859 5769
rect 4801 5729 4813 5763
rect 4847 5760 4859 5763
rect 4847 5732 5580 5760
rect 4847 5729 4859 5732
rect 4801 5723 4859 5729
rect 1673 5695 1731 5701
rect 1673 5661 1685 5695
rect 1719 5692 1731 5695
rect 2038 5692 2044 5704
rect 1719 5664 2044 5692
rect 1719 5661 1731 5664
rect 1673 5655 1731 5661
rect 2038 5652 2044 5664
rect 2096 5652 2102 5704
rect 2317 5695 2375 5701
rect 2317 5661 2329 5695
rect 2363 5692 2375 5695
rect 3145 5695 3203 5701
rect 2363 5664 2774 5692
rect 2363 5661 2375 5664
rect 2317 5655 2375 5661
rect 2746 5556 2774 5664
rect 3145 5661 3157 5695
rect 3191 5692 3203 5695
rect 4706 5692 4712 5704
rect 3191 5664 4712 5692
rect 3191 5661 3203 5664
rect 3145 5655 3203 5661
rect 4706 5652 4712 5664
rect 4764 5652 4770 5704
rect 5350 5652 5356 5704
rect 5408 5692 5414 5704
rect 5445 5695 5503 5701
rect 5445 5692 5457 5695
rect 5408 5664 5457 5692
rect 5408 5652 5414 5664
rect 5445 5661 5457 5664
rect 5491 5661 5503 5695
rect 5445 5655 5503 5661
rect 4154 5584 4160 5636
rect 4212 5624 4218 5636
rect 4341 5627 4399 5633
rect 4341 5624 4353 5627
rect 4212 5596 4353 5624
rect 4212 5584 4218 5596
rect 4341 5593 4353 5596
rect 4387 5593 4399 5627
rect 4341 5587 4399 5593
rect 4430 5584 4436 5636
rect 4488 5624 4494 5636
rect 5258 5624 5264 5636
rect 4488 5596 5264 5624
rect 4488 5584 4494 5596
rect 5258 5584 5264 5596
rect 5316 5584 5322 5636
rect 5552 5624 5580 5732
rect 5810 5720 5816 5772
rect 5868 5760 5874 5772
rect 5868 5732 7604 5760
rect 5868 5720 5874 5732
rect 5626 5652 5632 5704
rect 5684 5692 5690 5704
rect 6181 5695 6239 5701
rect 6181 5692 6193 5695
rect 5684 5664 6193 5692
rect 5684 5652 5690 5664
rect 6181 5661 6193 5664
rect 6227 5692 6239 5695
rect 6638 5692 6644 5704
rect 6227 5664 6644 5692
rect 6227 5661 6239 5664
rect 6181 5655 6239 5661
rect 6638 5652 6644 5664
rect 6696 5652 6702 5704
rect 7190 5692 7196 5704
rect 7151 5664 7196 5692
rect 7190 5652 7196 5664
rect 7248 5652 7254 5704
rect 7576 5692 7604 5732
rect 7834 5692 7840 5704
rect 7576 5664 7840 5692
rect 7834 5652 7840 5664
rect 7892 5692 7898 5704
rect 8110 5701 8116 5704
rect 8107 5692 8116 5701
rect 7892 5664 8116 5692
rect 7892 5652 7898 5664
rect 8107 5655 8116 5664
rect 8110 5652 8116 5655
rect 8168 5652 8174 5704
rect 5810 5624 5816 5636
rect 5552 5596 5816 5624
rect 5810 5584 5816 5596
rect 5868 5624 5874 5636
rect 5868 5596 6868 5624
rect 5868 5584 5874 5596
rect 3053 5559 3111 5565
rect 3053 5556 3065 5559
rect 2746 5528 3065 5556
rect 3053 5525 3065 5528
rect 3099 5556 3111 5559
rect 5902 5556 5908 5568
rect 3099 5528 5908 5556
rect 3099 5525 3111 5528
rect 3053 5519 3111 5525
rect 5902 5516 5908 5528
rect 5960 5516 5966 5568
rect 6730 5556 6736 5568
rect 6691 5528 6736 5556
rect 6730 5516 6736 5528
rect 6788 5516 6794 5568
rect 6840 5556 6868 5596
rect 7098 5584 7104 5636
rect 7156 5624 7162 5636
rect 7377 5627 7435 5633
rect 7377 5624 7389 5627
rect 7156 5596 7389 5624
rect 7156 5584 7162 5596
rect 7377 5593 7389 5596
rect 7423 5593 7435 5627
rect 7377 5587 7435 5593
rect 8202 5556 8208 5568
rect 6840 5528 8208 5556
rect 8202 5516 8208 5528
rect 8260 5516 8266 5568
rect 1104 5466 8832 5488
rect 1104 5414 3547 5466
rect 3599 5414 3611 5466
rect 3663 5414 3675 5466
rect 3727 5414 3739 5466
rect 3791 5414 3803 5466
rect 3855 5414 6144 5466
rect 6196 5414 6208 5466
rect 6260 5414 6272 5466
rect 6324 5414 6336 5466
rect 6388 5414 6400 5466
rect 6452 5414 8832 5466
rect 1104 5392 8832 5414
rect 1854 5312 1860 5364
rect 1912 5352 1918 5364
rect 1912 5324 2774 5352
rect 1912 5312 1918 5324
rect 2746 5284 2774 5324
rect 2958 5312 2964 5364
rect 3016 5352 3022 5364
rect 4430 5352 4436 5364
rect 3016 5324 4436 5352
rect 3016 5312 3022 5324
rect 4430 5312 4436 5324
rect 4488 5312 4494 5364
rect 4522 5312 4528 5364
rect 4580 5352 4586 5364
rect 5077 5355 5135 5361
rect 5077 5352 5089 5355
rect 4580 5324 5089 5352
rect 4580 5312 4586 5324
rect 5077 5321 5089 5324
rect 5123 5321 5135 5355
rect 5077 5315 5135 5321
rect 3786 5284 3792 5296
rect 2746 5256 3792 5284
rect 3786 5244 3792 5256
rect 3844 5244 3850 5296
rect 6822 5284 6828 5296
rect 3896 5256 6828 5284
rect 1664 5219 1722 5225
rect 1664 5185 1676 5219
rect 1710 5216 1722 5219
rect 1710 5188 2443 5216
rect 1710 5185 1722 5188
rect 1664 5179 1722 5185
rect 1394 5148 1400 5160
rect 1355 5120 1400 5148
rect 1394 5108 1400 5120
rect 1452 5108 1458 5160
rect 2415 5148 2443 5188
rect 2774 5176 2780 5228
rect 2832 5216 2838 5228
rect 3896 5216 3924 5256
rect 6822 5244 6828 5256
rect 6880 5244 6886 5296
rect 6914 5244 6920 5296
rect 6972 5244 6978 5296
rect 7374 5284 7380 5296
rect 7335 5256 7380 5284
rect 7374 5244 7380 5256
rect 7432 5244 7438 5296
rect 2832 5188 3924 5216
rect 3964 5219 4022 5225
rect 2832 5176 2838 5188
rect 3964 5185 3976 5219
rect 4010 5216 4022 5219
rect 6932 5216 6960 5244
rect 7926 5216 7932 5228
rect 4010 5188 5488 5216
rect 6932 5188 7932 5216
rect 4010 5185 4022 5188
rect 3964 5179 4022 5185
rect 5460 5157 5488 5188
rect 7926 5176 7932 5188
rect 7984 5176 7990 5228
rect 3145 5151 3203 5157
rect 3145 5148 3157 5151
rect 2415 5120 3157 5148
rect 3145 5117 3157 5120
rect 3191 5117 3203 5151
rect 3145 5111 3203 5117
rect 3697 5151 3755 5157
rect 3697 5117 3709 5151
rect 3743 5117 3755 5151
rect 3697 5111 3755 5117
rect 5445 5151 5503 5157
rect 5445 5117 5457 5151
rect 5491 5117 5503 5151
rect 6362 5148 6368 5160
rect 6323 5120 6368 5148
rect 5445 5111 5503 5117
rect 2777 5015 2835 5021
rect 2777 4981 2789 5015
rect 2823 5012 2835 5015
rect 3712 5012 3740 5111
rect 6362 5108 6368 5120
rect 6420 5108 6426 5160
rect 6546 5108 6552 5160
rect 6604 5148 6610 5160
rect 6917 5151 6975 5157
rect 6917 5148 6929 5151
rect 6604 5120 6929 5148
rect 6604 5108 6610 5120
rect 6917 5117 6929 5120
rect 6963 5117 6975 5151
rect 6917 5111 6975 5117
rect 5994 5040 6000 5092
rect 6052 5080 6058 5092
rect 6457 5083 6515 5089
rect 6457 5080 6469 5083
rect 6052 5052 6469 5080
rect 6052 5040 6058 5052
rect 6457 5049 6469 5052
rect 6503 5049 6515 5083
rect 6457 5043 6515 5049
rect 7190 5040 7196 5092
rect 7248 5080 7254 5092
rect 7469 5083 7527 5089
rect 7469 5080 7481 5083
rect 7248 5052 7481 5080
rect 7248 5040 7254 5052
rect 7469 5049 7481 5052
rect 7515 5049 7527 5083
rect 7469 5043 7527 5049
rect 2823 4984 3740 5012
rect 2823 4981 2835 4984
rect 2777 4975 2835 4981
rect 3878 4972 3884 5024
rect 3936 5012 3942 5024
rect 4430 5012 4436 5024
rect 3936 4984 4436 5012
rect 3936 4972 3942 4984
rect 4430 4972 4436 4984
rect 4488 4972 4494 5024
rect 1104 4922 8832 4944
rect 1104 4870 2248 4922
rect 2300 4870 2312 4922
rect 2364 4870 2376 4922
rect 2428 4870 2440 4922
rect 2492 4870 2504 4922
rect 2556 4870 4846 4922
rect 4898 4870 4910 4922
rect 4962 4870 4974 4922
rect 5026 4870 5038 4922
rect 5090 4870 5102 4922
rect 5154 4870 7443 4922
rect 7495 4870 7507 4922
rect 7559 4870 7571 4922
rect 7623 4870 7635 4922
rect 7687 4870 7699 4922
rect 7751 4870 8832 4922
rect 1104 4848 8832 4870
rect 1673 4811 1731 4817
rect 1673 4777 1685 4811
rect 1719 4808 1731 4811
rect 6362 4808 6368 4820
rect 1719 4780 6368 4808
rect 1719 4777 1731 4780
rect 1673 4771 1731 4777
rect 6362 4768 6368 4780
rect 6420 4768 6426 4820
rect 1780 4712 5948 4740
rect 1780 4613 1808 4712
rect 2038 4632 2044 4684
rect 2096 4672 2102 4684
rect 2225 4675 2283 4681
rect 2225 4672 2237 4675
rect 2096 4644 2237 4672
rect 2096 4632 2102 4644
rect 2225 4641 2237 4644
rect 2271 4641 2283 4675
rect 2225 4635 2283 4641
rect 5920 4672 5948 4712
rect 7377 4675 7435 4681
rect 7377 4672 7389 4675
rect 5920 4644 7389 4672
rect 1765 4607 1823 4613
rect 1765 4573 1777 4607
rect 1811 4573 1823 4607
rect 1765 4567 1823 4573
rect 2409 4607 2467 4613
rect 2409 4573 2421 4607
rect 2455 4604 2467 4607
rect 2774 4604 2780 4616
rect 2455 4576 2780 4604
rect 2455 4573 2467 4576
rect 2409 4567 2467 4573
rect 2774 4564 2780 4576
rect 2832 4564 2838 4616
rect 3068 4576 3280 4604
rect 2590 4496 2596 4548
rect 2648 4536 2654 4548
rect 3068 4536 3096 4576
rect 2648 4508 3096 4536
rect 3145 4539 3203 4545
rect 2648 4496 2654 4508
rect 3145 4505 3157 4539
rect 3191 4505 3203 4539
rect 3252 4536 3280 4576
rect 3970 4564 3976 4616
rect 4028 4604 4034 4616
rect 4341 4607 4399 4613
rect 4028 4576 4292 4604
rect 4028 4564 4034 4576
rect 3789 4539 3847 4545
rect 3789 4536 3801 4539
rect 3252 4508 3801 4536
rect 3145 4499 3203 4505
rect 3789 4505 3801 4508
rect 3835 4505 3847 4539
rect 3789 4499 3847 4505
rect 3881 4539 3939 4545
rect 3881 4505 3893 4539
rect 3927 4536 3939 4539
rect 4154 4536 4160 4548
rect 3927 4508 4160 4536
rect 3927 4505 3939 4508
rect 3881 4499 3939 4505
rect 2958 4428 2964 4480
rect 3016 4468 3022 4480
rect 3053 4471 3111 4477
rect 3053 4468 3065 4471
rect 3016 4440 3065 4468
rect 3016 4428 3022 4440
rect 3053 4437 3065 4440
rect 3099 4437 3111 4471
rect 3160 4468 3188 4499
rect 4154 4496 4160 4508
rect 4212 4496 4218 4548
rect 4264 4536 4292 4576
rect 4341 4573 4353 4607
rect 4387 4604 4399 4607
rect 4522 4604 4528 4616
rect 4387 4576 4528 4604
rect 4387 4573 4399 4576
rect 4341 4567 4399 4573
rect 4522 4564 4528 4576
rect 4580 4564 4586 4616
rect 5353 4607 5411 4613
rect 5353 4604 5365 4607
rect 4632 4576 5365 4604
rect 4632 4536 4660 4576
rect 5353 4573 5365 4576
rect 5399 4604 5411 4607
rect 5810 4604 5816 4616
rect 5399 4576 5816 4604
rect 5399 4573 5411 4576
rect 5353 4567 5411 4573
rect 5810 4564 5816 4576
rect 5868 4564 5874 4616
rect 5920 4604 5948 4644
rect 7377 4641 7389 4644
rect 7423 4641 7435 4675
rect 7377 4635 7435 4641
rect 6089 4607 6147 4613
rect 6089 4604 6101 4607
rect 5920 4576 6101 4604
rect 6089 4573 6101 4576
rect 6135 4573 6147 4607
rect 6822 4604 6828 4616
rect 6783 4576 6828 4604
rect 6089 4567 6147 4573
rect 6822 4564 6828 4576
rect 6880 4604 6886 4616
rect 7837 4607 7895 4613
rect 7837 4604 7849 4607
rect 6880 4576 7849 4604
rect 6880 4564 6886 4576
rect 7837 4573 7849 4576
rect 7883 4573 7895 4607
rect 7837 4567 7895 4573
rect 4798 4536 4804 4548
rect 4264 4508 4660 4536
rect 4759 4508 4804 4536
rect 4798 4496 4804 4508
rect 4856 4496 4862 4548
rect 4893 4539 4951 4545
rect 4893 4505 4905 4539
rect 4939 4505 4951 4539
rect 5902 4536 5908 4548
rect 5863 4508 5908 4536
rect 4893 4499 4951 4505
rect 4338 4468 4344 4480
rect 3160 4440 4344 4468
rect 3053 4431 3111 4437
rect 4338 4428 4344 4440
rect 4396 4468 4402 4480
rect 4908 4468 4936 4499
rect 5902 4496 5908 4508
rect 5960 4496 5966 4548
rect 7282 4536 7288 4548
rect 7243 4508 7288 4536
rect 7282 4496 7288 4508
rect 7340 4496 7346 4548
rect 4396 4440 4936 4468
rect 4396 4428 4402 4440
rect 1104 4378 8832 4400
rect 1104 4326 3547 4378
rect 3599 4326 3611 4378
rect 3663 4326 3675 4378
rect 3727 4326 3739 4378
rect 3791 4326 3803 4378
rect 3855 4326 6144 4378
rect 6196 4326 6208 4378
rect 6260 4326 6272 4378
rect 6324 4326 6336 4378
rect 6388 4326 6400 4378
rect 6452 4326 8832 4378
rect 1104 4304 8832 4326
rect 1673 4267 1731 4273
rect 1673 4233 1685 4267
rect 1719 4264 1731 4267
rect 4154 4264 4160 4276
rect 1719 4236 4160 4264
rect 1719 4233 1731 4236
rect 1673 4227 1731 4233
rect 4154 4224 4160 4236
rect 4212 4224 4218 4276
rect 4522 4224 4528 4276
rect 4580 4264 4586 4276
rect 4580 4236 5396 4264
rect 4580 4224 4586 4236
rect 1581 4199 1639 4205
rect 1581 4165 1593 4199
rect 1627 4196 1639 4199
rect 4798 4196 4804 4208
rect 1627 4168 4804 4196
rect 1627 4165 1639 4168
rect 1581 4159 1639 4165
rect 4798 4156 4804 4168
rect 4856 4156 4862 4208
rect 5368 4140 5396 4236
rect 2400 4131 2458 4137
rect 2400 4097 2412 4131
rect 2446 4128 2458 4131
rect 4430 4128 4436 4140
rect 2446 4100 3924 4128
rect 4391 4100 4436 4128
rect 2446 4097 2458 4100
rect 2400 4091 2458 4097
rect 1854 4020 1860 4072
rect 1912 4060 1918 4072
rect 3896 4069 3924 4100
rect 4430 4088 4436 4100
rect 4488 4088 4494 4140
rect 4617 4131 4675 4137
rect 4617 4097 4629 4131
rect 4663 4097 4675 4131
rect 5350 4128 5356 4140
rect 5263 4100 5356 4128
rect 4617 4091 4675 4097
rect 2133 4063 2191 4069
rect 2133 4060 2145 4063
rect 1912 4032 2145 4060
rect 1912 4020 1918 4032
rect 2133 4029 2145 4032
rect 2179 4029 2191 4063
rect 2133 4023 2191 4029
rect 3881 4063 3939 4069
rect 3881 4029 3893 4063
rect 3927 4029 3939 4063
rect 3881 4023 3939 4029
rect 4154 4020 4160 4072
rect 4212 4060 4218 4072
rect 4632 4060 4660 4091
rect 5350 4088 5356 4100
rect 5408 4088 5414 4140
rect 5902 4088 5908 4140
rect 5960 4128 5966 4140
rect 6457 4131 6515 4137
rect 6457 4128 6469 4131
rect 5960 4100 6469 4128
rect 5960 4088 5966 4100
rect 6457 4097 6469 4100
rect 6503 4097 6515 4131
rect 6457 4091 6515 4097
rect 6546 4088 6552 4140
rect 6604 4128 6610 4140
rect 7929 4131 7987 4137
rect 7929 4128 7941 4131
rect 6604 4100 7941 4128
rect 6604 4088 6610 4100
rect 7929 4097 7941 4100
rect 7975 4128 7987 4131
rect 8202 4128 8208 4140
rect 7975 4100 8208 4128
rect 7975 4097 7987 4100
rect 7929 4091 7987 4097
rect 8202 4088 8208 4100
rect 8260 4088 8266 4140
rect 4212 4032 4660 4060
rect 4212 4020 4218 4032
rect 5994 3992 6000 4004
rect 3436 3964 6000 3992
rect 2774 3884 2780 3936
rect 2832 3924 2838 3936
rect 3436 3924 3464 3964
rect 5994 3952 6000 3964
rect 6052 3992 6058 4004
rect 6457 3995 6515 4001
rect 6457 3992 6469 3995
rect 6052 3964 6469 3992
rect 6052 3952 6058 3964
rect 6457 3961 6469 3964
rect 6503 3961 6515 3995
rect 6457 3955 6515 3961
rect 2832 3896 3464 3924
rect 3513 3927 3571 3933
rect 2832 3884 2838 3896
rect 3513 3893 3525 3927
rect 3559 3924 3571 3927
rect 3970 3924 3976 3936
rect 3559 3896 3976 3924
rect 3559 3893 3571 3896
rect 3513 3887 3571 3893
rect 3970 3884 3976 3896
rect 4028 3884 4034 3936
rect 1104 3834 8832 3856
rect 1104 3782 2248 3834
rect 2300 3782 2312 3834
rect 2364 3782 2376 3834
rect 2428 3782 2440 3834
rect 2492 3782 2504 3834
rect 2556 3782 4846 3834
rect 4898 3782 4910 3834
rect 4962 3782 4974 3834
rect 5026 3782 5038 3834
rect 5090 3782 5102 3834
rect 5154 3782 7443 3834
rect 7495 3782 7507 3834
rect 7559 3782 7571 3834
rect 7623 3782 7635 3834
rect 7687 3782 7699 3834
rect 7751 3782 8832 3834
rect 1104 3760 8832 3782
rect 1854 3720 1860 3732
rect 1815 3692 1860 3720
rect 1854 3680 1860 3692
rect 1912 3680 1918 3732
rect 2038 3680 2044 3732
rect 2096 3720 2102 3732
rect 2096 3692 5948 3720
rect 2096 3680 2102 3692
rect 4338 3652 4344 3664
rect 4299 3624 4344 3652
rect 4338 3612 4344 3624
rect 4396 3612 4402 3664
rect 1489 3587 1547 3593
rect 1489 3553 1501 3587
rect 1535 3553 1547 3587
rect 1489 3547 1547 3553
rect 3237 3587 3295 3593
rect 3237 3553 3249 3587
rect 3283 3584 3295 3587
rect 3418 3584 3424 3596
rect 3283 3556 3424 3584
rect 3283 3553 3295 3556
rect 3237 3547 3295 3553
rect 1504 3516 1532 3547
rect 2970 3519 3028 3525
rect 2970 3516 2982 3519
rect 1504 3488 2982 3516
rect 2970 3485 2982 3488
rect 3016 3485 3028 3519
rect 2970 3479 3028 3485
rect 2682 3408 2688 3460
rect 2740 3448 2746 3460
rect 3252 3448 3280 3547
rect 3418 3544 3424 3556
rect 3476 3584 3482 3596
rect 4522 3584 4528 3596
rect 3476 3556 4528 3584
rect 3476 3544 3482 3556
rect 4522 3544 4528 3556
rect 4580 3544 4586 3596
rect 4430 3516 4436 3528
rect 4391 3488 4436 3516
rect 4430 3476 4436 3488
rect 4488 3476 4494 3528
rect 5810 3516 5816 3528
rect 5771 3488 5816 3516
rect 5810 3476 5816 3488
rect 5868 3476 5874 3528
rect 5920 3516 5948 3692
rect 6641 3519 6699 3525
rect 6641 3516 6653 3519
rect 5920 3488 6653 3516
rect 6641 3485 6653 3488
rect 6687 3516 6699 3519
rect 6914 3516 6920 3528
rect 6687 3488 6920 3516
rect 6687 3485 6699 3488
rect 6641 3479 6699 3485
rect 6914 3476 6920 3488
rect 6972 3476 6978 3528
rect 8113 3519 8171 3525
rect 8113 3485 8125 3519
rect 8159 3516 8171 3519
rect 8294 3516 8300 3528
rect 8159 3488 8300 3516
rect 8159 3485 8171 3488
rect 8113 3479 8171 3485
rect 8294 3476 8300 3488
rect 8352 3476 8358 3528
rect 6546 3448 6552 3460
rect 2740 3420 3280 3448
rect 6507 3420 6552 3448
rect 2740 3408 2746 3420
rect 6546 3408 6552 3420
rect 6604 3408 6610 3460
rect 1104 3290 8832 3312
rect 1104 3238 3547 3290
rect 3599 3238 3611 3290
rect 3663 3238 3675 3290
rect 3727 3238 3739 3290
rect 3791 3238 3803 3290
rect 3855 3238 6144 3290
rect 6196 3238 6208 3290
rect 6260 3238 6272 3290
rect 6324 3238 6336 3290
rect 6388 3238 6400 3290
rect 6452 3238 8832 3290
rect 1104 3216 8832 3238
rect 2866 3136 2872 3188
rect 2924 3176 2930 3188
rect 4338 3176 4344 3188
rect 2924 3148 4344 3176
rect 2924 3136 2930 3148
rect 4338 3136 4344 3148
rect 4396 3136 4402 3188
rect 5350 3136 5356 3188
rect 5408 3176 5414 3188
rect 6365 3179 6423 3185
rect 6365 3176 6377 3179
rect 5408 3148 6377 3176
rect 5408 3136 5414 3148
rect 6365 3145 6377 3148
rect 6411 3176 6423 3179
rect 6822 3176 6828 3188
rect 6411 3148 6828 3176
rect 6411 3145 6423 3148
rect 6365 3139 6423 3145
rect 6822 3136 6828 3148
rect 6880 3136 6886 3188
rect 1670 3068 1676 3120
rect 1728 3108 1734 3120
rect 1857 3111 1915 3117
rect 1857 3108 1869 3111
rect 1728 3080 1869 3108
rect 1728 3068 1734 3080
rect 1857 3077 1869 3080
rect 1903 3077 1915 3111
rect 1857 3071 1915 3077
rect 2041 3111 2099 3117
rect 2041 3077 2053 3111
rect 2087 3108 2099 3111
rect 6546 3108 6552 3120
rect 2087 3080 6552 3108
rect 2087 3077 2099 3080
rect 2041 3071 2099 3077
rect 6546 3068 6552 3080
rect 6604 3068 6610 3120
rect 6914 3108 6920 3120
rect 6875 3080 6920 3108
rect 6914 3068 6920 3080
rect 6972 3068 6978 3120
rect 7190 3108 7196 3120
rect 7151 3080 7196 3108
rect 7190 3068 7196 3080
rect 7248 3068 7254 3120
rect 2593 3043 2651 3049
rect 2593 3009 2605 3043
rect 2639 3040 2651 3043
rect 2682 3040 2688 3052
rect 2639 3012 2688 3040
rect 2639 3009 2651 3012
rect 2593 3003 2651 3009
rect 2682 3000 2688 3012
rect 2740 3000 2746 3052
rect 2860 3043 2918 3049
rect 2860 3009 2872 3043
rect 2906 3040 2918 3043
rect 4893 3043 4951 3049
rect 2906 3012 4384 3040
rect 2906 3009 2918 3012
rect 2860 3003 2918 3009
rect 4356 2981 4384 3012
rect 4893 3009 4905 3043
rect 4939 3040 4951 3043
rect 5258 3040 5264 3052
rect 4939 3012 5264 3040
rect 4939 3009 4951 3012
rect 4893 3003 4951 3009
rect 5258 3000 5264 3012
rect 5316 3000 5322 3052
rect 7837 3043 7895 3049
rect 7837 3009 7849 3043
rect 7883 3040 7895 3043
rect 7926 3040 7932 3052
rect 7883 3012 7932 3040
rect 7883 3009 7895 3012
rect 7837 3003 7895 3009
rect 7926 3000 7932 3012
rect 7984 3000 7990 3052
rect 4341 2975 4399 2981
rect 4341 2941 4353 2975
rect 4387 2941 4399 2975
rect 4341 2935 4399 2941
rect 5721 2975 5779 2981
rect 5721 2941 5733 2975
rect 5767 2972 5779 2975
rect 5767 2944 6960 2972
rect 5767 2941 5779 2944
rect 5721 2935 5779 2941
rect 6932 2916 6960 2944
rect 3602 2864 3608 2916
rect 3660 2904 3666 2916
rect 4430 2904 4436 2916
rect 3660 2876 4436 2904
rect 3660 2864 3666 2876
rect 4430 2864 4436 2876
rect 4488 2864 4494 2916
rect 6914 2864 6920 2916
rect 6972 2864 6978 2916
rect 934 2796 940 2848
rect 992 2836 998 2848
rect 1946 2836 1952 2848
rect 992 2808 1952 2836
rect 992 2796 998 2808
rect 1946 2796 1952 2808
rect 2004 2836 2010 2848
rect 3878 2836 3884 2848
rect 2004 2808 3884 2836
rect 2004 2796 2010 2808
rect 3878 2796 3884 2808
rect 3936 2796 3942 2848
rect 3973 2839 4031 2845
rect 3973 2805 3985 2839
rect 4019 2836 4031 2839
rect 4706 2836 4712 2848
rect 4019 2808 4712 2836
rect 4019 2805 4031 2808
rect 3973 2799 4031 2805
rect 4706 2796 4712 2808
rect 4764 2796 4770 2848
rect 6638 2796 6644 2848
rect 6696 2836 6702 2848
rect 6822 2836 6828 2848
rect 6696 2808 6828 2836
rect 6696 2796 6702 2808
rect 6822 2796 6828 2808
rect 6880 2796 6886 2848
rect 1104 2746 8832 2768
rect 1104 2694 2248 2746
rect 2300 2694 2312 2746
rect 2364 2694 2376 2746
rect 2428 2694 2440 2746
rect 2492 2694 2504 2746
rect 2556 2694 4846 2746
rect 4898 2694 4910 2746
rect 4962 2694 4974 2746
rect 5026 2694 5038 2746
rect 5090 2694 5102 2746
rect 5154 2694 7443 2746
rect 7495 2694 7507 2746
rect 7559 2694 7571 2746
rect 7623 2694 7635 2746
rect 7687 2694 7699 2746
rect 7751 2694 8832 2746
rect 1104 2672 8832 2694
rect 2501 2635 2559 2641
rect 2501 2601 2513 2635
rect 2547 2632 2559 2635
rect 2590 2632 2596 2644
rect 2547 2604 2596 2632
rect 2547 2601 2559 2604
rect 2501 2595 2559 2601
rect 2590 2592 2596 2604
rect 2648 2592 2654 2644
rect 5258 2632 5264 2644
rect 5219 2604 5264 2632
rect 5258 2592 5264 2604
rect 5316 2592 5322 2644
rect 6546 2592 6552 2644
rect 6604 2632 6610 2644
rect 6604 2604 7696 2632
rect 6604 2592 6610 2604
rect 6641 2567 6699 2573
rect 6641 2533 6653 2567
rect 6687 2564 6699 2567
rect 7006 2564 7012 2576
rect 6687 2536 7012 2564
rect 6687 2533 6699 2536
rect 6641 2527 6699 2533
rect 7006 2524 7012 2536
rect 7064 2524 7070 2576
rect 7668 2573 7696 2604
rect 7653 2567 7711 2573
rect 7653 2533 7665 2567
rect 7699 2533 7711 2567
rect 7653 2527 7711 2533
rect 1765 2499 1823 2505
rect 1765 2465 1777 2499
rect 1811 2496 1823 2499
rect 1811 2468 3740 2496
rect 1811 2465 1823 2468
rect 1765 2459 1823 2465
rect 2317 2431 2375 2437
rect 2317 2397 2329 2431
rect 2363 2428 2375 2431
rect 3602 2428 3608 2440
rect 2363 2400 3608 2428
rect 2363 2397 2375 2400
rect 2317 2391 2375 2397
rect 3602 2388 3608 2400
rect 3660 2388 3666 2440
rect 3050 2360 3056 2372
rect 3011 2332 3056 2360
rect 3050 2320 3056 2332
rect 3108 2320 3114 2372
rect 1854 2252 1860 2304
rect 1912 2292 1918 2304
rect 3142 2292 3148 2304
rect 1912 2264 1957 2292
rect 3103 2264 3148 2292
rect 1912 2252 1918 2264
rect 3142 2252 3148 2264
rect 3200 2252 3206 2304
rect 3712 2292 3740 2468
rect 3878 2456 3884 2508
rect 3936 2456 3942 2508
rect 5718 2456 5724 2508
rect 5776 2496 5782 2508
rect 6549 2499 6607 2505
rect 6549 2496 6561 2499
rect 5776 2468 6561 2496
rect 5776 2456 5782 2468
rect 6549 2465 6561 2468
rect 6595 2465 6607 2499
rect 6549 2459 6607 2465
rect 7101 2499 7159 2505
rect 7101 2465 7113 2499
rect 7147 2496 7159 2499
rect 7834 2496 7840 2508
rect 7147 2468 7840 2496
rect 7147 2465 7159 2468
rect 7101 2459 7159 2465
rect 7834 2456 7840 2468
rect 7892 2456 7898 2508
rect 8113 2499 8171 2505
rect 8113 2465 8125 2499
rect 8159 2496 8171 2499
rect 8294 2496 8300 2508
rect 8159 2468 8300 2496
rect 8159 2465 8171 2468
rect 8113 2459 8171 2465
rect 8294 2456 8300 2468
rect 8352 2456 8358 2508
rect 4338 2428 4344 2440
rect 4299 2400 4344 2428
rect 4338 2388 4344 2400
rect 4396 2388 4402 2440
rect 4706 2428 4712 2440
rect 4667 2400 4712 2428
rect 4706 2388 4712 2400
rect 4764 2388 4770 2440
rect 3970 2360 3976 2372
rect 3931 2332 3976 2360
rect 3970 2320 3976 2332
rect 4028 2320 4034 2372
rect 4246 2360 4252 2372
rect 4207 2332 4252 2360
rect 4246 2320 4252 2332
rect 4304 2320 4310 2372
rect 4522 2320 4528 2372
rect 4580 2360 4586 2372
rect 5077 2363 5135 2369
rect 5077 2360 5089 2363
rect 4580 2332 5089 2360
rect 4580 2320 4586 2332
rect 5077 2329 5089 2332
rect 5123 2329 5135 2363
rect 5077 2323 5135 2329
rect 7561 2363 7619 2369
rect 7561 2329 7573 2363
rect 7607 2329 7619 2363
rect 7561 2323 7619 2329
rect 7576 2292 7604 2323
rect 3712 2264 7604 2292
rect 1104 2202 8832 2224
rect 1104 2150 3547 2202
rect 3599 2150 3611 2202
rect 3663 2150 3675 2202
rect 3727 2150 3739 2202
rect 3791 2150 3803 2202
rect 3855 2150 6144 2202
rect 6196 2150 6208 2202
rect 6260 2150 6272 2202
rect 6324 2150 6336 2202
rect 6388 2150 6400 2202
rect 6452 2150 8832 2202
rect 1104 2128 8832 2150
rect 1854 2048 1860 2100
rect 1912 2088 1918 2100
rect 1912 2060 2774 2088
rect 1912 2048 1918 2060
rect 2746 2020 2774 2060
rect 3142 2048 3148 2100
rect 3200 2088 3206 2100
rect 5626 2088 5632 2100
rect 3200 2060 5632 2088
rect 3200 2048 3206 2060
rect 5626 2048 5632 2060
rect 5684 2048 5690 2100
rect 7190 2020 7196 2032
rect 2746 1992 7196 2020
rect 7190 1980 7196 1992
rect 7248 1980 7254 2032
rect 3050 1708 3056 1760
rect 3108 1748 3114 1760
rect 8938 1748 8944 1760
rect 3108 1720 8944 1748
rect 3108 1708 3114 1720
rect 8938 1708 8944 1720
rect 8996 1708 9002 1760
rect 4062 1300 4068 1352
rect 4120 1340 4126 1352
rect 6546 1340 6552 1352
rect 4120 1312 6552 1340
rect 4120 1300 4126 1312
rect 6546 1300 6552 1312
rect 6604 1300 6610 1352
<< via1 >>
rect 2248 27718 2300 27770
rect 2312 27718 2364 27770
rect 2376 27718 2428 27770
rect 2440 27718 2492 27770
rect 2504 27718 2556 27770
rect 4846 27718 4898 27770
rect 4910 27718 4962 27770
rect 4974 27718 5026 27770
rect 5038 27718 5090 27770
rect 5102 27718 5154 27770
rect 7443 27718 7495 27770
rect 7507 27718 7559 27770
rect 7571 27718 7623 27770
rect 7635 27718 7687 27770
rect 7699 27718 7751 27770
rect 2596 27548 2648 27600
rect 5816 27548 5868 27600
rect 2044 27480 2096 27532
rect 5540 27480 5592 27532
rect 4068 27412 4120 27464
rect 4160 27412 4212 27464
rect 7840 27455 7892 27464
rect 7840 27421 7849 27455
rect 7849 27421 7883 27455
rect 7883 27421 7892 27455
rect 7840 27412 7892 27421
rect 3884 27344 3936 27396
rect 4528 27387 4580 27396
rect 4528 27353 4537 27387
rect 4537 27353 4571 27387
rect 4571 27353 4580 27387
rect 4528 27344 4580 27353
rect 5448 27344 5500 27396
rect 6828 27344 6880 27396
rect 7380 27387 7432 27396
rect 7380 27353 7389 27387
rect 7389 27353 7423 27387
rect 7423 27353 7432 27387
rect 7380 27344 7432 27353
rect 2688 27319 2740 27328
rect 2688 27285 2697 27319
rect 2697 27285 2731 27319
rect 2731 27285 2740 27319
rect 2688 27276 2740 27285
rect 3976 27319 4028 27328
rect 3976 27285 3985 27319
rect 3985 27285 4019 27319
rect 4019 27285 4028 27319
rect 3976 27276 4028 27285
rect 5632 27319 5684 27328
rect 5632 27285 5641 27319
rect 5641 27285 5675 27319
rect 5675 27285 5684 27319
rect 5632 27276 5684 27285
rect 6920 27276 6972 27328
rect 3547 27174 3599 27226
rect 3611 27174 3663 27226
rect 3675 27174 3727 27226
rect 3739 27174 3791 27226
rect 3803 27174 3855 27226
rect 6144 27174 6196 27226
rect 6208 27174 6260 27226
rect 6272 27174 6324 27226
rect 6336 27174 6388 27226
rect 6400 27174 6452 27226
rect 2044 27115 2096 27124
rect 2044 27081 2053 27115
rect 2053 27081 2087 27115
rect 2087 27081 2096 27115
rect 2044 27072 2096 27081
rect 7380 27072 7432 27124
rect 5448 27004 5500 27056
rect 6460 27004 6512 27056
rect 3240 26979 3292 26988
rect 3240 26945 3249 26979
rect 3249 26945 3283 26979
rect 3283 26945 3292 26979
rect 3240 26936 3292 26945
rect 3424 26936 3476 26988
rect 4528 26979 4580 26988
rect 4528 26945 4537 26979
rect 4537 26945 4571 26979
rect 4571 26945 4580 26979
rect 4528 26936 4580 26945
rect 5540 26936 5592 26988
rect 5816 26936 5868 26988
rect 7932 26936 7984 26988
rect 7196 26868 7248 26920
rect 5908 26800 5960 26852
rect 6828 26800 6880 26852
rect 2780 26732 2832 26784
rect 5172 26732 5224 26784
rect 8208 26868 8260 26920
rect 2248 26630 2300 26682
rect 2312 26630 2364 26682
rect 2376 26630 2428 26682
rect 2440 26630 2492 26682
rect 2504 26630 2556 26682
rect 4846 26630 4898 26682
rect 4910 26630 4962 26682
rect 4974 26630 5026 26682
rect 5038 26630 5090 26682
rect 5102 26630 5154 26682
rect 7443 26630 7495 26682
rect 7507 26630 7559 26682
rect 7571 26630 7623 26682
rect 7635 26630 7687 26682
rect 7699 26630 7751 26682
rect 2596 26571 2648 26580
rect 2596 26537 2605 26571
rect 2605 26537 2639 26571
rect 2639 26537 2648 26571
rect 2596 26528 2648 26537
rect 2780 26528 2832 26580
rect 3240 26460 3292 26512
rect 3976 26435 4028 26444
rect 3976 26401 3985 26435
rect 3985 26401 4019 26435
rect 4019 26401 4028 26435
rect 3976 26392 4028 26401
rect 4160 26324 4212 26376
rect 4068 26256 4120 26308
rect 5908 26367 5960 26376
rect 5908 26333 5917 26367
rect 5917 26333 5951 26367
rect 5951 26333 5960 26367
rect 5908 26324 5960 26333
rect 6460 26503 6512 26512
rect 6460 26469 6469 26503
rect 6469 26469 6503 26503
rect 6503 26469 6512 26503
rect 6460 26460 6512 26469
rect 6920 26324 6972 26376
rect 7932 26367 7984 26376
rect 7932 26333 7941 26367
rect 7941 26333 7975 26367
rect 7975 26333 7984 26367
rect 7932 26324 7984 26333
rect 5264 26188 5316 26240
rect 5908 26188 5960 26240
rect 6644 26188 6696 26240
rect 3547 26086 3599 26138
rect 3611 26086 3663 26138
rect 3675 26086 3727 26138
rect 3739 26086 3791 26138
rect 3803 26086 3855 26138
rect 6144 26086 6196 26138
rect 6208 26086 6260 26138
rect 6272 26086 6324 26138
rect 6336 26086 6388 26138
rect 6400 26086 6452 26138
rect 2044 25984 2096 26036
rect 2688 25916 2740 25968
rect 4068 25916 4120 25968
rect 3424 25848 3476 25900
rect 4160 25848 4212 25900
rect 7196 25984 7248 26036
rect 7012 25959 7064 25968
rect 7012 25925 7021 25959
rect 7021 25925 7055 25959
rect 7055 25925 7064 25959
rect 7012 25916 7064 25925
rect 7288 25959 7340 25968
rect 7288 25925 7297 25959
rect 7297 25925 7331 25959
rect 7331 25925 7340 25959
rect 7288 25916 7340 25925
rect 5264 25891 5316 25900
rect 5264 25857 5273 25891
rect 5273 25857 5307 25891
rect 5307 25857 5316 25891
rect 5264 25848 5316 25857
rect 6920 25848 6972 25900
rect 7840 25848 7892 25900
rect 5724 25780 5776 25832
rect 5264 25712 5316 25764
rect 2248 25542 2300 25594
rect 2312 25542 2364 25594
rect 2376 25542 2428 25594
rect 2440 25542 2492 25594
rect 2504 25542 2556 25594
rect 4846 25542 4898 25594
rect 4910 25542 4962 25594
rect 4974 25542 5026 25594
rect 5038 25542 5090 25594
rect 5102 25542 5154 25594
rect 7443 25542 7495 25594
rect 7507 25542 7559 25594
rect 7571 25542 7623 25594
rect 7635 25542 7687 25594
rect 7699 25542 7751 25594
rect 2044 25483 2096 25492
rect 2044 25449 2053 25483
rect 2053 25449 2087 25483
rect 2087 25449 2096 25483
rect 2044 25440 2096 25449
rect 5264 25415 5316 25424
rect 5264 25381 5273 25415
rect 5273 25381 5307 25415
rect 5307 25381 5316 25415
rect 5264 25372 5316 25381
rect 6828 25415 6880 25424
rect 6828 25381 6837 25415
rect 6837 25381 6871 25415
rect 6871 25381 6880 25415
rect 6828 25372 6880 25381
rect 5172 25347 5224 25356
rect 5172 25313 5181 25347
rect 5181 25313 5215 25347
rect 5215 25313 5224 25347
rect 5172 25304 5224 25313
rect 5724 25347 5776 25356
rect 5724 25313 5733 25347
rect 5733 25313 5767 25347
rect 5767 25313 5776 25347
rect 5724 25304 5776 25313
rect 4528 25236 4580 25288
rect 6000 25236 6052 25288
rect 7196 25279 7248 25288
rect 7196 25245 7205 25279
rect 7205 25245 7239 25279
rect 7239 25245 7248 25279
rect 7196 25236 7248 25245
rect 4252 25211 4304 25220
rect 4252 25177 4261 25211
rect 4261 25177 4295 25211
rect 4295 25177 4304 25211
rect 4252 25168 4304 25177
rect 8208 25236 8260 25288
rect 3547 24998 3599 25050
rect 3611 24998 3663 25050
rect 3675 24998 3727 25050
rect 3739 24998 3791 25050
rect 3803 24998 3855 25050
rect 6144 24998 6196 25050
rect 6208 24998 6260 25050
rect 6272 24998 6324 25050
rect 6336 24998 6388 25050
rect 6400 24998 6452 25050
rect 6552 24896 6604 24948
rect 3424 24803 3476 24812
rect 3424 24769 3433 24803
rect 3433 24769 3467 24803
rect 3467 24769 3476 24803
rect 6000 24828 6052 24880
rect 6092 24828 6144 24880
rect 3424 24760 3476 24769
rect 5724 24760 5776 24812
rect 6552 24803 6604 24812
rect 6552 24769 6561 24803
rect 6561 24769 6595 24803
rect 6595 24769 6604 24803
rect 6552 24760 6604 24769
rect 6736 24760 6788 24812
rect 7840 24760 7892 24812
rect 3884 24624 3936 24676
rect 4252 24624 4304 24676
rect 7288 24624 7340 24676
rect 2964 24599 3016 24608
rect 2964 24565 2973 24599
rect 2973 24565 3007 24599
rect 3007 24565 3016 24599
rect 2964 24556 3016 24565
rect 2248 24454 2300 24506
rect 2312 24454 2364 24506
rect 2376 24454 2428 24506
rect 2440 24454 2492 24506
rect 2504 24454 2556 24506
rect 4846 24454 4898 24506
rect 4910 24454 4962 24506
rect 4974 24454 5026 24506
rect 5038 24454 5090 24506
rect 5102 24454 5154 24506
rect 7443 24454 7495 24506
rect 7507 24454 7559 24506
rect 7571 24454 7623 24506
rect 7635 24454 7687 24506
rect 7699 24454 7751 24506
rect 6552 24284 6604 24336
rect 6920 24284 6972 24336
rect 7380 24284 7432 24336
rect 4160 24216 4212 24268
rect 5356 24216 5408 24268
rect 8116 24259 8168 24268
rect 8116 24225 8125 24259
rect 8125 24225 8159 24259
rect 8159 24225 8168 24259
rect 8116 24216 8168 24225
rect 5632 24191 5684 24200
rect 2964 24080 3016 24132
rect 2136 24055 2188 24064
rect 2136 24021 2145 24055
rect 2145 24021 2179 24055
rect 2179 24021 2188 24055
rect 2136 24012 2188 24021
rect 3240 24055 3292 24064
rect 3240 24021 3249 24055
rect 3249 24021 3283 24055
rect 3283 24021 3292 24055
rect 3240 24012 3292 24021
rect 3976 24055 4028 24064
rect 3976 24021 3985 24055
rect 3985 24021 4019 24055
rect 4019 24021 4028 24055
rect 3976 24012 4028 24021
rect 4160 24080 4212 24132
rect 5632 24157 5641 24191
rect 5641 24157 5675 24191
rect 5675 24157 5684 24191
rect 5632 24148 5684 24157
rect 6644 24148 6696 24200
rect 6736 24080 6788 24132
rect 7564 24123 7616 24132
rect 7564 24089 7573 24123
rect 7573 24089 7607 24123
rect 7607 24089 7616 24123
rect 7564 24080 7616 24089
rect 3547 23910 3599 23962
rect 3611 23910 3663 23962
rect 3675 23910 3727 23962
rect 3739 23910 3791 23962
rect 3803 23910 3855 23962
rect 6144 23910 6196 23962
rect 6208 23910 6260 23962
rect 6272 23910 6324 23962
rect 6336 23910 6388 23962
rect 6400 23910 6452 23962
rect 3976 23808 4028 23860
rect 4160 23851 4212 23860
rect 4160 23817 4169 23851
rect 4169 23817 4203 23851
rect 4203 23817 4212 23851
rect 4160 23808 4212 23817
rect 7564 23808 7616 23860
rect 5356 23783 5408 23792
rect 5356 23749 5365 23783
rect 5365 23749 5399 23783
rect 5399 23749 5408 23783
rect 5356 23740 5408 23749
rect 7196 23783 7248 23792
rect 7196 23749 7205 23783
rect 7205 23749 7239 23783
rect 7239 23749 7248 23783
rect 7196 23740 7248 23749
rect 7380 23783 7432 23792
rect 7380 23749 7389 23783
rect 7389 23749 7423 23783
rect 7423 23749 7432 23783
rect 7380 23740 7432 23749
rect 6644 23715 6696 23724
rect 6644 23681 6653 23715
rect 6653 23681 6687 23715
rect 6687 23681 6696 23715
rect 6644 23672 6696 23681
rect 8116 23715 8168 23724
rect 8116 23681 8125 23715
rect 8125 23681 8159 23715
rect 8159 23681 8168 23715
rect 8116 23672 8168 23681
rect 5632 23604 5684 23656
rect 5816 23647 5868 23656
rect 5816 23613 5825 23647
rect 5825 23613 5859 23647
rect 5859 23613 5868 23647
rect 5816 23604 5868 23613
rect 6552 23604 6604 23656
rect 2136 23536 2188 23588
rect 3240 23536 3292 23588
rect 5816 23468 5868 23520
rect 2248 23366 2300 23418
rect 2312 23366 2364 23418
rect 2376 23366 2428 23418
rect 2440 23366 2492 23418
rect 2504 23366 2556 23418
rect 4846 23366 4898 23418
rect 4910 23366 4962 23418
rect 4974 23366 5026 23418
rect 5038 23366 5090 23418
rect 5102 23366 5154 23418
rect 7443 23366 7495 23418
rect 7507 23366 7559 23418
rect 7571 23366 7623 23418
rect 7635 23366 7687 23418
rect 7699 23366 7751 23418
rect 3056 23264 3108 23316
rect 6644 23196 6696 23248
rect 2596 23060 2648 23112
rect 5908 23060 5960 23112
rect 6736 23060 6788 23112
rect 8116 23060 8168 23112
rect 4620 22992 4672 23044
rect 5172 22992 5224 23044
rect 5264 22992 5316 23044
rect 3240 22967 3292 22976
rect 3240 22933 3249 22967
rect 3249 22933 3283 22967
rect 3283 22933 3292 22967
rect 3240 22924 3292 22933
rect 7012 22992 7064 23044
rect 3547 22822 3599 22874
rect 3611 22822 3663 22874
rect 3675 22822 3727 22874
rect 3739 22822 3791 22874
rect 3803 22822 3855 22874
rect 6144 22822 6196 22874
rect 6208 22822 6260 22874
rect 6272 22822 6324 22874
rect 6336 22822 6388 22874
rect 6400 22822 6452 22874
rect 3056 22763 3108 22772
rect 3056 22729 3065 22763
rect 3065 22729 3099 22763
rect 3099 22729 3108 22763
rect 3056 22720 3108 22729
rect 5264 22720 5316 22772
rect 4252 22695 4304 22704
rect 4252 22661 4261 22695
rect 4261 22661 4295 22695
rect 4295 22661 4304 22695
rect 4252 22652 4304 22661
rect 6920 22584 6972 22636
rect 7288 22584 7340 22636
rect 8116 22627 8168 22636
rect 8116 22593 8125 22627
rect 8125 22593 8159 22627
rect 8159 22593 8168 22627
rect 8116 22584 8168 22593
rect 4160 22516 4212 22568
rect 4528 22448 4580 22500
rect 4712 22448 4764 22500
rect 2688 22380 2740 22432
rect 4068 22380 4120 22432
rect 6000 22516 6052 22568
rect 6644 22491 6696 22500
rect 6644 22457 6653 22491
rect 6653 22457 6687 22491
rect 6687 22457 6696 22491
rect 6644 22448 6696 22457
rect 2248 22278 2300 22330
rect 2312 22278 2364 22330
rect 2376 22278 2428 22330
rect 2440 22278 2492 22330
rect 2504 22278 2556 22330
rect 4846 22278 4898 22330
rect 4910 22278 4962 22330
rect 4974 22278 5026 22330
rect 5038 22278 5090 22330
rect 5102 22278 5154 22330
rect 7443 22278 7495 22330
rect 7507 22278 7559 22330
rect 7571 22278 7623 22330
rect 7635 22278 7687 22330
rect 7699 22278 7751 22330
rect 3240 22219 3292 22228
rect 3240 22185 3249 22219
rect 3249 22185 3283 22219
rect 3283 22185 3292 22219
rect 3240 22176 3292 22185
rect 6736 22176 6788 22228
rect 2688 22151 2740 22160
rect 2688 22117 2697 22151
rect 2697 22117 2731 22151
rect 2731 22117 2740 22151
rect 2688 22108 2740 22117
rect 4068 22108 4120 22160
rect 4252 22108 4304 22160
rect 4712 22151 4764 22160
rect 4712 22117 4721 22151
rect 4721 22117 4755 22151
rect 4755 22117 4764 22151
rect 4712 22108 4764 22117
rect 4160 22040 4212 22092
rect 6644 22040 6696 22092
rect 4528 21972 4580 22024
rect 4896 22015 4948 22024
rect 4896 21981 4905 22015
rect 4905 21981 4939 22015
rect 4939 21981 4948 22015
rect 4896 21972 4948 21981
rect 6000 22015 6052 22024
rect 6000 21981 6009 22015
rect 6009 21981 6043 22015
rect 6043 21981 6052 22015
rect 6000 21972 6052 21981
rect 7012 22015 7064 22024
rect 7012 21981 7021 22015
rect 7021 21981 7055 22015
rect 7055 21981 7064 22015
rect 7012 21972 7064 21981
rect 6920 21904 6972 21956
rect 5080 21836 5132 21888
rect 3547 21734 3599 21786
rect 3611 21734 3663 21786
rect 3675 21734 3727 21786
rect 3739 21734 3791 21786
rect 3803 21734 3855 21786
rect 6144 21734 6196 21786
rect 6208 21734 6260 21786
rect 6272 21734 6324 21786
rect 6336 21734 6388 21786
rect 6400 21734 6452 21786
rect 2596 21675 2648 21684
rect 2596 21641 2605 21675
rect 2605 21641 2639 21675
rect 2639 21641 2648 21675
rect 2596 21632 2648 21641
rect 4620 21632 4672 21684
rect 4896 21607 4948 21616
rect 4896 21573 4905 21607
rect 4905 21573 4939 21607
rect 4939 21573 4948 21607
rect 4896 21564 4948 21573
rect 5080 21607 5132 21616
rect 5080 21573 5089 21607
rect 5089 21573 5123 21607
rect 5123 21573 5132 21607
rect 5080 21564 5132 21573
rect 5908 21496 5960 21548
rect 6552 21496 6604 21548
rect 4344 21428 4396 21480
rect 6644 21403 6696 21412
rect 3148 21335 3200 21344
rect 3148 21301 3157 21335
rect 3157 21301 3191 21335
rect 3191 21301 3200 21335
rect 3148 21292 3200 21301
rect 3240 21292 3292 21344
rect 5816 21292 5868 21344
rect 6644 21369 6653 21403
rect 6653 21369 6687 21403
rect 6687 21369 6696 21403
rect 6644 21360 6696 21369
rect 7288 21360 7340 21412
rect 8116 21292 8168 21344
rect 2248 21190 2300 21242
rect 2312 21190 2364 21242
rect 2376 21190 2428 21242
rect 2440 21190 2492 21242
rect 2504 21190 2556 21242
rect 4846 21190 4898 21242
rect 4910 21190 4962 21242
rect 4974 21190 5026 21242
rect 5038 21190 5090 21242
rect 5102 21190 5154 21242
rect 7443 21190 7495 21242
rect 7507 21190 7559 21242
rect 7571 21190 7623 21242
rect 7635 21190 7687 21242
rect 7699 21190 7751 21242
rect 3240 21131 3292 21140
rect 3240 21097 3249 21131
rect 3249 21097 3283 21131
rect 3283 21097 3292 21131
rect 3240 21088 3292 21097
rect 2596 21020 2648 21072
rect 6736 21088 6788 21140
rect 7840 21063 7892 21072
rect 7840 21029 7849 21063
rect 7849 21029 7883 21063
rect 7883 21029 7892 21063
rect 7840 21020 7892 21029
rect 5816 20952 5868 21004
rect 4160 20927 4212 20936
rect 4160 20893 4169 20927
rect 4169 20893 4203 20927
rect 4203 20893 4212 20927
rect 4160 20884 4212 20893
rect 5632 20859 5684 20868
rect 5632 20825 5641 20859
rect 5641 20825 5675 20859
rect 5675 20825 5684 20859
rect 5632 20816 5684 20825
rect 6736 20884 6788 20936
rect 6828 20884 6880 20936
rect 7012 20816 7064 20868
rect 2596 20791 2648 20800
rect 2596 20757 2605 20791
rect 2605 20757 2639 20791
rect 2639 20757 2648 20791
rect 2596 20748 2648 20757
rect 4068 20748 4120 20800
rect 6828 20748 6880 20800
rect 3547 20646 3599 20698
rect 3611 20646 3663 20698
rect 3675 20646 3727 20698
rect 3739 20646 3791 20698
rect 3803 20646 3855 20698
rect 6144 20646 6196 20698
rect 6208 20646 6260 20698
rect 6272 20646 6324 20698
rect 6336 20646 6388 20698
rect 6400 20646 6452 20698
rect 4344 20544 4396 20596
rect 4068 20476 4120 20528
rect 5632 20476 5684 20528
rect 4160 20408 4212 20460
rect 5816 20451 5868 20460
rect 5816 20417 5825 20451
rect 5825 20417 5859 20451
rect 5859 20417 5868 20451
rect 5816 20408 5868 20417
rect 6644 20451 6696 20460
rect 6644 20417 6653 20451
rect 6653 20417 6687 20451
rect 6687 20417 6696 20451
rect 6644 20408 6696 20417
rect 7196 20408 7248 20460
rect 6460 20315 6512 20324
rect 2688 20204 2740 20256
rect 4252 20204 4304 20256
rect 6000 20204 6052 20256
rect 6460 20281 6469 20315
rect 6469 20281 6503 20315
rect 6503 20281 6512 20315
rect 6460 20272 6512 20281
rect 7288 20204 7340 20256
rect 2248 20102 2300 20154
rect 2312 20102 2364 20154
rect 2376 20102 2428 20154
rect 2440 20102 2492 20154
rect 2504 20102 2556 20154
rect 4846 20102 4898 20154
rect 4910 20102 4962 20154
rect 4974 20102 5026 20154
rect 5038 20102 5090 20154
rect 5102 20102 5154 20154
rect 7443 20102 7495 20154
rect 7507 20102 7559 20154
rect 7571 20102 7623 20154
rect 7635 20102 7687 20154
rect 7699 20102 7751 20154
rect 3148 20000 3200 20052
rect 4344 20000 4396 20052
rect 4068 19864 4120 19916
rect 2964 19796 3016 19848
rect 5540 19796 5592 19848
rect 6552 19864 6604 19916
rect 6828 19796 6880 19848
rect 7288 19796 7340 19848
rect 8116 19839 8168 19848
rect 8116 19805 8125 19839
rect 8125 19805 8159 19839
rect 8159 19805 8168 19839
rect 8116 19796 8168 19805
rect 6460 19728 6512 19780
rect 6644 19728 6696 19780
rect 1584 19703 1636 19712
rect 1584 19669 1593 19703
rect 1593 19669 1627 19703
rect 1627 19669 1636 19703
rect 1584 19660 1636 19669
rect 2044 19703 2096 19712
rect 2044 19669 2053 19703
rect 2053 19669 2087 19703
rect 2087 19669 2096 19703
rect 2044 19660 2096 19669
rect 3547 19558 3599 19610
rect 3611 19558 3663 19610
rect 3675 19558 3727 19610
rect 3739 19558 3791 19610
rect 3803 19558 3855 19610
rect 6144 19558 6196 19610
rect 6208 19558 6260 19610
rect 6272 19558 6324 19610
rect 6336 19558 6388 19610
rect 6400 19558 6452 19610
rect 2964 19499 3016 19508
rect 2964 19465 2973 19499
rect 2973 19465 3007 19499
rect 3007 19465 3016 19499
rect 2964 19456 3016 19465
rect 4068 19499 4120 19508
rect 4068 19465 4077 19499
rect 4077 19465 4111 19499
rect 4111 19465 4120 19499
rect 4068 19456 4120 19465
rect 4252 19456 4304 19508
rect 6552 19388 6604 19440
rect 4436 19320 4488 19372
rect 2596 19252 2648 19304
rect 4712 19295 4764 19304
rect 4712 19261 4721 19295
rect 4721 19261 4755 19295
rect 4755 19261 4764 19295
rect 4712 19252 4764 19261
rect 1584 19184 1636 19236
rect 3240 19184 3292 19236
rect 5540 19320 5592 19372
rect 5632 19252 5684 19304
rect 6736 19320 6788 19372
rect 5724 19184 5776 19236
rect 7840 19252 7892 19304
rect 5540 19116 5592 19168
rect 5816 19159 5868 19168
rect 5816 19125 5825 19159
rect 5825 19125 5859 19159
rect 5859 19125 5868 19159
rect 5816 19116 5868 19125
rect 6828 19116 6880 19168
rect 2248 19014 2300 19066
rect 2312 19014 2364 19066
rect 2376 19014 2428 19066
rect 2440 19014 2492 19066
rect 2504 19014 2556 19066
rect 4846 19014 4898 19066
rect 4910 19014 4962 19066
rect 4974 19014 5026 19066
rect 5038 19014 5090 19066
rect 5102 19014 5154 19066
rect 7443 19014 7495 19066
rect 7507 19014 7559 19066
rect 7571 19014 7623 19066
rect 7635 19014 7687 19066
rect 7699 19014 7751 19066
rect 2688 18955 2740 18964
rect 2688 18921 2697 18955
rect 2697 18921 2731 18955
rect 2731 18921 2740 18955
rect 2688 18912 2740 18921
rect 7196 18912 7248 18964
rect 3240 18887 3292 18896
rect 3240 18853 3249 18887
rect 3249 18853 3283 18887
rect 3283 18853 3292 18887
rect 3240 18844 3292 18853
rect 4436 18887 4488 18896
rect 4436 18853 4445 18887
rect 4445 18853 4479 18887
rect 4479 18853 4488 18887
rect 4436 18844 4488 18853
rect 6644 18844 6696 18896
rect 6000 18776 6052 18828
rect 8024 18776 8076 18828
rect 4436 18751 4488 18760
rect 4436 18717 4445 18751
rect 4445 18717 4479 18751
rect 4479 18717 4488 18751
rect 4436 18708 4488 18717
rect 5724 18751 5776 18760
rect 5724 18717 5733 18751
rect 5733 18717 5767 18751
rect 5767 18717 5776 18751
rect 5724 18708 5776 18717
rect 6552 18708 6604 18760
rect 7196 18708 7248 18760
rect 7288 18708 7340 18760
rect 2044 18640 2096 18692
rect 2780 18640 2832 18692
rect 7104 18640 7156 18692
rect 2136 18615 2188 18624
rect 2136 18581 2145 18615
rect 2145 18581 2179 18615
rect 2179 18581 2188 18615
rect 2136 18572 2188 18581
rect 3547 18470 3599 18522
rect 3611 18470 3663 18522
rect 3675 18470 3727 18522
rect 3739 18470 3791 18522
rect 3803 18470 3855 18522
rect 6144 18470 6196 18522
rect 6208 18470 6260 18522
rect 6272 18470 6324 18522
rect 6336 18470 6388 18522
rect 6400 18470 6452 18522
rect 4712 18368 4764 18420
rect 4620 18300 4672 18352
rect 4436 18232 4488 18284
rect 5816 18368 5868 18420
rect 5172 18300 5224 18352
rect 5724 18232 5776 18284
rect 6920 18275 6972 18284
rect 6920 18241 6929 18275
rect 6929 18241 6963 18275
rect 6963 18241 6972 18275
rect 6920 18232 6972 18241
rect 7840 18232 7892 18284
rect 8208 18232 8260 18284
rect 5540 18164 5592 18216
rect 7012 18164 7064 18216
rect 5356 18096 5408 18148
rect 1676 18028 1728 18080
rect 2044 18071 2096 18080
rect 2044 18037 2053 18071
rect 2053 18037 2087 18071
rect 2087 18037 2096 18071
rect 2044 18028 2096 18037
rect 2596 18071 2648 18080
rect 2596 18037 2605 18071
rect 2605 18037 2639 18071
rect 2639 18037 2648 18071
rect 2596 18028 2648 18037
rect 5632 18028 5684 18080
rect 5908 18028 5960 18080
rect 2248 17926 2300 17978
rect 2312 17926 2364 17978
rect 2376 17926 2428 17978
rect 2440 17926 2492 17978
rect 2504 17926 2556 17978
rect 4846 17926 4898 17978
rect 4910 17926 4962 17978
rect 4974 17926 5026 17978
rect 5038 17926 5090 17978
rect 5102 17926 5154 17978
rect 7443 17926 7495 17978
rect 7507 17926 7559 17978
rect 7571 17926 7623 17978
rect 7635 17926 7687 17978
rect 7699 17926 7751 17978
rect 2596 17867 2648 17876
rect 2596 17833 2605 17867
rect 2605 17833 2639 17867
rect 2639 17833 2648 17867
rect 2596 17824 2648 17833
rect 3976 17824 4028 17876
rect 5816 17824 5868 17876
rect 2044 17756 2096 17808
rect 2596 17688 2648 17740
rect 4528 17688 4580 17740
rect 4620 17731 4672 17740
rect 4620 17697 4629 17731
rect 4629 17697 4663 17731
rect 4663 17697 4672 17731
rect 4620 17688 4672 17697
rect 4804 17688 4856 17740
rect 7012 17756 7064 17808
rect 3976 17620 4028 17672
rect 5356 17663 5408 17672
rect 1676 17552 1728 17604
rect 4436 17552 4488 17604
rect 5356 17629 5365 17663
rect 5365 17629 5399 17663
rect 5399 17629 5408 17663
rect 5356 17620 5408 17629
rect 6920 17620 6972 17672
rect 7196 17663 7248 17672
rect 7196 17629 7205 17663
rect 7205 17629 7239 17663
rect 7239 17629 7248 17663
rect 7196 17620 7248 17629
rect 8208 17620 8260 17672
rect 5080 17552 5132 17604
rect 5264 17552 5316 17604
rect 7932 17552 7984 17604
rect 1584 17527 1636 17536
rect 1584 17493 1593 17527
rect 1593 17493 1627 17527
rect 1627 17493 1636 17527
rect 1584 17484 1636 17493
rect 4804 17484 4856 17536
rect 3547 17382 3599 17434
rect 3611 17382 3663 17434
rect 3675 17382 3727 17434
rect 3739 17382 3791 17434
rect 3803 17382 3855 17434
rect 6144 17382 6196 17434
rect 6208 17382 6260 17434
rect 6272 17382 6324 17434
rect 6336 17382 6388 17434
rect 6400 17382 6452 17434
rect 1676 17323 1728 17332
rect 1676 17289 1685 17323
rect 1685 17289 1719 17323
rect 1719 17289 1728 17323
rect 1676 17280 1728 17289
rect 4804 17323 4856 17332
rect 4804 17289 4813 17323
rect 4813 17289 4847 17323
rect 4847 17289 4856 17323
rect 4804 17280 4856 17289
rect 2872 17187 2924 17196
rect 2872 17153 2881 17187
rect 2881 17153 2915 17187
rect 2915 17153 2924 17187
rect 2872 17144 2924 17153
rect 4344 17212 4396 17264
rect 4436 17212 4488 17264
rect 4068 17144 4120 17196
rect 5632 17144 5684 17196
rect 6368 17187 6420 17196
rect 6368 17153 6377 17187
rect 6377 17153 6411 17187
rect 6411 17153 6420 17187
rect 6368 17144 6420 17153
rect 6736 17144 6788 17196
rect 7840 17144 7892 17196
rect 5172 17076 5224 17128
rect 2596 17008 2648 17060
rect 5356 17076 5408 17128
rect 7196 17008 7248 17060
rect 5540 16940 5592 16992
rect 2248 16838 2300 16890
rect 2312 16838 2364 16890
rect 2376 16838 2428 16890
rect 2440 16838 2492 16890
rect 2504 16838 2556 16890
rect 4846 16838 4898 16890
rect 4910 16838 4962 16890
rect 4974 16838 5026 16890
rect 5038 16838 5090 16890
rect 5102 16838 5154 16890
rect 7443 16838 7495 16890
rect 7507 16838 7559 16890
rect 7571 16838 7623 16890
rect 7635 16838 7687 16890
rect 7699 16838 7751 16890
rect 2596 16779 2648 16788
rect 2596 16745 2605 16779
rect 2605 16745 2639 16779
rect 2639 16745 2648 16779
rect 2596 16736 2648 16745
rect 2872 16736 2924 16788
rect 7288 16736 7340 16788
rect 1584 16668 1636 16720
rect 6736 16668 6788 16720
rect 4068 16600 4120 16652
rect 3976 16532 4028 16584
rect 4344 16600 4396 16652
rect 4436 16575 4488 16584
rect 4436 16541 4445 16575
rect 4445 16541 4479 16575
rect 4479 16541 4488 16575
rect 4436 16532 4488 16541
rect 4528 16532 4580 16584
rect 5724 16532 5776 16584
rect 6000 16532 6052 16584
rect 6368 16532 6420 16584
rect 3884 16464 3936 16516
rect 5540 16464 5592 16516
rect 5908 16464 5960 16516
rect 7840 16464 7892 16516
rect 2596 16396 2648 16448
rect 7104 16396 7156 16448
rect 3547 16294 3599 16346
rect 3611 16294 3663 16346
rect 3675 16294 3727 16346
rect 3739 16294 3791 16346
rect 3803 16294 3855 16346
rect 6144 16294 6196 16346
rect 6208 16294 6260 16346
rect 6272 16294 6324 16346
rect 6336 16294 6388 16346
rect 6400 16294 6452 16346
rect 2596 16235 2648 16244
rect 2596 16201 2605 16235
rect 2605 16201 2639 16235
rect 2639 16201 2648 16235
rect 2596 16192 2648 16201
rect 3884 16235 3936 16244
rect 3516 16124 3568 16176
rect 3884 16201 3893 16235
rect 3893 16201 3927 16235
rect 3927 16201 3936 16235
rect 3884 16192 3936 16201
rect 3976 16192 4028 16244
rect 4712 16124 4764 16176
rect 5632 16124 5684 16176
rect 7196 16167 7248 16176
rect 7196 16133 7205 16167
rect 7205 16133 7239 16167
rect 7239 16133 7248 16167
rect 7196 16124 7248 16133
rect 7288 16124 7340 16176
rect 4528 16099 4580 16108
rect 4528 16065 4537 16099
rect 4537 16065 4571 16099
rect 4571 16065 4580 16099
rect 4528 16056 4580 16065
rect 4620 16056 4672 16108
rect 7012 16056 7064 16108
rect 8024 16056 8076 16108
rect 2688 15920 2740 15972
rect 5540 16031 5592 16040
rect 5540 15997 5549 16031
rect 5549 15997 5583 16031
rect 5583 15997 5592 16031
rect 5540 15988 5592 15997
rect 1952 15852 2004 15904
rect 2136 15895 2188 15904
rect 2136 15861 2145 15895
rect 2145 15861 2179 15895
rect 2179 15861 2188 15895
rect 2136 15852 2188 15861
rect 3148 15852 3200 15904
rect 3516 15852 3568 15904
rect 6000 15852 6052 15904
rect 2248 15750 2300 15802
rect 2312 15750 2364 15802
rect 2376 15750 2428 15802
rect 2440 15750 2492 15802
rect 2504 15750 2556 15802
rect 4846 15750 4898 15802
rect 4910 15750 4962 15802
rect 4974 15750 5026 15802
rect 5038 15750 5090 15802
rect 5102 15750 5154 15802
rect 7443 15750 7495 15802
rect 7507 15750 7559 15802
rect 7571 15750 7623 15802
rect 7635 15750 7687 15802
rect 7699 15750 7751 15802
rect 2688 15691 2740 15700
rect 2688 15657 2697 15691
rect 2697 15657 2731 15691
rect 2731 15657 2740 15691
rect 2688 15648 2740 15657
rect 5724 15648 5776 15700
rect 6000 15648 6052 15700
rect 3148 15580 3200 15632
rect 7012 15580 7064 15632
rect 7840 15580 7892 15632
rect 4068 15512 4120 15564
rect 4712 15487 4764 15496
rect 4712 15453 4721 15487
rect 4721 15453 4755 15487
rect 4755 15453 4764 15487
rect 4712 15444 4764 15453
rect 5540 15444 5592 15496
rect 6644 15444 6696 15496
rect 4620 15376 4672 15428
rect 5632 15376 5684 15428
rect 6552 15376 6604 15428
rect 1860 15308 1912 15360
rect 1952 15308 2004 15360
rect 2872 15308 2924 15360
rect 3056 15308 3108 15360
rect 8116 15376 8168 15428
rect 3547 15206 3599 15258
rect 3611 15206 3663 15258
rect 3675 15206 3727 15258
rect 3739 15206 3791 15258
rect 3803 15206 3855 15258
rect 6144 15206 6196 15258
rect 6208 15206 6260 15258
rect 6272 15206 6324 15258
rect 6336 15206 6388 15258
rect 6400 15206 6452 15258
rect 3056 15147 3108 15156
rect 3056 15113 3065 15147
rect 3065 15113 3099 15147
rect 3099 15113 3108 15147
rect 3056 15104 3108 15113
rect 6736 15104 6788 15156
rect 4528 15036 4580 15088
rect 4712 15011 4764 15020
rect 4712 14977 4721 15011
rect 4721 14977 4755 15011
rect 4755 14977 4764 15011
rect 4712 14968 4764 14977
rect 5724 14968 5776 15020
rect 6092 14968 6144 15020
rect 8116 14968 8168 15020
rect 5540 14900 5592 14952
rect 6552 14900 6604 14952
rect 6828 14900 6880 14952
rect 6092 14832 6144 14884
rect 1860 14807 1912 14816
rect 1860 14773 1869 14807
rect 1869 14773 1903 14807
rect 1903 14773 1912 14807
rect 1860 14764 1912 14773
rect 2596 14764 2648 14816
rect 3608 14807 3660 14816
rect 3608 14773 3617 14807
rect 3617 14773 3651 14807
rect 3651 14773 3660 14807
rect 3608 14764 3660 14773
rect 4252 14807 4304 14816
rect 4252 14773 4261 14807
rect 4261 14773 4295 14807
rect 4295 14773 4304 14807
rect 4252 14764 4304 14773
rect 4344 14764 4396 14816
rect 8208 14764 8260 14816
rect 2248 14662 2300 14714
rect 2312 14662 2364 14714
rect 2376 14662 2428 14714
rect 2440 14662 2492 14714
rect 2504 14662 2556 14714
rect 4846 14662 4898 14714
rect 4910 14662 4962 14714
rect 4974 14662 5026 14714
rect 5038 14662 5090 14714
rect 5102 14662 5154 14714
rect 7443 14662 7495 14714
rect 7507 14662 7559 14714
rect 7571 14662 7623 14714
rect 7635 14662 7687 14714
rect 7699 14662 7751 14714
rect 3608 14492 3660 14544
rect 5724 14492 5776 14544
rect 4252 14424 4304 14476
rect 5172 14467 5224 14476
rect 5172 14433 5181 14467
rect 5181 14433 5215 14467
rect 5215 14433 5224 14467
rect 5172 14424 5224 14433
rect 3884 14399 3936 14408
rect 3884 14365 3893 14399
rect 3893 14365 3927 14399
rect 3927 14365 3936 14399
rect 3884 14356 3936 14365
rect 4344 14356 4396 14408
rect 5540 14356 5592 14408
rect 5724 14356 5776 14408
rect 6092 14399 6144 14408
rect 6092 14365 6101 14399
rect 6101 14365 6135 14399
rect 6135 14365 6144 14399
rect 6092 14356 6144 14365
rect 6828 14356 6880 14408
rect 8208 14356 8260 14408
rect 2596 14288 2648 14340
rect 4804 14288 4856 14340
rect 6920 14288 6972 14340
rect 7656 14331 7708 14340
rect 7656 14297 7665 14331
rect 7665 14297 7699 14331
rect 7699 14297 7708 14331
rect 7656 14288 7708 14297
rect 1584 14263 1636 14272
rect 1584 14229 1593 14263
rect 1593 14229 1627 14263
rect 1627 14229 1636 14263
rect 1584 14220 1636 14229
rect 2688 14263 2740 14272
rect 2688 14229 2697 14263
rect 2697 14229 2731 14263
rect 2731 14229 2740 14263
rect 2688 14220 2740 14229
rect 5448 14220 5500 14272
rect 5724 14220 5776 14272
rect 6828 14220 6880 14272
rect 3547 14118 3599 14170
rect 3611 14118 3663 14170
rect 3675 14118 3727 14170
rect 3739 14118 3791 14170
rect 3803 14118 3855 14170
rect 6144 14118 6196 14170
rect 6208 14118 6260 14170
rect 6272 14118 6324 14170
rect 6336 14118 6388 14170
rect 6400 14118 6452 14170
rect 3884 14016 3936 14068
rect 5172 14016 5224 14068
rect 5632 13948 5684 14000
rect 7656 13948 7708 14000
rect 1584 13880 1636 13932
rect 2964 13880 3016 13932
rect 4804 13923 4856 13932
rect 4804 13889 4813 13923
rect 4813 13889 4847 13923
rect 4847 13889 4856 13923
rect 4804 13880 4856 13889
rect 5356 13880 5408 13932
rect 7012 13923 7064 13932
rect 7012 13889 7021 13923
rect 7021 13889 7055 13923
rect 7055 13889 7064 13923
rect 7012 13880 7064 13889
rect 8208 13880 8260 13932
rect 5540 13855 5592 13864
rect 1584 13676 1636 13728
rect 2688 13676 2740 13728
rect 5540 13821 5549 13855
rect 5549 13821 5583 13855
rect 5583 13821 5592 13855
rect 5540 13812 5592 13821
rect 4712 13676 4764 13728
rect 2248 13574 2300 13626
rect 2312 13574 2364 13626
rect 2376 13574 2428 13626
rect 2440 13574 2492 13626
rect 2504 13574 2556 13626
rect 4846 13574 4898 13626
rect 4910 13574 4962 13626
rect 4974 13574 5026 13626
rect 5038 13574 5090 13626
rect 5102 13574 5154 13626
rect 7443 13574 7495 13626
rect 7507 13574 7559 13626
rect 7571 13574 7623 13626
rect 7635 13574 7687 13626
rect 7699 13574 7751 13626
rect 1768 13472 1820 13524
rect 5816 13472 5868 13524
rect 6092 13472 6144 13524
rect 8392 13472 8444 13524
rect 6000 13404 6052 13456
rect 7012 13336 7064 13388
rect 5448 13311 5500 13320
rect 2412 13200 2464 13252
rect 4528 13243 4580 13252
rect 4528 13209 4537 13243
rect 4537 13209 4571 13243
rect 4571 13209 4580 13243
rect 5448 13277 5457 13311
rect 5457 13277 5491 13311
rect 5491 13277 5500 13311
rect 5448 13268 5500 13277
rect 5816 13268 5868 13320
rect 7104 13268 7156 13320
rect 7932 13268 7984 13320
rect 8116 13311 8168 13320
rect 8116 13277 8125 13311
rect 8125 13277 8159 13311
rect 8159 13277 8168 13311
rect 8116 13268 8168 13277
rect 4528 13200 4580 13209
rect 7012 13200 7064 13252
rect 7380 13243 7432 13252
rect 7380 13209 7389 13243
rect 7389 13209 7423 13243
rect 7423 13209 7432 13243
rect 7380 13200 7432 13209
rect 1584 13175 1636 13184
rect 1584 13141 1593 13175
rect 1593 13141 1627 13175
rect 1627 13141 1636 13175
rect 1584 13132 1636 13141
rect 3056 13132 3108 13184
rect 7564 13132 7616 13184
rect 3547 13030 3599 13082
rect 3611 13030 3663 13082
rect 3675 13030 3727 13082
rect 3739 13030 3791 13082
rect 3803 13030 3855 13082
rect 6144 13030 6196 13082
rect 6208 13030 6260 13082
rect 6272 13030 6324 13082
rect 6336 13030 6388 13082
rect 6400 13030 6452 13082
rect 1768 12971 1820 12980
rect 1768 12937 1777 12971
rect 1777 12937 1811 12971
rect 1811 12937 1820 12971
rect 1768 12928 1820 12937
rect 2412 12971 2464 12980
rect 2412 12937 2421 12971
rect 2421 12937 2455 12971
rect 2455 12937 2464 12971
rect 2412 12928 2464 12937
rect 2872 12928 2924 12980
rect 5632 12928 5684 12980
rect 6920 12928 6972 12980
rect 4528 12860 4580 12912
rect 7380 12860 7432 12912
rect 3700 12835 3752 12844
rect 3700 12801 3709 12835
rect 3709 12801 3743 12835
rect 3743 12801 3752 12835
rect 3700 12792 3752 12801
rect 4252 12835 4304 12844
rect 4252 12801 4261 12835
rect 4261 12801 4295 12835
rect 4295 12801 4304 12835
rect 4252 12792 4304 12801
rect 7564 12835 7616 12844
rect 7564 12801 7573 12835
rect 7573 12801 7607 12835
rect 7607 12801 7616 12835
rect 7564 12792 7616 12801
rect 8116 12835 8168 12844
rect 8116 12801 8125 12835
rect 8125 12801 8159 12835
rect 8159 12801 8168 12835
rect 8116 12792 8168 12801
rect 5816 12724 5868 12776
rect 4344 12656 4396 12708
rect 4160 12588 4212 12640
rect 7012 12724 7064 12776
rect 7288 12656 7340 12708
rect 2248 12486 2300 12538
rect 2312 12486 2364 12538
rect 2376 12486 2428 12538
rect 2440 12486 2492 12538
rect 2504 12486 2556 12538
rect 4846 12486 4898 12538
rect 4910 12486 4962 12538
rect 4974 12486 5026 12538
rect 5038 12486 5090 12538
rect 5102 12486 5154 12538
rect 7443 12486 7495 12538
rect 7507 12486 7559 12538
rect 7571 12486 7623 12538
rect 7635 12486 7687 12538
rect 7699 12486 7751 12538
rect 4160 12384 4212 12436
rect 3700 12316 3752 12368
rect 4712 12359 4764 12368
rect 4712 12325 4721 12359
rect 4721 12325 4755 12359
rect 4755 12325 4764 12359
rect 4712 12316 4764 12325
rect 5448 12384 5500 12436
rect 5540 12316 5592 12368
rect 5356 12248 5408 12300
rect 5448 12180 5500 12232
rect 5816 12180 5868 12232
rect 6552 12223 6604 12232
rect 1952 12087 2004 12096
rect 1952 12053 1961 12087
rect 1961 12053 1995 12087
rect 1995 12053 2004 12087
rect 1952 12044 2004 12053
rect 5908 12112 5960 12164
rect 6552 12189 6561 12223
rect 6561 12189 6595 12223
rect 6595 12189 6604 12223
rect 6552 12180 6604 12189
rect 6736 12180 6788 12232
rect 6644 12112 6696 12164
rect 3884 12087 3936 12096
rect 3884 12053 3893 12087
rect 3893 12053 3927 12087
rect 3927 12053 3936 12087
rect 3884 12044 3936 12053
rect 7104 12044 7156 12096
rect 7288 12044 7340 12096
rect 3547 11942 3599 11994
rect 3611 11942 3663 11994
rect 3675 11942 3727 11994
rect 3739 11942 3791 11994
rect 3803 11942 3855 11994
rect 6144 11942 6196 11994
rect 6208 11942 6260 11994
rect 6272 11942 6324 11994
rect 6336 11942 6388 11994
rect 6400 11942 6452 11994
rect 3148 11840 3200 11892
rect 3976 11840 4028 11892
rect 5540 11772 5592 11824
rect 4252 11747 4304 11756
rect 4252 11713 4261 11747
rect 4261 11713 4295 11747
rect 4295 11713 4304 11747
rect 4252 11704 4304 11713
rect 5264 11704 5316 11756
rect 6000 11840 6052 11892
rect 6552 11772 6604 11824
rect 7104 11815 7156 11824
rect 7104 11781 7113 11815
rect 7113 11781 7147 11815
rect 7147 11781 7156 11815
rect 7104 11772 7156 11781
rect 7012 11704 7064 11756
rect 7840 11747 7892 11756
rect 7840 11713 7849 11747
rect 7849 11713 7883 11747
rect 7883 11713 7892 11747
rect 7840 11704 7892 11713
rect 3240 11636 3292 11688
rect 6736 11636 6788 11688
rect 4160 11611 4212 11620
rect 4160 11577 4169 11611
rect 4169 11577 4203 11611
rect 4203 11577 4212 11611
rect 4160 11568 4212 11577
rect 1676 11543 1728 11552
rect 1676 11509 1685 11543
rect 1685 11509 1719 11543
rect 1719 11509 1728 11543
rect 1676 11500 1728 11509
rect 1860 11500 1912 11552
rect 5448 11500 5500 11552
rect 2248 11398 2300 11450
rect 2312 11398 2364 11450
rect 2376 11398 2428 11450
rect 2440 11398 2492 11450
rect 2504 11398 2556 11450
rect 4846 11398 4898 11450
rect 4910 11398 4962 11450
rect 4974 11398 5026 11450
rect 5038 11398 5090 11450
rect 5102 11398 5154 11450
rect 7443 11398 7495 11450
rect 7507 11398 7559 11450
rect 7571 11398 7623 11450
rect 7635 11398 7687 11450
rect 7699 11398 7751 11450
rect 3240 11339 3292 11348
rect 3240 11305 3249 11339
rect 3249 11305 3283 11339
rect 3283 11305 3292 11339
rect 3240 11296 3292 11305
rect 3884 11296 3936 11348
rect 7932 11339 7984 11348
rect 4160 11228 4212 11280
rect 5356 11228 5408 11280
rect 3976 11160 4028 11212
rect 4344 11203 4396 11212
rect 4344 11169 4353 11203
rect 4353 11169 4387 11203
rect 4387 11169 4396 11203
rect 4344 11160 4396 11169
rect 5448 11203 5500 11212
rect 5448 11169 5457 11203
rect 5457 11169 5491 11203
rect 5491 11169 5500 11203
rect 5448 11160 5500 11169
rect 7932 11305 7941 11339
rect 7941 11305 7975 11339
rect 7975 11305 7984 11339
rect 7932 11296 7984 11305
rect 1676 11092 1728 11144
rect 5264 11092 5316 11144
rect 1952 11024 2004 11076
rect 2136 10999 2188 11008
rect 2136 10965 2145 10999
rect 2145 10965 2179 10999
rect 2179 10965 2188 10999
rect 2136 10956 2188 10965
rect 4712 11024 4764 11076
rect 5816 11024 5868 11076
rect 6736 11092 6788 11144
rect 7380 11135 7432 11144
rect 7380 11101 7389 11135
rect 7389 11101 7423 11135
rect 7423 11101 7432 11135
rect 7380 11092 7432 11101
rect 7840 11024 7892 11076
rect 8208 10956 8260 11008
rect 8392 10956 8444 11008
rect 3547 10854 3599 10906
rect 3611 10854 3663 10906
rect 3675 10854 3727 10906
rect 3739 10854 3791 10906
rect 3803 10854 3855 10906
rect 6144 10854 6196 10906
rect 6208 10854 6260 10906
rect 6272 10854 6324 10906
rect 6336 10854 6388 10906
rect 6400 10854 6452 10906
rect 3056 10752 3108 10804
rect 4620 10795 4672 10804
rect 4620 10761 4629 10795
rect 4629 10761 4663 10795
rect 4663 10761 4672 10795
rect 4620 10752 4672 10761
rect 5540 10752 5592 10804
rect 6092 10684 6144 10736
rect 6920 10752 6972 10804
rect 4712 10659 4764 10668
rect 4712 10625 4721 10659
rect 4721 10625 4755 10659
rect 4755 10625 4764 10659
rect 4712 10616 4764 10625
rect 5908 10616 5960 10668
rect 7196 10616 7248 10668
rect 4344 10548 4396 10600
rect 5816 10591 5868 10600
rect 5816 10557 5825 10591
rect 5825 10557 5859 10591
rect 5859 10557 5868 10591
rect 5816 10548 5868 10557
rect 6552 10548 6604 10600
rect 8208 10548 8260 10600
rect 2044 10480 2096 10532
rect 1860 10412 1912 10464
rect 2780 10412 2832 10464
rect 4620 10480 4672 10532
rect 5448 10480 5500 10532
rect 7840 10480 7892 10532
rect 7288 10412 7340 10464
rect 2248 10310 2300 10362
rect 2312 10310 2364 10362
rect 2376 10310 2428 10362
rect 2440 10310 2492 10362
rect 2504 10310 2556 10362
rect 4846 10310 4898 10362
rect 4910 10310 4962 10362
rect 4974 10310 5026 10362
rect 5038 10310 5090 10362
rect 5102 10310 5154 10362
rect 7443 10310 7495 10362
rect 7507 10310 7559 10362
rect 7571 10310 7623 10362
rect 7635 10310 7687 10362
rect 7699 10310 7751 10362
rect 2780 10208 2832 10260
rect 4436 10208 4488 10260
rect 4712 10208 4764 10260
rect 6552 10140 6604 10192
rect 7288 10115 7340 10124
rect 2872 10004 2924 10056
rect 4160 10004 4212 10056
rect 7288 10081 7297 10115
rect 7297 10081 7331 10115
rect 7331 10081 7340 10115
rect 7288 10072 7340 10081
rect 6092 10047 6144 10056
rect 3056 9936 3108 9988
rect 4252 9979 4304 9988
rect 4252 9945 4261 9979
rect 4261 9945 4295 9979
rect 4295 9945 4304 9979
rect 4252 9936 4304 9945
rect 6092 10013 6101 10047
rect 6101 10013 6135 10047
rect 6135 10013 6144 10047
rect 6092 10004 6144 10013
rect 6644 10004 6696 10056
rect 6828 10047 6880 10056
rect 6828 10013 6837 10047
rect 6837 10013 6871 10047
rect 6871 10013 6880 10047
rect 6828 10004 6880 10013
rect 7932 10004 7984 10056
rect 5540 9936 5592 9988
rect 5908 9979 5960 9988
rect 5908 9945 5917 9979
rect 5917 9945 5951 9979
rect 5951 9945 5960 9979
rect 5908 9936 5960 9945
rect 7380 9979 7432 9988
rect 7380 9945 7389 9979
rect 7389 9945 7423 9979
rect 7423 9945 7432 9979
rect 7380 9936 7432 9945
rect 2136 9868 2188 9920
rect 2596 9868 2648 9920
rect 5448 9868 5500 9920
rect 3547 9766 3599 9818
rect 3611 9766 3663 9818
rect 3675 9766 3727 9818
rect 3739 9766 3791 9818
rect 3803 9766 3855 9818
rect 6144 9766 6196 9818
rect 6208 9766 6260 9818
rect 6272 9766 6324 9818
rect 6336 9766 6388 9818
rect 6400 9766 6452 9818
rect 4252 9664 4304 9716
rect 4436 9664 4488 9716
rect 6552 9664 6604 9716
rect 7380 9596 7432 9648
rect 1952 9367 2004 9376
rect 1952 9333 1961 9367
rect 1961 9333 1995 9367
rect 1995 9333 2004 9367
rect 1952 9324 2004 9333
rect 4344 9528 4396 9580
rect 4528 9528 4580 9580
rect 5540 9571 5592 9580
rect 5540 9537 5549 9571
rect 5549 9537 5583 9571
rect 5583 9537 5592 9571
rect 5540 9528 5592 9537
rect 5908 9528 5960 9580
rect 7932 9571 7984 9580
rect 7932 9537 7941 9571
rect 7941 9537 7975 9571
rect 7975 9537 7984 9571
rect 7932 9528 7984 9537
rect 4160 9460 4212 9512
rect 4620 9460 4672 9512
rect 5356 9503 5408 9512
rect 5356 9469 5365 9503
rect 5365 9469 5399 9503
rect 5399 9469 5408 9503
rect 5356 9460 5408 9469
rect 7196 9392 7248 9444
rect 3884 9367 3936 9376
rect 3884 9333 3893 9367
rect 3893 9333 3927 9367
rect 3927 9333 3936 9367
rect 3884 9324 3936 9333
rect 5816 9324 5868 9376
rect 8116 9324 8168 9376
rect 2248 9222 2300 9274
rect 2312 9222 2364 9274
rect 2376 9222 2428 9274
rect 2440 9222 2492 9274
rect 2504 9222 2556 9274
rect 4846 9222 4898 9274
rect 4910 9222 4962 9274
rect 4974 9222 5026 9274
rect 5038 9222 5090 9274
rect 5102 9222 5154 9274
rect 7443 9222 7495 9274
rect 7507 9222 7559 9274
rect 7571 9222 7623 9274
rect 7635 9222 7687 9274
rect 7699 9222 7751 9274
rect 2044 9163 2096 9172
rect 2044 9129 2053 9163
rect 2053 9129 2087 9163
rect 2087 9129 2096 9163
rect 2044 9120 2096 9129
rect 4160 9163 4212 9172
rect 4160 9129 4169 9163
rect 4169 9129 4203 9163
rect 4203 9129 4212 9163
rect 4160 9120 4212 9129
rect 6000 9052 6052 9104
rect 7840 9095 7892 9104
rect 7840 9061 7849 9095
rect 7849 9061 7883 9095
rect 7883 9061 7892 9095
rect 7840 9052 7892 9061
rect 6644 8984 6696 9036
rect 4528 8916 4580 8968
rect 5356 8916 5408 8968
rect 6828 8916 6880 8968
rect 7196 8916 7248 8968
rect 3148 8848 3200 8900
rect 5908 8848 5960 8900
rect 6184 8848 6236 8900
rect 8300 8848 8352 8900
rect 1492 8823 1544 8832
rect 1492 8789 1501 8823
rect 1501 8789 1535 8823
rect 1535 8789 1544 8823
rect 1492 8780 1544 8789
rect 2044 8780 2096 8832
rect 4252 8780 4304 8832
rect 3547 8678 3599 8730
rect 3611 8678 3663 8730
rect 3675 8678 3727 8730
rect 3739 8678 3791 8730
rect 3803 8678 3855 8730
rect 6144 8678 6196 8730
rect 6208 8678 6260 8730
rect 6272 8678 6324 8730
rect 6336 8678 6388 8730
rect 6400 8678 6452 8730
rect 1492 8619 1544 8628
rect 1492 8585 1501 8619
rect 1501 8585 1535 8619
rect 1535 8585 1544 8619
rect 3148 8619 3200 8628
rect 1492 8576 1544 8585
rect 3148 8585 3157 8619
rect 3157 8585 3191 8619
rect 3191 8585 3200 8619
rect 3148 8576 3200 8585
rect 5448 8576 5500 8628
rect 3884 8508 3936 8560
rect 4712 8508 4764 8560
rect 7196 8551 7248 8560
rect 7196 8517 7205 8551
rect 7205 8517 7239 8551
rect 7239 8517 7248 8551
rect 7196 8508 7248 8517
rect 3884 8372 3936 8424
rect 4160 8440 4212 8492
rect 5448 8440 5500 8492
rect 8116 8483 8168 8492
rect 8116 8449 8125 8483
rect 8125 8449 8159 8483
rect 8159 8449 8168 8483
rect 8116 8440 8168 8449
rect 4528 8415 4580 8424
rect 4528 8381 4537 8415
rect 4537 8381 4571 8415
rect 4571 8381 4580 8415
rect 4528 8372 4580 8381
rect 5724 8372 5776 8424
rect 5356 8347 5408 8356
rect 5356 8313 5365 8347
rect 5365 8313 5399 8347
rect 5399 8313 5408 8347
rect 5356 8304 5408 8313
rect 3976 8236 4028 8288
rect 6184 8236 6236 8288
rect 7288 8236 7340 8288
rect 2248 8134 2300 8186
rect 2312 8134 2364 8186
rect 2376 8134 2428 8186
rect 2440 8134 2492 8186
rect 2504 8134 2556 8186
rect 4846 8134 4898 8186
rect 4910 8134 4962 8186
rect 4974 8134 5026 8186
rect 5038 8134 5090 8186
rect 5102 8134 5154 8186
rect 7443 8134 7495 8186
rect 7507 8134 7559 8186
rect 7571 8134 7623 8186
rect 7635 8134 7687 8186
rect 7699 8134 7751 8186
rect 1860 8032 1912 8084
rect 2044 8032 2096 8084
rect 3424 7964 3476 8016
rect 4528 7964 4580 8016
rect 5172 7964 5224 8016
rect 5908 7964 5960 8016
rect 1492 7896 1544 7948
rect 2412 7871 2464 7880
rect 2412 7837 2421 7871
rect 2421 7837 2455 7871
rect 2455 7837 2464 7871
rect 2412 7828 2464 7837
rect 4528 7828 4580 7880
rect 4344 7803 4396 7812
rect 4344 7769 4353 7803
rect 4353 7769 4387 7803
rect 4387 7769 4396 7803
rect 4344 7760 4396 7769
rect 4436 7803 4488 7812
rect 4436 7769 4445 7803
rect 4445 7769 4479 7803
rect 4479 7769 4488 7803
rect 4436 7760 4488 7769
rect 2596 7735 2648 7744
rect 2596 7701 2605 7735
rect 2605 7701 2639 7735
rect 2639 7701 2648 7735
rect 2596 7692 2648 7701
rect 3240 7735 3292 7744
rect 3240 7701 3249 7735
rect 3249 7701 3283 7735
rect 3283 7701 3292 7735
rect 3240 7692 3292 7701
rect 3976 7692 4028 7744
rect 5264 7828 5316 7880
rect 6184 7871 6236 7880
rect 6184 7837 6193 7871
rect 6193 7837 6227 7871
rect 6227 7837 6236 7871
rect 6184 7828 6236 7837
rect 7012 7828 7064 7880
rect 7840 7828 7892 7880
rect 6736 7803 6788 7812
rect 6736 7769 6745 7803
rect 6745 7769 6779 7803
rect 6779 7769 6788 7803
rect 6736 7760 6788 7769
rect 6920 7803 6972 7812
rect 6920 7769 6929 7803
rect 6929 7769 6963 7803
rect 6963 7769 6972 7803
rect 6920 7760 6972 7769
rect 3547 7590 3599 7642
rect 3611 7590 3663 7642
rect 3675 7590 3727 7642
rect 3739 7590 3791 7642
rect 3803 7590 3855 7642
rect 6144 7590 6196 7642
rect 6208 7590 6260 7642
rect 6272 7590 6324 7642
rect 6336 7590 6388 7642
rect 6400 7590 6452 7642
rect 2596 7420 2648 7472
rect 6920 7488 6972 7540
rect 4068 7420 4120 7472
rect 4252 7463 4304 7472
rect 4252 7429 4261 7463
rect 4261 7429 4295 7463
rect 4295 7429 4304 7463
rect 4252 7420 4304 7429
rect 4436 7463 4488 7472
rect 4436 7429 4445 7463
rect 4445 7429 4479 7463
rect 4479 7429 4488 7463
rect 4436 7420 4488 7429
rect 4160 7352 4212 7404
rect 3792 7327 3844 7336
rect 3792 7293 3801 7327
rect 3801 7293 3835 7327
rect 3835 7293 3844 7327
rect 3792 7284 3844 7293
rect 3976 7284 4028 7336
rect 5356 7352 5408 7404
rect 6736 7395 6788 7404
rect 6736 7361 6745 7395
rect 6745 7361 6779 7395
rect 6779 7361 6788 7395
rect 6736 7352 6788 7361
rect 7288 7352 7340 7404
rect 7932 7395 7984 7404
rect 7932 7361 7941 7395
rect 7941 7361 7975 7395
rect 7975 7361 7984 7395
rect 7932 7352 7984 7361
rect 2412 7216 2464 7268
rect 2044 7148 2096 7200
rect 4252 7148 4304 7200
rect 5172 7148 5224 7200
rect 2248 7046 2300 7098
rect 2312 7046 2364 7098
rect 2376 7046 2428 7098
rect 2440 7046 2492 7098
rect 2504 7046 2556 7098
rect 4846 7046 4898 7098
rect 4910 7046 4962 7098
rect 4974 7046 5026 7098
rect 5038 7046 5090 7098
rect 5102 7046 5154 7098
rect 7443 7046 7495 7098
rect 7507 7046 7559 7098
rect 7571 7046 7623 7098
rect 7635 7046 7687 7098
rect 7699 7046 7751 7098
rect 1492 6987 1544 6996
rect 1492 6953 1501 6987
rect 1501 6953 1535 6987
rect 1535 6953 1544 6987
rect 1492 6944 1544 6953
rect 4436 6944 4488 6996
rect 4712 6944 4764 6996
rect 5448 6876 5500 6928
rect 3240 6851 3292 6860
rect 3240 6817 3249 6851
rect 3249 6817 3283 6851
rect 3283 6817 3292 6851
rect 3240 6808 3292 6817
rect 3332 6808 3384 6860
rect 2044 6783 2096 6792
rect 2044 6749 2053 6783
rect 2053 6749 2087 6783
rect 2087 6749 2096 6783
rect 2044 6740 2096 6749
rect 2596 6740 2648 6792
rect 4252 6783 4304 6792
rect 4252 6749 4261 6783
rect 4261 6749 4295 6783
rect 4295 6749 4304 6783
rect 4252 6740 4304 6749
rect 4712 6808 4764 6860
rect 5264 6808 5316 6860
rect 5356 6672 5408 6724
rect 5724 6740 5776 6792
rect 7104 6808 7156 6860
rect 4344 6604 4396 6656
rect 4528 6604 4580 6656
rect 5264 6604 5316 6656
rect 7012 6740 7064 6792
rect 8024 6740 8076 6792
rect 6736 6604 6788 6656
rect 3547 6502 3599 6554
rect 3611 6502 3663 6554
rect 3675 6502 3727 6554
rect 3739 6502 3791 6554
rect 3803 6502 3855 6554
rect 6144 6502 6196 6554
rect 6208 6502 6260 6554
rect 6272 6502 6324 6554
rect 6336 6502 6388 6554
rect 6400 6502 6452 6554
rect 3240 6400 3292 6452
rect 1676 6264 1728 6316
rect 5172 6332 5224 6384
rect 7196 6264 7248 6316
rect 8208 6264 8260 6316
rect 4528 6239 4580 6248
rect 4528 6205 4537 6239
rect 4537 6205 4571 6239
rect 4571 6205 4580 6239
rect 4528 6196 4580 6205
rect 5448 6196 5500 6248
rect 5724 6196 5776 6248
rect 6736 6196 6788 6248
rect 1584 6103 1636 6112
rect 1584 6069 1593 6103
rect 1593 6069 1627 6103
rect 1627 6069 1636 6103
rect 1584 6060 1636 6069
rect 2136 6103 2188 6112
rect 2136 6069 2145 6103
rect 2145 6069 2179 6103
rect 2179 6069 2188 6103
rect 2136 6060 2188 6069
rect 4252 6060 4304 6112
rect 4344 6060 4396 6112
rect 2248 5958 2300 6010
rect 2312 5958 2364 6010
rect 2376 5958 2428 6010
rect 2440 5958 2492 6010
rect 2504 5958 2556 6010
rect 4846 5958 4898 6010
rect 4910 5958 4962 6010
rect 4974 5958 5026 6010
rect 5038 5958 5090 6010
rect 5102 5958 5154 6010
rect 7443 5958 7495 6010
rect 7507 5958 7559 6010
rect 7571 5958 7623 6010
rect 7635 5958 7687 6010
rect 7699 5958 7751 6010
rect 7288 5856 7340 5908
rect 7380 5788 7432 5840
rect 2136 5720 2188 5772
rect 2044 5652 2096 5704
rect 4712 5652 4764 5704
rect 5356 5652 5408 5704
rect 4160 5584 4212 5636
rect 4436 5584 4488 5636
rect 5264 5627 5316 5636
rect 5264 5593 5273 5627
rect 5273 5593 5307 5627
rect 5307 5593 5316 5627
rect 5264 5584 5316 5593
rect 5816 5720 5868 5772
rect 5632 5652 5684 5704
rect 6644 5652 6696 5704
rect 7196 5695 7248 5704
rect 7196 5661 7205 5695
rect 7205 5661 7239 5695
rect 7239 5661 7248 5695
rect 7196 5652 7248 5661
rect 7840 5652 7892 5704
rect 8116 5695 8168 5704
rect 8116 5661 8119 5695
rect 8119 5661 8153 5695
rect 8153 5661 8168 5695
rect 8116 5652 8168 5661
rect 5816 5584 5868 5636
rect 5908 5516 5960 5568
rect 6736 5559 6788 5568
rect 6736 5525 6745 5559
rect 6745 5525 6779 5559
rect 6779 5525 6788 5559
rect 6736 5516 6788 5525
rect 7104 5584 7156 5636
rect 8208 5516 8260 5568
rect 3547 5414 3599 5466
rect 3611 5414 3663 5466
rect 3675 5414 3727 5466
rect 3739 5414 3791 5466
rect 3803 5414 3855 5466
rect 6144 5414 6196 5466
rect 6208 5414 6260 5466
rect 6272 5414 6324 5466
rect 6336 5414 6388 5466
rect 6400 5414 6452 5466
rect 1860 5312 1912 5364
rect 2964 5312 3016 5364
rect 4436 5312 4488 5364
rect 4528 5312 4580 5364
rect 3792 5244 3844 5296
rect 1400 5151 1452 5160
rect 1400 5117 1409 5151
rect 1409 5117 1443 5151
rect 1443 5117 1452 5151
rect 1400 5108 1452 5117
rect 2780 5176 2832 5228
rect 6828 5244 6880 5296
rect 6920 5244 6972 5296
rect 7380 5287 7432 5296
rect 7380 5253 7389 5287
rect 7389 5253 7423 5287
rect 7423 5253 7432 5287
rect 7380 5244 7432 5253
rect 7932 5219 7984 5228
rect 7932 5185 7941 5219
rect 7941 5185 7975 5219
rect 7975 5185 7984 5219
rect 7932 5176 7984 5185
rect 6368 5151 6420 5160
rect 6368 5117 6377 5151
rect 6377 5117 6411 5151
rect 6411 5117 6420 5151
rect 6368 5108 6420 5117
rect 6552 5108 6604 5160
rect 6000 5040 6052 5092
rect 7196 5040 7248 5092
rect 3884 4972 3936 5024
rect 4436 4972 4488 5024
rect 2248 4870 2300 4922
rect 2312 4870 2364 4922
rect 2376 4870 2428 4922
rect 2440 4870 2492 4922
rect 2504 4870 2556 4922
rect 4846 4870 4898 4922
rect 4910 4870 4962 4922
rect 4974 4870 5026 4922
rect 5038 4870 5090 4922
rect 5102 4870 5154 4922
rect 7443 4870 7495 4922
rect 7507 4870 7559 4922
rect 7571 4870 7623 4922
rect 7635 4870 7687 4922
rect 7699 4870 7751 4922
rect 6368 4768 6420 4820
rect 2044 4632 2096 4684
rect 2780 4564 2832 4616
rect 2596 4496 2648 4548
rect 3976 4564 4028 4616
rect 2964 4428 3016 4480
rect 4160 4496 4212 4548
rect 4528 4564 4580 4616
rect 5816 4564 5868 4616
rect 6828 4607 6880 4616
rect 6828 4573 6837 4607
rect 6837 4573 6871 4607
rect 6871 4573 6880 4607
rect 6828 4564 6880 4573
rect 4804 4539 4856 4548
rect 4804 4505 4813 4539
rect 4813 4505 4847 4539
rect 4847 4505 4856 4539
rect 4804 4496 4856 4505
rect 5908 4539 5960 4548
rect 4344 4428 4396 4480
rect 5908 4505 5917 4539
rect 5917 4505 5951 4539
rect 5951 4505 5960 4539
rect 5908 4496 5960 4505
rect 7288 4539 7340 4548
rect 7288 4505 7297 4539
rect 7297 4505 7331 4539
rect 7331 4505 7340 4539
rect 7288 4496 7340 4505
rect 3547 4326 3599 4378
rect 3611 4326 3663 4378
rect 3675 4326 3727 4378
rect 3739 4326 3791 4378
rect 3803 4326 3855 4378
rect 6144 4326 6196 4378
rect 6208 4326 6260 4378
rect 6272 4326 6324 4378
rect 6336 4326 6388 4378
rect 6400 4326 6452 4378
rect 4160 4224 4212 4276
rect 4528 4224 4580 4276
rect 4804 4156 4856 4208
rect 4436 4131 4488 4140
rect 1860 4020 1912 4072
rect 4436 4097 4445 4131
rect 4445 4097 4479 4131
rect 4479 4097 4488 4131
rect 4436 4088 4488 4097
rect 5356 4131 5408 4140
rect 4160 4020 4212 4072
rect 5356 4097 5365 4131
rect 5365 4097 5399 4131
rect 5399 4097 5408 4131
rect 5356 4088 5408 4097
rect 5908 4088 5960 4140
rect 6552 4088 6604 4140
rect 8208 4088 8260 4140
rect 2780 3884 2832 3936
rect 6000 3952 6052 4004
rect 3976 3884 4028 3936
rect 2248 3782 2300 3834
rect 2312 3782 2364 3834
rect 2376 3782 2428 3834
rect 2440 3782 2492 3834
rect 2504 3782 2556 3834
rect 4846 3782 4898 3834
rect 4910 3782 4962 3834
rect 4974 3782 5026 3834
rect 5038 3782 5090 3834
rect 5102 3782 5154 3834
rect 7443 3782 7495 3834
rect 7507 3782 7559 3834
rect 7571 3782 7623 3834
rect 7635 3782 7687 3834
rect 7699 3782 7751 3834
rect 1860 3723 1912 3732
rect 1860 3689 1869 3723
rect 1869 3689 1903 3723
rect 1903 3689 1912 3723
rect 1860 3680 1912 3689
rect 2044 3680 2096 3732
rect 4344 3655 4396 3664
rect 4344 3621 4353 3655
rect 4353 3621 4387 3655
rect 4387 3621 4396 3655
rect 4344 3612 4396 3621
rect 2688 3408 2740 3460
rect 3424 3544 3476 3596
rect 4528 3544 4580 3596
rect 4436 3519 4488 3528
rect 4436 3485 4445 3519
rect 4445 3485 4479 3519
rect 4479 3485 4488 3519
rect 4436 3476 4488 3485
rect 5816 3519 5868 3528
rect 5816 3485 5825 3519
rect 5825 3485 5859 3519
rect 5859 3485 5868 3519
rect 5816 3476 5868 3485
rect 6920 3476 6972 3528
rect 8300 3476 8352 3528
rect 6552 3451 6604 3460
rect 6552 3417 6561 3451
rect 6561 3417 6595 3451
rect 6595 3417 6604 3451
rect 6552 3408 6604 3417
rect 3547 3238 3599 3290
rect 3611 3238 3663 3290
rect 3675 3238 3727 3290
rect 3739 3238 3791 3290
rect 3803 3238 3855 3290
rect 6144 3238 6196 3290
rect 6208 3238 6260 3290
rect 6272 3238 6324 3290
rect 6336 3238 6388 3290
rect 6400 3238 6452 3290
rect 2872 3136 2924 3188
rect 4344 3136 4396 3188
rect 5356 3136 5408 3188
rect 6828 3136 6880 3188
rect 1676 3068 1728 3120
rect 6552 3068 6604 3120
rect 6920 3111 6972 3120
rect 6920 3077 6929 3111
rect 6929 3077 6963 3111
rect 6963 3077 6972 3111
rect 6920 3068 6972 3077
rect 7196 3111 7248 3120
rect 7196 3077 7205 3111
rect 7205 3077 7239 3111
rect 7239 3077 7248 3111
rect 7196 3068 7248 3077
rect 2688 3000 2740 3052
rect 5264 3000 5316 3052
rect 7932 3000 7984 3052
rect 3608 2864 3660 2916
rect 4436 2864 4488 2916
rect 6920 2864 6972 2916
rect 940 2796 992 2848
rect 1952 2796 2004 2848
rect 3884 2796 3936 2848
rect 4712 2796 4764 2848
rect 6644 2796 6696 2848
rect 6828 2796 6880 2848
rect 2248 2694 2300 2746
rect 2312 2694 2364 2746
rect 2376 2694 2428 2746
rect 2440 2694 2492 2746
rect 2504 2694 2556 2746
rect 4846 2694 4898 2746
rect 4910 2694 4962 2746
rect 4974 2694 5026 2746
rect 5038 2694 5090 2746
rect 5102 2694 5154 2746
rect 7443 2694 7495 2746
rect 7507 2694 7559 2746
rect 7571 2694 7623 2746
rect 7635 2694 7687 2746
rect 7699 2694 7751 2746
rect 2596 2592 2648 2644
rect 5264 2635 5316 2644
rect 5264 2601 5273 2635
rect 5273 2601 5307 2635
rect 5307 2601 5316 2635
rect 5264 2592 5316 2601
rect 6552 2592 6604 2644
rect 7012 2524 7064 2576
rect 3608 2388 3660 2440
rect 3056 2363 3108 2372
rect 3056 2329 3065 2363
rect 3065 2329 3099 2363
rect 3099 2329 3108 2363
rect 3056 2320 3108 2329
rect 1860 2295 1912 2304
rect 1860 2261 1869 2295
rect 1869 2261 1903 2295
rect 1903 2261 1912 2295
rect 3148 2295 3200 2304
rect 1860 2252 1912 2261
rect 3148 2261 3157 2295
rect 3157 2261 3191 2295
rect 3191 2261 3200 2295
rect 3148 2252 3200 2261
rect 3884 2456 3936 2508
rect 5724 2456 5776 2508
rect 7840 2456 7892 2508
rect 8300 2456 8352 2508
rect 4344 2431 4396 2440
rect 4344 2397 4353 2431
rect 4353 2397 4387 2431
rect 4387 2397 4396 2431
rect 4344 2388 4396 2397
rect 4712 2431 4764 2440
rect 4712 2397 4721 2431
rect 4721 2397 4755 2431
rect 4755 2397 4764 2431
rect 4712 2388 4764 2397
rect 3976 2363 4028 2372
rect 3976 2329 3985 2363
rect 3985 2329 4019 2363
rect 4019 2329 4028 2363
rect 3976 2320 4028 2329
rect 4252 2363 4304 2372
rect 4252 2329 4261 2363
rect 4261 2329 4295 2363
rect 4295 2329 4304 2363
rect 4252 2320 4304 2329
rect 4528 2320 4580 2372
rect 3547 2150 3599 2202
rect 3611 2150 3663 2202
rect 3675 2150 3727 2202
rect 3739 2150 3791 2202
rect 3803 2150 3855 2202
rect 6144 2150 6196 2202
rect 6208 2150 6260 2202
rect 6272 2150 6324 2202
rect 6336 2150 6388 2202
rect 6400 2150 6452 2202
rect 1860 2048 1912 2100
rect 3148 2048 3200 2100
rect 5632 2048 5684 2100
rect 7196 1980 7248 2032
rect 3056 1708 3108 1760
rect 8944 1708 8996 1760
rect 4068 1300 4120 1352
rect 6552 1300 6604 1352
<< metal2 >>
rect 6642 29744 6698 29753
rect 6642 29679 6698 29688
rect 6550 29200 6606 29209
rect 6550 29135 6606 29144
rect 5538 28656 5594 28665
rect 5538 28591 5594 28600
rect 2248 27772 2556 27792
rect 2248 27770 2254 27772
rect 2310 27770 2334 27772
rect 2390 27770 2414 27772
rect 2470 27770 2494 27772
rect 2550 27770 2556 27772
rect 2310 27718 2312 27770
rect 2492 27718 2494 27770
rect 2248 27716 2254 27718
rect 2310 27716 2334 27718
rect 2390 27716 2414 27718
rect 2470 27716 2494 27718
rect 2550 27716 2556 27718
rect 2248 27696 2556 27716
rect 4846 27772 5154 27792
rect 4846 27770 4852 27772
rect 4908 27770 4932 27772
rect 4988 27770 5012 27772
rect 5068 27770 5092 27772
rect 5148 27770 5154 27772
rect 4908 27718 4910 27770
rect 5090 27718 5092 27770
rect 4846 27716 4852 27718
rect 4908 27716 4932 27718
rect 4988 27716 5012 27718
rect 5068 27716 5092 27718
rect 5148 27716 5154 27718
rect 4846 27696 5154 27716
rect 2596 27600 2648 27606
rect 2596 27542 2648 27548
rect 2044 27532 2096 27538
rect 2044 27474 2096 27480
rect 2056 27130 2084 27474
rect 2044 27124 2096 27130
rect 2044 27066 2096 27072
rect 2248 26684 2556 26704
rect 2248 26682 2254 26684
rect 2310 26682 2334 26684
rect 2390 26682 2414 26684
rect 2470 26682 2494 26684
rect 2550 26682 2556 26684
rect 2310 26630 2312 26682
rect 2492 26630 2494 26682
rect 2248 26628 2254 26630
rect 2310 26628 2334 26630
rect 2390 26628 2414 26630
rect 2470 26628 2494 26630
rect 2550 26628 2556 26630
rect 2248 26608 2556 26628
rect 2608 26586 2636 27542
rect 5552 27538 5580 28591
rect 5998 28112 6054 28121
rect 5998 28047 6054 28056
rect 5816 27600 5868 27606
rect 5816 27542 5868 27548
rect 5906 27568 5962 27577
rect 5540 27532 5592 27538
rect 5540 27474 5592 27480
rect 4068 27464 4120 27470
rect 4068 27406 4120 27412
rect 4160 27464 4212 27470
rect 4160 27406 4212 27412
rect 3884 27396 3936 27402
rect 3884 27338 3936 27344
rect 2688 27328 2740 27334
rect 2688 27270 2740 27276
rect 2596 26580 2648 26586
rect 2596 26522 2648 26528
rect 2044 26036 2096 26042
rect 2044 25978 2096 25984
rect 2056 25498 2084 25978
rect 2700 25974 2728 27270
rect 3547 27228 3855 27248
rect 3547 27226 3553 27228
rect 3609 27226 3633 27228
rect 3689 27226 3713 27228
rect 3769 27226 3793 27228
rect 3849 27226 3855 27228
rect 3609 27174 3611 27226
rect 3791 27174 3793 27226
rect 3547 27172 3553 27174
rect 3609 27172 3633 27174
rect 3689 27172 3713 27174
rect 3769 27172 3793 27174
rect 3849 27172 3855 27174
rect 3547 27152 3855 27172
rect 3240 26988 3292 26994
rect 3240 26930 3292 26936
rect 3424 26988 3476 26994
rect 3424 26930 3476 26936
rect 2780 26784 2832 26790
rect 2780 26726 2832 26732
rect 2792 26586 2820 26726
rect 2780 26580 2832 26586
rect 2780 26522 2832 26528
rect 3252 26518 3280 26930
rect 3240 26512 3292 26518
rect 3240 26454 3292 26460
rect 2688 25968 2740 25974
rect 2688 25910 2740 25916
rect 3436 25906 3464 26930
rect 3547 26140 3855 26160
rect 3547 26138 3553 26140
rect 3609 26138 3633 26140
rect 3689 26138 3713 26140
rect 3769 26138 3793 26140
rect 3849 26138 3855 26140
rect 3609 26086 3611 26138
rect 3791 26086 3793 26138
rect 3547 26084 3553 26086
rect 3609 26084 3633 26086
rect 3689 26084 3713 26086
rect 3769 26084 3793 26086
rect 3849 26084 3855 26086
rect 3547 26064 3855 26084
rect 3424 25900 3476 25906
rect 3424 25842 3476 25848
rect 2248 25596 2556 25616
rect 2248 25594 2254 25596
rect 2310 25594 2334 25596
rect 2390 25594 2414 25596
rect 2470 25594 2494 25596
rect 2550 25594 2556 25596
rect 2310 25542 2312 25594
rect 2492 25542 2494 25594
rect 2248 25540 2254 25542
rect 2310 25540 2334 25542
rect 2390 25540 2414 25542
rect 2470 25540 2494 25542
rect 2550 25540 2556 25542
rect 2248 25520 2556 25540
rect 2044 25492 2096 25498
rect 2044 25434 2096 25440
rect 3436 24818 3464 25842
rect 3547 25052 3855 25072
rect 3547 25050 3553 25052
rect 3609 25050 3633 25052
rect 3689 25050 3713 25052
rect 3769 25050 3793 25052
rect 3849 25050 3855 25052
rect 3609 24998 3611 25050
rect 3791 24998 3793 25050
rect 3547 24996 3553 24998
rect 3609 24996 3633 24998
rect 3689 24996 3713 24998
rect 3769 24996 3793 24998
rect 3849 24996 3855 24998
rect 3547 24976 3855 24996
rect 3424 24812 3476 24818
rect 3424 24754 3476 24760
rect 3896 24682 3924 27338
rect 3976 27328 4028 27334
rect 3976 27270 4028 27276
rect 3988 26450 4016 27270
rect 3976 26444 4028 26450
rect 3976 26386 4028 26392
rect 4080 26314 4108 27406
rect 4172 26382 4200 27406
rect 4528 27396 4580 27402
rect 4528 27338 4580 27344
rect 5448 27396 5500 27402
rect 5448 27338 5500 27344
rect 4540 26994 4568 27338
rect 5460 27062 5488 27338
rect 5448 27056 5500 27062
rect 5448 26998 5500 27004
rect 5552 26994 5580 27474
rect 5632 27328 5684 27334
rect 5632 27270 5684 27276
rect 4528 26988 4580 26994
rect 4528 26930 4580 26936
rect 5540 26988 5592 26994
rect 5540 26930 5592 26936
rect 4160 26376 4212 26382
rect 4160 26318 4212 26324
rect 4068 26308 4120 26314
rect 4068 26250 4120 26256
rect 4080 25974 4108 26250
rect 4068 25968 4120 25974
rect 4068 25910 4120 25916
rect 4160 25900 4212 25906
rect 4160 25842 4212 25848
rect 3884 24676 3936 24682
rect 3884 24618 3936 24624
rect 2964 24608 3016 24614
rect 2964 24550 3016 24556
rect 2248 24508 2556 24528
rect 2248 24506 2254 24508
rect 2310 24506 2334 24508
rect 2390 24506 2414 24508
rect 2470 24506 2494 24508
rect 2550 24506 2556 24508
rect 2310 24454 2312 24506
rect 2492 24454 2494 24506
rect 2248 24452 2254 24454
rect 2310 24452 2334 24454
rect 2390 24452 2414 24454
rect 2470 24452 2494 24454
rect 2550 24452 2556 24454
rect 2248 24432 2556 24452
rect 2976 24138 3004 24550
rect 4172 24274 4200 25842
rect 4540 25294 4568 26930
rect 5172 26784 5224 26790
rect 5172 26726 5224 26732
rect 4846 26684 5154 26704
rect 4846 26682 4852 26684
rect 4908 26682 4932 26684
rect 4988 26682 5012 26684
rect 5068 26682 5092 26684
rect 5148 26682 5154 26684
rect 4908 26630 4910 26682
rect 5090 26630 5092 26682
rect 4846 26628 4852 26630
rect 4908 26628 4932 26630
rect 4988 26628 5012 26630
rect 5068 26628 5092 26630
rect 5148 26628 5154 26630
rect 4846 26608 5154 26628
rect 4846 25596 5154 25616
rect 4846 25594 4852 25596
rect 4908 25594 4932 25596
rect 4988 25594 5012 25596
rect 5068 25594 5092 25596
rect 5148 25594 5154 25596
rect 4908 25542 4910 25594
rect 5090 25542 5092 25594
rect 4846 25540 4852 25542
rect 4908 25540 4932 25542
rect 4988 25540 5012 25542
rect 5068 25540 5092 25542
rect 5148 25540 5154 25542
rect 4846 25520 5154 25540
rect 5184 25362 5212 26726
rect 5264 26240 5316 26246
rect 5264 26182 5316 26188
rect 5276 25906 5304 26182
rect 5264 25900 5316 25906
rect 5264 25842 5316 25848
rect 5264 25764 5316 25770
rect 5264 25706 5316 25712
rect 5276 25430 5304 25706
rect 5264 25424 5316 25430
rect 5264 25366 5316 25372
rect 5172 25356 5224 25362
rect 5172 25298 5224 25304
rect 4528 25288 4580 25294
rect 4528 25230 4580 25236
rect 4252 25220 4304 25226
rect 4252 25162 4304 25168
rect 4264 24682 4292 25162
rect 5644 24834 5672 27270
rect 5722 27024 5778 27033
rect 5828 26994 5856 27542
rect 5906 27503 5962 27512
rect 5722 26959 5778 26968
rect 5816 26988 5868 26994
rect 5736 25838 5764 26959
rect 5816 26930 5868 26936
rect 5920 26858 5948 27503
rect 5908 26852 5960 26858
rect 5908 26794 5960 26800
rect 5920 26382 5948 26794
rect 5908 26376 5960 26382
rect 5908 26318 5960 26324
rect 5908 26240 5960 26246
rect 5908 26182 5960 26188
rect 5724 25832 5776 25838
rect 5724 25774 5776 25780
rect 5736 25362 5764 25774
rect 5724 25356 5776 25362
rect 5724 25298 5776 25304
rect 5644 24818 5764 24834
rect 5644 24812 5776 24818
rect 5644 24806 5724 24812
rect 4252 24676 4304 24682
rect 4252 24618 4304 24624
rect 4160 24268 4212 24274
rect 4160 24210 4212 24216
rect 2964 24132 3016 24138
rect 2964 24074 3016 24080
rect 4160 24132 4212 24138
rect 4160 24074 4212 24080
rect 2136 24064 2188 24070
rect 2136 24006 2188 24012
rect 3240 24064 3292 24070
rect 3240 24006 3292 24012
rect 3976 24064 4028 24070
rect 3976 24006 4028 24012
rect 2148 23594 2176 24006
rect 3252 23594 3280 24006
rect 3547 23964 3855 23984
rect 3547 23962 3553 23964
rect 3609 23962 3633 23964
rect 3689 23962 3713 23964
rect 3769 23962 3793 23964
rect 3849 23962 3855 23964
rect 3609 23910 3611 23962
rect 3791 23910 3793 23962
rect 3547 23908 3553 23910
rect 3609 23908 3633 23910
rect 3689 23908 3713 23910
rect 3769 23908 3793 23910
rect 3849 23908 3855 23910
rect 3547 23888 3855 23908
rect 3988 23866 4016 24006
rect 4172 23866 4200 24074
rect 3976 23860 4028 23866
rect 3976 23802 4028 23808
rect 4160 23860 4212 23866
rect 4160 23802 4212 23808
rect 2136 23588 2188 23594
rect 2136 23530 2188 23536
rect 3240 23588 3292 23594
rect 3240 23530 3292 23536
rect 2248 23420 2556 23440
rect 2248 23418 2254 23420
rect 2310 23418 2334 23420
rect 2390 23418 2414 23420
rect 2470 23418 2494 23420
rect 2550 23418 2556 23420
rect 2310 23366 2312 23418
rect 2492 23366 2494 23418
rect 2248 23364 2254 23366
rect 2310 23364 2334 23366
rect 2390 23364 2414 23366
rect 2470 23364 2494 23366
rect 2550 23364 2556 23366
rect 2248 23344 2556 23364
rect 3056 23316 3108 23322
rect 3056 23258 3108 23264
rect 2596 23112 2648 23118
rect 2596 23054 2648 23060
rect 2248 22332 2556 22352
rect 2248 22330 2254 22332
rect 2310 22330 2334 22332
rect 2390 22330 2414 22332
rect 2470 22330 2494 22332
rect 2550 22330 2556 22332
rect 2310 22278 2312 22330
rect 2492 22278 2494 22330
rect 2248 22276 2254 22278
rect 2310 22276 2334 22278
rect 2390 22276 2414 22278
rect 2470 22276 2494 22278
rect 2550 22276 2556 22278
rect 2248 22256 2556 22276
rect 2608 21690 2636 23054
rect 3068 22778 3096 23258
rect 3240 22976 3292 22982
rect 3240 22918 3292 22924
rect 3056 22772 3108 22778
rect 3056 22714 3108 22720
rect 2688 22432 2740 22438
rect 2688 22374 2740 22380
rect 2700 22166 2728 22374
rect 3252 22234 3280 22918
rect 3547 22876 3855 22896
rect 3547 22874 3553 22876
rect 3609 22874 3633 22876
rect 3689 22874 3713 22876
rect 3769 22874 3793 22876
rect 3849 22874 3855 22876
rect 3609 22822 3611 22874
rect 3791 22822 3793 22874
rect 3547 22820 3553 22822
rect 3609 22820 3633 22822
rect 3689 22820 3713 22822
rect 3769 22820 3793 22822
rect 3849 22820 3855 22822
rect 3547 22800 3855 22820
rect 4264 22710 4292 24618
rect 4846 24508 5154 24528
rect 4846 24506 4852 24508
rect 4908 24506 4932 24508
rect 4988 24506 5012 24508
rect 5068 24506 5092 24508
rect 5148 24506 5154 24508
rect 4908 24454 4910 24506
rect 5090 24454 5092 24506
rect 4846 24452 4852 24454
rect 4908 24452 4932 24454
rect 4988 24452 5012 24454
rect 5068 24452 5092 24454
rect 5148 24452 5154 24454
rect 4846 24432 5154 24452
rect 5356 24268 5408 24274
rect 5356 24210 5408 24216
rect 5368 23798 5396 24210
rect 5644 24206 5672 24806
rect 5724 24754 5776 24760
rect 5632 24200 5684 24206
rect 5632 24142 5684 24148
rect 5356 23792 5408 23798
rect 5356 23734 5408 23740
rect 5644 23662 5672 24142
rect 5632 23656 5684 23662
rect 5632 23598 5684 23604
rect 5816 23656 5868 23662
rect 5816 23598 5868 23604
rect 5828 23526 5856 23598
rect 5816 23520 5868 23526
rect 5816 23462 5868 23468
rect 4846 23420 5154 23440
rect 4846 23418 4852 23420
rect 4908 23418 4932 23420
rect 4988 23418 5012 23420
rect 5068 23418 5092 23420
rect 5148 23418 5154 23420
rect 4908 23366 4910 23418
rect 5090 23366 5092 23418
rect 4846 23364 4852 23366
rect 4908 23364 4932 23366
rect 4988 23364 5012 23366
rect 5068 23364 5092 23366
rect 5148 23364 5154 23366
rect 4846 23344 5154 23364
rect 5920 23118 5948 26182
rect 6012 25294 6040 28047
rect 6144 27228 6452 27248
rect 6144 27226 6150 27228
rect 6206 27226 6230 27228
rect 6286 27226 6310 27228
rect 6366 27226 6390 27228
rect 6446 27226 6452 27228
rect 6206 27174 6208 27226
rect 6388 27174 6390 27226
rect 6144 27172 6150 27174
rect 6206 27172 6230 27174
rect 6286 27172 6310 27174
rect 6366 27172 6390 27174
rect 6446 27172 6452 27174
rect 6144 27152 6452 27172
rect 6460 27056 6512 27062
rect 6460 26998 6512 27004
rect 6472 26518 6500 26998
rect 6460 26512 6512 26518
rect 6460 26454 6512 26460
rect 6144 26140 6452 26160
rect 6144 26138 6150 26140
rect 6206 26138 6230 26140
rect 6286 26138 6310 26140
rect 6366 26138 6390 26140
rect 6446 26138 6452 26140
rect 6206 26086 6208 26138
rect 6388 26086 6390 26138
rect 6144 26084 6150 26086
rect 6206 26084 6230 26086
rect 6286 26084 6310 26086
rect 6366 26084 6390 26086
rect 6446 26084 6452 26086
rect 6144 26064 6452 26084
rect 6000 25288 6052 25294
rect 6000 25230 6052 25236
rect 6012 24886 6040 25230
rect 6144 25052 6452 25072
rect 6144 25050 6150 25052
rect 6206 25050 6230 25052
rect 6286 25050 6310 25052
rect 6366 25050 6390 25052
rect 6446 25050 6452 25052
rect 6206 24998 6208 25050
rect 6388 24998 6390 25050
rect 6144 24996 6150 24998
rect 6206 24996 6230 24998
rect 6286 24996 6310 24998
rect 6366 24996 6390 24998
rect 6446 24996 6452 24998
rect 6144 24976 6452 24996
rect 6564 24954 6592 29135
rect 6656 26246 6684 29679
rect 7443 27772 7751 27792
rect 7443 27770 7449 27772
rect 7505 27770 7529 27772
rect 7585 27770 7609 27772
rect 7665 27770 7689 27772
rect 7745 27770 7751 27772
rect 7505 27718 7507 27770
rect 7687 27718 7689 27770
rect 7443 27716 7449 27718
rect 7505 27716 7529 27718
rect 7585 27716 7609 27718
rect 7665 27716 7689 27718
rect 7745 27716 7751 27718
rect 7443 27696 7751 27716
rect 7840 27464 7892 27470
rect 7840 27406 7892 27412
rect 6828 27396 6880 27402
rect 6828 27338 6880 27344
rect 7380 27396 7432 27402
rect 7380 27338 7432 27344
rect 6840 26858 6868 27338
rect 6920 27328 6972 27334
rect 6920 27270 6972 27276
rect 6828 26852 6880 26858
rect 6828 26794 6880 26800
rect 6734 26480 6790 26489
rect 6734 26415 6790 26424
rect 6644 26240 6696 26246
rect 6644 26182 6696 26188
rect 6642 25936 6698 25945
rect 6642 25871 6698 25880
rect 6552 24948 6604 24954
rect 6552 24890 6604 24896
rect 6000 24880 6052 24886
rect 6000 24822 6052 24828
rect 6092 24880 6144 24886
rect 6092 24822 6144 24828
rect 6104 24154 6132 24822
rect 6552 24812 6604 24818
rect 6552 24754 6604 24760
rect 6564 24342 6592 24754
rect 6552 24336 6604 24342
rect 6552 24278 6604 24284
rect 6656 24206 6684 25871
rect 6748 24818 6776 26415
rect 6840 25430 6868 26794
rect 6932 26382 6960 27270
rect 7392 27130 7420 27338
rect 7380 27124 7432 27130
rect 7380 27066 7432 27072
rect 7196 26920 7248 26926
rect 7392 26874 7420 27066
rect 7196 26862 7248 26868
rect 6920 26376 6972 26382
rect 6972 26324 7052 26330
rect 6920 26318 7052 26324
rect 6932 26302 7052 26318
rect 7024 25974 7052 26302
rect 7208 26042 7236 26862
rect 7300 26846 7420 26874
rect 7196 26036 7248 26042
rect 7196 25978 7248 25984
rect 7300 25974 7328 26846
rect 7443 26684 7751 26704
rect 7443 26682 7449 26684
rect 7505 26682 7529 26684
rect 7585 26682 7609 26684
rect 7665 26682 7689 26684
rect 7745 26682 7751 26684
rect 7505 26630 7507 26682
rect 7687 26630 7689 26682
rect 7443 26628 7449 26630
rect 7505 26628 7529 26630
rect 7585 26628 7609 26630
rect 7665 26628 7689 26630
rect 7745 26628 7751 26630
rect 7443 26608 7751 26628
rect 7012 25968 7064 25974
rect 7012 25910 7064 25916
rect 7288 25968 7340 25974
rect 7288 25910 7340 25916
rect 7852 25906 7880 27406
rect 7932 26988 7984 26994
rect 7932 26930 7984 26936
rect 7944 26382 7972 26930
rect 8208 26920 8260 26926
rect 8208 26862 8260 26868
rect 7932 26376 7984 26382
rect 7932 26318 7984 26324
rect 6920 25900 6972 25906
rect 6920 25842 6972 25848
rect 7840 25900 7892 25906
rect 7840 25842 7892 25848
rect 6828 25424 6880 25430
rect 6828 25366 6880 25372
rect 6736 24812 6788 24818
rect 6736 24754 6788 24760
rect 6012 24126 6132 24154
rect 6644 24200 6696 24206
rect 6644 24142 6696 24148
rect 5908 23112 5960 23118
rect 5908 23054 5960 23060
rect 4620 23044 4672 23050
rect 4620 22986 4672 22992
rect 5172 23044 5224 23050
rect 5172 22986 5224 22992
rect 5264 23044 5316 23050
rect 5264 22986 5316 22992
rect 4252 22704 4304 22710
rect 4252 22646 4304 22652
rect 4160 22568 4212 22574
rect 4160 22510 4212 22516
rect 4068 22432 4120 22438
rect 4068 22374 4120 22380
rect 3240 22228 3292 22234
rect 3240 22170 3292 22176
rect 4080 22166 4108 22374
rect 2688 22160 2740 22166
rect 2688 22102 2740 22108
rect 4068 22160 4120 22166
rect 4068 22102 4120 22108
rect 4172 22098 4200 22510
rect 4528 22500 4580 22506
rect 4528 22442 4580 22448
rect 4252 22160 4304 22166
rect 4252 22102 4304 22108
rect 4160 22092 4212 22098
rect 4160 22034 4212 22040
rect 3547 21788 3855 21808
rect 3547 21786 3553 21788
rect 3609 21786 3633 21788
rect 3689 21786 3713 21788
rect 3769 21786 3793 21788
rect 3849 21786 3855 21788
rect 3609 21734 3611 21786
rect 3791 21734 3793 21786
rect 3547 21732 3553 21734
rect 3609 21732 3633 21734
rect 3689 21732 3713 21734
rect 3769 21732 3793 21734
rect 3849 21732 3855 21734
rect 3547 21712 3855 21732
rect 2596 21684 2648 21690
rect 2596 21626 2648 21632
rect 3148 21344 3200 21350
rect 3148 21286 3200 21292
rect 3240 21344 3292 21350
rect 3240 21286 3292 21292
rect 2248 21244 2556 21264
rect 2248 21242 2254 21244
rect 2310 21242 2334 21244
rect 2390 21242 2414 21244
rect 2470 21242 2494 21244
rect 2550 21242 2556 21244
rect 2310 21190 2312 21242
rect 2492 21190 2494 21242
rect 2248 21188 2254 21190
rect 2310 21188 2334 21190
rect 2390 21188 2414 21190
rect 2470 21188 2494 21190
rect 2550 21188 2556 21190
rect 2248 21168 2556 21188
rect 2596 21072 2648 21078
rect 2596 21014 2648 21020
rect 2608 20806 2636 21014
rect 2596 20800 2648 20806
rect 2596 20742 2648 20748
rect 2248 20156 2556 20176
rect 2248 20154 2254 20156
rect 2310 20154 2334 20156
rect 2390 20154 2414 20156
rect 2470 20154 2494 20156
rect 2550 20154 2556 20156
rect 2310 20102 2312 20154
rect 2492 20102 2494 20154
rect 2248 20100 2254 20102
rect 2310 20100 2334 20102
rect 2390 20100 2414 20102
rect 2470 20100 2494 20102
rect 2550 20100 2556 20102
rect 2248 20080 2556 20100
rect 1584 19712 1636 19718
rect 1584 19654 1636 19660
rect 2044 19712 2096 19718
rect 2044 19654 2096 19660
rect 1596 19242 1624 19654
rect 1584 19236 1636 19242
rect 1584 19178 1636 19184
rect 2056 18698 2084 19654
rect 2608 19310 2636 20742
rect 2688 20256 2740 20262
rect 2688 20198 2740 20204
rect 2596 19304 2648 19310
rect 2596 19246 2648 19252
rect 2248 19068 2556 19088
rect 2248 19066 2254 19068
rect 2310 19066 2334 19068
rect 2390 19066 2414 19068
rect 2470 19066 2494 19068
rect 2550 19066 2556 19068
rect 2310 19014 2312 19066
rect 2492 19014 2494 19066
rect 2248 19012 2254 19014
rect 2310 19012 2334 19014
rect 2390 19012 2414 19014
rect 2470 19012 2494 19014
rect 2550 19012 2556 19014
rect 2248 18992 2556 19012
rect 2700 18970 2728 20198
rect 3160 20058 3188 21286
rect 3252 21146 3280 21286
rect 3240 21140 3292 21146
rect 3240 21082 3292 21088
rect 4160 20936 4212 20942
rect 4160 20878 4212 20884
rect 4068 20800 4120 20806
rect 4068 20742 4120 20748
rect 3547 20700 3855 20720
rect 3547 20698 3553 20700
rect 3609 20698 3633 20700
rect 3689 20698 3713 20700
rect 3769 20698 3793 20700
rect 3849 20698 3855 20700
rect 3609 20646 3611 20698
rect 3791 20646 3793 20698
rect 3547 20644 3553 20646
rect 3609 20644 3633 20646
rect 3689 20644 3713 20646
rect 3769 20644 3793 20646
rect 3849 20644 3855 20646
rect 3547 20624 3855 20644
rect 4080 20534 4108 20742
rect 4068 20528 4120 20534
rect 4068 20470 4120 20476
rect 4172 20466 4200 20878
rect 4160 20460 4212 20466
rect 4160 20402 4212 20408
rect 4264 20346 4292 22102
rect 4540 22030 4568 22442
rect 4528 22024 4580 22030
rect 4528 21966 4580 21972
rect 4632 21690 4660 22986
rect 4712 22500 4764 22506
rect 4712 22442 4764 22448
rect 4724 22166 4752 22442
rect 4846 22332 5154 22352
rect 4846 22330 4852 22332
rect 4908 22330 4932 22332
rect 4988 22330 5012 22332
rect 5068 22330 5092 22332
rect 5148 22330 5154 22332
rect 4908 22278 4910 22330
rect 5090 22278 5092 22330
rect 4846 22276 4852 22278
rect 4908 22276 4932 22278
rect 4988 22276 5012 22278
rect 5068 22276 5092 22278
rect 5148 22276 5154 22278
rect 4846 22256 5154 22276
rect 4712 22160 4764 22166
rect 4712 22102 4764 22108
rect 5184 22094 5212 22986
rect 5276 22778 5304 22986
rect 5264 22772 5316 22778
rect 5264 22714 5316 22720
rect 5092 22066 5212 22094
rect 4896 22024 4948 22030
rect 4896 21966 4948 21972
rect 4620 21684 4672 21690
rect 4620 21626 4672 21632
rect 4908 21622 4936 21966
rect 5092 21894 5120 22066
rect 5080 21888 5132 21894
rect 5080 21830 5132 21836
rect 5092 21622 5120 21830
rect 4896 21616 4948 21622
rect 4896 21558 4948 21564
rect 5080 21616 5132 21622
rect 5080 21558 5132 21564
rect 5920 21554 5948 23054
rect 6012 22574 6040 24126
rect 6144 23964 6452 23984
rect 6144 23962 6150 23964
rect 6206 23962 6230 23964
rect 6286 23962 6310 23964
rect 6366 23962 6390 23964
rect 6446 23962 6452 23964
rect 6206 23910 6208 23962
rect 6388 23910 6390 23962
rect 6144 23908 6150 23910
rect 6206 23908 6230 23910
rect 6286 23908 6310 23910
rect 6366 23908 6390 23910
rect 6446 23908 6452 23910
rect 6144 23888 6452 23908
rect 6656 23882 6684 24142
rect 6748 24138 6776 24754
rect 6932 24342 6960 25842
rect 7443 25596 7751 25616
rect 7443 25594 7449 25596
rect 7505 25594 7529 25596
rect 7585 25594 7609 25596
rect 7665 25594 7689 25596
rect 7745 25594 7751 25596
rect 7505 25542 7507 25594
rect 7687 25542 7689 25594
rect 7443 25540 7449 25542
rect 7505 25540 7529 25542
rect 7585 25540 7609 25542
rect 7665 25540 7689 25542
rect 7745 25540 7751 25542
rect 7443 25520 7751 25540
rect 7852 25401 7880 25842
rect 7838 25392 7894 25401
rect 7838 25327 7894 25336
rect 7196 25288 7248 25294
rect 7196 25230 7248 25236
rect 6920 24336 6972 24342
rect 6920 24278 6972 24284
rect 6736 24132 6788 24138
rect 6736 24074 6788 24080
rect 6564 23854 6684 23882
rect 6564 23662 6592 23854
rect 7208 23798 7236 25230
rect 7944 24857 7972 26318
rect 8220 25294 8248 26862
rect 8208 25288 8260 25294
rect 8208 25230 8260 25236
rect 7930 24848 7986 24857
rect 7840 24812 7892 24818
rect 7930 24783 7986 24792
rect 7840 24754 7892 24760
rect 7288 24676 7340 24682
rect 7288 24618 7340 24624
rect 7196 23792 7248 23798
rect 7196 23734 7248 23740
rect 6644 23724 6696 23730
rect 6644 23666 6696 23672
rect 6552 23656 6604 23662
rect 6552 23598 6604 23604
rect 6656 23254 6684 23666
rect 6644 23248 6696 23254
rect 6644 23190 6696 23196
rect 6734 23216 6790 23225
rect 6144 22876 6452 22896
rect 6144 22874 6150 22876
rect 6206 22874 6230 22876
rect 6286 22874 6310 22876
rect 6366 22874 6390 22876
rect 6446 22874 6452 22876
rect 6206 22822 6208 22874
rect 6388 22822 6390 22874
rect 6144 22820 6150 22822
rect 6206 22820 6230 22822
rect 6286 22820 6310 22822
rect 6366 22820 6390 22822
rect 6446 22820 6452 22822
rect 6144 22800 6452 22820
rect 6000 22568 6052 22574
rect 6000 22510 6052 22516
rect 6012 22030 6040 22510
rect 6656 22506 6684 23190
rect 6734 23151 6790 23160
rect 6748 23118 6776 23151
rect 6736 23112 6788 23118
rect 6736 23054 6788 23060
rect 6644 22500 6696 22506
rect 6644 22442 6696 22448
rect 6748 22234 6776 23054
rect 7012 23044 7064 23050
rect 7012 22986 7064 22992
rect 6920 22636 6972 22642
rect 6920 22578 6972 22584
rect 6736 22228 6788 22234
rect 6736 22170 6788 22176
rect 6644 22094 6696 22098
rect 6748 22094 6776 22170
rect 6644 22092 6776 22094
rect 6696 22066 6776 22092
rect 6644 22034 6696 22040
rect 6000 22024 6052 22030
rect 6000 21966 6052 21972
rect 6932 21962 6960 22578
rect 7024 22030 7052 22986
rect 7300 22642 7328 24618
rect 7443 24508 7751 24528
rect 7443 24506 7449 24508
rect 7505 24506 7529 24508
rect 7585 24506 7609 24508
rect 7665 24506 7689 24508
rect 7745 24506 7751 24508
rect 7505 24454 7507 24506
rect 7687 24454 7689 24506
rect 7443 24452 7449 24454
rect 7505 24452 7529 24454
rect 7585 24452 7609 24454
rect 7665 24452 7689 24454
rect 7745 24452 7751 24454
rect 7443 24432 7751 24452
rect 7380 24336 7432 24342
rect 7380 24278 7432 24284
rect 7392 23798 7420 24278
rect 7564 24132 7616 24138
rect 7564 24074 7616 24080
rect 7576 23866 7604 24074
rect 7564 23860 7616 23866
rect 7564 23802 7616 23808
rect 7380 23792 7432 23798
rect 7380 23734 7432 23740
rect 7443 23420 7751 23440
rect 7443 23418 7449 23420
rect 7505 23418 7529 23420
rect 7585 23418 7609 23420
rect 7665 23418 7689 23420
rect 7745 23418 7751 23420
rect 7505 23366 7507 23418
rect 7687 23366 7689 23418
rect 7443 23364 7449 23366
rect 7505 23364 7529 23366
rect 7585 23364 7609 23366
rect 7665 23364 7689 23366
rect 7745 23364 7751 23366
rect 7443 23344 7751 23364
rect 7288 22636 7340 22642
rect 7288 22578 7340 22584
rect 7443 22332 7751 22352
rect 7443 22330 7449 22332
rect 7505 22330 7529 22332
rect 7585 22330 7609 22332
rect 7665 22330 7689 22332
rect 7745 22330 7751 22332
rect 7505 22278 7507 22330
rect 7687 22278 7689 22330
rect 7443 22276 7449 22278
rect 7505 22276 7529 22278
rect 7585 22276 7609 22278
rect 7665 22276 7689 22278
rect 7745 22276 7751 22278
rect 7443 22256 7751 22276
rect 7012 22024 7064 22030
rect 7012 21966 7064 21972
rect 6920 21956 6972 21962
rect 6920 21898 6972 21904
rect 6144 21788 6452 21808
rect 6144 21786 6150 21788
rect 6206 21786 6230 21788
rect 6286 21786 6310 21788
rect 6366 21786 6390 21788
rect 6446 21786 6452 21788
rect 6206 21734 6208 21786
rect 6388 21734 6390 21786
rect 6144 21732 6150 21734
rect 6206 21732 6230 21734
rect 6286 21732 6310 21734
rect 6366 21732 6390 21734
rect 6446 21732 6452 21734
rect 6144 21712 6452 21732
rect 6734 21584 6790 21593
rect 5908 21548 5960 21554
rect 5908 21490 5960 21496
rect 6552 21548 6604 21554
rect 6734 21519 6790 21528
rect 6552 21490 6604 21496
rect 4344 21480 4396 21486
rect 4344 21422 4396 21428
rect 4356 20602 4384 21422
rect 5816 21344 5868 21350
rect 5816 21286 5868 21292
rect 4846 21244 5154 21264
rect 4846 21242 4852 21244
rect 4908 21242 4932 21244
rect 4988 21242 5012 21244
rect 5068 21242 5092 21244
rect 5148 21242 5154 21244
rect 4908 21190 4910 21242
rect 5090 21190 5092 21242
rect 4846 21188 4852 21190
rect 4908 21188 4932 21190
rect 4988 21188 5012 21190
rect 5068 21188 5092 21190
rect 5148 21188 5154 21190
rect 4846 21168 5154 21188
rect 5828 21010 5856 21286
rect 5816 21004 5868 21010
rect 5816 20946 5868 20952
rect 5632 20868 5684 20874
rect 5632 20810 5684 20816
rect 4344 20596 4396 20602
rect 4344 20538 4396 20544
rect 5644 20534 5672 20810
rect 5632 20528 5684 20534
rect 5632 20470 5684 20476
rect 5828 20466 5856 20946
rect 6144 20700 6452 20720
rect 6144 20698 6150 20700
rect 6206 20698 6230 20700
rect 6286 20698 6310 20700
rect 6366 20698 6390 20700
rect 6446 20698 6452 20700
rect 6206 20646 6208 20698
rect 6388 20646 6390 20698
rect 6144 20644 6150 20646
rect 6206 20644 6230 20646
rect 6286 20644 6310 20646
rect 6366 20644 6390 20646
rect 6446 20644 6452 20646
rect 6144 20624 6452 20644
rect 5816 20460 5868 20466
rect 5816 20402 5868 20408
rect 4172 20318 4292 20346
rect 3148 20052 3200 20058
rect 3148 19994 3200 20000
rect 4068 19916 4120 19922
rect 4068 19858 4120 19864
rect 2964 19848 3016 19854
rect 2964 19790 3016 19796
rect 2976 19514 3004 19790
rect 3547 19612 3855 19632
rect 3547 19610 3553 19612
rect 3609 19610 3633 19612
rect 3689 19610 3713 19612
rect 3769 19610 3793 19612
rect 3849 19610 3855 19612
rect 3609 19558 3611 19610
rect 3791 19558 3793 19610
rect 3547 19556 3553 19558
rect 3609 19556 3633 19558
rect 3689 19556 3713 19558
rect 3769 19556 3793 19558
rect 3849 19556 3855 19558
rect 3547 19536 3855 19556
rect 4080 19514 4108 19858
rect 2964 19508 3016 19514
rect 2964 19450 3016 19456
rect 4068 19508 4120 19514
rect 4068 19450 4120 19456
rect 3240 19236 3292 19242
rect 3240 19178 3292 19184
rect 2688 18964 2740 18970
rect 2688 18906 2740 18912
rect 3252 18902 3280 19178
rect 3240 18896 3292 18902
rect 3240 18838 3292 18844
rect 2044 18692 2096 18698
rect 2044 18634 2096 18640
rect 2780 18692 2832 18698
rect 2780 18634 2832 18640
rect 2136 18624 2188 18630
rect 2136 18566 2188 18572
rect 1676 18080 1728 18086
rect 1676 18022 1728 18028
rect 2044 18080 2096 18086
rect 2044 18022 2096 18028
rect 1688 17610 1716 18022
rect 2056 17814 2084 18022
rect 2044 17808 2096 17814
rect 2044 17750 2096 17756
rect 1676 17604 1728 17610
rect 1676 17546 1728 17552
rect 1584 17536 1636 17542
rect 1584 17478 1636 17484
rect 1596 16726 1624 17478
rect 1688 17338 1716 17546
rect 1676 17332 1728 17338
rect 1676 17274 1728 17280
rect 1584 16720 1636 16726
rect 1584 16662 1636 16668
rect 2148 15910 2176 18566
rect 2596 18080 2648 18086
rect 2596 18022 2648 18028
rect 2248 17980 2556 18000
rect 2248 17978 2254 17980
rect 2310 17978 2334 17980
rect 2390 17978 2414 17980
rect 2470 17978 2494 17980
rect 2550 17978 2556 17980
rect 2310 17926 2312 17978
rect 2492 17926 2494 17978
rect 2248 17924 2254 17926
rect 2310 17924 2334 17926
rect 2390 17924 2414 17926
rect 2470 17924 2494 17926
rect 2550 17924 2556 17926
rect 2248 17904 2556 17924
rect 2608 17882 2636 18022
rect 2596 17876 2648 17882
rect 2596 17818 2648 17824
rect 2608 17746 2636 17818
rect 2596 17740 2648 17746
rect 2596 17682 2648 17688
rect 2594 17096 2650 17105
rect 2594 17031 2596 17040
rect 2648 17031 2650 17040
rect 2596 17002 2648 17008
rect 2248 16892 2556 16912
rect 2248 16890 2254 16892
rect 2310 16890 2334 16892
rect 2390 16890 2414 16892
rect 2470 16890 2494 16892
rect 2550 16890 2556 16892
rect 2310 16838 2312 16890
rect 2492 16838 2494 16890
rect 2248 16836 2254 16838
rect 2310 16836 2334 16838
rect 2390 16836 2414 16838
rect 2470 16836 2494 16838
rect 2550 16836 2556 16838
rect 2248 16816 2556 16836
rect 2608 16794 2636 17002
rect 2596 16788 2648 16794
rect 2596 16730 2648 16736
rect 2596 16448 2648 16454
rect 2596 16390 2648 16396
rect 2608 16250 2636 16390
rect 2596 16244 2648 16250
rect 2596 16186 2648 16192
rect 2688 15972 2740 15978
rect 2688 15914 2740 15920
rect 1952 15904 2004 15910
rect 1952 15846 2004 15852
rect 2136 15904 2188 15910
rect 2136 15846 2188 15852
rect 1964 15366 1992 15846
rect 2248 15804 2556 15824
rect 2248 15802 2254 15804
rect 2310 15802 2334 15804
rect 2390 15802 2414 15804
rect 2470 15802 2494 15804
rect 2550 15802 2556 15804
rect 2310 15750 2312 15802
rect 2492 15750 2494 15802
rect 2248 15748 2254 15750
rect 2310 15748 2334 15750
rect 2390 15748 2414 15750
rect 2470 15748 2494 15750
rect 2550 15748 2556 15750
rect 2248 15728 2556 15748
rect 2700 15706 2728 15914
rect 2688 15700 2740 15706
rect 2688 15642 2740 15648
rect 1860 15360 1912 15366
rect 1860 15302 1912 15308
rect 1952 15360 2004 15366
rect 1952 15302 2004 15308
rect 1872 14822 1900 15302
rect 1860 14816 1912 14822
rect 1860 14758 1912 14764
rect 2596 14816 2648 14822
rect 2596 14758 2648 14764
rect 1584 14272 1636 14278
rect 1584 14214 1636 14220
rect 1596 13938 1624 14214
rect 1584 13932 1636 13938
rect 1584 13874 1636 13880
rect 1584 13728 1636 13734
rect 1584 13670 1636 13676
rect 1596 13190 1624 13670
rect 1768 13524 1820 13530
rect 1768 13466 1820 13472
rect 1584 13184 1636 13190
rect 1584 13126 1636 13132
rect 1596 10033 1624 13126
rect 1780 12986 1808 13466
rect 1768 12980 1820 12986
rect 1768 12922 1820 12928
rect 1872 11642 1900 14758
rect 2248 14716 2556 14736
rect 2248 14714 2254 14716
rect 2310 14714 2334 14716
rect 2390 14714 2414 14716
rect 2470 14714 2494 14716
rect 2550 14714 2556 14716
rect 2310 14662 2312 14714
rect 2492 14662 2494 14714
rect 2248 14660 2254 14662
rect 2310 14660 2334 14662
rect 2390 14660 2414 14662
rect 2470 14660 2494 14662
rect 2550 14660 2556 14662
rect 2248 14640 2556 14660
rect 2608 14346 2636 14758
rect 2596 14340 2648 14346
rect 2596 14282 2648 14288
rect 2248 13628 2556 13648
rect 2248 13626 2254 13628
rect 2310 13626 2334 13628
rect 2390 13626 2414 13628
rect 2470 13626 2494 13628
rect 2550 13626 2556 13628
rect 2310 13574 2312 13626
rect 2492 13574 2494 13626
rect 2248 13572 2254 13574
rect 2310 13572 2334 13574
rect 2390 13572 2414 13574
rect 2470 13572 2494 13574
rect 2550 13572 2556 13574
rect 2248 13552 2556 13572
rect 2412 13252 2464 13258
rect 2412 13194 2464 13200
rect 2424 12986 2452 13194
rect 2412 12980 2464 12986
rect 2412 12922 2464 12928
rect 2248 12540 2556 12560
rect 2248 12538 2254 12540
rect 2310 12538 2334 12540
rect 2390 12538 2414 12540
rect 2470 12538 2494 12540
rect 2550 12538 2556 12540
rect 2310 12486 2312 12538
rect 2492 12486 2494 12538
rect 2248 12484 2254 12486
rect 2310 12484 2334 12486
rect 2390 12484 2414 12486
rect 2470 12484 2494 12486
rect 2550 12484 2556 12486
rect 2248 12464 2556 12484
rect 1952 12096 2004 12102
rect 1952 12038 2004 12044
rect 1780 11614 1900 11642
rect 1676 11552 1728 11558
rect 1676 11494 1728 11500
rect 1688 11150 1716 11494
rect 1676 11144 1728 11150
rect 1676 11086 1728 11092
rect 1582 10024 1638 10033
rect 1582 9959 1638 9968
rect 1492 8832 1544 8838
rect 1492 8774 1544 8780
rect 1504 8634 1532 8774
rect 1492 8628 1544 8634
rect 1492 8570 1544 8576
rect 1492 7948 1544 7954
rect 1492 7890 1544 7896
rect 1504 7002 1532 7890
rect 1780 7313 1808 11614
rect 1860 11552 1912 11558
rect 1860 11494 1912 11500
rect 1872 10470 1900 11494
rect 1964 11082 1992 12038
rect 2248 11452 2556 11472
rect 2248 11450 2254 11452
rect 2310 11450 2334 11452
rect 2390 11450 2414 11452
rect 2470 11450 2494 11452
rect 2550 11450 2556 11452
rect 2310 11398 2312 11450
rect 2492 11398 2494 11450
rect 2248 11396 2254 11398
rect 2310 11396 2334 11398
rect 2390 11396 2414 11398
rect 2470 11396 2494 11398
rect 2550 11396 2556 11398
rect 2248 11376 2556 11396
rect 1952 11076 2004 11082
rect 1952 11018 2004 11024
rect 2136 11008 2188 11014
rect 2136 10950 2188 10956
rect 2044 10532 2096 10538
rect 2044 10474 2096 10480
rect 1860 10464 1912 10470
rect 1860 10406 1912 10412
rect 1952 9376 2004 9382
rect 1952 9318 2004 9324
rect 1860 8084 1912 8090
rect 1860 8026 1912 8032
rect 1766 7304 1822 7313
rect 1766 7239 1822 7248
rect 1492 6996 1544 7002
rect 1492 6938 1544 6944
rect 1676 6316 1728 6322
rect 1676 6258 1728 6264
rect 1584 6112 1636 6118
rect 1584 6054 1636 6060
rect 1596 5681 1624 6054
rect 1582 5672 1638 5681
rect 1582 5607 1638 5616
rect 1400 5160 1452 5166
rect 1398 5128 1400 5137
rect 1452 5128 1454 5137
rect 1398 5063 1454 5072
rect 1688 3126 1716 6258
rect 1872 5370 1900 8026
rect 1860 5364 1912 5370
rect 1860 5306 1912 5312
rect 1860 4072 1912 4078
rect 1860 4014 1912 4020
rect 1872 3738 1900 4014
rect 1860 3732 1912 3738
rect 1860 3674 1912 3680
rect 1676 3120 1728 3126
rect 1676 3062 1728 3068
rect 1964 2854 1992 9318
rect 2056 9178 2084 10474
rect 2148 9926 2176 10950
rect 2248 10364 2556 10384
rect 2248 10362 2254 10364
rect 2310 10362 2334 10364
rect 2390 10362 2414 10364
rect 2470 10362 2494 10364
rect 2550 10362 2556 10364
rect 2310 10310 2312 10362
rect 2492 10310 2494 10362
rect 2248 10308 2254 10310
rect 2310 10308 2334 10310
rect 2390 10308 2414 10310
rect 2470 10308 2494 10310
rect 2550 10308 2556 10310
rect 2248 10288 2556 10308
rect 2608 10169 2636 14282
rect 2688 14272 2740 14278
rect 2688 14214 2740 14220
rect 2700 13734 2728 14214
rect 2688 13728 2740 13734
rect 2688 13670 2740 13676
rect 2700 10577 2728 13670
rect 2792 10713 2820 18634
rect 3547 18524 3855 18544
rect 3547 18522 3553 18524
rect 3609 18522 3633 18524
rect 3689 18522 3713 18524
rect 3769 18522 3793 18524
rect 3849 18522 3855 18524
rect 3609 18470 3611 18522
rect 3791 18470 3793 18522
rect 3547 18468 3553 18470
rect 3609 18468 3633 18470
rect 3689 18468 3713 18470
rect 3769 18468 3793 18470
rect 3849 18468 3855 18470
rect 3547 18448 3855 18468
rect 3976 17876 4028 17882
rect 3976 17818 4028 17824
rect 3988 17678 4016 17818
rect 3976 17672 4028 17678
rect 3976 17614 4028 17620
rect 4080 17513 4108 19450
rect 4066 17504 4122 17513
rect 3547 17436 3855 17456
rect 4066 17439 4122 17448
rect 3547 17434 3553 17436
rect 3609 17434 3633 17436
rect 3689 17434 3713 17436
rect 3769 17434 3793 17436
rect 3849 17434 3855 17436
rect 3609 17382 3611 17434
rect 3791 17382 3793 17434
rect 3547 17380 3553 17382
rect 3609 17380 3633 17382
rect 3689 17380 3713 17382
rect 3769 17380 3793 17382
rect 3849 17380 3855 17382
rect 3547 17360 3855 17380
rect 4080 17202 4108 17439
rect 2872 17196 2924 17202
rect 2872 17138 2924 17144
rect 4068 17196 4120 17202
rect 4068 17138 4120 17144
rect 2884 16794 2912 17138
rect 2872 16788 2924 16794
rect 2872 16730 2924 16736
rect 4068 16652 4120 16658
rect 4068 16594 4120 16600
rect 3976 16584 4028 16590
rect 3976 16526 4028 16532
rect 3884 16516 3936 16522
rect 3884 16458 3936 16464
rect 3547 16348 3855 16368
rect 3547 16346 3553 16348
rect 3609 16346 3633 16348
rect 3689 16346 3713 16348
rect 3769 16346 3793 16348
rect 3849 16346 3855 16348
rect 3609 16294 3611 16346
rect 3791 16294 3793 16346
rect 3547 16292 3553 16294
rect 3609 16292 3633 16294
rect 3689 16292 3713 16294
rect 3769 16292 3793 16294
rect 3849 16292 3855 16294
rect 3547 16272 3855 16292
rect 3896 16250 3924 16458
rect 3988 16250 4016 16526
rect 3884 16244 3936 16250
rect 3884 16186 3936 16192
rect 3976 16244 4028 16250
rect 3976 16186 4028 16192
rect 3516 16176 3568 16182
rect 3516 16118 3568 16124
rect 3528 15910 3556 16118
rect 3148 15904 3200 15910
rect 3148 15846 3200 15852
rect 3516 15904 3568 15910
rect 3516 15846 3568 15852
rect 3160 15638 3188 15846
rect 3148 15632 3200 15638
rect 3148 15574 3200 15580
rect 4080 15570 4108 16594
rect 4068 15564 4120 15570
rect 4068 15506 4120 15512
rect 4172 15450 4200 20318
rect 4252 20256 4304 20262
rect 4252 20198 4304 20204
rect 4264 19514 4292 20198
rect 4846 20156 5154 20176
rect 4846 20154 4852 20156
rect 4908 20154 4932 20156
rect 4988 20154 5012 20156
rect 5068 20154 5092 20156
rect 5148 20154 5154 20156
rect 4908 20102 4910 20154
rect 5090 20102 5092 20154
rect 4846 20100 4852 20102
rect 4908 20100 4932 20102
rect 4988 20100 5012 20102
rect 5068 20100 5092 20102
rect 5148 20100 5154 20102
rect 4846 20080 5154 20100
rect 4344 20052 4396 20058
rect 4344 19994 4396 20000
rect 4252 19508 4304 19514
rect 4252 19450 4304 19456
rect 4356 17270 4384 19994
rect 5540 19848 5592 19854
rect 5540 19790 5592 19796
rect 5552 19378 5580 19790
rect 4436 19372 4488 19378
rect 4436 19314 4488 19320
rect 5540 19372 5592 19378
rect 5540 19314 5592 19320
rect 4448 18902 4476 19314
rect 4712 19304 4764 19310
rect 4712 19246 4764 19252
rect 5632 19304 5684 19310
rect 5828 19281 5856 20402
rect 6460 20324 6512 20330
rect 6460 20266 6512 20272
rect 6000 20256 6052 20262
rect 6000 20198 6052 20204
rect 5632 19246 5684 19252
rect 5814 19272 5870 19281
rect 4436 18896 4488 18902
rect 4436 18838 4488 18844
rect 4436 18760 4488 18766
rect 4436 18702 4488 18708
rect 4448 18290 4476 18702
rect 4724 18426 4752 19246
rect 5540 19168 5592 19174
rect 5540 19110 5592 19116
rect 4846 19068 5154 19088
rect 4846 19066 4852 19068
rect 4908 19066 4932 19068
rect 4988 19066 5012 19068
rect 5068 19066 5092 19068
rect 5148 19066 5154 19068
rect 4908 19014 4910 19066
rect 5090 19014 5092 19066
rect 4846 19012 4852 19014
rect 4908 19012 4932 19014
rect 4988 19012 5012 19014
rect 5068 19012 5092 19014
rect 5148 19012 5154 19014
rect 4846 18992 5154 19012
rect 4712 18420 4764 18426
rect 4712 18362 4764 18368
rect 4620 18352 4672 18358
rect 4620 18294 4672 18300
rect 5172 18352 5224 18358
rect 5552 18306 5580 19110
rect 5172 18294 5224 18300
rect 4436 18284 4488 18290
rect 4436 18226 4488 18232
rect 4632 17746 4660 18294
rect 4846 17980 5154 18000
rect 4846 17978 4852 17980
rect 4908 17978 4932 17980
rect 4988 17978 5012 17980
rect 5068 17978 5092 17980
rect 5148 17978 5154 17980
rect 4908 17926 4910 17978
rect 5090 17926 5092 17978
rect 4846 17924 4852 17926
rect 4908 17924 4932 17926
rect 4988 17924 5012 17926
rect 5068 17924 5092 17926
rect 5148 17924 5154 17926
rect 4846 17904 5154 17924
rect 4528 17740 4580 17746
rect 4528 17682 4580 17688
rect 4620 17740 4672 17746
rect 4620 17682 4672 17688
rect 4804 17740 4856 17746
rect 4804 17682 4856 17688
rect 4434 17640 4490 17649
rect 4540 17626 4568 17682
rect 4816 17626 4844 17682
rect 4540 17598 4844 17626
rect 5080 17604 5132 17610
rect 4434 17575 4436 17584
rect 4488 17575 4490 17584
rect 4436 17546 4488 17552
rect 5080 17546 5132 17552
rect 4804 17536 4856 17542
rect 5092 17513 5120 17546
rect 4804 17478 4856 17484
rect 5078 17504 5134 17513
rect 4816 17338 4844 17478
rect 5078 17439 5134 17448
rect 4804 17332 4856 17338
rect 4804 17274 4856 17280
rect 4344 17264 4396 17270
rect 4344 17206 4396 17212
rect 4436 17264 4488 17270
rect 4436 17206 4488 17212
rect 4356 16658 4384 17206
rect 4344 16652 4396 16658
rect 4344 16594 4396 16600
rect 4448 16590 4476 17206
rect 5184 17134 5212 18294
rect 5460 18278 5580 18306
rect 5356 18148 5408 18154
rect 5356 18090 5408 18096
rect 5368 17678 5396 18090
rect 5356 17672 5408 17678
rect 5262 17640 5318 17649
rect 5356 17614 5408 17620
rect 5262 17575 5264 17584
rect 5316 17575 5318 17584
rect 5264 17546 5316 17552
rect 5172 17128 5224 17134
rect 5356 17128 5408 17134
rect 5172 17070 5224 17076
rect 5354 17096 5356 17105
rect 5408 17096 5410 17105
rect 5354 17031 5410 17040
rect 4846 16892 5154 16912
rect 4846 16890 4852 16892
rect 4908 16890 4932 16892
rect 4988 16890 5012 16892
rect 5068 16890 5092 16892
rect 5148 16890 5154 16892
rect 4908 16838 4910 16890
rect 5090 16838 5092 16890
rect 4846 16836 4852 16838
rect 4908 16836 4932 16838
rect 4988 16836 5012 16838
rect 5068 16836 5092 16838
rect 5148 16836 5154 16838
rect 4846 16816 5154 16836
rect 5460 16810 5488 18278
rect 5540 18216 5592 18222
rect 5540 18158 5592 18164
rect 5552 16998 5580 18158
rect 5644 18086 5672 19246
rect 5724 19236 5776 19242
rect 5814 19207 5870 19216
rect 5724 19178 5776 19184
rect 5736 18766 5764 19178
rect 5816 19168 5868 19174
rect 5816 19110 5868 19116
rect 5724 18760 5776 18766
rect 5724 18702 5776 18708
rect 5828 18426 5856 19110
rect 6012 18834 6040 20198
rect 6472 19786 6500 20266
rect 6564 19922 6592 21490
rect 6644 21412 6696 21418
rect 6644 21354 6696 21360
rect 6656 20466 6684 21354
rect 6748 21146 6776 21519
rect 7288 21412 7340 21418
rect 7288 21354 7340 21360
rect 6736 21140 6788 21146
rect 6736 21082 6788 21088
rect 6748 20942 6776 21082
rect 6736 20936 6788 20942
rect 6736 20878 6788 20884
rect 6828 20936 6880 20942
rect 6828 20878 6880 20884
rect 6644 20460 6696 20466
rect 6644 20402 6696 20408
rect 6552 19916 6604 19922
rect 6552 19858 6604 19864
rect 6460 19780 6512 19786
rect 6460 19722 6512 19728
rect 6144 19612 6452 19632
rect 6144 19610 6150 19612
rect 6206 19610 6230 19612
rect 6286 19610 6310 19612
rect 6366 19610 6390 19612
rect 6446 19610 6452 19612
rect 6206 19558 6208 19610
rect 6388 19558 6390 19610
rect 6144 19556 6150 19558
rect 6206 19556 6230 19558
rect 6286 19556 6310 19558
rect 6366 19556 6390 19558
rect 6446 19556 6452 19558
rect 6144 19536 6452 19556
rect 6564 19446 6592 19858
rect 6644 19780 6696 19786
rect 6644 19722 6696 19728
rect 6552 19440 6604 19446
rect 6090 19408 6146 19417
rect 6552 19382 6604 19388
rect 6090 19343 6146 19352
rect 6000 18828 6052 18834
rect 6000 18770 6052 18776
rect 6104 18714 6132 19343
rect 6656 18902 6684 19722
rect 6748 19378 6776 20878
rect 6840 20806 6868 20878
rect 7012 20868 7064 20874
rect 7012 20810 7064 20816
rect 6828 20800 6880 20806
rect 6828 20742 6880 20748
rect 6840 19854 6868 20742
rect 6828 19848 6880 19854
rect 6828 19790 6880 19796
rect 6826 19680 6882 19689
rect 6826 19615 6882 19624
rect 6736 19372 6788 19378
rect 6736 19314 6788 19320
rect 6840 19258 6868 19615
rect 6748 19230 6868 19258
rect 6644 18896 6696 18902
rect 6644 18838 6696 18844
rect 6012 18686 6132 18714
rect 6552 18760 6604 18766
rect 6552 18702 6604 18708
rect 5816 18420 5868 18426
rect 5816 18362 5868 18368
rect 5724 18284 5776 18290
rect 5724 18226 5776 18232
rect 5632 18080 5684 18086
rect 5632 18022 5684 18028
rect 5736 17898 5764 18226
rect 5644 17870 5764 17898
rect 5828 17882 5856 18362
rect 5908 18080 5960 18086
rect 5908 18022 5960 18028
rect 5816 17876 5868 17882
rect 5644 17202 5672 17870
rect 5816 17818 5868 17824
rect 5632 17196 5684 17202
rect 5632 17138 5684 17144
rect 5540 16992 5592 16998
rect 5540 16934 5592 16940
rect 5460 16782 5580 16810
rect 4436 16584 4488 16590
rect 4436 16526 4488 16532
rect 4528 16584 4580 16590
rect 4528 16526 4580 16532
rect 4540 16114 4568 16526
rect 5552 16522 5580 16782
rect 5540 16516 5592 16522
rect 5540 16458 5592 16464
rect 5644 16182 5672 17138
rect 5828 17105 5856 17818
rect 5814 17096 5870 17105
rect 5814 17031 5870 17040
rect 5920 16674 5948 18022
rect 5736 16646 5948 16674
rect 5736 16590 5764 16646
rect 6012 16590 6040 18686
rect 6144 18524 6452 18544
rect 6144 18522 6150 18524
rect 6206 18522 6230 18524
rect 6286 18522 6310 18524
rect 6366 18522 6390 18524
rect 6446 18522 6452 18524
rect 6206 18470 6208 18522
rect 6388 18470 6390 18522
rect 6144 18468 6150 18470
rect 6206 18468 6230 18470
rect 6286 18468 6310 18470
rect 6366 18468 6390 18470
rect 6446 18468 6452 18470
rect 6144 18448 6452 18468
rect 6144 17436 6452 17456
rect 6144 17434 6150 17436
rect 6206 17434 6230 17436
rect 6286 17434 6310 17436
rect 6366 17434 6390 17436
rect 6446 17434 6452 17436
rect 6206 17382 6208 17434
rect 6388 17382 6390 17434
rect 6144 17380 6150 17382
rect 6206 17380 6230 17382
rect 6286 17380 6310 17382
rect 6366 17380 6390 17382
rect 6446 17380 6452 17382
rect 6144 17360 6452 17380
rect 6368 17196 6420 17202
rect 6368 17138 6420 17144
rect 6380 16590 6408 17138
rect 5724 16584 5776 16590
rect 5724 16526 5776 16532
rect 6000 16584 6052 16590
rect 6000 16526 6052 16532
rect 6368 16584 6420 16590
rect 6368 16526 6420 16532
rect 4712 16176 4764 16182
rect 4712 16118 4764 16124
rect 5632 16176 5684 16182
rect 5632 16118 5684 16124
rect 4528 16108 4580 16114
rect 4528 16050 4580 16056
rect 4620 16108 4672 16114
rect 4620 16050 4672 16056
rect 4172 15422 4476 15450
rect 2872 15360 2924 15366
rect 2872 15302 2924 15308
rect 3056 15360 3108 15366
rect 3056 15302 3108 15308
rect 2884 12986 2912 15302
rect 3068 15162 3096 15302
rect 3547 15260 3855 15280
rect 3547 15258 3553 15260
rect 3609 15258 3633 15260
rect 3689 15258 3713 15260
rect 3769 15258 3793 15260
rect 3849 15258 3855 15260
rect 3609 15206 3611 15258
rect 3791 15206 3793 15258
rect 3547 15204 3553 15206
rect 3609 15204 3633 15206
rect 3689 15204 3713 15206
rect 3769 15204 3793 15206
rect 3849 15204 3855 15206
rect 3547 15184 3855 15204
rect 3056 15156 3108 15162
rect 3056 15098 3108 15104
rect 3608 14816 3660 14822
rect 3608 14758 3660 14764
rect 4252 14816 4304 14822
rect 4252 14758 4304 14764
rect 4344 14816 4396 14822
rect 4344 14758 4396 14764
rect 3620 14550 3648 14758
rect 3608 14544 3660 14550
rect 3608 14486 3660 14492
rect 4264 14482 4292 14758
rect 4252 14476 4304 14482
rect 4252 14418 4304 14424
rect 4356 14414 4384 14758
rect 3884 14408 3936 14414
rect 3884 14350 3936 14356
rect 4344 14408 4396 14414
rect 4344 14350 4396 14356
rect 3547 14172 3855 14192
rect 3547 14170 3553 14172
rect 3609 14170 3633 14172
rect 3689 14170 3713 14172
rect 3769 14170 3793 14172
rect 3849 14170 3855 14172
rect 3609 14118 3611 14170
rect 3791 14118 3793 14170
rect 3547 14116 3553 14118
rect 3609 14116 3633 14118
rect 3689 14116 3713 14118
rect 3769 14116 3793 14118
rect 3849 14116 3855 14118
rect 3547 14096 3855 14116
rect 3896 14074 3924 14350
rect 3884 14068 3936 14074
rect 3884 14010 3936 14016
rect 2964 13932 3016 13938
rect 2964 13874 3016 13880
rect 2872 12980 2924 12986
rect 2872 12922 2924 12928
rect 2976 12866 3004 13874
rect 3056 13184 3108 13190
rect 3108 13132 3188 13138
rect 3056 13126 3188 13132
rect 3068 13110 3188 13126
rect 3054 12880 3110 12889
rect 2976 12838 3054 12866
rect 3054 12815 3110 12824
rect 3068 10810 3096 12815
rect 3160 11898 3188 13110
rect 3547 13084 3855 13104
rect 3547 13082 3553 13084
rect 3609 13082 3633 13084
rect 3689 13082 3713 13084
rect 3769 13082 3793 13084
rect 3849 13082 3855 13084
rect 3609 13030 3611 13082
rect 3791 13030 3793 13082
rect 3547 13028 3553 13030
rect 3609 13028 3633 13030
rect 3689 13028 3713 13030
rect 3769 13028 3793 13030
rect 3849 13028 3855 13030
rect 3547 13008 3855 13028
rect 3700 12844 3752 12850
rect 3700 12786 3752 12792
rect 4252 12844 4304 12850
rect 4252 12786 4304 12792
rect 3712 12374 3740 12786
rect 4160 12640 4212 12646
rect 4160 12582 4212 12588
rect 4172 12442 4200 12582
rect 4160 12436 4212 12442
rect 4160 12378 4212 12384
rect 3700 12368 3752 12374
rect 3700 12310 3752 12316
rect 3884 12096 3936 12102
rect 3884 12038 3936 12044
rect 3547 11996 3855 12016
rect 3547 11994 3553 11996
rect 3609 11994 3633 11996
rect 3689 11994 3713 11996
rect 3769 11994 3793 11996
rect 3849 11994 3855 11996
rect 3609 11942 3611 11994
rect 3791 11942 3793 11994
rect 3547 11940 3553 11942
rect 3609 11940 3633 11942
rect 3689 11940 3713 11942
rect 3769 11940 3793 11942
rect 3849 11940 3855 11942
rect 3547 11920 3855 11940
rect 3148 11892 3200 11898
rect 3148 11834 3200 11840
rect 3240 11688 3292 11694
rect 3240 11630 3292 11636
rect 3252 11354 3280 11630
rect 3896 11354 3924 12038
rect 3976 11892 4028 11898
rect 3976 11834 4028 11840
rect 3240 11348 3292 11354
rect 3240 11290 3292 11296
rect 3884 11348 3936 11354
rect 3884 11290 3936 11296
rect 3988 11218 4016 11834
rect 4264 11762 4292 12786
rect 4344 12708 4396 12714
rect 4344 12650 4396 12656
rect 4252 11756 4304 11762
rect 4252 11698 4304 11704
rect 4160 11620 4212 11626
rect 4160 11562 4212 11568
rect 4172 11286 4200 11562
rect 4160 11280 4212 11286
rect 4160 11222 4212 11228
rect 3976 11212 4028 11218
rect 3976 11154 4028 11160
rect 3547 10908 3855 10928
rect 3547 10906 3553 10908
rect 3609 10906 3633 10908
rect 3689 10906 3713 10908
rect 3769 10906 3793 10908
rect 3849 10906 3855 10908
rect 3609 10854 3611 10906
rect 3791 10854 3793 10906
rect 3547 10852 3553 10854
rect 3609 10852 3633 10854
rect 3689 10852 3713 10854
rect 3769 10852 3793 10854
rect 3849 10852 3855 10854
rect 3547 10832 3855 10852
rect 3056 10804 3108 10810
rect 3056 10746 3108 10752
rect 2778 10704 2834 10713
rect 2778 10639 2834 10648
rect 2686 10568 2742 10577
rect 2686 10503 2742 10512
rect 2780 10464 2832 10470
rect 2780 10406 2832 10412
rect 2792 10266 2820 10406
rect 2780 10260 2832 10266
rect 2780 10202 2832 10208
rect 2594 10160 2650 10169
rect 2594 10095 2650 10104
rect 4172 10062 4200 11222
rect 4356 11218 4384 12650
rect 4448 12434 4476 15422
rect 4540 15094 4568 16050
rect 4632 15434 4660 16050
rect 4724 15502 4752 16118
rect 5540 16040 5592 16046
rect 5540 15982 5592 15988
rect 4846 15804 5154 15824
rect 4846 15802 4852 15804
rect 4908 15802 4932 15804
rect 4988 15802 5012 15804
rect 5068 15802 5092 15804
rect 5148 15802 5154 15804
rect 4908 15750 4910 15802
rect 5090 15750 5092 15802
rect 4846 15748 4852 15750
rect 4908 15748 4932 15750
rect 4988 15748 5012 15750
rect 5068 15748 5092 15750
rect 5148 15748 5154 15750
rect 4846 15728 5154 15748
rect 5552 15502 5580 15982
rect 5736 15706 5764 16526
rect 5908 16516 5960 16522
rect 5908 16458 5960 16464
rect 5724 15700 5776 15706
rect 5724 15642 5776 15648
rect 5736 15609 5764 15642
rect 5722 15600 5778 15609
rect 5920 15586 5948 16458
rect 6012 15910 6040 16526
rect 6144 16348 6452 16368
rect 6144 16346 6150 16348
rect 6206 16346 6230 16348
rect 6286 16346 6310 16348
rect 6366 16346 6390 16348
rect 6446 16346 6452 16348
rect 6206 16294 6208 16346
rect 6388 16294 6390 16346
rect 6144 16292 6150 16294
rect 6206 16292 6230 16294
rect 6286 16292 6310 16294
rect 6366 16292 6390 16294
rect 6446 16292 6452 16294
rect 6144 16272 6452 16292
rect 6564 16289 6592 18702
rect 6748 17202 6776 19230
rect 6828 19168 6880 19174
rect 6828 19110 6880 19116
rect 6840 17377 6868 19110
rect 6920 18284 6972 18290
rect 6920 18226 6972 18232
rect 6932 17678 6960 18226
rect 7024 18222 7052 20810
rect 7196 20460 7248 20466
rect 7196 20402 7248 20408
rect 7208 18970 7236 20402
rect 7300 20262 7328 21354
rect 7443 21244 7751 21264
rect 7443 21242 7449 21244
rect 7505 21242 7529 21244
rect 7585 21242 7609 21244
rect 7665 21242 7689 21244
rect 7745 21242 7751 21244
rect 7505 21190 7507 21242
rect 7687 21190 7689 21242
rect 7443 21188 7449 21190
rect 7505 21188 7529 21190
rect 7585 21188 7609 21190
rect 7665 21188 7689 21190
rect 7745 21188 7751 21190
rect 7443 21168 7751 21188
rect 7852 21078 7880 24754
rect 8114 24304 8170 24313
rect 8114 24239 8116 24248
rect 8168 24239 8170 24248
rect 8116 24210 8168 24216
rect 8128 23730 8156 24210
rect 8220 23769 8248 25230
rect 8206 23760 8262 23769
rect 8116 23724 8168 23730
rect 8206 23695 8262 23704
rect 8116 23666 8168 23672
rect 8116 23112 8168 23118
rect 8116 23054 8168 23060
rect 8128 22681 8156 23054
rect 8114 22672 8170 22681
rect 8114 22607 8116 22616
rect 8168 22607 8170 22616
rect 8116 22578 8168 22584
rect 8114 22128 8170 22137
rect 8114 22063 8170 22072
rect 8128 21350 8156 22063
rect 8116 21344 8168 21350
rect 8116 21286 8168 21292
rect 7840 21072 7892 21078
rect 7840 21014 7892 21020
rect 8022 21040 8078 21049
rect 7288 20256 7340 20262
rect 7288 20198 7340 20204
rect 7300 19854 7328 20198
rect 7443 20156 7751 20176
rect 7443 20154 7449 20156
rect 7505 20154 7529 20156
rect 7585 20154 7609 20156
rect 7665 20154 7689 20156
rect 7745 20154 7751 20156
rect 7505 20102 7507 20154
rect 7687 20102 7689 20154
rect 7443 20100 7449 20102
rect 7505 20100 7529 20102
rect 7585 20100 7609 20102
rect 7665 20100 7689 20102
rect 7745 20100 7751 20102
rect 7443 20080 7751 20100
rect 7288 19848 7340 19854
rect 7288 19790 7340 19796
rect 7852 19310 7880 21014
rect 8022 20975 8078 20984
rect 7840 19304 7892 19310
rect 7840 19246 7892 19252
rect 7443 19068 7751 19088
rect 7443 19066 7449 19068
rect 7505 19066 7529 19068
rect 7585 19066 7609 19068
rect 7665 19066 7689 19068
rect 7745 19066 7751 19068
rect 7505 19014 7507 19066
rect 7687 19014 7689 19066
rect 7443 19012 7449 19014
rect 7505 19012 7529 19014
rect 7585 19012 7609 19014
rect 7665 19012 7689 19014
rect 7745 19012 7751 19014
rect 7443 18992 7751 19012
rect 7196 18964 7248 18970
rect 7196 18906 7248 18912
rect 7208 18766 7236 18906
rect 8036 18834 8064 20975
rect 8128 19854 8156 21286
rect 8206 20496 8262 20505
rect 8206 20431 8262 20440
rect 8116 19848 8168 19854
rect 8116 19790 8168 19796
rect 8024 18828 8076 18834
rect 8024 18770 8076 18776
rect 7196 18760 7248 18766
rect 7196 18702 7248 18708
rect 7288 18760 7340 18766
rect 7288 18702 7340 18708
rect 7104 18692 7156 18698
rect 7104 18634 7156 18640
rect 7012 18216 7064 18222
rect 7012 18158 7064 18164
rect 7024 17814 7052 18158
rect 7012 17808 7064 17814
rect 7012 17750 7064 17756
rect 6920 17672 6972 17678
rect 6920 17614 6972 17620
rect 6826 17368 6882 17377
rect 6826 17303 6882 17312
rect 6736 17196 6788 17202
rect 6736 17138 6788 17144
rect 6736 16720 6788 16726
rect 6736 16662 6788 16668
rect 6550 16280 6606 16289
rect 6550 16215 6606 16224
rect 6000 15904 6052 15910
rect 6000 15846 6052 15852
rect 6012 15706 6040 15846
rect 6000 15700 6052 15706
rect 6000 15642 6052 15648
rect 5920 15558 6040 15586
rect 5722 15535 5778 15544
rect 4712 15496 4764 15502
rect 4712 15438 4764 15444
rect 5540 15496 5592 15502
rect 5540 15438 5592 15444
rect 4620 15428 4672 15434
rect 4620 15370 4672 15376
rect 4528 15088 4580 15094
rect 4528 15030 4580 15036
rect 4724 15026 4752 15438
rect 5632 15428 5684 15434
rect 5632 15370 5684 15376
rect 4712 15020 4764 15026
rect 4712 14962 4764 14968
rect 4724 14770 4752 14962
rect 5540 14952 5592 14958
rect 5540 14894 5592 14900
rect 4632 14742 4752 14770
rect 4528 13252 4580 13258
rect 4528 13194 4580 13200
rect 4540 12918 4568 13194
rect 4528 12912 4580 12918
rect 4528 12854 4580 12860
rect 4448 12406 4568 12434
rect 4344 11212 4396 11218
rect 4344 11154 4396 11160
rect 4344 10600 4396 10606
rect 4344 10542 4396 10548
rect 2872 10056 2924 10062
rect 2872 9998 2924 10004
rect 4160 10056 4212 10062
rect 4160 9998 4212 10004
rect 2136 9920 2188 9926
rect 2136 9862 2188 9868
rect 2596 9920 2648 9926
rect 2596 9862 2648 9868
rect 2248 9276 2556 9296
rect 2248 9274 2254 9276
rect 2310 9274 2334 9276
rect 2390 9274 2414 9276
rect 2470 9274 2494 9276
rect 2550 9274 2556 9276
rect 2310 9222 2312 9274
rect 2492 9222 2494 9274
rect 2248 9220 2254 9222
rect 2310 9220 2334 9222
rect 2390 9220 2414 9222
rect 2470 9220 2494 9222
rect 2550 9220 2556 9222
rect 2248 9200 2556 9220
rect 2044 9172 2096 9178
rect 2044 9114 2096 9120
rect 2056 8922 2084 9114
rect 2056 8894 2176 8922
rect 2044 8832 2096 8838
rect 2044 8774 2096 8780
rect 2056 8090 2084 8774
rect 2044 8084 2096 8090
rect 2044 8026 2096 8032
rect 2044 7200 2096 7206
rect 2044 7142 2096 7148
rect 2056 6798 2084 7142
rect 2148 6914 2176 8894
rect 2248 8188 2556 8208
rect 2248 8186 2254 8188
rect 2310 8186 2334 8188
rect 2390 8186 2414 8188
rect 2470 8186 2494 8188
rect 2550 8186 2556 8188
rect 2310 8134 2312 8186
rect 2492 8134 2494 8186
rect 2248 8132 2254 8134
rect 2310 8132 2334 8134
rect 2390 8132 2414 8134
rect 2470 8132 2494 8134
rect 2550 8132 2556 8134
rect 2248 8112 2556 8132
rect 2608 7970 2636 9862
rect 2516 7942 2636 7970
rect 2412 7880 2464 7886
rect 2412 7822 2464 7828
rect 2424 7274 2452 7822
rect 2516 7290 2544 7942
rect 2596 7744 2648 7750
rect 2596 7686 2648 7692
rect 2608 7478 2636 7686
rect 2596 7472 2648 7478
rect 2596 7414 2648 7420
rect 2412 7268 2464 7274
rect 2516 7262 2636 7290
rect 2412 7210 2464 7216
rect 2248 7100 2556 7120
rect 2248 7098 2254 7100
rect 2310 7098 2334 7100
rect 2390 7098 2414 7100
rect 2470 7098 2494 7100
rect 2550 7098 2556 7100
rect 2310 7046 2312 7098
rect 2492 7046 2494 7098
rect 2248 7044 2254 7046
rect 2310 7044 2334 7046
rect 2390 7044 2414 7046
rect 2470 7044 2494 7046
rect 2550 7044 2556 7046
rect 2248 7024 2556 7044
rect 2608 7018 2636 7262
rect 2608 6990 2728 7018
rect 2148 6886 2636 6914
rect 2608 6798 2636 6886
rect 2044 6792 2096 6798
rect 2044 6734 2096 6740
rect 2596 6792 2648 6798
rect 2596 6734 2648 6740
rect 2608 6225 2636 6734
rect 2594 6216 2650 6225
rect 2594 6151 2650 6160
rect 2136 6112 2188 6118
rect 2136 6054 2188 6060
rect 2148 5778 2176 6054
rect 2248 6012 2556 6032
rect 2248 6010 2254 6012
rect 2310 6010 2334 6012
rect 2390 6010 2414 6012
rect 2470 6010 2494 6012
rect 2550 6010 2556 6012
rect 2310 5958 2312 6010
rect 2492 5958 2494 6010
rect 2248 5956 2254 5958
rect 2310 5956 2334 5958
rect 2390 5956 2414 5958
rect 2470 5956 2494 5958
rect 2550 5956 2556 5958
rect 2248 5936 2556 5956
rect 2136 5772 2188 5778
rect 2136 5714 2188 5720
rect 2044 5704 2096 5710
rect 2044 5646 2096 5652
rect 2056 4690 2084 5646
rect 2700 5080 2728 6990
rect 2780 5228 2832 5234
rect 2780 5170 2832 5176
rect 2792 5080 2820 5170
rect 2700 5052 2820 5080
rect 2248 4924 2556 4944
rect 2248 4922 2254 4924
rect 2310 4922 2334 4924
rect 2390 4922 2414 4924
rect 2470 4922 2494 4924
rect 2550 4922 2556 4924
rect 2310 4870 2312 4922
rect 2492 4870 2494 4922
rect 2248 4868 2254 4870
rect 2310 4868 2334 4870
rect 2390 4868 2414 4870
rect 2470 4868 2494 4870
rect 2550 4868 2556 4870
rect 2248 4848 2556 4868
rect 2044 4684 2096 4690
rect 2044 4626 2096 4632
rect 2056 3738 2084 4626
rect 2780 4616 2832 4622
rect 2780 4558 2832 4564
rect 2596 4548 2648 4554
rect 2596 4490 2648 4496
rect 2248 3836 2556 3856
rect 2248 3834 2254 3836
rect 2310 3834 2334 3836
rect 2390 3834 2414 3836
rect 2470 3834 2494 3836
rect 2550 3834 2556 3836
rect 2310 3782 2312 3834
rect 2492 3782 2494 3834
rect 2248 3780 2254 3782
rect 2310 3780 2334 3782
rect 2390 3780 2414 3782
rect 2470 3780 2494 3782
rect 2550 3780 2556 3782
rect 2248 3760 2556 3780
rect 2044 3732 2096 3738
rect 2044 3674 2096 3680
rect 940 2848 992 2854
rect 940 2790 992 2796
rect 1952 2848 2004 2854
rect 1952 2790 2004 2796
rect 952 800 980 2790
rect 2248 2748 2556 2768
rect 2248 2746 2254 2748
rect 2310 2746 2334 2748
rect 2390 2746 2414 2748
rect 2470 2746 2494 2748
rect 2550 2746 2556 2748
rect 2310 2694 2312 2746
rect 2492 2694 2494 2746
rect 2248 2692 2254 2694
rect 2310 2692 2334 2694
rect 2390 2692 2414 2694
rect 2470 2692 2494 2694
rect 2550 2692 2556 2694
rect 2248 2672 2556 2692
rect 2608 2650 2636 4490
rect 2792 3942 2820 4558
rect 2780 3936 2832 3942
rect 2780 3878 2832 3884
rect 2688 3460 2740 3466
rect 2688 3402 2740 3408
rect 2700 3058 2728 3402
rect 2884 3194 2912 9998
rect 3056 9988 3108 9994
rect 3056 9930 3108 9936
rect 4252 9988 4304 9994
rect 4252 9930 4304 9936
rect 2964 5364 3016 5370
rect 2964 5306 3016 5312
rect 2976 4486 3004 5306
rect 2964 4480 3016 4486
rect 2964 4422 3016 4428
rect 2872 3188 2924 3194
rect 2872 3130 2924 3136
rect 2688 3052 2740 3058
rect 2688 2994 2740 3000
rect 2596 2644 2648 2650
rect 2596 2586 2648 2592
rect 1860 2304 1912 2310
rect 1860 2246 1912 2252
rect 1872 2106 1900 2246
rect 1860 2100 1912 2106
rect 1860 2042 1912 2048
rect 2884 800 2912 3130
rect 3068 2378 3096 9930
rect 3547 9820 3855 9840
rect 3547 9818 3553 9820
rect 3609 9818 3633 9820
rect 3689 9818 3713 9820
rect 3769 9818 3793 9820
rect 3849 9818 3855 9820
rect 3609 9766 3611 9818
rect 3791 9766 3793 9818
rect 3547 9764 3553 9766
rect 3609 9764 3633 9766
rect 3689 9764 3713 9766
rect 3769 9764 3793 9766
rect 3849 9764 3855 9766
rect 3547 9744 3855 9764
rect 4264 9722 4292 9930
rect 4252 9716 4304 9722
rect 4252 9658 4304 9664
rect 4356 9586 4384 10542
rect 4436 10260 4488 10266
rect 4436 10202 4488 10208
rect 4448 9722 4476 10202
rect 4436 9716 4488 9722
rect 4436 9658 4488 9664
rect 4540 9586 4568 12406
rect 4632 10810 4660 14742
rect 4846 14716 5154 14736
rect 4846 14714 4852 14716
rect 4908 14714 4932 14716
rect 4988 14714 5012 14716
rect 5068 14714 5092 14716
rect 5148 14714 5154 14716
rect 4908 14662 4910 14714
rect 5090 14662 5092 14714
rect 4846 14660 4852 14662
rect 4908 14660 4932 14662
rect 4988 14660 5012 14662
rect 5068 14660 5092 14662
rect 5148 14660 5154 14662
rect 4846 14640 5154 14660
rect 5172 14476 5224 14482
rect 5172 14418 5224 14424
rect 4804 14340 4856 14346
rect 4804 14282 4856 14288
rect 4816 13938 4844 14282
rect 5184 14074 5212 14418
rect 5552 14414 5580 14894
rect 5540 14408 5592 14414
rect 5540 14350 5592 14356
rect 5448 14272 5500 14278
rect 5448 14214 5500 14220
rect 5172 14068 5224 14074
rect 5172 14010 5224 14016
rect 5262 13968 5318 13977
rect 4804 13932 4856 13938
rect 5262 13903 5318 13912
rect 5356 13932 5408 13938
rect 4804 13874 4856 13880
rect 4712 13728 4764 13734
rect 4712 13670 4764 13676
rect 4724 12434 4752 13670
rect 4846 13628 5154 13648
rect 4846 13626 4852 13628
rect 4908 13626 4932 13628
rect 4988 13626 5012 13628
rect 5068 13626 5092 13628
rect 5148 13626 5154 13628
rect 4908 13574 4910 13626
rect 5090 13574 5092 13626
rect 4846 13572 4852 13574
rect 4908 13572 4932 13574
rect 4988 13572 5012 13574
rect 5068 13572 5092 13574
rect 5148 13572 5154 13574
rect 4846 13552 5154 13572
rect 4846 12540 5154 12560
rect 4846 12538 4852 12540
rect 4908 12538 4932 12540
rect 4988 12538 5012 12540
rect 5068 12538 5092 12540
rect 5148 12538 5154 12540
rect 4908 12486 4910 12538
rect 5090 12486 5092 12538
rect 4846 12484 4852 12486
rect 4908 12484 4932 12486
rect 4988 12484 5012 12486
rect 5068 12484 5092 12486
rect 5148 12484 5154 12486
rect 4846 12464 5154 12484
rect 4724 12406 5212 12434
rect 4712 12368 4764 12374
rect 4712 12310 4764 12316
rect 4724 11082 4752 12310
rect 4846 11452 5154 11472
rect 4846 11450 4852 11452
rect 4908 11450 4932 11452
rect 4988 11450 5012 11452
rect 5068 11450 5092 11452
rect 5148 11450 5154 11452
rect 4908 11398 4910 11450
rect 5090 11398 5092 11450
rect 4846 11396 4852 11398
rect 4908 11396 4932 11398
rect 4988 11396 5012 11398
rect 5068 11396 5092 11398
rect 5148 11396 5154 11398
rect 4846 11376 5154 11396
rect 4712 11076 4764 11082
rect 4712 11018 4764 11024
rect 4620 10804 4672 10810
rect 4620 10746 4672 10752
rect 4712 10668 4764 10674
rect 4712 10610 4764 10616
rect 4620 10532 4672 10538
rect 4620 10474 4672 10480
rect 4344 9580 4396 9586
rect 4344 9522 4396 9528
rect 4528 9580 4580 9586
rect 4528 9522 4580 9528
rect 4160 9512 4212 9518
rect 4160 9454 4212 9460
rect 3884 9376 3936 9382
rect 3884 9318 3936 9324
rect 3148 8900 3200 8906
rect 3148 8842 3200 8848
rect 3160 8634 3188 8842
rect 3547 8732 3855 8752
rect 3547 8730 3553 8732
rect 3609 8730 3633 8732
rect 3689 8730 3713 8732
rect 3769 8730 3793 8732
rect 3849 8730 3855 8732
rect 3609 8678 3611 8730
rect 3791 8678 3793 8730
rect 3547 8676 3553 8678
rect 3609 8676 3633 8678
rect 3689 8676 3713 8678
rect 3769 8676 3793 8678
rect 3849 8676 3855 8678
rect 3547 8656 3855 8676
rect 3148 8628 3200 8634
rect 3148 8570 3200 8576
rect 3896 8566 3924 9318
rect 4172 9178 4200 9454
rect 4160 9172 4212 9178
rect 4160 9114 4212 9120
rect 4540 8974 4568 9522
rect 4632 9518 4660 10474
rect 4724 10266 4752 10610
rect 4846 10364 5154 10384
rect 4846 10362 4852 10364
rect 4908 10362 4932 10364
rect 4988 10362 5012 10364
rect 5068 10362 5092 10364
rect 5148 10362 5154 10364
rect 4908 10310 4910 10362
rect 5090 10310 5092 10362
rect 4846 10308 4852 10310
rect 4908 10308 4932 10310
rect 4988 10308 5012 10310
rect 5068 10308 5092 10310
rect 5148 10308 5154 10310
rect 4846 10288 5154 10308
rect 4712 10260 4764 10266
rect 4712 10202 4764 10208
rect 4620 9512 4672 9518
rect 4620 9454 4672 9460
rect 4528 8968 4580 8974
rect 4528 8910 4580 8916
rect 4252 8832 4304 8838
rect 4252 8774 4304 8780
rect 3884 8560 3936 8566
rect 3884 8502 3936 8508
rect 4160 8492 4212 8498
rect 4160 8434 4212 8440
rect 3884 8424 3936 8430
rect 3884 8366 3936 8372
rect 3424 8016 3476 8022
rect 3424 7958 3476 7964
rect 3240 7744 3292 7750
rect 3240 7686 3292 7692
rect 3252 6866 3280 7686
rect 3240 6860 3292 6866
rect 3240 6802 3292 6808
rect 3332 6860 3384 6866
rect 3332 6802 3384 6808
rect 3344 6746 3372 6802
rect 3252 6718 3372 6746
rect 3252 6458 3280 6718
rect 3240 6452 3292 6458
rect 3240 6394 3292 6400
rect 3436 5137 3464 7958
rect 3547 7644 3855 7664
rect 3547 7642 3553 7644
rect 3609 7642 3633 7644
rect 3689 7642 3713 7644
rect 3769 7642 3793 7644
rect 3849 7642 3855 7644
rect 3609 7590 3611 7642
rect 3791 7590 3793 7642
rect 3547 7588 3553 7590
rect 3609 7588 3633 7590
rect 3689 7588 3713 7590
rect 3769 7588 3793 7590
rect 3849 7588 3855 7590
rect 3547 7568 3855 7588
rect 3792 7336 3844 7342
rect 3790 7304 3792 7313
rect 3844 7304 3846 7313
rect 3790 7239 3846 7248
rect 3547 6556 3855 6576
rect 3547 6554 3553 6556
rect 3609 6554 3633 6556
rect 3689 6554 3713 6556
rect 3769 6554 3793 6556
rect 3849 6554 3855 6556
rect 3609 6502 3611 6554
rect 3791 6502 3793 6554
rect 3547 6500 3553 6502
rect 3609 6500 3633 6502
rect 3689 6500 3713 6502
rect 3769 6500 3793 6502
rect 3849 6500 3855 6502
rect 3547 6480 3855 6500
rect 3547 5468 3855 5488
rect 3547 5466 3553 5468
rect 3609 5466 3633 5468
rect 3689 5466 3713 5468
rect 3769 5466 3793 5468
rect 3849 5466 3855 5468
rect 3609 5414 3611 5466
rect 3791 5414 3793 5466
rect 3547 5412 3553 5414
rect 3609 5412 3633 5414
rect 3689 5412 3713 5414
rect 3769 5412 3793 5414
rect 3849 5412 3855 5414
rect 3547 5392 3855 5412
rect 3792 5296 3844 5302
rect 3792 5238 3844 5244
rect 3422 5128 3478 5137
rect 3422 5063 3478 5072
rect 3436 3602 3464 5063
rect 3804 4706 3832 5238
rect 3896 5030 3924 8366
rect 3976 8288 4028 8294
rect 3976 8230 4028 8236
rect 3988 7750 4016 8230
rect 3976 7744 4028 7750
rect 3976 7686 4028 7692
rect 3988 7342 4016 7686
rect 4068 7472 4120 7478
rect 4068 7414 4120 7420
rect 3976 7336 4028 7342
rect 3976 7278 4028 7284
rect 4080 7290 4108 7414
rect 4172 7410 4200 8434
rect 4264 7478 4292 8774
rect 4528 8424 4580 8430
rect 4528 8366 4580 8372
rect 4540 8022 4568 8366
rect 4528 8016 4580 8022
rect 4528 7958 4580 7964
rect 4528 7880 4580 7886
rect 4528 7822 4580 7828
rect 4344 7812 4396 7818
rect 4344 7754 4396 7760
rect 4436 7812 4488 7818
rect 4436 7754 4488 7760
rect 4252 7472 4304 7478
rect 4252 7414 4304 7420
rect 4160 7404 4212 7410
rect 4160 7346 4212 7352
rect 3988 7154 4016 7278
rect 4080 7262 4200 7290
rect 3988 7126 4108 7154
rect 3884 5024 3936 5030
rect 3884 4966 3936 4972
rect 3804 4678 4016 4706
rect 3988 4622 4016 4678
rect 3976 4616 4028 4622
rect 3976 4558 4028 4564
rect 3547 4380 3855 4400
rect 3547 4378 3553 4380
rect 3609 4378 3633 4380
rect 3689 4378 3713 4380
rect 3769 4378 3793 4380
rect 3849 4378 3855 4380
rect 3609 4326 3611 4378
rect 3791 4326 3793 4378
rect 3547 4324 3553 4326
rect 3609 4324 3633 4326
rect 3689 4324 3713 4326
rect 3769 4324 3793 4326
rect 3849 4324 3855 4326
rect 3547 4304 3855 4324
rect 3976 3936 4028 3942
rect 3976 3878 4028 3884
rect 3424 3596 3476 3602
rect 3424 3538 3476 3544
rect 3547 3292 3855 3312
rect 3547 3290 3553 3292
rect 3609 3290 3633 3292
rect 3689 3290 3713 3292
rect 3769 3290 3793 3292
rect 3849 3290 3855 3292
rect 3609 3238 3611 3290
rect 3791 3238 3793 3290
rect 3547 3236 3553 3238
rect 3609 3236 3633 3238
rect 3689 3236 3713 3238
rect 3769 3236 3793 3238
rect 3849 3236 3855 3238
rect 3547 3216 3855 3236
rect 3608 2916 3660 2922
rect 3608 2858 3660 2864
rect 3620 2446 3648 2858
rect 3884 2848 3936 2854
rect 3884 2790 3936 2796
rect 3896 2514 3924 2790
rect 3884 2508 3936 2514
rect 3884 2450 3936 2456
rect 3608 2440 3660 2446
rect 3608 2382 3660 2388
rect 3988 2378 4016 3878
rect 3056 2372 3108 2378
rect 3056 2314 3108 2320
rect 3976 2372 4028 2378
rect 3976 2314 4028 2320
rect 3068 1766 3096 2314
rect 3148 2304 3200 2310
rect 3148 2246 3200 2252
rect 3160 2106 3188 2246
rect 3547 2204 3855 2224
rect 3547 2202 3553 2204
rect 3609 2202 3633 2204
rect 3689 2202 3713 2204
rect 3769 2202 3793 2204
rect 3849 2202 3855 2204
rect 3609 2150 3611 2202
rect 3791 2150 3793 2202
rect 3547 2148 3553 2150
rect 3609 2148 3633 2150
rect 3689 2148 3713 2150
rect 3769 2148 3793 2150
rect 3849 2148 3855 2150
rect 3547 2128 3855 2148
rect 3148 2100 3200 2106
rect 3148 2042 3200 2048
rect 3056 1760 3108 1766
rect 3056 1702 3108 1708
rect 4080 1358 4108 7126
rect 4172 6202 4200 7262
rect 4264 7206 4292 7414
rect 4252 7200 4304 7206
rect 4252 7142 4304 7148
rect 4264 6798 4292 7142
rect 4252 6792 4304 6798
rect 4252 6734 4304 6740
rect 4356 6662 4384 7754
rect 4448 7478 4476 7754
rect 4436 7472 4488 7478
rect 4436 7414 4488 7420
rect 4436 6996 4488 7002
rect 4436 6938 4488 6944
rect 4344 6656 4396 6662
rect 4344 6598 4396 6604
rect 4172 6174 4384 6202
rect 4172 5642 4200 6174
rect 4356 6118 4384 6174
rect 4252 6112 4304 6118
rect 4252 6054 4304 6060
rect 4344 6112 4396 6118
rect 4344 6054 4396 6060
rect 4160 5636 4212 5642
rect 4160 5578 4212 5584
rect 4160 4548 4212 4554
rect 4160 4490 4212 4496
rect 4172 4282 4200 4490
rect 4160 4276 4212 4282
rect 4160 4218 4212 4224
rect 4172 4078 4200 4218
rect 4160 4072 4212 4078
rect 4160 4014 4212 4020
rect 4264 2378 4292 6054
rect 4448 5794 4476 6938
rect 4540 6662 4568 7822
rect 4528 6656 4580 6662
rect 4528 6598 4580 6604
rect 4528 6248 4580 6254
rect 4528 6190 4580 6196
rect 4356 5766 4476 5794
rect 4356 4706 4384 5766
rect 4436 5636 4488 5642
rect 4436 5578 4488 5584
rect 4448 5370 4476 5578
rect 4540 5370 4568 6190
rect 4436 5364 4488 5370
rect 4436 5306 4488 5312
rect 4528 5364 4580 5370
rect 4528 5306 4580 5312
rect 4436 5024 4488 5030
rect 4436 4966 4488 4972
rect 4448 4842 4476 4966
rect 4448 4814 4568 4842
rect 4356 4678 4476 4706
rect 4344 4480 4396 4486
rect 4344 4422 4396 4428
rect 4356 3670 4384 4422
rect 4448 4146 4476 4678
rect 4540 4622 4568 4814
rect 4528 4616 4580 4622
rect 4528 4558 4580 4564
rect 4540 4282 4568 4558
rect 4528 4276 4580 4282
rect 4528 4218 4580 4224
rect 4436 4140 4488 4146
rect 4436 4082 4488 4088
rect 4344 3664 4396 3670
rect 4344 3606 4396 3612
rect 4448 3534 4476 4082
rect 4528 3596 4580 3602
rect 4528 3538 4580 3544
rect 4436 3528 4488 3534
rect 4436 3470 4488 3476
rect 4344 3188 4396 3194
rect 4344 3130 4396 3136
rect 4356 2446 4384 3130
rect 4448 2922 4476 3470
rect 4436 2916 4488 2922
rect 4436 2858 4488 2864
rect 4344 2440 4396 2446
rect 4344 2382 4396 2388
rect 4540 2378 4568 3538
rect 4252 2372 4304 2378
rect 4252 2314 4304 2320
rect 4528 2372 4580 2378
rect 4528 2314 4580 2320
rect 4068 1352 4120 1358
rect 4068 1294 4120 1300
rect 938 0 994 800
rect 2870 0 2926 800
rect 4632 762 4660 9454
rect 4846 9276 5154 9296
rect 4846 9274 4852 9276
rect 4908 9274 4932 9276
rect 4988 9274 5012 9276
rect 5068 9274 5092 9276
rect 5148 9274 5154 9276
rect 4908 9222 4910 9274
rect 5090 9222 5092 9274
rect 4846 9220 4852 9222
rect 4908 9220 4932 9222
rect 4988 9220 5012 9222
rect 5068 9220 5092 9222
rect 5148 9220 5154 9222
rect 4846 9200 5154 9220
rect 4712 8560 4764 8566
rect 4712 8502 4764 8508
rect 4724 7002 4752 8502
rect 4846 8188 5154 8208
rect 4846 8186 4852 8188
rect 4908 8186 4932 8188
rect 4988 8186 5012 8188
rect 5068 8186 5092 8188
rect 5148 8186 5154 8188
rect 4908 8134 4910 8186
rect 5090 8134 5092 8186
rect 4846 8132 4852 8134
rect 4908 8132 4932 8134
rect 4988 8132 5012 8134
rect 5068 8132 5092 8134
rect 5148 8132 5154 8134
rect 4846 8112 5154 8132
rect 5184 8022 5212 12406
rect 5276 11762 5304 13903
rect 5356 13874 5408 13880
rect 5368 12306 5396 13874
rect 5460 13326 5488 14214
rect 5644 14006 5672 15370
rect 5736 15026 5764 15535
rect 5724 15020 5776 15026
rect 5724 14962 5776 14968
rect 5724 14544 5776 14550
rect 5724 14486 5776 14492
rect 5814 14512 5870 14521
rect 5736 14414 5764 14486
rect 5814 14447 5870 14456
rect 5724 14408 5776 14414
rect 5724 14350 5776 14356
rect 5736 14278 5764 14350
rect 5724 14272 5776 14278
rect 5724 14214 5776 14220
rect 5632 14000 5684 14006
rect 5632 13942 5684 13948
rect 5540 13864 5592 13870
rect 5540 13806 5592 13812
rect 5448 13320 5500 13326
rect 5448 13262 5500 13268
rect 5460 12442 5488 13262
rect 5448 12436 5500 12442
rect 5448 12378 5500 12384
rect 5356 12300 5408 12306
rect 5356 12242 5408 12248
rect 5264 11756 5316 11762
rect 5264 11698 5316 11704
rect 5276 11150 5304 11698
rect 5368 11286 5396 12242
rect 5460 12238 5488 12378
rect 5552 12374 5580 13806
rect 5828 13530 5856 14447
rect 6012 13988 6040 15558
rect 6644 15496 6696 15502
rect 6644 15438 6696 15444
rect 6552 15428 6604 15434
rect 6552 15370 6604 15376
rect 6144 15260 6452 15280
rect 6144 15258 6150 15260
rect 6206 15258 6230 15260
rect 6286 15258 6310 15260
rect 6366 15258 6390 15260
rect 6446 15258 6452 15260
rect 6206 15206 6208 15258
rect 6388 15206 6390 15258
rect 6144 15204 6150 15206
rect 6206 15204 6230 15206
rect 6286 15204 6310 15206
rect 6366 15204 6390 15206
rect 6446 15204 6452 15206
rect 6144 15184 6452 15204
rect 6092 15020 6144 15026
rect 6092 14962 6144 14968
rect 6104 14890 6132 14962
rect 6564 14958 6592 15370
rect 6656 15201 6684 15438
rect 6642 15192 6698 15201
rect 6748 15162 6776 16662
rect 7116 16454 7144 18634
rect 7208 18465 7236 18702
rect 7194 18456 7250 18465
rect 7194 18391 7250 18400
rect 7196 17672 7248 17678
rect 7196 17614 7248 17620
rect 7208 17066 7236 17614
rect 7196 17060 7248 17066
rect 7196 17002 7248 17008
rect 7104 16448 7156 16454
rect 7104 16390 7156 16396
rect 7208 16182 7236 17002
rect 7300 16794 7328 18702
rect 7840 18284 7892 18290
rect 7840 18226 7892 18232
rect 7443 17980 7751 18000
rect 7443 17978 7449 17980
rect 7505 17978 7529 17980
rect 7585 17978 7609 17980
rect 7665 17978 7689 17980
rect 7745 17978 7751 17980
rect 7505 17926 7507 17978
rect 7687 17926 7689 17978
rect 7443 17924 7449 17926
rect 7505 17924 7529 17926
rect 7585 17924 7609 17926
rect 7665 17924 7689 17926
rect 7745 17924 7751 17926
rect 7443 17904 7751 17924
rect 7852 17921 7880 18226
rect 7838 17912 7894 17921
rect 7838 17847 7894 17856
rect 7932 17604 7984 17610
rect 7932 17546 7984 17552
rect 7840 17196 7892 17202
rect 7840 17138 7892 17144
rect 7443 16892 7751 16912
rect 7443 16890 7449 16892
rect 7505 16890 7529 16892
rect 7585 16890 7609 16892
rect 7665 16890 7689 16892
rect 7745 16890 7751 16892
rect 7505 16838 7507 16890
rect 7687 16838 7689 16890
rect 7443 16836 7449 16838
rect 7505 16836 7529 16838
rect 7585 16836 7609 16838
rect 7665 16836 7689 16838
rect 7745 16836 7751 16838
rect 7443 16816 7751 16836
rect 7288 16788 7340 16794
rect 7288 16730 7340 16736
rect 7300 16182 7328 16730
rect 7852 16522 7880 17138
rect 7840 16516 7892 16522
rect 7840 16458 7892 16464
rect 7196 16176 7248 16182
rect 7196 16118 7248 16124
rect 7288 16176 7340 16182
rect 7288 16118 7340 16124
rect 7012 16108 7064 16114
rect 7012 16050 7064 16056
rect 7024 15638 7052 16050
rect 7443 15804 7751 15824
rect 7443 15802 7449 15804
rect 7505 15802 7529 15804
rect 7585 15802 7609 15804
rect 7665 15802 7689 15804
rect 7745 15802 7751 15804
rect 7505 15750 7507 15802
rect 7687 15750 7689 15802
rect 7443 15748 7449 15750
rect 7505 15748 7529 15750
rect 7585 15748 7609 15750
rect 7665 15748 7689 15750
rect 7745 15748 7751 15750
rect 7443 15728 7751 15748
rect 7852 15638 7880 16458
rect 7944 15994 7972 17546
rect 8036 16114 8064 18770
rect 8220 18290 8248 20431
rect 8208 18284 8260 18290
rect 8208 18226 8260 18232
rect 8220 17678 8248 18226
rect 8208 17672 8260 17678
rect 8208 17614 8260 17620
rect 8024 16108 8076 16114
rect 8024 16050 8076 16056
rect 7944 15966 8064 15994
rect 7012 15632 7064 15638
rect 7012 15574 7064 15580
rect 7840 15632 7892 15638
rect 7840 15574 7892 15580
rect 6642 15127 6698 15136
rect 6736 15156 6788 15162
rect 6736 15098 6788 15104
rect 6552 14952 6604 14958
rect 6552 14894 6604 14900
rect 6828 14952 6880 14958
rect 6828 14894 6880 14900
rect 6092 14884 6144 14890
rect 6092 14826 6144 14832
rect 6104 14414 6132 14826
rect 6840 14804 6868 14894
rect 6748 14776 6868 14804
rect 6092 14408 6144 14414
rect 6092 14350 6144 14356
rect 6144 14172 6452 14192
rect 6144 14170 6150 14172
rect 6206 14170 6230 14172
rect 6286 14170 6310 14172
rect 6366 14170 6390 14172
rect 6446 14170 6452 14172
rect 6206 14118 6208 14170
rect 6388 14118 6390 14170
rect 6144 14116 6150 14118
rect 6206 14116 6230 14118
rect 6286 14116 6310 14118
rect 6366 14116 6390 14118
rect 6446 14116 6452 14118
rect 6144 14096 6452 14116
rect 6012 13960 6132 13988
rect 6104 13530 6132 13960
rect 5816 13524 5868 13530
rect 5816 13466 5868 13472
rect 6092 13524 6144 13530
rect 6092 13466 6144 13472
rect 5828 13326 5856 13466
rect 6000 13456 6052 13462
rect 6000 13398 6052 13404
rect 5816 13320 5868 13326
rect 5816 13262 5868 13268
rect 5632 12980 5684 12986
rect 5632 12922 5684 12928
rect 5540 12368 5592 12374
rect 5540 12310 5592 12316
rect 5448 12232 5500 12238
rect 5448 12174 5500 12180
rect 5540 11824 5592 11830
rect 5540 11766 5592 11772
rect 5448 11552 5500 11558
rect 5448 11494 5500 11500
rect 5356 11280 5408 11286
rect 5356 11222 5408 11228
rect 5460 11218 5488 11494
rect 5448 11212 5500 11218
rect 5448 11154 5500 11160
rect 5264 11144 5316 11150
rect 5264 11086 5316 11092
rect 5552 10810 5580 11766
rect 5540 10804 5592 10810
rect 5540 10746 5592 10752
rect 5644 10690 5672 12922
rect 5828 12782 5856 13262
rect 5816 12776 5868 12782
rect 5816 12718 5868 12724
rect 5816 12232 5868 12238
rect 5816 12174 5868 12180
rect 5828 11082 5856 12174
rect 5908 12164 5960 12170
rect 5908 12106 5960 12112
rect 5816 11076 5868 11082
rect 5816 11018 5868 11024
rect 5814 10704 5870 10713
rect 5644 10662 5764 10690
rect 5448 10532 5500 10538
rect 5448 10474 5500 10480
rect 5460 9926 5488 10474
rect 5630 10160 5686 10169
rect 5630 10095 5686 10104
rect 5540 9988 5592 9994
rect 5540 9930 5592 9936
rect 5448 9920 5500 9926
rect 5448 9862 5500 9868
rect 5356 9512 5408 9518
rect 5356 9454 5408 9460
rect 5368 8974 5396 9454
rect 5356 8968 5408 8974
rect 5356 8910 5408 8916
rect 5460 8634 5488 9862
rect 5552 9586 5580 9930
rect 5540 9580 5592 9586
rect 5540 9522 5592 9528
rect 5448 8628 5500 8634
rect 5448 8570 5500 8576
rect 5448 8492 5500 8498
rect 5448 8434 5500 8440
rect 5356 8356 5408 8362
rect 5356 8298 5408 8304
rect 5172 8016 5224 8022
rect 5172 7958 5224 7964
rect 5264 7880 5316 7886
rect 5264 7822 5316 7828
rect 5172 7200 5224 7206
rect 5172 7142 5224 7148
rect 4846 7100 5154 7120
rect 4846 7098 4852 7100
rect 4908 7098 4932 7100
rect 4988 7098 5012 7100
rect 5068 7098 5092 7100
rect 5148 7098 5154 7100
rect 4908 7046 4910 7098
rect 5090 7046 5092 7098
rect 4846 7044 4852 7046
rect 4908 7044 4932 7046
rect 4988 7044 5012 7046
rect 5068 7044 5092 7046
rect 5148 7044 5154 7046
rect 4846 7024 5154 7044
rect 4712 6996 4764 7002
rect 4712 6938 4764 6944
rect 4712 6860 4764 6866
rect 4712 6802 4764 6808
rect 4724 5710 4752 6802
rect 5184 6390 5212 7142
rect 5276 6866 5304 7822
rect 5368 7410 5396 8298
rect 5356 7404 5408 7410
rect 5356 7346 5408 7352
rect 5460 6934 5488 8434
rect 5448 6928 5500 6934
rect 5448 6870 5500 6876
rect 5264 6860 5316 6866
rect 5264 6802 5316 6808
rect 5356 6724 5408 6730
rect 5356 6666 5408 6672
rect 5264 6656 5316 6662
rect 5264 6598 5316 6604
rect 5172 6384 5224 6390
rect 5172 6326 5224 6332
rect 4846 6012 5154 6032
rect 4846 6010 4852 6012
rect 4908 6010 4932 6012
rect 4988 6010 5012 6012
rect 5068 6010 5092 6012
rect 5148 6010 5154 6012
rect 4908 5958 4910 6010
rect 5090 5958 5092 6010
rect 4846 5956 4852 5958
rect 4908 5956 4932 5958
rect 4988 5956 5012 5958
rect 5068 5956 5092 5958
rect 5148 5956 5154 5958
rect 4846 5936 5154 5956
rect 4712 5704 4764 5710
rect 4712 5646 4764 5652
rect 5276 5642 5304 6598
rect 5368 5710 5396 6666
rect 5460 6254 5488 6870
rect 5448 6248 5500 6254
rect 5448 6190 5500 6196
rect 5356 5704 5408 5710
rect 5356 5646 5408 5652
rect 5264 5636 5316 5642
rect 5264 5578 5316 5584
rect 4846 4924 5154 4944
rect 4846 4922 4852 4924
rect 4908 4922 4932 4924
rect 4988 4922 5012 4924
rect 5068 4922 5092 4924
rect 5148 4922 5154 4924
rect 4908 4870 4910 4922
rect 5090 4870 5092 4922
rect 4846 4868 4852 4870
rect 4908 4868 4932 4870
rect 4988 4868 5012 4870
rect 5068 4868 5092 4870
rect 5148 4868 5154 4870
rect 4846 4848 5154 4868
rect 4804 4548 4856 4554
rect 4804 4490 4856 4496
rect 4816 4214 4844 4490
rect 4804 4208 4856 4214
rect 4804 4150 4856 4156
rect 5356 4140 5408 4146
rect 5356 4082 5408 4088
rect 4846 3836 5154 3856
rect 4846 3834 4852 3836
rect 4908 3834 4932 3836
rect 4988 3834 5012 3836
rect 5068 3834 5092 3836
rect 5148 3834 5154 3836
rect 4908 3782 4910 3834
rect 5090 3782 5092 3834
rect 4846 3780 4852 3782
rect 4908 3780 4932 3782
rect 4988 3780 5012 3782
rect 5068 3780 5092 3782
rect 5148 3780 5154 3782
rect 4846 3760 5154 3780
rect 5368 3194 5396 4082
rect 5356 3188 5408 3194
rect 5356 3130 5408 3136
rect 5264 3052 5316 3058
rect 5264 2994 5316 3000
rect 4712 2848 4764 2854
rect 4712 2790 4764 2796
rect 4724 2446 4752 2790
rect 4846 2748 5154 2768
rect 4846 2746 4852 2748
rect 4908 2746 4932 2748
rect 4988 2746 5012 2748
rect 5068 2746 5092 2748
rect 5148 2746 5154 2748
rect 4908 2694 4910 2746
rect 5090 2694 5092 2746
rect 4846 2692 4852 2694
rect 4908 2692 4932 2694
rect 4988 2692 5012 2694
rect 5068 2692 5092 2694
rect 5148 2692 5154 2694
rect 4846 2672 5154 2692
rect 5276 2650 5304 2994
rect 5552 2774 5580 9522
rect 5644 6882 5672 10095
rect 5736 8430 5764 10662
rect 5920 10674 5948 12106
rect 6012 11898 6040 13398
rect 6144 13084 6452 13104
rect 6144 13082 6150 13084
rect 6206 13082 6230 13084
rect 6286 13082 6310 13084
rect 6366 13082 6390 13084
rect 6446 13082 6452 13084
rect 6206 13030 6208 13082
rect 6388 13030 6390 13082
rect 6144 13028 6150 13030
rect 6206 13028 6230 13030
rect 6286 13028 6310 13030
rect 6366 13028 6390 13030
rect 6446 13028 6452 13030
rect 6144 13008 6452 13028
rect 6642 13016 6698 13025
rect 6642 12951 6698 12960
rect 6552 12232 6604 12238
rect 6552 12174 6604 12180
rect 6144 11996 6452 12016
rect 6144 11994 6150 11996
rect 6206 11994 6230 11996
rect 6286 11994 6310 11996
rect 6366 11994 6390 11996
rect 6446 11994 6452 11996
rect 6206 11942 6208 11994
rect 6388 11942 6390 11994
rect 6144 11940 6150 11942
rect 6206 11940 6230 11942
rect 6286 11940 6310 11942
rect 6366 11940 6390 11942
rect 6446 11940 6452 11942
rect 6144 11920 6452 11940
rect 6000 11892 6052 11898
rect 6000 11834 6052 11840
rect 6564 11830 6592 12174
rect 6656 12170 6684 12951
rect 6748 12594 6776 14776
rect 7443 14716 7751 14736
rect 7443 14714 7449 14716
rect 7505 14714 7529 14716
rect 7585 14714 7609 14716
rect 7665 14714 7689 14716
rect 7745 14714 7751 14716
rect 7505 14662 7507 14714
rect 7687 14662 7689 14714
rect 7443 14660 7449 14662
rect 7505 14660 7529 14662
rect 7585 14660 7609 14662
rect 7665 14660 7689 14662
rect 7745 14660 7751 14662
rect 7443 14640 7751 14660
rect 6828 14408 6880 14414
rect 6828 14350 6880 14356
rect 6840 14278 6868 14350
rect 6920 14340 6972 14346
rect 6920 14282 6972 14288
rect 7656 14340 7708 14346
rect 7656 14282 7708 14288
rect 6828 14272 6880 14278
rect 6828 14214 6880 14220
rect 6840 12753 6868 14214
rect 6932 12986 6960 14282
rect 7668 14006 7696 14282
rect 7656 14000 7708 14006
rect 7656 13942 7708 13948
rect 7012 13932 7064 13938
rect 7012 13874 7064 13880
rect 7024 13394 7052 13874
rect 7443 13628 7751 13648
rect 7443 13626 7449 13628
rect 7505 13626 7529 13628
rect 7585 13626 7609 13628
rect 7665 13626 7689 13628
rect 7745 13626 7751 13628
rect 7505 13574 7507 13626
rect 7687 13574 7689 13626
rect 7443 13572 7449 13574
rect 7505 13572 7529 13574
rect 7585 13572 7609 13574
rect 7665 13572 7689 13574
rect 7745 13572 7751 13574
rect 7443 13552 7751 13572
rect 7194 13424 7250 13433
rect 7012 13388 7064 13394
rect 7194 13359 7250 13368
rect 7012 13330 7064 13336
rect 7104 13320 7156 13326
rect 7208 13274 7236 13359
rect 7156 13268 7236 13274
rect 7104 13262 7236 13268
rect 7932 13320 7984 13326
rect 7932 13262 7984 13268
rect 7012 13252 7064 13258
rect 7116 13246 7236 13262
rect 7012 13194 7064 13200
rect 6920 12980 6972 12986
rect 6920 12922 6972 12928
rect 7024 12866 7052 13194
rect 7208 12889 7236 13246
rect 7380 13252 7432 13258
rect 7380 13194 7432 13200
rect 7392 12918 7420 13194
rect 7564 13184 7616 13190
rect 7564 13126 7616 13132
rect 7380 12912 7432 12918
rect 6932 12838 7052 12866
rect 7194 12880 7250 12889
rect 6826 12744 6882 12753
rect 6826 12679 6882 12688
rect 6748 12566 6868 12594
rect 6736 12232 6788 12238
rect 6736 12174 6788 12180
rect 6644 12164 6696 12170
rect 6644 12106 6696 12112
rect 6552 11824 6604 11830
rect 6552 11766 6604 11772
rect 6748 11694 6776 12174
rect 6736 11688 6788 11694
rect 6736 11630 6788 11636
rect 6748 11150 6776 11630
rect 6736 11144 6788 11150
rect 6736 11086 6788 11092
rect 6144 10908 6452 10928
rect 6144 10906 6150 10908
rect 6206 10906 6230 10908
rect 6286 10906 6310 10908
rect 6366 10906 6390 10908
rect 6446 10906 6452 10908
rect 6206 10854 6208 10906
rect 6388 10854 6390 10906
rect 6144 10852 6150 10854
rect 6206 10852 6230 10854
rect 6286 10852 6310 10854
rect 6366 10852 6390 10854
rect 6446 10852 6452 10854
rect 6144 10832 6452 10852
rect 6092 10736 6144 10742
rect 6092 10678 6144 10684
rect 5814 10639 5870 10648
rect 5908 10668 5960 10674
rect 5828 10606 5856 10639
rect 5908 10610 5960 10616
rect 5816 10600 5868 10606
rect 5816 10542 5868 10548
rect 5828 9382 5856 10542
rect 6104 10062 6132 10678
rect 6552 10600 6604 10606
rect 6552 10542 6604 10548
rect 6734 10568 6790 10577
rect 6564 10198 6592 10542
rect 6734 10503 6790 10512
rect 6552 10192 6604 10198
rect 6552 10134 6604 10140
rect 6092 10056 6144 10062
rect 6092 9998 6144 10004
rect 6644 10056 6696 10062
rect 6644 9998 6696 10004
rect 5908 9988 5960 9994
rect 5908 9930 5960 9936
rect 5920 9586 5948 9930
rect 6104 9908 6132 9998
rect 6012 9880 6132 9908
rect 5908 9580 5960 9586
rect 5908 9522 5960 9528
rect 5816 9376 5868 9382
rect 5816 9318 5868 9324
rect 5920 8906 5948 9522
rect 6012 9110 6040 9880
rect 6144 9820 6452 9840
rect 6144 9818 6150 9820
rect 6206 9818 6230 9820
rect 6286 9818 6310 9820
rect 6366 9818 6390 9820
rect 6446 9818 6452 9820
rect 6206 9766 6208 9818
rect 6388 9766 6390 9818
rect 6144 9764 6150 9766
rect 6206 9764 6230 9766
rect 6286 9764 6310 9766
rect 6366 9764 6390 9766
rect 6446 9764 6452 9766
rect 6144 9744 6452 9764
rect 6552 9716 6604 9722
rect 6182 9688 6238 9697
rect 6552 9658 6604 9664
rect 6182 9623 6238 9632
rect 6000 9104 6052 9110
rect 6000 9046 6052 9052
rect 6196 8906 6224 9623
rect 5908 8900 5960 8906
rect 5908 8842 5960 8848
rect 6184 8900 6236 8906
rect 6184 8842 6236 8848
rect 6144 8732 6452 8752
rect 6144 8730 6150 8732
rect 6206 8730 6230 8732
rect 6286 8730 6310 8732
rect 6366 8730 6390 8732
rect 6446 8730 6452 8732
rect 6206 8678 6208 8730
rect 6388 8678 6390 8730
rect 6144 8676 6150 8678
rect 6206 8676 6230 8678
rect 6286 8676 6310 8678
rect 6366 8676 6390 8678
rect 6446 8676 6452 8678
rect 6144 8656 6452 8676
rect 5724 8424 5776 8430
rect 5724 8366 5776 8372
rect 6184 8288 6236 8294
rect 6184 8230 6236 8236
rect 5908 8016 5960 8022
rect 5908 7958 5960 7964
rect 5644 6854 5856 6882
rect 5724 6792 5776 6798
rect 5724 6734 5776 6740
rect 5736 6254 5764 6734
rect 5724 6248 5776 6254
rect 5630 6216 5686 6225
rect 5724 6190 5776 6196
rect 5630 6151 5686 6160
rect 5644 5710 5672 6151
rect 5828 5778 5856 6854
rect 5816 5772 5868 5778
rect 5816 5714 5868 5720
rect 5632 5704 5684 5710
rect 5632 5646 5684 5652
rect 5722 5672 5778 5681
rect 5920 5658 5948 7958
rect 6196 7886 6224 8230
rect 6184 7880 6236 7886
rect 6184 7822 6236 7828
rect 6144 7644 6452 7664
rect 6144 7642 6150 7644
rect 6206 7642 6230 7644
rect 6286 7642 6310 7644
rect 6366 7642 6390 7644
rect 6446 7642 6452 7644
rect 6206 7590 6208 7642
rect 6388 7590 6390 7642
rect 6144 7588 6150 7590
rect 6206 7588 6230 7590
rect 6286 7588 6310 7590
rect 6366 7588 6390 7590
rect 6446 7588 6452 7590
rect 6144 7568 6452 7588
rect 6144 6556 6452 6576
rect 6144 6554 6150 6556
rect 6206 6554 6230 6556
rect 6286 6554 6310 6556
rect 6366 6554 6390 6556
rect 6446 6554 6452 6556
rect 6206 6502 6208 6554
rect 6388 6502 6390 6554
rect 6144 6500 6150 6502
rect 6206 6500 6230 6502
rect 6286 6500 6310 6502
rect 6366 6500 6390 6502
rect 6446 6500 6452 6502
rect 6144 6480 6452 6500
rect 6564 6474 6592 9658
rect 6656 9042 6684 9998
rect 6644 9036 6696 9042
rect 6644 8978 6696 8984
rect 6656 7993 6684 8978
rect 6642 7984 6698 7993
rect 6748 7970 6776 10503
rect 6840 10062 6868 12566
rect 6932 10810 6960 12838
rect 7380 12854 7432 12860
rect 7576 12850 7604 13126
rect 7194 12815 7250 12824
rect 7564 12844 7616 12850
rect 7012 12776 7064 12782
rect 7012 12718 7064 12724
rect 7024 11762 7052 12718
rect 7104 12096 7156 12102
rect 7104 12038 7156 12044
rect 7116 11830 7144 12038
rect 7104 11824 7156 11830
rect 7104 11766 7156 11772
rect 7012 11756 7064 11762
rect 7012 11698 7064 11704
rect 6920 10804 6972 10810
rect 6920 10746 6972 10752
rect 7208 10674 7236 12815
rect 7564 12786 7616 12792
rect 7288 12708 7340 12714
rect 7288 12650 7340 12656
rect 7300 12102 7328 12650
rect 7443 12540 7751 12560
rect 7443 12538 7449 12540
rect 7505 12538 7529 12540
rect 7585 12538 7609 12540
rect 7665 12538 7689 12540
rect 7745 12538 7751 12540
rect 7505 12486 7507 12538
rect 7687 12486 7689 12538
rect 7443 12484 7449 12486
rect 7505 12484 7529 12486
rect 7585 12484 7609 12486
rect 7665 12484 7689 12486
rect 7745 12484 7751 12486
rect 7443 12464 7751 12484
rect 7288 12096 7340 12102
rect 7288 12038 7340 12044
rect 7840 11756 7892 11762
rect 7840 11698 7892 11704
rect 7443 11452 7751 11472
rect 7443 11450 7449 11452
rect 7505 11450 7529 11452
rect 7585 11450 7609 11452
rect 7665 11450 7689 11452
rect 7745 11450 7751 11452
rect 7505 11398 7507 11450
rect 7687 11398 7689 11450
rect 7443 11396 7449 11398
rect 7505 11396 7529 11398
rect 7585 11396 7609 11398
rect 7665 11396 7689 11398
rect 7745 11396 7751 11398
rect 7443 11376 7751 11396
rect 7852 11393 7880 11698
rect 7838 11384 7894 11393
rect 7944 11354 7972 13262
rect 7838 11319 7894 11328
rect 7932 11348 7984 11354
rect 7932 11290 7984 11296
rect 7380 11144 7432 11150
rect 7380 11086 7432 11092
rect 7392 10849 7420 11086
rect 7840 11076 7892 11082
rect 7840 11018 7892 11024
rect 7378 10840 7434 10849
rect 7378 10775 7434 10784
rect 7196 10668 7248 10674
rect 7196 10610 7248 10616
rect 7852 10538 7880 11018
rect 7840 10532 7892 10538
rect 7840 10474 7892 10480
rect 7288 10464 7340 10470
rect 7288 10406 7340 10412
rect 7300 10130 7328 10406
rect 7443 10364 7751 10384
rect 7443 10362 7449 10364
rect 7505 10362 7529 10364
rect 7585 10362 7609 10364
rect 7665 10362 7689 10364
rect 7745 10362 7751 10364
rect 7505 10310 7507 10362
rect 7687 10310 7689 10362
rect 7443 10308 7449 10310
rect 7505 10308 7529 10310
rect 7585 10308 7609 10310
rect 7665 10308 7689 10310
rect 7745 10308 7751 10310
rect 7443 10288 7751 10308
rect 7288 10124 7340 10130
rect 7288 10066 7340 10072
rect 6828 10056 6880 10062
rect 6828 9998 6880 10004
rect 7380 9988 7432 9994
rect 7380 9930 7432 9936
rect 7392 9654 7420 9930
rect 7380 9648 7432 9654
rect 7380 9590 7432 9596
rect 7196 9444 7248 9450
rect 7196 9386 7248 9392
rect 7208 8974 7236 9386
rect 7443 9276 7751 9296
rect 7443 9274 7449 9276
rect 7505 9274 7529 9276
rect 7585 9274 7609 9276
rect 7665 9274 7689 9276
rect 7745 9274 7751 9276
rect 7505 9222 7507 9274
rect 7687 9222 7689 9274
rect 7443 9220 7449 9222
rect 7505 9220 7529 9222
rect 7585 9220 7609 9222
rect 7665 9220 7689 9222
rect 7745 9220 7751 9222
rect 7443 9200 7751 9220
rect 7852 9110 7880 10474
rect 8036 10146 8064 15966
rect 8116 15428 8168 15434
rect 8116 15370 8168 15376
rect 8128 15026 8156 15370
rect 8116 15020 8168 15026
rect 8116 14962 8168 14968
rect 8128 13682 8156 14962
rect 8208 14816 8260 14822
rect 8208 14758 8260 14764
rect 8220 14414 8248 14758
rect 8208 14408 8260 14414
rect 8208 14350 8260 14356
rect 8220 13938 8248 14350
rect 8208 13932 8260 13938
rect 8208 13874 8260 13880
rect 8220 13818 8248 13874
rect 8220 13790 8340 13818
rect 8128 13654 8248 13682
rect 8116 13320 8168 13326
rect 8116 13262 8168 13268
rect 8128 12850 8156 13262
rect 8116 12844 8168 12850
rect 8116 12786 8168 12792
rect 8128 10305 8156 12786
rect 8220 11937 8248 13654
rect 8206 11928 8262 11937
rect 8206 11863 8262 11872
rect 8208 11008 8260 11014
rect 8208 10950 8260 10956
rect 8220 10606 8248 10950
rect 8208 10600 8260 10606
rect 8208 10542 8260 10548
rect 8114 10296 8170 10305
rect 8114 10231 8170 10240
rect 7944 10118 8064 10146
rect 7944 10062 7972 10118
rect 7932 10056 7984 10062
rect 7932 9998 7984 10004
rect 7944 9586 7972 9998
rect 7932 9580 7984 9586
rect 7932 9522 7984 9528
rect 7840 9104 7892 9110
rect 7840 9046 7892 9052
rect 6828 8968 6880 8974
rect 6828 8910 6880 8916
rect 7196 8968 7248 8974
rect 7196 8910 7248 8916
rect 6840 8809 6868 8910
rect 6826 8800 6882 8809
rect 6826 8735 6882 8744
rect 7208 8566 7236 8910
rect 7196 8560 7248 8566
rect 7196 8502 7248 8508
rect 7288 8288 7340 8294
rect 7288 8230 7340 8236
rect 6748 7942 6868 7970
rect 6642 7919 6698 7928
rect 6736 7812 6788 7818
rect 6736 7754 6788 7760
rect 6748 7410 6776 7754
rect 6736 7404 6788 7410
rect 6736 7346 6788 7352
rect 6736 6656 6788 6662
rect 6736 6598 6788 6604
rect 6564 6446 6684 6474
rect 6656 5794 6684 6446
rect 6748 6254 6776 6598
rect 6736 6248 6788 6254
rect 6736 6190 6788 6196
rect 5828 5642 5948 5658
rect 5722 5607 5778 5616
rect 5816 5636 5948 5642
rect 5552 2746 5672 2774
rect 5264 2644 5316 2650
rect 5264 2586 5316 2592
rect 4712 2440 4764 2446
rect 4712 2382 4764 2388
rect 5644 2106 5672 2746
rect 5736 2514 5764 5607
rect 5868 5630 5948 5636
rect 6564 5766 6684 5794
rect 5816 5578 5868 5584
rect 5908 5568 5960 5574
rect 5908 5510 5960 5516
rect 5816 4616 5868 4622
rect 5816 4558 5868 4564
rect 5828 3534 5856 4558
rect 5920 4554 5948 5510
rect 6144 5468 6452 5488
rect 6144 5466 6150 5468
rect 6206 5466 6230 5468
rect 6286 5466 6310 5468
rect 6366 5466 6390 5468
rect 6446 5466 6452 5468
rect 6206 5414 6208 5466
rect 6388 5414 6390 5466
rect 6144 5412 6150 5414
rect 6206 5412 6230 5414
rect 6286 5412 6310 5414
rect 6366 5412 6390 5414
rect 6446 5412 6452 5414
rect 6144 5392 6452 5412
rect 6564 5166 6592 5766
rect 6644 5704 6696 5710
rect 6644 5646 6696 5652
rect 6368 5160 6420 5166
rect 6368 5102 6420 5108
rect 6552 5160 6604 5166
rect 6552 5102 6604 5108
rect 6000 5092 6052 5098
rect 6000 5034 6052 5040
rect 5908 4548 5960 4554
rect 5908 4490 5960 4496
rect 5920 4146 5948 4490
rect 5908 4140 5960 4146
rect 5908 4082 5960 4088
rect 6012 4010 6040 5034
rect 6380 4826 6408 5102
rect 6368 4820 6420 4826
rect 6368 4762 6420 4768
rect 6144 4380 6452 4400
rect 6144 4378 6150 4380
rect 6206 4378 6230 4380
rect 6286 4378 6310 4380
rect 6366 4378 6390 4380
rect 6446 4378 6452 4380
rect 6206 4326 6208 4378
rect 6388 4326 6390 4378
rect 6144 4324 6150 4326
rect 6206 4324 6230 4326
rect 6286 4324 6310 4326
rect 6366 4324 6390 4326
rect 6446 4324 6452 4326
rect 6144 4304 6452 4324
rect 6564 4146 6592 5102
rect 6552 4140 6604 4146
rect 6552 4082 6604 4088
rect 6000 4004 6052 4010
rect 6000 3946 6052 3952
rect 5816 3528 5868 3534
rect 5816 3470 5868 3476
rect 5828 2774 5856 3470
rect 6552 3460 6604 3466
rect 6552 3402 6604 3408
rect 6144 3292 6452 3312
rect 6144 3290 6150 3292
rect 6206 3290 6230 3292
rect 6286 3290 6310 3292
rect 6366 3290 6390 3292
rect 6446 3290 6452 3292
rect 6206 3238 6208 3290
rect 6388 3238 6390 3290
rect 6144 3236 6150 3238
rect 6206 3236 6230 3238
rect 6286 3236 6310 3238
rect 6366 3236 6390 3238
rect 6446 3236 6452 3238
rect 6144 3216 6452 3236
rect 6564 3126 6592 3402
rect 6552 3120 6604 3126
rect 6552 3062 6604 3068
rect 5828 2746 6040 2774
rect 5724 2508 5776 2514
rect 5724 2450 5776 2456
rect 5632 2100 5684 2106
rect 5632 2042 5684 2048
rect 6012 1193 6040 2746
rect 6564 2650 6592 3062
rect 6656 2961 6684 5646
rect 6748 5574 6776 6190
rect 6736 5568 6788 5574
rect 6736 5510 6788 5516
rect 6642 2952 6698 2961
rect 6642 2887 6698 2896
rect 6644 2848 6696 2854
rect 6644 2790 6696 2796
rect 6552 2644 6604 2650
rect 6552 2586 6604 2592
rect 6144 2204 6452 2224
rect 6144 2202 6150 2204
rect 6206 2202 6230 2204
rect 6286 2202 6310 2204
rect 6366 2202 6390 2204
rect 6446 2202 6452 2204
rect 6206 2150 6208 2202
rect 6388 2150 6390 2202
rect 6144 2148 6150 2150
rect 6206 2148 6230 2150
rect 6286 2148 6310 2150
rect 6366 2148 6390 2150
rect 6446 2148 6452 2150
rect 6144 2128 6452 2148
rect 6656 1737 6684 2790
rect 6642 1728 6698 1737
rect 6642 1663 6698 1672
rect 6552 1352 6604 1358
rect 6552 1294 6604 1300
rect 5998 1184 6054 1193
rect 5998 1119 6054 1128
rect 4816 870 4936 898
rect 4816 762 4844 870
rect 4908 800 4936 870
rect 4632 734 4844 762
rect 4894 0 4950 800
rect 6564 649 6592 1294
rect 6550 640 6606 649
rect 6550 575 6606 584
rect 6642 232 6698 241
rect 6748 218 6776 5510
rect 6840 5386 6868 7942
rect 7012 7880 7064 7886
rect 7012 7822 7064 7828
rect 6920 7812 6972 7818
rect 6920 7754 6972 7760
rect 6932 7546 6960 7754
rect 6920 7540 6972 7546
rect 6920 7482 6972 7488
rect 7024 6798 7052 7822
rect 7300 7410 7328 8230
rect 7443 8188 7751 8208
rect 7443 8186 7449 8188
rect 7505 8186 7529 8188
rect 7585 8186 7609 8188
rect 7665 8186 7689 8188
rect 7745 8186 7751 8188
rect 7505 8134 7507 8186
rect 7687 8134 7689 8186
rect 7443 8132 7449 8134
rect 7505 8132 7529 8134
rect 7585 8132 7609 8134
rect 7665 8132 7689 8134
rect 7745 8132 7751 8134
rect 7443 8112 7751 8132
rect 7840 7880 7892 7886
rect 7840 7822 7892 7828
rect 7288 7404 7340 7410
rect 7288 7346 7340 7352
rect 7852 7177 7880 7822
rect 7944 7721 7972 9522
rect 8128 9382 8156 9413
rect 8116 9376 8168 9382
rect 8114 9344 8116 9353
rect 8168 9344 8170 9353
rect 8114 9279 8170 9288
rect 8128 8498 8156 9279
rect 8220 8809 8248 10542
rect 8312 9897 8340 13790
rect 8392 13524 8444 13530
rect 8392 13466 8444 13472
rect 8404 11014 8432 13466
rect 8392 11008 8444 11014
rect 8392 10950 8444 10956
rect 8298 9888 8354 9897
rect 8298 9823 8354 9832
rect 8300 8900 8352 8906
rect 8300 8842 8352 8848
rect 8206 8800 8262 8809
rect 8206 8735 8262 8744
rect 8116 8492 8168 8498
rect 8116 8434 8168 8440
rect 7930 7712 7986 7721
rect 7930 7647 7986 7656
rect 7932 7404 7984 7410
rect 7932 7346 7984 7352
rect 7838 7168 7894 7177
rect 7443 7100 7751 7120
rect 7838 7103 7894 7112
rect 7443 7098 7449 7100
rect 7505 7098 7529 7100
rect 7585 7098 7609 7100
rect 7665 7098 7689 7100
rect 7745 7098 7751 7100
rect 7505 7046 7507 7098
rect 7687 7046 7689 7098
rect 7443 7044 7449 7046
rect 7505 7044 7529 7046
rect 7585 7044 7609 7046
rect 7665 7044 7689 7046
rect 7745 7044 7751 7046
rect 7443 7024 7751 7044
rect 7104 6860 7156 6866
rect 7104 6802 7156 6808
rect 7012 6792 7064 6798
rect 7012 6734 7064 6740
rect 7116 5642 7144 6802
rect 7944 6633 7972 7346
rect 8024 6792 8076 6798
rect 8024 6734 8076 6740
rect 7930 6624 7986 6633
rect 7930 6559 7986 6568
rect 7196 6316 7248 6322
rect 7196 6258 7248 6264
rect 7208 5710 7236 6258
rect 7443 6012 7751 6032
rect 7443 6010 7449 6012
rect 7505 6010 7529 6012
rect 7585 6010 7609 6012
rect 7665 6010 7689 6012
rect 7745 6010 7751 6012
rect 7505 5958 7507 6010
rect 7687 5958 7689 6010
rect 7443 5956 7449 5958
rect 7505 5956 7529 5958
rect 7585 5956 7609 5958
rect 7665 5956 7689 5958
rect 7745 5956 7751 5958
rect 7443 5936 7751 5956
rect 7288 5908 7340 5914
rect 7288 5850 7340 5856
rect 7196 5704 7248 5710
rect 7196 5646 7248 5652
rect 7104 5636 7156 5642
rect 7104 5578 7156 5584
rect 6840 5358 6960 5386
rect 6932 5302 6960 5358
rect 6828 5296 6880 5302
rect 6828 5238 6880 5244
rect 6920 5296 6972 5302
rect 6920 5238 6972 5244
rect 6840 4622 6868 5238
rect 7116 4978 7144 5578
rect 7196 5092 7248 5098
rect 7196 5034 7248 5040
rect 7024 4950 7144 4978
rect 6828 4616 6880 4622
rect 6828 4558 6880 4564
rect 6840 4049 6868 4558
rect 6826 4040 6882 4049
rect 6826 3975 6882 3984
rect 6920 3528 6972 3534
rect 6920 3470 6972 3476
rect 6828 3188 6880 3194
rect 6828 3130 6880 3136
rect 6840 2854 6868 3130
rect 6932 3126 6960 3470
rect 6920 3120 6972 3126
rect 6920 3062 6972 3068
rect 6920 2916 6972 2922
rect 6920 2858 6972 2864
rect 6828 2848 6880 2854
rect 6828 2790 6880 2796
rect 6932 800 6960 2858
rect 7024 2582 7052 4950
rect 7208 3126 7236 5034
rect 7300 4554 7328 5850
rect 7380 5840 7432 5846
rect 7380 5782 7432 5788
rect 7392 5302 7420 5782
rect 7840 5704 7892 5710
rect 7840 5646 7892 5652
rect 7380 5296 7432 5302
rect 7380 5238 7432 5244
rect 7443 4924 7751 4944
rect 7443 4922 7449 4924
rect 7505 4922 7529 4924
rect 7585 4922 7609 4924
rect 7665 4922 7689 4924
rect 7745 4922 7751 4924
rect 7505 4870 7507 4922
rect 7687 4870 7689 4922
rect 7443 4868 7449 4870
rect 7505 4868 7529 4870
rect 7585 4868 7609 4870
rect 7665 4868 7689 4870
rect 7745 4868 7751 4870
rect 7443 4848 7751 4868
rect 7288 4548 7340 4554
rect 7288 4490 7340 4496
rect 7443 3836 7751 3856
rect 7443 3834 7449 3836
rect 7505 3834 7529 3836
rect 7585 3834 7609 3836
rect 7665 3834 7689 3836
rect 7745 3834 7751 3836
rect 7505 3782 7507 3834
rect 7687 3782 7689 3834
rect 7443 3780 7449 3782
rect 7505 3780 7529 3782
rect 7585 3780 7609 3782
rect 7665 3780 7689 3782
rect 7745 3780 7751 3782
rect 7443 3760 7751 3780
rect 7196 3120 7248 3126
rect 7196 3062 7248 3068
rect 7012 2576 7064 2582
rect 7012 2518 7064 2524
rect 7208 2038 7236 3062
rect 7443 2748 7751 2768
rect 7443 2746 7449 2748
rect 7505 2746 7529 2748
rect 7585 2746 7609 2748
rect 7665 2746 7689 2748
rect 7745 2746 7751 2748
rect 7505 2694 7507 2746
rect 7687 2694 7689 2746
rect 7443 2692 7449 2694
rect 7505 2692 7529 2694
rect 7585 2692 7609 2694
rect 7665 2692 7689 2694
rect 7745 2692 7751 2694
rect 7443 2672 7751 2692
rect 7852 2514 7880 5646
rect 7932 5228 7984 5234
rect 7932 5170 7984 5176
rect 7944 5001 7972 5170
rect 7930 4992 7986 5001
rect 7930 4927 7986 4936
rect 7944 3058 7972 4927
rect 7932 3052 7984 3058
rect 7932 2994 7984 3000
rect 7840 2508 7892 2514
rect 7840 2450 7892 2456
rect 8036 2281 8064 6734
rect 8208 6316 8260 6322
rect 8208 6258 8260 6264
rect 8114 6080 8170 6089
rect 8114 6015 8170 6024
rect 8128 5710 8156 6015
rect 8116 5704 8168 5710
rect 8116 5646 8168 5652
rect 8220 5574 8248 6258
rect 8208 5568 8260 5574
rect 8206 5536 8208 5545
rect 8260 5536 8262 5545
rect 8206 5471 8262 5480
rect 8220 5445 8248 5471
rect 8312 4457 8340 8842
rect 8298 4448 8354 4457
rect 8298 4383 8354 4392
rect 8208 4140 8260 4146
rect 8208 4082 8260 4088
rect 8220 3369 8248 4082
rect 8312 3534 8340 4383
rect 8300 3528 8352 3534
rect 8300 3470 8352 3476
rect 8206 3360 8262 3369
rect 8206 3295 8262 3304
rect 8312 2514 8340 3470
rect 8300 2508 8352 2514
rect 8300 2450 8352 2456
rect 8022 2272 8078 2281
rect 8022 2207 8078 2216
rect 7196 2032 7248 2038
rect 7196 1974 7248 1980
rect 8944 1760 8996 1766
rect 8944 1702 8996 1708
rect 8956 800 8984 1702
rect 6698 190 6776 218
rect 6642 167 6698 176
rect 6918 0 6974 800
rect 8942 0 8998 800
<< via2 >>
rect 6642 29688 6698 29744
rect 6550 29144 6606 29200
rect 5538 28600 5594 28656
rect 2254 27770 2310 27772
rect 2334 27770 2390 27772
rect 2414 27770 2470 27772
rect 2494 27770 2550 27772
rect 2254 27718 2300 27770
rect 2300 27718 2310 27770
rect 2334 27718 2364 27770
rect 2364 27718 2376 27770
rect 2376 27718 2390 27770
rect 2414 27718 2428 27770
rect 2428 27718 2440 27770
rect 2440 27718 2470 27770
rect 2494 27718 2504 27770
rect 2504 27718 2550 27770
rect 2254 27716 2310 27718
rect 2334 27716 2390 27718
rect 2414 27716 2470 27718
rect 2494 27716 2550 27718
rect 4852 27770 4908 27772
rect 4932 27770 4988 27772
rect 5012 27770 5068 27772
rect 5092 27770 5148 27772
rect 4852 27718 4898 27770
rect 4898 27718 4908 27770
rect 4932 27718 4962 27770
rect 4962 27718 4974 27770
rect 4974 27718 4988 27770
rect 5012 27718 5026 27770
rect 5026 27718 5038 27770
rect 5038 27718 5068 27770
rect 5092 27718 5102 27770
rect 5102 27718 5148 27770
rect 4852 27716 4908 27718
rect 4932 27716 4988 27718
rect 5012 27716 5068 27718
rect 5092 27716 5148 27718
rect 2254 26682 2310 26684
rect 2334 26682 2390 26684
rect 2414 26682 2470 26684
rect 2494 26682 2550 26684
rect 2254 26630 2300 26682
rect 2300 26630 2310 26682
rect 2334 26630 2364 26682
rect 2364 26630 2376 26682
rect 2376 26630 2390 26682
rect 2414 26630 2428 26682
rect 2428 26630 2440 26682
rect 2440 26630 2470 26682
rect 2494 26630 2504 26682
rect 2504 26630 2550 26682
rect 2254 26628 2310 26630
rect 2334 26628 2390 26630
rect 2414 26628 2470 26630
rect 2494 26628 2550 26630
rect 5998 28056 6054 28112
rect 3553 27226 3609 27228
rect 3633 27226 3689 27228
rect 3713 27226 3769 27228
rect 3793 27226 3849 27228
rect 3553 27174 3599 27226
rect 3599 27174 3609 27226
rect 3633 27174 3663 27226
rect 3663 27174 3675 27226
rect 3675 27174 3689 27226
rect 3713 27174 3727 27226
rect 3727 27174 3739 27226
rect 3739 27174 3769 27226
rect 3793 27174 3803 27226
rect 3803 27174 3849 27226
rect 3553 27172 3609 27174
rect 3633 27172 3689 27174
rect 3713 27172 3769 27174
rect 3793 27172 3849 27174
rect 3553 26138 3609 26140
rect 3633 26138 3689 26140
rect 3713 26138 3769 26140
rect 3793 26138 3849 26140
rect 3553 26086 3599 26138
rect 3599 26086 3609 26138
rect 3633 26086 3663 26138
rect 3663 26086 3675 26138
rect 3675 26086 3689 26138
rect 3713 26086 3727 26138
rect 3727 26086 3739 26138
rect 3739 26086 3769 26138
rect 3793 26086 3803 26138
rect 3803 26086 3849 26138
rect 3553 26084 3609 26086
rect 3633 26084 3689 26086
rect 3713 26084 3769 26086
rect 3793 26084 3849 26086
rect 2254 25594 2310 25596
rect 2334 25594 2390 25596
rect 2414 25594 2470 25596
rect 2494 25594 2550 25596
rect 2254 25542 2300 25594
rect 2300 25542 2310 25594
rect 2334 25542 2364 25594
rect 2364 25542 2376 25594
rect 2376 25542 2390 25594
rect 2414 25542 2428 25594
rect 2428 25542 2440 25594
rect 2440 25542 2470 25594
rect 2494 25542 2504 25594
rect 2504 25542 2550 25594
rect 2254 25540 2310 25542
rect 2334 25540 2390 25542
rect 2414 25540 2470 25542
rect 2494 25540 2550 25542
rect 3553 25050 3609 25052
rect 3633 25050 3689 25052
rect 3713 25050 3769 25052
rect 3793 25050 3849 25052
rect 3553 24998 3599 25050
rect 3599 24998 3609 25050
rect 3633 24998 3663 25050
rect 3663 24998 3675 25050
rect 3675 24998 3689 25050
rect 3713 24998 3727 25050
rect 3727 24998 3739 25050
rect 3739 24998 3769 25050
rect 3793 24998 3803 25050
rect 3803 24998 3849 25050
rect 3553 24996 3609 24998
rect 3633 24996 3689 24998
rect 3713 24996 3769 24998
rect 3793 24996 3849 24998
rect 2254 24506 2310 24508
rect 2334 24506 2390 24508
rect 2414 24506 2470 24508
rect 2494 24506 2550 24508
rect 2254 24454 2300 24506
rect 2300 24454 2310 24506
rect 2334 24454 2364 24506
rect 2364 24454 2376 24506
rect 2376 24454 2390 24506
rect 2414 24454 2428 24506
rect 2428 24454 2440 24506
rect 2440 24454 2470 24506
rect 2494 24454 2504 24506
rect 2504 24454 2550 24506
rect 2254 24452 2310 24454
rect 2334 24452 2390 24454
rect 2414 24452 2470 24454
rect 2494 24452 2550 24454
rect 4852 26682 4908 26684
rect 4932 26682 4988 26684
rect 5012 26682 5068 26684
rect 5092 26682 5148 26684
rect 4852 26630 4898 26682
rect 4898 26630 4908 26682
rect 4932 26630 4962 26682
rect 4962 26630 4974 26682
rect 4974 26630 4988 26682
rect 5012 26630 5026 26682
rect 5026 26630 5038 26682
rect 5038 26630 5068 26682
rect 5092 26630 5102 26682
rect 5102 26630 5148 26682
rect 4852 26628 4908 26630
rect 4932 26628 4988 26630
rect 5012 26628 5068 26630
rect 5092 26628 5148 26630
rect 4852 25594 4908 25596
rect 4932 25594 4988 25596
rect 5012 25594 5068 25596
rect 5092 25594 5148 25596
rect 4852 25542 4898 25594
rect 4898 25542 4908 25594
rect 4932 25542 4962 25594
rect 4962 25542 4974 25594
rect 4974 25542 4988 25594
rect 5012 25542 5026 25594
rect 5026 25542 5038 25594
rect 5038 25542 5068 25594
rect 5092 25542 5102 25594
rect 5102 25542 5148 25594
rect 4852 25540 4908 25542
rect 4932 25540 4988 25542
rect 5012 25540 5068 25542
rect 5092 25540 5148 25542
rect 5722 26968 5778 27024
rect 5906 27512 5962 27568
rect 3553 23962 3609 23964
rect 3633 23962 3689 23964
rect 3713 23962 3769 23964
rect 3793 23962 3849 23964
rect 3553 23910 3599 23962
rect 3599 23910 3609 23962
rect 3633 23910 3663 23962
rect 3663 23910 3675 23962
rect 3675 23910 3689 23962
rect 3713 23910 3727 23962
rect 3727 23910 3739 23962
rect 3739 23910 3769 23962
rect 3793 23910 3803 23962
rect 3803 23910 3849 23962
rect 3553 23908 3609 23910
rect 3633 23908 3689 23910
rect 3713 23908 3769 23910
rect 3793 23908 3849 23910
rect 2254 23418 2310 23420
rect 2334 23418 2390 23420
rect 2414 23418 2470 23420
rect 2494 23418 2550 23420
rect 2254 23366 2300 23418
rect 2300 23366 2310 23418
rect 2334 23366 2364 23418
rect 2364 23366 2376 23418
rect 2376 23366 2390 23418
rect 2414 23366 2428 23418
rect 2428 23366 2440 23418
rect 2440 23366 2470 23418
rect 2494 23366 2504 23418
rect 2504 23366 2550 23418
rect 2254 23364 2310 23366
rect 2334 23364 2390 23366
rect 2414 23364 2470 23366
rect 2494 23364 2550 23366
rect 2254 22330 2310 22332
rect 2334 22330 2390 22332
rect 2414 22330 2470 22332
rect 2494 22330 2550 22332
rect 2254 22278 2300 22330
rect 2300 22278 2310 22330
rect 2334 22278 2364 22330
rect 2364 22278 2376 22330
rect 2376 22278 2390 22330
rect 2414 22278 2428 22330
rect 2428 22278 2440 22330
rect 2440 22278 2470 22330
rect 2494 22278 2504 22330
rect 2504 22278 2550 22330
rect 2254 22276 2310 22278
rect 2334 22276 2390 22278
rect 2414 22276 2470 22278
rect 2494 22276 2550 22278
rect 3553 22874 3609 22876
rect 3633 22874 3689 22876
rect 3713 22874 3769 22876
rect 3793 22874 3849 22876
rect 3553 22822 3599 22874
rect 3599 22822 3609 22874
rect 3633 22822 3663 22874
rect 3663 22822 3675 22874
rect 3675 22822 3689 22874
rect 3713 22822 3727 22874
rect 3727 22822 3739 22874
rect 3739 22822 3769 22874
rect 3793 22822 3803 22874
rect 3803 22822 3849 22874
rect 3553 22820 3609 22822
rect 3633 22820 3689 22822
rect 3713 22820 3769 22822
rect 3793 22820 3849 22822
rect 4852 24506 4908 24508
rect 4932 24506 4988 24508
rect 5012 24506 5068 24508
rect 5092 24506 5148 24508
rect 4852 24454 4898 24506
rect 4898 24454 4908 24506
rect 4932 24454 4962 24506
rect 4962 24454 4974 24506
rect 4974 24454 4988 24506
rect 5012 24454 5026 24506
rect 5026 24454 5038 24506
rect 5038 24454 5068 24506
rect 5092 24454 5102 24506
rect 5102 24454 5148 24506
rect 4852 24452 4908 24454
rect 4932 24452 4988 24454
rect 5012 24452 5068 24454
rect 5092 24452 5148 24454
rect 4852 23418 4908 23420
rect 4932 23418 4988 23420
rect 5012 23418 5068 23420
rect 5092 23418 5148 23420
rect 4852 23366 4898 23418
rect 4898 23366 4908 23418
rect 4932 23366 4962 23418
rect 4962 23366 4974 23418
rect 4974 23366 4988 23418
rect 5012 23366 5026 23418
rect 5026 23366 5038 23418
rect 5038 23366 5068 23418
rect 5092 23366 5102 23418
rect 5102 23366 5148 23418
rect 4852 23364 4908 23366
rect 4932 23364 4988 23366
rect 5012 23364 5068 23366
rect 5092 23364 5148 23366
rect 6150 27226 6206 27228
rect 6230 27226 6286 27228
rect 6310 27226 6366 27228
rect 6390 27226 6446 27228
rect 6150 27174 6196 27226
rect 6196 27174 6206 27226
rect 6230 27174 6260 27226
rect 6260 27174 6272 27226
rect 6272 27174 6286 27226
rect 6310 27174 6324 27226
rect 6324 27174 6336 27226
rect 6336 27174 6366 27226
rect 6390 27174 6400 27226
rect 6400 27174 6446 27226
rect 6150 27172 6206 27174
rect 6230 27172 6286 27174
rect 6310 27172 6366 27174
rect 6390 27172 6446 27174
rect 6150 26138 6206 26140
rect 6230 26138 6286 26140
rect 6310 26138 6366 26140
rect 6390 26138 6446 26140
rect 6150 26086 6196 26138
rect 6196 26086 6206 26138
rect 6230 26086 6260 26138
rect 6260 26086 6272 26138
rect 6272 26086 6286 26138
rect 6310 26086 6324 26138
rect 6324 26086 6336 26138
rect 6336 26086 6366 26138
rect 6390 26086 6400 26138
rect 6400 26086 6446 26138
rect 6150 26084 6206 26086
rect 6230 26084 6286 26086
rect 6310 26084 6366 26086
rect 6390 26084 6446 26086
rect 6150 25050 6206 25052
rect 6230 25050 6286 25052
rect 6310 25050 6366 25052
rect 6390 25050 6446 25052
rect 6150 24998 6196 25050
rect 6196 24998 6206 25050
rect 6230 24998 6260 25050
rect 6260 24998 6272 25050
rect 6272 24998 6286 25050
rect 6310 24998 6324 25050
rect 6324 24998 6336 25050
rect 6336 24998 6366 25050
rect 6390 24998 6400 25050
rect 6400 24998 6446 25050
rect 6150 24996 6206 24998
rect 6230 24996 6286 24998
rect 6310 24996 6366 24998
rect 6390 24996 6446 24998
rect 7449 27770 7505 27772
rect 7529 27770 7585 27772
rect 7609 27770 7665 27772
rect 7689 27770 7745 27772
rect 7449 27718 7495 27770
rect 7495 27718 7505 27770
rect 7529 27718 7559 27770
rect 7559 27718 7571 27770
rect 7571 27718 7585 27770
rect 7609 27718 7623 27770
rect 7623 27718 7635 27770
rect 7635 27718 7665 27770
rect 7689 27718 7699 27770
rect 7699 27718 7745 27770
rect 7449 27716 7505 27718
rect 7529 27716 7585 27718
rect 7609 27716 7665 27718
rect 7689 27716 7745 27718
rect 6734 26424 6790 26480
rect 6642 25880 6698 25936
rect 7449 26682 7505 26684
rect 7529 26682 7585 26684
rect 7609 26682 7665 26684
rect 7689 26682 7745 26684
rect 7449 26630 7495 26682
rect 7495 26630 7505 26682
rect 7529 26630 7559 26682
rect 7559 26630 7571 26682
rect 7571 26630 7585 26682
rect 7609 26630 7623 26682
rect 7623 26630 7635 26682
rect 7635 26630 7665 26682
rect 7689 26630 7699 26682
rect 7699 26630 7745 26682
rect 7449 26628 7505 26630
rect 7529 26628 7585 26630
rect 7609 26628 7665 26630
rect 7689 26628 7745 26630
rect 3553 21786 3609 21788
rect 3633 21786 3689 21788
rect 3713 21786 3769 21788
rect 3793 21786 3849 21788
rect 3553 21734 3599 21786
rect 3599 21734 3609 21786
rect 3633 21734 3663 21786
rect 3663 21734 3675 21786
rect 3675 21734 3689 21786
rect 3713 21734 3727 21786
rect 3727 21734 3739 21786
rect 3739 21734 3769 21786
rect 3793 21734 3803 21786
rect 3803 21734 3849 21786
rect 3553 21732 3609 21734
rect 3633 21732 3689 21734
rect 3713 21732 3769 21734
rect 3793 21732 3849 21734
rect 2254 21242 2310 21244
rect 2334 21242 2390 21244
rect 2414 21242 2470 21244
rect 2494 21242 2550 21244
rect 2254 21190 2300 21242
rect 2300 21190 2310 21242
rect 2334 21190 2364 21242
rect 2364 21190 2376 21242
rect 2376 21190 2390 21242
rect 2414 21190 2428 21242
rect 2428 21190 2440 21242
rect 2440 21190 2470 21242
rect 2494 21190 2504 21242
rect 2504 21190 2550 21242
rect 2254 21188 2310 21190
rect 2334 21188 2390 21190
rect 2414 21188 2470 21190
rect 2494 21188 2550 21190
rect 2254 20154 2310 20156
rect 2334 20154 2390 20156
rect 2414 20154 2470 20156
rect 2494 20154 2550 20156
rect 2254 20102 2300 20154
rect 2300 20102 2310 20154
rect 2334 20102 2364 20154
rect 2364 20102 2376 20154
rect 2376 20102 2390 20154
rect 2414 20102 2428 20154
rect 2428 20102 2440 20154
rect 2440 20102 2470 20154
rect 2494 20102 2504 20154
rect 2504 20102 2550 20154
rect 2254 20100 2310 20102
rect 2334 20100 2390 20102
rect 2414 20100 2470 20102
rect 2494 20100 2550 20102
rect 2254 19066 2310 19068
rect 2334 19066 2390 19068
rect 2414 19066 2470 19068
rect 2494 19066 2550 19068
rect 2254 19014 2300 19066
rect 2300 19014 2310 19066
rect 2334 19014 2364 19066
rect 2364 19014 2376 19066
rect 2376 19014 2390 19066
rect 2414 19014 2428 19066
rect 2428 19014 2440 19066
rect 2440 19014 2470 19066
rect 2494 19014 2504 19066
rect 2504 19014 2550 19066
rect 2254 19012 2310 19014
rect 2334 19012 2390 19014
rect 2414 19012 2470 19014
rect 2494 19012 2550 19014
rect 3553 20698 3609 20700
rect 3633 20698 3689 20700
rect 3713 20698 3769 20700
rect 3793 20698 3849 20700
rect 3553 20646 3599 20698
rect 3599 20646 3609 20698
rect 3633 20646 3663 20698
rect 3663 20646 3675 20698
rect 3675 20646 3689 20698
rect 3713 20646 3727 20698
rect 3727 20646 3739 20698
rect 3739 20646 3769 20698
rect 3793 20646 3803 20698
rect 3803 20646 3849 20698
rect 3553 20644 3609 20646
rect 3633 20644 3689 20646
rect 3713 20644 3769 20646
rect 3793 20644 3849 20646
rect 4852 22330 4908 22332
rect 4932 22330 4988 22332
rect 5012 22330 5068 22332
rect 5092 22330 5148 22332
rect 4852 22278 4898 22330
rect 4898 22278 4908 22330
rect 4932 22278 4962 22330
rect 4962 22278 4974 22330
rect 4974 22278 4988 22330
rect 5012 22278 5026 22330
rect 5026 22278 5038 22330
rect 5038 22278 5068 22330
rect 5092 22278 5102 22330
rect 5102 22278 5148 22330
rect 4852 22276 4908 22278
rect 4932 22276 4988 22278
rect 5012 22276 5068 22278
rect 5092 22276 5148 22278
rect 6150 23962 6206 23964
rect 6230 23962 6286 23964
rect 6310 23962 6366 23964
rect 6390 23962 6446 23964
rect 6150 23910 6196 23962
rect 6196 23910 6206 23962
rect 6230 23910 6260 23962
rect 6260 23910 6272 23962
rect 6272 23910 6286 23962
rect 6310 23910 6324 23962
rect 6324 23910 6336 23962
rect 6336 23910 6366 23962
rect 6390 23910 6400 23962
rect 6400 23910 6446 23962
rect 6150 23908 6206 23910
rect 6230 23908 6286 23910
rect 6310 23908 6366 23910
rect 6390 23908 6446 23910
rect 7449 25594 7505 25596
rect 7529 25594 7585 25596
rect 7609 25594 7665 25596
rect 7689 25594 7745 25596
rect 7449 25542 7495 25594
rect 7495 25542 7505 25594
rect 7529 25542 7559 25594
rect 7559 25542 7571 25594
rect 7571 25542 7585 25594
rect 7609 25542 7623 25594
rect 7623 25542 7635 25594
rect 7635 25542 7665 25594
rect 7689 25542 7699 25594
rect 7699 25542 7745 25594
rect 7449 25540 7505 25542
rect 7529 25540 7585 25542
rect 7609 25540 7665 25542
rect 7689 25540 7745 25542
rect 7838 25336 7894 25392
rect 7930 24792 7986 24848
rect 6150 22874 6206 22876
rect 6230 22874 6286 22876
rect 6310 22874 6366 22876
rect 6390 22874 6446 22876
rect 6150 22822 6196 22874
rect 6196 22822 6206 22874
rect 6230 22822 6260 22874
rect 6260 22822 6272 22874
rect 6272 22822 6286 22874
rect 6310 22822 6324 22874
rect 6324 22822 6336 22874
rect 6336 22822 6366 22874
rect 6390 22822 6400 22874
rect 6400 22822 6446 22874
rect 6150 22820 6206 22822
rect 6230 22820 6286 22822
rect 6310 22820 6366 22822
rect 6390 22820 6446 22822
rect 6734 23160 6790 23216
rect 7449 24506 7505 24508
rect 7529 24506 7585 24508
rect 7609 24506 7665 24508
rect 7689 24506 7745 24508
rect 7449 24454 7495 24506
rect 7495 24454 7505 24506
rect 7529 24454 7559 24506
rect 7559 24454 7571 24506
rect 7571 24454 7585 24506
rect 7609 24454 7623 24506
rect 7623 24454 7635 24506
rect 7635 24454 7665 24506
rect 7689 24454 7699 24506
rect 7699 24454 7745 24506
rect 7449 24452 7505 24454
rect 7529 24452 7585 24454
rect 7609 24452 7665 24454
rect 7689 24452 7745 24454
rect 7449 23418 7505 23420
rect 7529 23418 7585 23420
rect 7609 23418 7665 23420
rect 7689 23418 7745 23420
rect 7449 23366 7495 23418
rect 7495 23366 7505 23418
rect 7529 23366 7559 23418
rect 7559 23366 7571 23418
rect 7571 23366 7585 23418
rect 7609 23366 7623 23418
rect 7623 23366 7635 23418
rect 7635 23366 7665 23418
rect 7689 23366 7699 23418
rect 7699 23366 7745 23418
rect 7449 23364 7505 23366
rect 7529 23364 7585 23366
rect 7609 23364 7665 23366
rect 7689 23364 7745 23366
rect 7449 22330 7505 22332
rect 7529 22330 7585 22332
rect 7609 22330 7665 22332
rect 7689 22330 7745 22332
rect 7449 22278 7495 22330
rect 7495 22278 7505 22330
rect 7529 22278 7559 22330
rect 7559 22278 7571 22330
rect 7571 22278 7585 22330
rect 7609 22278 7623 22330
rect 7623 22278 7635 22330
rect 7635 22278 7665 22330
rect 7689 22278 7699 22330
rect 7699 22278 7745 22330
rect 7449 22276 7505 22278
rect 7529 22276 7585 22278
rect 7609 22276 7665 22278
rect 7689 22276 7745 22278
rect 6150 21786 6206 21788
rect 6230 21786 6286 21788
rect 6310 21786 6366 21788
rect 6390 21786 6446 21788
rect 6150 21734 6196 21786
rect 6196 21734 6206 21786
rect 6230 21734 6260 21786
rect 6260 21734 6272 21786
rect 6272 21734 6286 21786
rect 6310 21734 6324 21786
rect 6324 21734 6336 21786
rect 6336 21734 6366 21786
rect 6390 21734 6400 21786
rect 6400 21734 6446 21786
rect 6150 21732 6206 21734
rect 6230 21732 6286 21734
rect 6310 21732 6366 21734
rect 6390 21732 6446 21734
rect 6734 21528 6790 21584
rect 4852 21242 4908 21244
rect 4932 21242 4988 21244
rect 5012 21242 5068 21244
rect 5092 21242 5148 21244
rect 4852 21190 4898 21242
rect 4898 21190 4908 21242
rect 4932 21190 4962 21242
rect 4962 21190 4974 21242
rect 4974 21190 4988 21242
rect 5012 21190 5026 21242
rect 5026 21190 5038 21242
rect 5038 21190 5068 21242
rect 5092 21190 5102 21242
rect 5102 21190 5148 21242
rect 4852 21188 4908 21190
rect 4932 21188 4988 21190
rect 5012 21188 5068 21190
rect 5092 21188 5148 21190
rect 6150 20698 6206 20700
rect 6230 20698 6286 20700
rect 6310 20698 6366 20700
rect 6390 20698 6446 20700
rect 6150 20646 6196 20698
rect 6196 20646 6206 20698
rect 6230 20646 6260 20698
rect 6260 20646 6272 20698
rect 6272 20646 6286 20698
rect 6310 20646 6324 20698
rect 6324 20646 6336 20698
rect 6336 20646 6366 20698
rect 6390 20646 6400 20698
rect 6400 20646 6446 20698
rect 6150 20644 6206 20646
rect 6230 20644 6286 20646
rect 6310 20644 6366 20646
rect 6390 20644 6446 20646
rect 3553 19610 3609 19612
rect 3633 19610 3689 19612
rect 3713 19610 3769 19612
rect 3793 19610 3849 19612
rect 3553 19558 3599 19610
rect 3599 19558 3609 19610
rect 3633 19558 3663 19610
rect 3663 19558 3675 19610
rect 3675 19558 3689 19610
rect 3713 19558 3727 19610
rect 3727 19558 3739 19610
rect 3739 19558 3769 19610
rect 3793 19558 3803 19610
rect 3803 19558 3849 19610
rect 3553 19556 3609 19558
rect 3633 19556 3689 19558
rect 3713 19556 3769 19558
rect 3793 19556 3849 19558
rect 2254 17978 2310 17980
rect 2334 17978 2390 17980
rect 2414 17978 2470 17980
rect 2494 17978 2550 17980
rect 2254 17926 2300 17978
rect 2300 17926 2310 17978
rect 2334 17926 2364 17978
rect 2364 17926 2376 17978
rect 2376 17926 2390 17978
rect 2414 17926 2428 17978
rect 2428 17926 2440 17978
rect 2440 17926 2470 17978
rect 2494 17926 2504 17978
rect 2504 17926 2550 17978
rect 2254 17924 2310 17926
rect 2334 17924 2390 17926
rect 2414 17924 2470 17926
rect 2494 17924 2550 17926
rect 2594 17060 2650 17096
rect 2594 17040 2596 17060
rect 2596 17040 2648 17060
rect 2648 17040 2650 17060
rect 2254 16890 2310 16892
rect 2334 16890 2390 16892
rect 2414 16890 2470 16892
rect 2494 16890 2550 16892
rect 2254 16838 2300 16890
rect 2300 16838 2310 16890
rect 2334 16838 2364 16890
rect 2364 16838 2376 16890
rect 2376 16838 2390 16890
rect 2414 16838 2428 16890
rect 2428 16838 2440 16890
rect 2440 16838 2470 16890
rect 2494 16838 2504 16890
rect 2504 16838 2550 16890
rect 2254 16836 2310 16838
rect 2334 16836 2390 16838
rect 2414 16836 2470 16838
rect 2494 16836 2550 16838
rect 2254 15802 2310 15804
rect 2334 15802 2390 15804
rect 2414 15802 2470 15804
rect 2494 15802 2550 15804
rect 2254 15750 2300 15802
rect 2300 15750 2310 15802
rect 2334 15750 2364 15802
rect 2364 15750 2376 15802
rect 2376 15750 2390 15802
rect 2414 15750 2428 15802
rect 2428 15750 2440 15802
rect 2440 15750 2470 15802
rect 2494 15750 2504 15802
rect 2504 15750 2550 15802
rect 2254 15748 2310 15750
rect 2334 15748 2390 15750
rect 2414 15748 2470 15750
rect 2494 15748 2550 15750
rect 2254 14714 2310 14716
rect 2334 14714 2390 14716
rect 2414 14714 2470 14716
rect 2494 14714 2550 14716
rect 2254 14662 2300 14714
rect 2300 14662 2310 14714
rect 2334 14662 2364 14714
rect 2364 14662 2376 14714
rect 2376 14662 2390 14714
rect 2414 14662 2428 14714
rect 2428 14662 2440 14714
rect 2440 14662 2470 14714
rect 2494 14662 2504 14714
rect 2504 14662 2550 14714
rect 2254 14660 2310 14662
rect 2334 14660 2390 14662
rect 2414 14660 2470 14662
rect 2494 14660 2550 14662
rect 2254 13626 2310 13628
rect 2334 13626 2390 13628
rect 2414 13626 2470 13628
rect 2494 13626 2550 13628
rect 2254 13574 2300 13626
rect 2300 13574 2310 13626
rect 2334 13574 2364 13626
rect 2364 13574 2376 13626
rect 2376 13574 2390 13626
rect 2414 13574 2428 13626
rect 2428 13574 2440 13626
rect 2440 13574 2470 13626
rect 2494 13574 2504 13626
rect 2504 13574 2550 13626
rect 2254 13572 2310 13574
rect 2334 13572 2390 13574
rect 2414 13572 2470 13574
rect 2494 13572 2550 13574
rect 2254 12538 2310 12540
rect 2334 12538 2390 12540
rect 2414 12538 2470 12540
rect 2494 12538 2550 12540
rect 2254 12486 2300 12538
rect 2300 12486 2310 12538
rect 2334 12486 2364 12538
rect 2364 12486 2376 12538
rect 2376 12486 2390 12538
rect 2414 12486 2428 12538
rect 2428 12486 2440 12538
rect 2440 12486 2470 12538
rect 2494 12486 2504 12538
rect 2504 12486 2550 12538
rect 2254 12484 2310 12486
rect 2334 12484 2390 12486
rect 2414 12484 2470 12486
rect 2494 12484 2550 12486
rect 1582 9968 1638 10024
rect 2254 11450 2310 11452
rect 2334 11450 2390 11452
rect 2414 11450 2470 11452
rect 2494 11450 2550 11452
rect 2254 11398 2300 11450
rect 2300 11398 2310 11450
rect 2334 11398 2364 11450
rect 2364 11398 2376 11450
rect 2376 11398 2390 11450
rect 2414 11398 2428 11450
rect 2428 11398 2440 11450
rect 2440 11398 2470 11450
rect 2494 11398 2504 11450
rect 2504 11398 2550 11450
rect 2254 11396 2310 11398
rect 2334 11396 2390 11398
rect 2414 11396 2470 11398
rect 2494 11396 2550 11398
rect 1766 7248 1822 7304
rect 1582 5616 1638 5672
rect 1398 5108 1400 5128
rect 1400 5108 1452 5128
rect 1452 5108 1454 5128
rect 1398 5072 1454 5108
rect 2254 10362 2310 10364
rect 2334 10362 2390 10364
rect 2414 10362 2470 10364
rect 2494 10362 2550 10364
rect 2254 10310 2300 10362
rect 2300 10310 2310 10362
rect 2334 10310 2364 10362
rect 2364 10310 2376 10362
rect 2376 10310 2390 10362
rect 2414 10310 2428 10362
rect 2428 10310 2440 10362
rect 2440 10310 2470 10362
rect 2494 10310 2504 10362
rect 2504 10310 2550 10362
rect 2254 10308 2310 10310
rect 2334 10308 2390 10310
rect 2414 10308 2470 10310
rect 2494 10308 2550 10310
rect 3553 18522 3609 18524
rect 3633 18522 3689 18524
rect 3713 18522 3769 18524
rect 3793 18522 3849 18524
rect 3553 18470 3599 18522
rect 3599 18470 3609 18522
rect 3633 18470 3663 18522
rect 3663 18470 3675 18522
rect 3675 18470 3689 18522
rect 3713 18470 3727 18522
rect 3727 18470 3739 18522
rect 3739 18470 3769 18522
rect 3793 18470 3803 18522
rect 3803 18470 3849 18522
rect 3553 18468 3609 18470
rect 3633 18468 3689 18470
rect 3713 18468 3769 18470
rect 3793 18468 3849 18470
rect 4066 17448 4122 17504
rect 3553 17434 3609 17436
rect 3633 17434 3689 17436
rect 3713 17434 3769 17436
rect 3793 17434 3849 17436
rect 3553 17382 3599 17434
rect 3599 17382 3609 17434
rect 3633 17382 3663 17434
rect 3663 17382 3675 17434
rect 3675 17382 3689 17434
rect 3713 17382 3727 17434
rect 3727 17382 3739 17434
rect 3739 17382 3769 17434
rect 3793 17382 3803 17434
rect 3803 17382 3849 17434
rect 3553 17380 3609 17382
rect 3633 17380 3689 17382
rect 3713 17380 3769 17382
rect 3793 17380 3849 17382
rect 3553 16346 3609 16348
rect 3633 16346 3689 16348
rect 3713 16346 3769 16348
rect 3793 16346 3849 16348
rect 3553 16294 3599 16346
rect 3599 16294 3609 16346
rect 3633 16294 3663 16346
rect 3663 16294 3675 16346
rect 3675 16294 3689 16346
rect 3713 16294 3727 16346
rect 3727 16294 3739 16346
rect 3739 16294 3769 16346
rect 3793 16294 3803 16346
rect 3803 16294 3849 16346
rect 3553 16292 3609 16294
rect 3633 16292 3689 16294
rect 3713 16292 3769 16294
rect 3793 16292 3849 16294
rect 4852 20154 4908 20156
rect 4932 20154 4988 20156
rect 5012 20154 5068 20156
rect 5092 20154 5148 20156
rect 4852 20102 4898 20154
rect 4898 20102 4908 20154
rect 4932 20102 4962 20154
rect 4962 20102 4974 20154
rect 4974 20102 4988 20154
rect 5012 20102 5026 20154
rect 5026 20102 5038 20154
rect 5038 20102 5068 20154
rect 5092 20102 5102 20154
rect 5102 20102 5148 20154
rect 4852 20100 4908 20102
rect 4932 20100 4988 20102
rect 5012 20100 5068 20102
rect 5092 20100 5148 20102
rect 4852 19066 4908 19068
rect 4932 19066 4988 19068
rect 5012 19066 5068 19068
rect 5092 19066 5148 19068
rect 4852 19014 4898 19066
rect 4898 19014 4908 19066
rect 4932 19014 4962 19066
rect 4962 19014 4974 19066
rect 4974 19014 4988 19066
rect 5012 19014 5026 19066
rect 5026 19014 5038 19066
rect 5038 19014 5068 19066
rect 5092 19014 5102 19066
rect 5102 19014 5148 19066
rect 4852 19012 4908 19014
rect 4932 19012 4988 19014
rect 5012 19012 5068 19014
rect 5092 19012 5148 19014
rect 4852 17978 4908 17980
rect 4932 17978 4988 17980
rect 5012 17978 5068 17980
rect 5092 17978 5148 17980
rect 4852 17926 4898 17978
rect 4898 17926 4908 17978
rect 4932 17926 4962 17978
rect 4962 17926 4974 17978
rect 4974 17926 4988 17978
rect 5012 17926 5026 17978
rect 5026 17926 5038 17978
rect 5038 17926 5068 17978
rect 5092 17926 5102 17978
rect 5102 17926 5148 17978
rect 4852 17924 4908 17926
rect 4932 17924 4988 17926
rect 5012 17924 5068 17926
rect 5092 17924 5148 17926
rect 4434 17604 4490 17640
rect 4434 17584 4436 17604
rect 4436 17584 4488 17604
rect 4488 17584 4490 17604
rect 5078 17448 5134 17504
rect 5262 17604 5318 17640
rect 5262 17584 5264 17604
rect 5264 17584 5316 17604
rect 5316 17584 5318 17604
rect 5354 17076 5356 17096
rect 5356 17076 5408 17096
rect 5408 17076 5410 17096
rect 5354 17040 5410 17076
rect 4852 16890 4908 16892
rect 4932 16890 4988 16892
rect 5012 16890 5068 16892
rect 5092 16890 5148 16892
rect 4852 16838 4898 16890
rect 4898 16838 4908 16890
rect 4932 16838 4962 16890
rect 4962 16838 4974 16890
rect 4974 16838 4988 16890
rect 5012 16838 5026 16890
rect 5026 16838 5038 16890
rect 5038 16838 5068 16890
rect 5092 16838 5102 16890
rect 5102 16838 5148 16890
rect 4852 16836 4908 16838
rect 4932 16836 4988 16838
rect 5012 16836 5068 16838
rect 5092 16836 5148 16838
rect 5814 19216 5870 19272
rect 6150 19610 6206 19612
rect 6230 19610 6286 19612
rect 6310 19610 6366 19612
rect 6390 19610 6446 19612
rect 6150 19558 6196 19610
rect 6196 19558 6206 19610
rect 6230 19558 6260 19610
rect 6260 19558 6272 19610
rect 6272 19558 6286 19610
rect 6310 19558 6324 19610
rect 6324 19558 6336 19610
rect 6336 19558 6366 19610
rect 6390 19558 6400 19610
rect 6400 19558 6446 19610
rect 6150 19556 6206 19558
rect 6230 19556 6286 19558
rect 6310 19556 6366 19558
rect 6390 19556 6446 19558
rect 6090 19352 6146 19408
rect 6826 19624 6882 19680
rect 5814 17040 5870 17096
rect 6150 18522 6206 18524
rect 6230 18522 6286 18524
rect 6310 18522 6366 18524
rect 6390 18522 6446 18524
rect 6150 18470 6196 18522
rect 6196 18470 6206 18522
rect 6230 18470 6260 18522
rect 6260 18470 6272 18522
rect 6272 18470 6286 18522
rect 6310 18470 6324 18522
rect 6324 18470 6336 18522
rect 6336 18470 6366 18522
rect 6390 18470 6400 18522
rect 6400 18470 6446 18522
rect 6150 18468 6206 18470
rect 6230 18468 6286 18470
rect 6310 18468 6366 18470
rect 6390 18468 6446 18470
rect 6150 17434 6206 17436
rect 6230 17434 6286 17436
rect 6310 17434 6366 17436
rect 6390 17434 6446 17436
rect 6150 17382 6196 17434
rect 6196 17382 6206 17434
rect 6230 17382 6260 17434
rect 6260 17382 6272 17434
rect 6272 17382 6286 17434
rect 6310 17382 6324 17434
rect 6324 17382 6336 17434
rect 6336 17382 6366 17434
rect 6390 17382 6400 17434
rect 6400 17382 6446 17434
rect 6150 17380 6206 17382
rect 6230 17380 6286 17382
rect 6310 17380 6366 17382
rect 6390 17380 6446 17382
rect 3553 15258 3609 15260
rect 3633 15258 3689 15260
rect 3713 15258 3769 15260
rect 3793 15258 3849 15260
rect 3553 15206 3599 15258
rect 3599 15206 3609 15258
rect 3633 15206 3663 15258
rect 3663 15206 3675 15258
rect 3675 15206 3689 15258
rect 3713 15206 3727 15258
rect 3727 15206 3739 15258
rect 3739 15206 3769 15258
rect 3793 15206 3803 15258
rect 3803 15206 3849 15258
rect 3553 15204 3609 15206
rect 3633 15204 3689 15206
rect 3713 15204 3769 15206
rect 3793 15204 3849 15206
rect 3553 14170 3609 14172
rect 3633 14170 3689 14172
rect 3713 14170 3769 14172
rect 3793 14170 3849 14172
rect 3553 14118 3599 14170
rect 3599 14118 3609 14170
rect 3633 14118 3663 14170
rect 3663 14118 3675 14170
rect 3675 14118 3689 14170
rect 3713 14118 3727 14170
rect 3727 14118 3739 14170
rect 3739 14118 3769 14170
rect 3793 14118 3803 14170
rect 3803 14118 3849 14170
rect 3553 14116 3609 14118
rect 3633 14116 3689 14118
rect 3713 14116 3769 14118
rect 3793 14116 3849 14118
rect 3054 12824 3110 12880
rect 3553 13082 3609 13084
rect 3633 13082 3689 13084
rect 3713 13082 3769 13084
rect 3793 13082 3849 13084
rect 3553 13030 3599 13082
rect 3599 13030 3609 13082
rect 3633 13030 3663 13082
rect 3663 13030 3675 13082
rect 3675 13030 3689 13082
rect 3713 13030 3727 13082
rect 3727 13030 3739 13082
rect 3739 13030 3769 13082
rect 3793 13030 3803 13082
rect 3803 13030 3849 13082
rect 3553 13028 3609 13030
rect 3633 13028 3689 13030
rect 3713 13028 3769 13030
rect 3793 13028 3849 13030
rect 3553 11994 3609 11996
rect 3633 11994 3689 11996
rect 3713 11994 3769 11996
rect 3793 11994 3849 11996
rect 3553 11942 3599 11994
rect 3599 11942 3609 11994
rect 3633 11942 3663 11994
rect 3663 11942 3675 11994
rect 3675 11942 3689 11994
rect 3713 11942 3727 11994
rect 3727 11942 3739 11994
rect 3739 11942 3769 11994
rect 3793 11942 3803 11994
rect 3803 11942 3849 11994
rect 3553 11940 3609 11942
rect 3633 11940 3689 11942
rect 3713 11940 3769 11942
rect 3793 11940 3849 11942
rect 3553 10906 3609 10908
rect 3633 10906 3689 10908
rect 3713 10906 3769 10908
rect 3793 10906 3849 10908
rect 3553 10854 3599 10906
rect 3599 10854 3609 10906
rect 3633 10854 3663 10906
rect 3663 10854 3675 10906
rect 3675 10854 3689 10906
rect 3713 10854 3727 10906
rect 3727 10854 3739 10906
rect 3739 10854 3769 10906
rect 3793 10854 3803 10906
rect 3803 10854 3849 10906
rect 3553 10852 3609 10854
rect 3633 10852 3689 10854
rect 3713 10852 3769 10854
rect 3793 10852 3849 10854
rect 2778 10648 2834 10704
rect 2686 10512 2742 10568
rect 2594 10104 2650 10160
rect 4852 15802 4908 15804
rect 4932 15802 4988 15804
rect 5012 15802 5068 15804
rect 5092 15802 5148 15804
rect 4852 15750 4898 15802
rect 4898 15750 4908 15802
rect 4932 15750 4962 15802
rect 4962 15750 4974 15802
rect 4974 15750 4988 15802
rect 5012 15750 5026 15802
rect 5026 15750 5038 15802
rect 5038 15750 5068 15802
rect 5092 15750 5102 15802
rect 5102 15750 5148 15802
rect 4852 15748 4908 15750
rect 4932 15748 4988 15750
rect 5012 15748 5068 15750
rect 5092 15748 5148 15750
rect 5722 15544 5778 15600
rect 6150 16346 6206 16348
rect 6230 16346 6286 16348
rect 6310 16346 6366 16348
rect 6390 16346 6446 16348
rect 6150 16294 6196 16346
rect 6196 16294 6206 16346
rect 6230 16294 6260 16346
rect 6260 16294 6272 16346
rect 6272 16294 6286 16346
rect 6310 16294 6324 16346
rect 6324 16294 6336 16346
rect 6336 16294 6366 16346
rect 6390 16294 6400 16346
rect 6400 16294 6446 16346
rect 6150 16292 6206 16294
rect 6230 16292 6286 16294
rect 6310 16292 6366 16294
rect 6390 16292 6446 16294
rect 7449 21242 7505 21244
rect 7529 21242 7585 21244
rect 7609 21242 7665 21244
rect 7689 21242 7745 21244
rect 7449 21190 7495 21242
rect 7495 21190 7505 21242
rect 7529 21190 7559 21242
rect 7559 21190 7571 21242
rect 7571 21190 7585 21242
rect 7609 21190 7623 21242
rect 7623 21190 7635 21242
rect 7635 21190 7665 21242
rect 7689 21190 7699 21242
rect 7699 21190 7745 21242
rect 7449 21188 7505 21190
rect 7529 21188 7585 21190
rect 7609 21188 7665 21190
rect 7689 21188 7745 21190
rect 8114 24268 8170 24304
rect 8114 24248 8116 24268
rect 8116 24248 8168 24268
rect 8168 24248 8170 24268
rect 8206 23704 8262 23760
rect 8114 22636 8170 22672
rect 8114 22616 8116 22636
rect 8116 22616 8168 22636
rect 8168 22616 8170 22636
rect 8114 22072 8170 22128
rect 7449 20154 7505 20156
rect 7529 20154 7585 20156
rect 7609 20154 7665 20156
rect 7689 20154 7745 20156
rect 7449 20102 7495 20154
rect 7495 20102 7505 20154
rect 7529 20102 7559 20154
rect 7559 20102 7571 20154
rect 7571 20102 7585 20154
rect 7609 20102 7623 20154
rect 7623 20102 7635 20154
rect 7635 20102 7665 20154
rect 7689 20102 7699 20154
rect 7699 20102 7745 20154
rect 7449 20100 7505 20102
rect 7529 20100 7585 20102
rect 7609 20100 7665 20102
rect 7689 20100 7745 20102
rect 8022 20984 8078 21040
rect 7449 19066 7505 19068
rect 7529 19066 7585 19068
rect 7609 19066 7665 19068
rect 7689 19066 7745 19068
rect 7449 19014 7495 19066
rect 7495 19014 7505 19066
rect 7529 19014 7559 19066
rect 7559 19014 7571 19066
rect 7571 19014 7585 19066
rect 7609 19014 7623 19066
rect 7623 19014 7635 19066
rect 7635 19014 7665 19066
rect 7689 19014 7699 19066
rect 7699 19014 7745 19066
rect 7449 19012 7505 19014
rect 7529 19012 7585 19014
rect 7609 19012 7665 19014
rect 7689 19012 7745 19014
rect 8206 20440 8262 20496
rect 6826 17312 6882 17368
rect 6550 16224 6606 16280
rect 2254 9274 2310 9276
rect 2334 9274 2390 9276
rect 2414 9274 2470 9276
rect 2494 9274 2550 9276
rect 2254 9222 2300 9274
rect 2300 9222 2310 9274
rect 2334 9222 2364 9274
rect 2364 9222 2376 9274
rect 2376 9222 2390 9274
rect 2414 9222 2428 9274
rect 2428 9222 2440 9274
rect 2440 9222 2470 9274
rect 2494 9222 2504 9274
rect 2504 9222 2550 9274
rect 2254 9220 2310 9222
rect 2334 9220 2390 9222
rect 2414 9220 2470 9222
rect 2494 9220 2550 9222
rect 2254 8186 2310 8188
rect 2334 8186 2390 8188
rect 2414 8186 2470 8188
rect 2494 8186 2550 8188
rect 2254 8134 2300 8186
rect 2300 8134 2310 8186
rect 2334 8134 2364 8186
rect 2364 8134 2376 8186
rect 2376 8134 2390 8186
rect 2414 8134 2428 8186
rect 2428 8134 2440 8186
rect 2440 8134 2470 8186
rect 2494 8134 2504 8186
rect 2504 8134 2550 8186
rect 2254 8132 2310 8134
rect 2334 8132 2390 8134
rect 2414 8132 2470 8134
rect 2494 8132 2550 8134
rect 2254 7098 2310 7100
rect 2334 7098 2390 7100
rect 2414 7098 2470 7100
rect 2494 7098 2550 7100
rect 2254 7046 2300 7098
rect 2300 7046 2310 7098
rect 2334 7046 2364 7098
rect 2364 7046 2376 7098
rect 2376 7046 2390 7098
rect 2414 7046 2428 7098
rect 2428 7046 2440 7098
rect 2440 7046 2470 7098
rect 2494 7046 2504 7098
rect 2504 7046 2550 7098
rect 2254 7044 2310 7046
rect 2334 7044 2390 7046
rect 2414 7044 2470 7046
rect 2494 7044 2550 7046
rect 2594 6160 2650 6216
rect 2254 6010 2310 6012
rect 2334 6010 2390 6012
rect 2414 6010 2470 6012
rect 2494 6010 2550 6012
rect 2254 5958 2300 6010
rect 2300 5958 2310 6010
rect 2334 5958 2364 6010
rect 2364 5958 2376 6010
rect 2376 5958 2390 6010
rect 2414 5958 2428 6010
rect 2428 5958 2440 6010
rect 2440 5958 2470 6010
rect 2494 5958 2504 6010
rect 2504 5958 2550 6010
rect 2254 5956 2310 5958
rect 2334 5956 2390 5958
rect 2414 5956 2470 5958
rect 2494 5956 2550 5958
rect 2254 4922 2310 4924
rect 2334 4922 2390 4924
rect 2414 4922 2470 4924
rect 2494 4922 2550 4924
rect 2254 4870 2300 4922
rect 2300 4870 2310 4922
rect 2334 4870 2364 4922
rect 2364 4870 2376 4922
rect 2376 4870 2390 4922
rect 2414 4870 2428 4922
rect 2428 4870 2440 4922
rect 2440 4870 2470 4922
rect 2494 4870 2504 4922
rect 2504 4870 2550 4922
rect 2254 4868 2310 4870
rect 2334 4868 2390 4870
rect 2414 4868 2470 4870
rect 2494 4868 2550 4870
rect 2254 3834 2310 3836
rect 2334 3834 2390 3836
rect 2414 3834 2470 3836
rect 2494 3834 2550 3836
rect 2254 3782 2300 3834
rect 2300 3782 2310 3834
rect 2334 3782 2364 3834
rect 2364 3782 2376 3834
rect 2376 3782 2390 3834
rect 2414 3782 2428 3834
rect 2428 3782 2440 3834
rect 2440 3782 2470 3834
rect 2494 3782 2504 3834
rect 2504 3782 2550 3834
rect 2254 3780 2310 3782
rect 2334 3780 2390 3782
rect 2414 3780 2470 3782
rect 2494 3780 2550 3782
rect 2254 2746 2310 2748
rect 2334 2746 2390 2748
rect 2414 2746 2470 2748
rect 2494 2746 2550 2748
rect 2254 2694 2300 2746
rect 2300 2694 2310 2746
rect 2334 2694 2364 2746
rect 2364 2694 2376 2746
rect 2376 2694 2390 2746
rect 2414 2694 2428 2746
rect 2428 2694 2440 2746
rect 2440 2694 2470 2746
rect 2494 2694 2504 2746
rect 2504 2694 2550 2746
rect 2254 2692 2310 2694
rect 2334 2692 2390 2694
rect 2414 2692 2470 2694
rect 2494 2692 2550 2694
rect 3553 9818 3609 9820
rect 3633 9818 3689 9820
rect 3713 9818 3769 9820
rect 3793 9818 3849 9820
rect 3553 9766 3599 9818
rect 3599 9766 3609 9818
rect 3633 9766 3663 9818
rect 3663 9766 3675 9818
rect 3675 9766 3689 9818
rect 3713 9766 3727 9818
rect 3727 9766 3739 9818
rect 3739 9766 3769 9818
rect 3793 9766 3803 9818
rect 3803 9766 3849 9818
rect 3553 9764 3609 9766
rect 3633 9764 3689 9766
rect 3713 9764 3769 9766
rect 3793 9764 3849 9766
rect 4852 14714 4908 14716
rect 4932 14714 4988 14716
rect 5012 14714 5068 14716
rect 5092 14714 5148 14716
rect 4852 14662 4898 14714
rect 4898 14662 4908 14714
rect 4932 14662 4962 14714
rect 4962 14662 4974 14714
rect 4974 14662 4988 14714
rect 5012 14662 5026 14714
rect 5026 14662 5038 14714
rect 5038 14662 5068 14714
rect 5092 14662 5102 14714
rect 5102 14662 5148 14714
rect 4852 14660 4908 14662
rect 4932 14660 4988 14662
rect 5012 14660 5068 14662
rect 5092 14660 5148 14662
rect 5262 13912 5318 13968
rect 4852 13626 4908 13628
rect 4932 13626 4988 13628
rect 5012 13626 5068 13628
rect 5092 13626 5148 13628
rect 4852 13574 4898 13626
rect 4898 13574 4908 13626
rect 4932 13574 4962 13626
rect 4962 13574 4974 13626
rect 4974 13574 4988 13626
rect 5012 13574 5026 13626
rect 5026 13574 5038 13626
rect 5038 13574 5068 13626
rect 5092 13574 5102 13626
rect 5102 13574 5148 13626
rect 4852 13572 4908 13574
rect 4932 13572 4988 13574
rect 5012 13572 5068 13574
rect 5092 13572 5148 13574
rect 4852 12538 4908 12540
rect 4932 12538 4988 12540
rect 5012 12538 5068 12540
rect 5092 12538 5148 12540
rect 4852 12486 4898 12538
rect 4898 12486 4908 12538
rect 4932 12486 4962 12538
rect 4962 12486 4974 12538
rect 4974 12486 4988 12538
rect 5012 12486 5026 12538
rect 5026 12486 5038 12538
rect 5038 12486 5068 12538
rect 5092 12486 5102 12538
rect 5102 12486 5148 12538
rect 4852 12484 4908 12486
rect 4932 12484 4988 12486
rect 5012 12484 5068 12486
rect 5092 12484 5148 12486
rect 4852 11450 4908 11452
rect 4932 11450 4988 11452
rect 5012 11450 5068 11452
rect 5092 11450 5148 11452
rect 4852 11398 4898 11450
rect 4898 11398 4908 11450
rect 4932 11398 4962 11450
rect 4962 11398 4974 11450
rect 4974 11398 4988 11450
rect 5012 11398 5026 11450
rect 5026 11398 5038 11450
rect 5038 11398 5068 11450
rect 5092 11398 5102 11450
rect 5102 11398 5148 11450
rect 4852 11396 4908 11398
rect 4932 11396 4988 11398
rect 5012 11396 5068 11398
rect 5092 11396 5148 11398
rect 3553 8730 3609 8732
rect 3633 8730 3689 8732
rect 3713 8730 3769 8732
rect 3793 8730 3849 8732
rect 3553 8678 3599 8730
rect 3599 8678 3609 8730
rect 3633 8678 3663 8730
rect 3663 8678 3675 8730
rect 3675 8678 3689 8730
rect 3713 8678 3727 8730
rect 3727 8678 3739 8730
rect 3739 8678 3769 8730
rect 3793 8678 3803 8730
rect 3803 8678 3849 8730
rect 3553 8676 3609 8678
rect 3633 8676 3689 8678
rect 3713 8676 3769 8678
rect 3793 8676 3849 8678
rect 4852 10362 4908 10364
rect 4932 10362 4988 10364
rect 5012 10362 5068 10364
rect 5092 10362 5148 10364
rect 4852 10310 4898 10362
rect 4898 10310 4908 10362
rect 4932 10310 4962 10362
rect 4962 10310 4974 10362
rect 4974 10310 4988 10362
rect 5012 10310 5026 10362
rect 5026 10310 5038 10362
rect 5038 10310 5068 10362
rect 5092 10310 5102 10362
rect 5102 10310 5148 10362
rect 4852 10308 4908 10310
rect 4932 10308 4988 10310
rect 5012 10308 5068 10310
rect 5092 10308 5148 10310
rect 3553 7642 3609 7644
rect 3633 7642 3689 7644
rect 3713 7642 3769 7644
rect 3793 7642 3849 7644
rect 3553 7590 3599 7642
rect 3599 7590 3609 7642
rect 3633 7590 3663 7642
rect 3663 7590 3675 7642
rect 3675 7590 3689 7642
rect 3713 7590 3727 7642
rect 3727 7590 3739 7642
rect 3739 7590 3769 7642
rect 3793 7590 3803 7642
rect 3803 7590 3849 7642
rect 3553 7588 3609 7590
rect 3633 7588 3689 7590
rect 3713 7588 3769 7590
rect 3793 7588 3849 7590
rect 3790 7284 3792 7304
rect 3792 7284 3844 7304
rect 3844 7284 3846 7304
rect 3790 7248 3846 7284
rect 3553 6554 3609 6556
rect 3633 6554 3689 6556
rect 3713 6554 3769 6556
rect 3793 6554 3849 6556
rect 3553 6502 3599 6554
rect 3599 6502 3609 6554
rect 3633 6502 3663 6554
rect 3663 6502 3675 6554
rect 3675 6502 3689 6554
rect 3713 6502 3727 6554
rect 3727 6502 3739 6554
rect 3739 6502 3769 6554
rect 3793 6502 3803 6554
rect 3803 6502 3849 6554
rect 3553 6500 3609 6502
rect 3633 6500 3689 6502
rect 3713 6500 3769 6502
rect 3793 6500 3849 6502
rect 3553 5466 3609 5468
rect 3633 5466 3689 5468
rect 3713 5466 3769 5468
rect 3793 5466 3849 5468
rect 3553 5414 3599 5466
rect 3599 5414 3609 5466
rect 3633 5414 3663 5466
rect 3663 5414 3675 5466
rect 3675 5414 3689 5466
rect 3713 5414 3727 5466
rect 3727 5414 3739 5466
rect 3739 5414 3769 5466
rect 3793 5414 3803 5466
rect 3803 5414 3849 5466
rect 3553 5412 3609 5414
rect 3633 5412 3689 5414
rect 3713 5412 3769 5414
rect 3793 5412 3849 5414
rect 3422 5072 3478 5128
rect 3553 4378 3609 4380
rect 3633 4378 3689 4380
rect 3713 4378 3769 4380
rect 3793 4378 3849 4380
rect 3553 4326 3599 4378
rect 3599 4326 3609 4378
rect 3633 4326 3663 4378
rect 3663 4326 3675 4378
rect 3675 4326 3689 4378
rect 3713 4326 3727 4378
rect 3727 4326 3739 4378
rect 3739 4326 3769 4378
rect 3793 4326 3803 4378
rect 3803 4326 3849 4378
rect 3553 4324 3609 4326
rect 3633 4324 3689 4326
rect 3713 4324 3769 4326
rect 3793 4324 3849 4326
rect 3553 3290 3609 3292
rect 3633 3290 3689 3292
rect 3713 3290 3769 3292
rect 3793 3290 3849 3292
rect 3553 3238 3599 3290
rect 3599 3238 3609 3290
rect 3633 3238 3663 3290
rect 3663 3238 3675 3290
rect 3675 3238 3689 3290
rect 3713 3238 3727 3290
rect 3727 3238 3739 3290
rect 3739 3238 3769 3290
rect 3793 3238 3803 3290
rect 3803 3238 3849 3290
rect 3553 3236 3609 3238
rect 3633 3236 3689 3238
rect 3713 3236 3769 3238
rect 3793 3236 3849 3238
rect 3553 2202 3609 2204
rect 3633 2202 3689 2204
rect 3713 2202 3769 2204
rect 3793 2202 3849 2204
rect 3553 2150 3599 2202
rect 3599 2150 3609 2202
rect 3633 2150 3663 2202
rect 3663 2150 3675 2202
rect 3675 2150 3689 2202
rect 3713 2150 3727 2202
rect 3727 2150 3739 2202
rect 3739 2150 3769 2202
rect 3793 2150 3803 2202
rect 3803 2150 3849 2202
rect 3553 2148 3609 2150
rect 3633 2148 3689 2150
rect 3713 2148 3769 2150
rect 3793 2148 3849 2150
rect 4852 9274 4908 9276
rect 4932 9274 4988 9276
rect 5012 9274 5068 9276
rect 5092 9274 5148 9276
rect 4852 9222 4898 9274
rect 4898 9222 4908 9274
rect 4932 9222 4962 9274
rect 4962 9222 4974 9274
rect 4974 9222 4988 9274
rect 5012 9222 5026 9274
rect 5026 9222 5038 9274
rect 5038 9222 5068 9274
rect 5092 9222 5102 9274
rect 5102 9222 5148 9274
rect 4852 9220 4908 9222
rect 4932 9220 4988 9222
rect 5012 9220 5068 9222
rect 5092 9220 5148 9222
rect 4852 8186 4908 8188
rect 4932 8186 4988 8188
rect 5012 8186 5068 8188
rect 5092 8186 5148 8188
rect 4852 8134 4898 8186
rect 4898 8134 4908 8186
rect 4932 8134 4962 8186
rect 4962 8134 4974 8186
rect 4974 8134 4988 8186
rect 5012 8134 5026 8186
rect 5026 8134 5038 8186
rect 5038 8134 5068 8186
rect 5092 8134 5102 8186
rect 5102 8134 5148 8186
rect 4852 8132 4908 8134
rect 4932 8132 4988 8134
rect 5012 8132 5068 8134
rect 5092 8132 5148 8134
rect 5814 14456 5870 14512
rect 6150 15258 6206 15260
rect 6230 15258 6286 15260
rect 6310 15258 6366 15260
rect 6390 15258 6446 15260
rect 6150 15206 6196 15258
rect 6196 15206 6206 15258
rect 6230 15206 6260 15258
rect 6260 15206 6272 15258
rect 6272 15206 6286 15258
rect 6310 15206 6324 15258
rect 6324 15206 6336 15258
rect 6336 15206 6366 15258
rect 6390 15206 6400 15258
rect 6400 15206 6446 15258
rect 6150 15204 6206 15206
rect 6230 15204 6286 15206
rect 6310 15204 6366 15206
rect 6390 15204 6446 15206
rect 6642 15136 6698 15192
rect 7194 18400 7250 18456
rect 7449 17978 7505 17980
rect 7529 17978 7585 17980
rect 7609 17978 7665 17980
rect 7689 17978 7745 17980
rect 7449 17926 7495 17978
rect 7495 17926 7505 17978
rect 7529 17926 7559 17978
rect 7559 17926 7571 17978
rect 7571 17926 7585 17978
rect 7609 17926 7623 17978
rect 7623 17926 7635 17978
rect 7635 17926 7665 17978
rect 7689 17926 7699 17978
rect 7699 17926 7745 17978
rect 7449 17924 7505 17926
rect 7529 17924 7585 17926
rect 7609 17924 7665 17926
rect 7689 17924 7745 17926
rect 7838 17856 7894 17912
rect 7449 16890 7505 16892
rect 7529 16890 7585 16892
rect 7609 16890 7665 16892
rect 7689 16890 7745 16892
rect 7449 16838 7495 16890
rect 7495 16838 7505 16890
rect 7529 16838 7559 16890
rect 7559 16838 7571 16890
rect 7571 16838 7585 16890
rect 7609 16838 7623 16890
rect 7623 16838 7635 16890
rect 7635 16838 7665 16890
rect 7689 16838 7699 16890
rect 7699 16838 7745 16890
rect 7449 16836 7505 16838
rect 7529 16836 7585 16838
rect 7609 16836 7665 16838
rect 7689 16836 7745 16838
rect 7449 15802 7505 15804
rect 7529 15802 7585 15804
rect 7609 15802 7665 15804
rect 7689 15802 7745 15804
rect 7449 15750 7495 15802
rect 7495 15750 7505 15802
rect 7529 15750 7559 15802
rect 7559 15750 7571 15802
rect 7571 15750 7585 15802
rect 7609 15750 7623 15802
rect 7623 15750 7635 15802
rect 7635 15750 7665 15802
rect 7689 15750 7699 15802
rect 7699 15750 7745 15802
rect 7449 15748 7505 15750
rect 7529 15748 7585 15750
rect 7609 15748 7665 15750
rect 7689 15748 7745 15750
rect 6150 14170 6206 14172
rect 6230 14170 6286 14172
rect 6310 14170 6366 14172
rect 6390 14170 6446 14172
rect 6150 14118 6196 14170
rect 6196 14118 6206 14170
rect 6230 14118 6260 14170
rect 6260 14118 6272 14170
rect 6272 14118 6286 14170
rect 6310 14118 6324 14170
rect 6324 14118 6336 14170
rect 6336 14118 6366 14170
rect 6390 14118 6400 14170
rect 6400 14118 6446 14170
rect 6150 14116 6206 14118
rect 6230 14116 6286 14118
rect 6310 14116 6366 14118
rect 6390 14116 6446 14118
rect 5630 10104 5686 10160
rect 4852 7098 4908 7100
rect 4932 7098 4988 7100
rect 5012 7098 5068 7100
rect 5092 7098 5148 7100
rect 4852 7046 4898 7098
rect 4898 7046 4908 7098
rect 4932 7046 4962 7098
rect 4962 7046 4974 7098
rect 4974 7046 4988 7098
rect 5012 7046 5026 7098
rect 5026 7046 5038 7098
rect 5038 7046 5068 7098
rect 5092 7046 5102 7098
rect 5102 7046 5148 7098
rect 4852 7044 4908 7046
rect 4932 7044 4988 7046
rect 5012 7044 5068 7046
rect 5092 7044 5148 7046
rect 4852 6010 4908 6012
rect 4932 6010 4988 6012
rect 5012 6010 5068 6012
rect 5092 6010 5148 6012
rect 4852 5958 4898 6010
rect 4898 5958 4908 6010
rect 4932 5958 4962 6010
rect 4962 5958 4974 6010
rect 4974 5958 4988 6010
rect 5012 5958 5026 6010
rect 5026 5958 5038 6010
rect 5038 5958 5068 6010
rect 5092 5958 5102 6010
rect 5102 5958 5148 6010
rect 4852 5956 4908 5958
rect 4932 5956 4988 5958
rect 5012 5956 5068 5958
rect 5092 5956 5148 5958
rect 4852 4922 4908 4924
rect 4932 4922 4988 4924
rect 5012 4922 5068 4924
rect 5092 4922 5148 4924
rect 4852 4870 4898 4922
rect 4898 4870 4908 4922
rect 4932 4870 4962 4922
rect 4962 4870 4974 4922
rect 4974 4870 4988 4922
rect 5012 4870 5026 4922
rect 5026 4870 5038 4922
rect 5038 4870 5068 4922
rect 5092 4870 5102 4922
rect 5102 4870 5148 4922
rect 4852 4868 4908 4870
rect 4932 4868 4988 4870
rect 5012 4868 5068 4870
rect 5092 4868 5148 4870
rect 4852 3834 4908 3836
rect 4932 3834 4988 3836
rect 5012 3834 5068 3836
rect 5092 3834 5148 3836
rect 4852 3782 4898 3834
rect 4898 3782 4908 3834
rect 4932 3782 4962 3834
rect 4962 3782 4974 3834
rect 4974 3782 4988 3834
rect 5012 3782 5026 3834
rect 5026 3782 5038 3834
rect 5038 3782 5068 3834
rect 5092 3782 5102 3834
rect 5102 3782 5148 3834
rect 4852 3780 4908 3782
rect 4932 3780 4988 3782
rect 5012 3780 5068 3782
rect 5092 3780 5148 3782
rect 4852 2746 4908 2748
rect 4932 2746 4988 2748
rect 5012 2746 5068 2748
rect 5092 2746 5148 2748
rect 4852 2694 4898 2746
rect 4898 2694 4908 2746
rect 4932 2694 4962 2746
rect 4962 2694 4974 2746
rect 4974 2694 4988 2746
rect 5012 2694 5026 2746
rect 5026 2694 5038 2746
rect 5038 2694 5068 2746
rect 5092 2694 5102 2746
rect 5102 2694 5148 2746
rect 4852 2692 4908 2694
rect 4932 2692 4988 2694
rect 5012 2692 5068 2694
rect 5092 2692 5148 2694
rect 5814 10648 5870 10704
rect 6150 13082 6206 13084
rect 6230 13082 6286 13084
rect 6310 13082 6366 13084
rect 6390 13082 6446 13084
rect 6150 13030 6196 13082
rect 6196 13030 6206 13082
rect 6230 13030 6260 13082
rect 6260 13030 6272 13082
rect 6272 13030 6286 13082
rect 6310 13030 6324 13082
rect 6324 13030 6336 13082
rect 6336 13030 6366 13082
rect 6390 13030 6400 13082
rect 6400 13030 6446 13082
rect 6150 13028 6206 13030
rect 6230 13028 6286 13030
rect 6310 13028 6366 13030
rect 6390 13028 6446 13030
rect 6642 12960 6698 13016
rect 6150 11994 6206 11996
rect 6230 11994 6286 11996
rect 6310 11994 6366 11996
rect 6390 11994 6446 11996
rect 6150 11942 6196 11994
rect 6196 11942 6206 11994
rect 6230 11942 6260 11994
rect 6260 11942 6272 11994
rect 6272 11942 6286 11994
rect 6310 11942 6324 11994
rect 6324 11942 6336 11994
rect 6336 11942 6366 11994
rect 6390 11942 6400 11994
rect 6400 11942 6446 11994
rect 6150 11940 6206 11942
rect 6230 11940 6286 11942
rect 6310 11940 6366 11942
rect 6390 11940 6446 11942
rect 7449 14714 7505 14716
rect 7529 14714 7585 14716
rect 7609 14714 7665 14716
rect 7689 14714 7745 14716
rect 7449 14662 7495 14714
rect 7495 14662 7505 14714
rect 7529 14662 7559 14714
rect 7559 14662 7571 14714
rect 7571 14662 7585 14714
rect 7609 14662 7623 14714
rect 7623 14662 7635 14714
rect 7635 14662 7665 14714
rect 7689 14662 7699 14714
rect 7699 14662 7745 14714
rect 7449 14660 7505 14662
rect 7529 14660 7585 14662
rect 7609 14660 7665 14662
rect 7689 14660 7745 14662
rect 7449 13626 7505 13628
rect 7529 13626 7585 13628
rect 7609 13626 7665 13628
rect 7689 13626 7745 13628
rect 7449 13574 7495 13626
rect 7495 13574 7505 13626
rect 7529 13574 7559 13626
rect 7559 13574 7571 13626
rect 7571 13574 7585 13626
rect 7609 13574 7623 13626
rect 7623 13574 7635 13626
rect 7635 13574 7665 13626
rect 7689 13574 7699 13626
rect 7699 13574 7745 13626
rect 7449 13572 7505 13574
rect 7529 13572 7585 13574
rect 7609 13572 7665 13574
rect 7689 13572 7745 13574
rect 7194 13368 7250 13424
rect 6826 12688 6882 12744
rect 6150 10906 6206 10908
rect 6230 10906 6286 10908
rect 6310 10906 6366 10908
rect 6390 10906 6446 10908
rect 6150 10854 6196 10906
rect 6196 10854 6206 10906
rect 6230 10854 6260 10906
rect 6260 10854 6272 10906
rect 6272 10854 6286 10906
rect 6310 10854 6324 10906
rect 6324 10854 6336 10906
rect 6336 10854 6366 10906
rect 6390 10854 6400 10906
rect 6400 10854 6446 10906
rect 6150 10852 6206 10854
rect 6230 10852 6286 10854
rect 6310 10852 6366 10854
rect 6390 10852 6446 10854
rect 6734 10512 6790 10568
rect 6150 9818 6206 9820
rect 6230 9818 6286 9820
rect 6310 9818 6366 9820
rect 6390 9818 6446 9820
rect 6150 9766 6196 9818
rect 6196 9766 6206 9818
rect 6230 9766 6260 9818
rect 6260 9766 6272 9818
rect 6272 9766 6286 9818
rect 6310 9766 6324 9818
rect 6324 9766 6336 9818
rect 6336 9766 6366 9818
rect 6390 9766 6400 9818
rect 6400 9766 6446 9818
rect 6150 9764 6206 9766
rect 6230 9764 6286 9766
rect 6310 9764 6366 9766
rect 6390 9764 6446 9766
rect 6182 9632 6238 9688
rect 6150 8730 6206 8732
rect 6230 8730 6286 8732
rect 6310 8730 6366 8732
rect 6390 8730 6446 8732
rect 6150 8678 6196 8730
rect 6196 8678 6206 8730
rect 6230 8678 6260 8730
rect 6260 8678 6272 8730
rect 6272 8678 6286 8730
rect 6310 8678 6324 8730
rect 6324 8678 6336 8730
rect 6336 8678 6366 8730
rect 6390 8678 6400 8730
rect 6400 8678 6446 8730
rect 6150 8676 6206 8678
rect 6230 8676 6286 8678
rect 6310 8676 6366 8678
rect 6390 8676 6446 8678
rect 5630 6160 5686 6216
rect 5722 5616 5778 5672
rect 6150 7642 6206 7644
rect 6230 7642 6286 7644
rect 6310 7642 6366 7644
rect 6390 7642 6446 7644
rect 6150 7590 6196 7642
rect 6196 7590 6206 7642
rect 6230 7590 6260 7642
rect 6260 7590 6272 7642
rect 6272 7590 6286 7642
rect 6310 7590 6324 7642
rect 6324 7590 6336 7642
rect 6336 7590 6366 7642
rect 6390 7590 6400 7642
rect 6400 7590 6446 7642
rect 6150 7588 6206 7590
rect 6230 7588 6286 7590
rect 6310 7588 6366 7590
rect 6390 7588 6446 7590
rect 6150 6554 6206 6556
rect 6230 6554 6286 6556
rect 6310 6554 6366 6556
rect 6390 6554 6446 6556
rect 6150 6502 6196 6554
rect 6196 6502 6206 6554
rect 6230 6502 6260 6554
rect 6260 6502 6272 6554
rect 6272 6502 6286 6554
rect 6310 6502 6324 6554
rect 6324 6502 6336 6554
rect 6336 6502 6366 6554
rect 6390 6502 6400 6554
rect 6400 6502 6446 6554
rect 6150 6500 6206 6502
rect 6230 6500 6286 6502
rect 6310 6500 6366 6502
rect 6390 6500 6446 6502
rect 6642 7928 6698 7984
rect 7194 12824 7250 12880
rect 7449 12538 7505 12540
rect 7529 12538 7585 12540
rect 7609 12538 7665 12540
rect 7689 12538 7745 12540
rect 7449 12486 7495 12538
rect 7495 12486 7505 12538
rect 7529 12486 7559 12538
rect 7559 12486 7571 12538
rect 7571 12486 7585 12538
rect 7609 12486 7623 12538
rect 7623 12486 7635 12538
rect 7635 12486 7665 12538
rect 7689 12486 7699 12538
rect 7699 12486 7745 12538
rect 7449 12484 7505 12486
rect 7529 12484 7585 12486
rect 7609 12484 7665 12486
rect 7689 12484 7745 12486
rect 7449 11450 7505 11452
rect 7529 11450 7585 11452
rect 7609 11450 7665 11452
rect 7689 11450 7745 11452
rect 7449 11398 7495 11450
rect 7495 11398 7505 11450
rect 7529 11398 7559 11450
rect 7559 11398 7571 11450
rect 7571 11398 7585 11450
rect 7609 11398 7623 11450
rect 7623 11398 7635 11450
rect 7635 11398 7665 11450
rect 7689 11398 7699 11450
rect 7699 11398 7745 11450
rect 7449 11396 7505 11398
rect 7529 11396 7585 11398
rect 7609 11396 7665 11398
rect 7689 11396 7745 11398
rect 7838 11328 7894 11384
rect 7378 10784 7434 10840
rect 7449 10362 7505 10364
rect 7529 10362 7585 10364
rect 7609 10362 7665 10364
rect 7689 10362 7745 10364
rect 7449 10310 7495 10362
rect 7495 10310 7505 10362
rect 7529 10310 7559 10362
rect 7559 10310 7571 10362
rect 7571 10310 7585 10362
rect 7609 10310 7623 10362
rect 7623 10310 7635 10362
rect 7635 10310 7665 10362
rect 7689 10310 7699 10362
rect 7699 10310 7745 10362
rect 7449 10308 7505 10310
rect 7529 10308 7585 10310
rect 7609 10308 7665 10310
rect 7689 10308 7745 10310
rect 7449 9274 7505 9276
rect 7529 9274 7585 9276
rect 7609 9274 7665 9276
rect 7689 9274 7745 9276
rect 7449 9222 7495 9274
rect 7495 9222 7505 9274
rect 7529 9222 7559 9274
rect 7559 9222 7571 9274
rect 7571 9222 7585 9274
rect 7609 9222 7623 9274
rect 7623 9222 7635 9274
rect 7635 9222 7665 9274
rect 7689 9222 7699 9274
rect 7699 9222 7745 9274
rect 7449 9220 7505 9222
rect 7529 9220 7585 9222
rect 7609 9220 7665 9222
rect 7689 9220 7745 9222
rect 8206 11872 8262 11928
rect 8114 10240 8170 10296
rect 6826 8744 6882 8800
rect 6150 5466 6206 5468
rect 6230 5466 6286 5468
rect 6310 5466 6366 5468
rect 6390 5466 6446 5468
rect 6150 5414 6196 5466
rect 6196 5414 6206 5466
rect 6230 5414 6260 5466
rect 6260 5414 6272 5466
rect 6272 5414 6286 5466
rect 6310 5414 6324 5466
rect 6324 5414 6336 5466
rect 6336 5414 6366 5466
rect 6390 5414 6400 5466
rect 6400 5414 6446 5466
rect 6150 5412 6206 5414
rect 6230 5412 6286 5414
rect 6310 5412 6366 5414
rect 6390 5412 6446 5414
rect 6150 4378 6206 4380
rect 6230 4378 6286 4380
rect 6310 4378 6366 4380
rect 6390 4378 6446 4380
rect 6150 4326 6196 4378
rect 6196 4326 6206 4378
rect 6230 4326 6260 4378
rect 6260 4326 6272 4378
rect 6272 4326 6286 4378
rect 6310 4326 6324 4378
rect 6324 4326 6336 4378
rect 6336 4326 6366 4378
rect 6390 4326 6400 4378
rect 6400 4326 6446 4378
rect 6150 4324 6206 4326
rect 6230 4324 6286 4326
rect 6310 4324 6366 4326
rect 6390 4324 6446 4326
rect 6150 3290 6206 3292
rect 6230 3290 6286 3292
rect 6310 3290 6366 3292
rect 6390 3290 6446 3292
rect 6150 3238 6196 3290
rect 6196 3238 6206 3290
rect 6230 3238 6260 3290
rect 6260 3238 6272 3290
rect 6272 3238 6286 3290
rect 6310 3238 6324 3290
rect 6324 3238 6336 3290
rect 6336 3238 6366 3290
rect 6390 3238 6400 3290
rect 6400 3238 6446 3290
rect 6150 3236 6206 3238
rect 6230 3236 6286 3238
rect 6310 3236 6366 3238
rect 6390 3236 6446 3238
rect 6642 2896 6698 2952
rect 6150 2202 6206 2204
rect 6230 2202 6286 2204
rect 6310 2202 6366 2204
rect 6390 2202 6446 2204
rect 6150 2150 6196 2202
rect 6196 2150 6206 2202
rect 6230 2150 6260 2202
rect 6260 2150 6272 2202
rect 6272 2150 6286 2202
rect 6310 2150 6324 2202
rect 6324 2150 6336 2202
rect 6336 2150 6366 2202
rect 6390 2150 6400 2202
rect 6400 2150 6446 2202
rect 6150 2148 6206 2150
rect 6230 2148 6286 2150
rect 6310 2148 6366 2150
rect 6390 2148 6446 2150
rect 6642 1672 6698 1728
rect 5998 1128 6054 1184
rect 6550 584 6606 640
rect 6642 176 6698 232
rect 7449 8186 7505 8188
rect 7529 8186 7585 8188
rect 7609 8186 7665 8188
rect 7689 8186 7745 8188
rect 7449 8134 7495 8186
rect 7495 8134 7505 8186
rect 7529 8134 7559 8186
rect 7559 8134 7571 8186
rect 7571 8134 7585 8186
rect 7609 8134 7623 8186
rect 7623 8134 7635 8186
rect 7635 8134 7665 8186
rect 7689 8134 7699 8186
rect 7699 8134 7745 8186
rect 7449 8132 7505 8134
rect 7529 8132 7585 8134
rect 7609 8132 7665 8134
rect 7689 8132 7745 8134
rect 8114 9324 8116 9344
rect 8116 9324 8168 9344
rect 8168 9324 8170 9344
rect 8114 9288 8170 9324
rect 8298 9832 8354 9888
rect 8206 8744 8262 8800
rect 7930 7656 7986 7712
rect 7838 7112 7894 7168
rect 7449 7098 7505 7100
rect 7529 7098 7585 7100
rect 7609 7098 7665 7100
rect 7689 7098 7745 7100
rect 7449 7046 7495 7098
rect 7495 7046 7505 7098
rect 7529 7046 7559 7098
rect 7559 7046 7571 7098
rect 7571 7046 7585 7098
rect 7609 7046 7623 7098
rect 7623 7046 7635 7098
rect 7635 7046 7665 7098
rect 7689 7046 7699 7098
rect 7699 7046 7745 7098
rect 7449 7044 7505 7046
rect 7529 7044 7585 7046
rect 7609 7044 7665 7046
rect 7689 7044 7745 7046
rect 7930 6568 7986 6624
rect 7449 6010 7505 6012
rect 7529 6010 7585 6012
rect 7609 6010 7665 6012
rect 7689 6010 7745 6012
rect 7449 5958 7495 6010
rect 7495 5958 7505 6010
rect 7529 5958 7559 6010
rect 7559 5958 7571 6010
rect 7571 5958 7585 6010
rect 7609 5958 7623 6010
rect 7623 5958 7635 6010
rect 7635 5958 7665 6010
rect 7689 5958 7699 6010
rect 7699 5958 7745 6010
rect 7449 5956 7505 5958
rect 7529 5956 7585 5958
rect 7609 5956 7665 5958
rect 7689 5956 7745 5958
rect 6826 3984 6882 4040
rect 7449 4922 7505 4924
rect 7529 4922 7585 4924
rect 7609 4922 7665 4924
rect 7689 4922 7745 4924
rect 7449 4870 7495 4922
rect 7495 4870 7505 4922
rect 7529 4870 7559 4922
rect 7559 4870 7571 4922
rect 7571 4870 7585 4922
rect 7609 4870 7623 4922
rect 7623 4870 7635 4922
rect 7635 4870 7665 4922
rect 7689 4870 7699 4922
rect 7699 4870 7745 4922
rect 7449 4868 7505 4870
rect 7529 4868 7585 4870
rect 7609 4868 7665 4870
rect 7689 4868 7745 4870
rect 7449 3834 7505 3836
rect 7529 3834 7585 3836
rect 7609 3834 7665 3836
rect 7689 3834 7745 3836
rect 7449 3782 7495 3834
rect 7495 3782 7505 3834
rect 7529 3782 7559 3834
rect 7559 3782 7571 3834
rect 7571 3782 7585 3834
rect 7609 3782 7623 3834
rect 7623 3782 7635 3834
rect 7635 3782 7665 3834
rect 7689 3782 7699 3834
rect 7699 3782 7745 3834
rect 7449 3780 7505 3782
rect 7529 3780 7585 3782
rect 7609 3780 7665 3782
rect 7689 3780 7745 3782
rect 7449 2746 7505 2748
rect 7529 2746 7585 2748
rect 7609 2746 7665 2748
rect 7689 2746 7745 2748
rect 7449 2694 7495 2746
rect 7495 2694 7505 2746
rect 7529 2694 7559 2746
rect 7559 2694 7571 2746
rect 7571 2694 7585 2746
rect 7609 2694 7623 2746
rect 7623 2694 7635 2746
rect 7635 2694 7665 2746
rect 7689 2694 7699 2746
rect 7699 2694 7745 2746
rect 7449 2692 7505 2694
rect 7529 2692 7585 2694
rect 7609 2692 7665 2694
rect 7689 2692 7745 2694
rect 7930 4936 7986 4992
rect 8114 6024 8170 6080
rect 8206 5516 8208 5536
rect 8208 5516 8260 5536
rect 8260 5516 8262 5536
rect 8206 5480 8262 5516
rect 8298 4392 8354 4448
rect 8206 3304 8262 3360
rect 8022 2216 8078 2272
<< metal3 >>
rect 6637 29746 6703 29749
rect 9200 29746 10000 29776
rect 6637 29744 10000 29746
rect 6637 29688 6642 29744
rect 6698 29688 10000 29744
rect 6637 29686 10000 29688
rect 6637 29683 6703 29686
rect 9200 29656 10000 29686
rect 6545 29202 6611 29205
rect 9200 29202 10000 29232
rect 6545 29200 10000 29202
rect 6545 29144 6550 29200
rect 6606 29144 10000 29200
rect 6545 29142 10000 29144
rect 6545 29139 6611 29142
rect 9200 29112 10000 29142
rect 5533 28658 5599 28661
rect 9200 28658 10000 28688
rect 5533 28656 10000 28658
rect 5533 28600 5538 28656
rect 5594 28600 10000 28656
rect 5533 28598 10000 28600
rect 5533 28595 5599 28598
rect 9200 28568 10000 28598
rect 5993 28114 6059 28117
rect 9200 28114 10000 28144
rect 5993 28112 10000 28114
rect 5993 28056 5998 28112
rect 6054 28056 10000 28112
rect 5993 28054 10000 28056
rect 5993 28051 6059 28054
rect 9200 28024 10000 28054
rect 2242 27776 2562 27777
rect 2242 27712 2250 27776
rect 2314 27712 2330 27776
rect 2394 27712 2410 27776
rect 2474 27712 2490 27776
rect 2554 27712 2562 27776
rect 2242 27711 2562 27712
rect 4840 27776 5160 27777
rect 4840 27712 4848 27776
rect 4912 27712 4928 27776
rect 4992 27712 5008 27776
rect 5072 27712 5088 27776
rect 5152 27712 5160 27776
rect 4840 27711 5160 27712
rect 7437 27776 7757 27777
rect 7437 27712 7445 27776
rect 7509 27712 7525 27776
rect 7589 27712 7605 27776
rect 7669 27712 7685 27776
rect 7749 27712 7757 27776
rect 7437 27711 7757 27712
rect 5901 27570 5967 27573
rect 9200 27570 10000 27600
rect 5901 27568 10000 27570
rect 5901 27512 5906 27568
rect 5962 27512 10000 27568
rect 5901 27510 10000 27512
rect 5901 27507 5967 27510
rect 9200 27480 10000 27510
rect 3541 27232 3861 27233
rect 3541 27168 3549 27232
rect 3613 27168 3629 27232
rect 3693 27168 3709 27232
rect 3773 27168 3789 27232
rect 3853 27168 3861 27232
rect 3541 27167 3861 27168
rect 6138 27232 6458 27233
rect 6138 27168 6146 27232
rect 6210 27168 6226 27232
rect 6290 27168 6306 27232
rect 6370 27168 6386 27232
rect 6450 27168 6458 27232
rect 6138 27167 6458 27168
rect 5717 27026 5783 27029
rect 9200 27026 10000 27056
rect 5717 27024 10000 27026
rect 5717 26968 5722 27024
rect 5778 26968 10000 27024
rect 5717 26966 10000 26968
rect 5717 26963 5783 26966
rect 9200 26936 10000 26966
rect 2242 26688 2562 26689
rect 2242 26624 2250 26688
rect 2314 26624 2330 26688
rect 2394 26624 2410 26688
rect 2474 26624 2490 26688
rect 2554 26624 2562 26688
rect 2242 26623 2562 26624
rect 4840 26688 5160 26689
rect 4840 26624 4848 26688
rect 4912 26624 4928 26688
rect 4992 26624 5008 26688
rect 5072 26624 5088 26688
rect 5152 26624 5160 26688
rect 4840 26623 5160 26624
rect 7437 26688 7757 26689
rect 7437 26624 7445 26688
rect 7509 26624 7525 26688
rect 7589 26624 7605 26688
rect 7669 26624 7685 26688
rect 7749 26624 7757 26688
rect 7437 26623 7757 26624
rect 6729 26482 6795 26485
rect 9200 26482 10000 26512
rect 6729 26480 10000 26482
rect 6729 26424 6734 26480
rect 6790 26424 10000 26480
rect 6729 26422 10000 26424
rect 6729 26419 6795 26422
rect 9200 26392 10000 26422
rect 3541 26144 3861 26145
rect 3541 26080 3549 26144
rect 3613 26080 3629 26144
rect 3693 26080 3709 26144
rect 3773 26080 3789 26144
rect 3853 26080 3861 26144
rect 3541 26079 3861 26080
rect 6138 26144 6458 26145
rect 6138 26080 6146 26144
rect 6210 26080 6226 26144
rect 6290 26080 6306 26144
rect 6370 26080 6386 26144
rect 6450 26080 6458 26144
rect 6138 26079 6458 26080
rect 6637 25938 6703 25941
rect 9200 25938 10000 25968
rect 6637 25936 10000 25938
rect 6637 25880 6642 25936
rect 6698 25880 10000 25936
rect 6637 25878 10000 25880
rect 6637 25875 6703 25878
rect 9200 25848 10000 25878
rect 2242 25600 2562 25601
rect 2242 25536 2250 25600
rect 2314 25536 2330 25600
rect 2394 25536 2410 25600
rect 2474 25536 2490 25600
rect 2554 25536 2562 25600
rect 2242 25535 2562 25536
rect 4840 25600 5160 25601
rect 4840 25536 4848 25600
rect 4912 25536 4928 25600
rect 4992 25536 5008 25600
rect 5072 25536 5088 25600
rect 5152 25536 5160 25600
rect 4840 25535 5160 25536
rect 7437 25600 7757 25601
rect 7437 25536 7445 25600
rect 7509 25536 7525 25600
rect 7589 25536 7605 25600
rect 7669 25536 7685 25600
rect 7749 25536 7757 25600
rect 7437 25535 7757 25536
rect 7833 25394 7899 25397
rect 9200 25394 10000 25424
rect 7833 25392 10000 25394
rect 7833 25336 7838 25392
rect 7894 25336 10000 25392
rect 7833 25334 10000 25336
rect 7833 25331 7899 25334
rect 9200 25304 10000 25334
rect 3541 25056 3861 25057
rect 3541 24992 3549 25056
rect 3613 24992 3629 25056
rect 3693 24992 3709 25056
rect 3773 24992 3789 25056
rect 3853 24992 3861 25056
rect 3541 24991 3861 24992
rect 6138 25056 6458 25057
rect 6138 24992 6146 25056
rect 6210 24992 6226 25056
rect 6290 24992 6306 25056
rect 6370 24992 6386 25056
rect 6450 24992 6458 25056
rect 6138 24991 6458 24992
rect 7925 24850 7991 24853
rect 9200 24850 10000 24880
rect 7925 24848 10000 24850
rect 7925 24792 7930 24848
rect 7986 24792 10000 24848
rect 7925 24790 10000 24792
rect 7925 24787 7991 24790
rect 9200 24760 10000 24790
rect 2242 24512 2562 24513
rect 2242 24448 2250 24512
rect 2314 24448 2330 24512
rect 2394 24448 2410 24512
rect 2474 24448 2490 24512
rect 2554 24448 2562 24512
rect 2242 24447 2562 24448
rect 4840 24512 5160 24513
rect 4840 24448 4848 24512
rect 4912 24448 4928 24512
rect 4992 24448 5008 24512
rect 5072 24448 5088 24512
rect 5152 24448 5160 24512
rect 4840 24447 5160 24448
rect 7437 24512 7757 24513
rect 7437 24448 7445 24512
rect 7509 24448 7525 24512
rect 7589 24448 7605 24512
rect 7669 24448 7685 24512
rect 7749 24448 7757 24512
rect 7437 24447 7757 24448
rect 8109 24306 8175 24309
rect 9200 24306 10000 24336
rect 8109 24304 10000 24306
rect 8109 24248 8114 24304
rect 8170 24248 10000 24304
rect 8109 24246 10000 24248
rect 8109 24243 8175 24246
rect 9200 24216 10000 24246
rect 3541 23968 3861 23969
rect 3541 23904 3549 23968
rect 3613 23904 3629 23968
rect 3693 23904 3709 23968
rect 3773 23904 3789 23968
rect 3853 23904 3861 23968
rect 3541 23903 3861 23904
rect 6138 23968 6458 23969
rect 6138 23904 6146 23968
rect 6210 23904 6226 23968
rect 6290 23904 6306 23968
rect 6370 23904 6386 23968
rect 6450 23904 6458 23968
rect 6138 23903 6458 23904
rect 8201 23762 8267 23765
rect 9200 23762 10000 23792
rect 8201 23760 10000 23762
rect 8201 23704 8206 23760
rect 8262 23704 10000 23760
rect 8201 23702 10000 23704
rect 8201 23699 8267 23702
rect 9200 23672 10000 23702
rect 2242 23424 2562 23425
rect 2242 23360 2250 23424
rect 2314 23360 2330 23424
rect 2394 23360 2410 23424
rect 2474 23360 2490 23424
rect 2554 23360 2562 23424
rect 2242 23359 2562 23360
rect 4840 23424 5160 23425
rect 4840 23360 4848 23424
rect 4912 23360 4928 23424
rect 4992 23360 5008 23424
rect 5072 23360 5088 23424
rect 5152 23360 5160 23424
rect 4840 23359 5160 23360
rect 7437 23424 7757 23425
rect 7437 23360 7445 23424
rect 7509 23360 7525 23424
rect 7589 23360 7605 23424
rect 7669 23360 7685 23424
rect 7749 23360 7757 23424
rect 7437 23359 7757 23360
rect 6729 23218 6795 23221
rect 9200 23218 10000 23248
rect 6729 23216 10000 23218
rect 6729 23160 6734 23216
rect 6790 23160 10000 23216
rect 6729 23158 10000 23160
rect 6729 23155 6795 23158
rect 9200 23128 10000 23158
rect 3541 22880 3861 22881
rect 3541 22816 3549 22880
rect 3613 22816 3629 22880
rect 3693 22816 3709 22880
rect 3773 22816 3789 22880
rect 3853 22816 3861 22880
rect 3541 22815 3861 22816
rect 6138 22880 6458 22881
rect 6138 22816 6146 22880
rect 6210 22816 6226 22880
rect 6290 22816 6306 22880
rect 6370 22816 6386 22880
rect 6450 22816 6458 22880
rect 6138 22815 6458 22816
rect 8109 22674 8175 22677
rect 9200 22674 10000 22704
rect 8109 22672 10000 22674
rect 8109 22616 8114 22672
rect 8170 22616 10000 22672
rect 8109 22614 10000 22616
rect 8109 22611 8175 22614
rect 9200 22584 10000 22614
rect 2242 22336 2562 22337
rect 2242 22272 2250 22336
rect 2314 22272 2330 22336
rect 2394 22272 2410 22336
rect 2474 22272 2490 22336
rect 2554 22272 2562 22336
rect 2242 22271 2562 22272
rect 4840 22336 5160 22337
rect 4840 22272 4848 22336
rect 4912 22272 4928 22336
rect 4992 22272 5008 22336
rect 5072 22272 5088 22336
rect 5152 22272 5160 22336
rect 4840 22271 5160 22272
rect 7437 22336 7757 22337
rect 7437 22272 7445 22336
rect 7509 22272 7525 22336
rect 7589 22272 7605 22336
rect 7669 22272 7685 22336
rect 7749 22272 7757 22336
rect 7437 22271 7757 22272
rect 8109 22130 8175 22133
rect 9200 22130 10000 22160
rect 8109 22128 10000 22130
rect 8109 22072 8114 22128
rect 8170 22072 10000 22128
rect 8109 22070 10000 22072
rect 8109 22067 8175 22070
rect 9200 22040 10000 22070
rect 3541 21792 3861 21793
rect 3541 21728 3549 21792
rect 3613 21728 3629 21792
rect 3693 21728 3709 21792
rect 3773 21728 3789 21792
rect 3853 21728 3861 21792
rect 3541 21727 3861 21728
rect 6138 21792 6458 21793
rect 6138 21728 6146 21792
rect 6210 21728 6226 21792
rect 6290 21728 6306 21792
rect 6370 21728 6386 21792
rect 6450 21728 6458 21792
rect 6138 21727 6458 21728
rect 6729 21586 6795 21589
rect 9200 21586 10000 21616
rect 6729 21584 10000 21586
rect 6729 21528 6734 21584
rect 6790 21528 10000 21584
rect 6729 21526 10000 21528
rect 6729 21523 6795 21526
rect 9200 21496 10000 21526
rect 2242 21248 2562 21249
rect 2242 21184 2250 21248
rect 2314 21184 2330 21248
rect 2394 21184 2410 21248
rect 2474 21184 2490 21248
rect 2554 21184 2562 21248
rect 2242 21183 2562 21184
rect 4840 21248 5160 21249
rect 4840 21184 4848 21248
rect 4912 21184 4928 21248
rect 4992 21184 5008 21248
rect 5072 21184 5088 21248
rect 5152 21184 5160 21248
rect 4840 21183 5160 21184
rect 7437 21248 7757 21249
rect 7437 21184 7445 21248
rect 7509 21184 7525 21248
rect 7589 21184 7605 21248
rect 7669 21184 7685 21248
rect 7749 21184 7757 21248
rect 7437 21183 7757 21184
rect 8017 21042 8083 21045
rect 9200 21042 10000 21072
rect 8017 21040 10000 21042
rect 8017 20984 8022 21040
rect 8078 20984 10000 21040
rect 8017 20982 10000 20984
rect 8017 20979 8083 20982
rect 9200 20952 10000 20982
rect 3541 20704 3861 20705
rect 3541 20640 3549 20704
rect 3613 20640 3629 20704
rect 3693 20640 3709 20704
rect 3773 20640 3789 20704
rect 3853 20640 3861 20704
rect 3541 20639 3861 20640
rect 6138 20704 6458 20705
rect 6138 20640 6146 20704
rect 6210 20640 6226 20704
rect 6290 20640 6306 20704
rect 6370 20640 6386 20704
rect 6450 20640 6458 20704
rect 6138 20639 6458 20640
rect 8201 20498 8267 20501
rect 9200 20498 10000 20528
rect 8201 20496 10000 20498
rect 8201 20440 8206 20496
rect 8262 20440 10000 20496
rect 8201 20438 10000 20440
rect 8201 20435 8267 20438
rect 9200 20408 10000 20438
rect 2242 20160 2562 20161
rect 2242 20096 2250 20160
rect 2314 20096 2330 20160
rect 2394 20096 2410 20160
rect 2474 20096 2490 20160
rect 2554 20096 2562 20160
rect 2242 20095 2562 20096
rect 4840 20160 5160 20161
rect 4840 20096 4848 20160
rect 4912 20096 4928 20160
rect 4992 20096 5008 20160
rect 5072 20096 5088 20160
rect 5152 20096 5160 20160
rect 4840 20095 5160 20096
rect 7437 20160 7757 20161
rect 7437 20096 7445 20160
rect 7509 20096 7525 20160
rect 7589 20096 7605 20160
rect 7669 20096 7685 20160
rect 7749 20096 7757 20160
rect 7437 20095 7757 20096
rect 9200 20090 10000 20120
rect 7974 20030 10000 20090
rect 6821 19682 6887 19685
rect 7974 19682 8034 20030
rect 9200 20000 10000 20030
rect 6821 19680 8034 19682
rect 6821 19624 6826 19680
rect 6882 19624 8034 19680
rect 6821 19622 8034 19624
rect 6821 19619 6887 19622
rect 3541 19616 3861 19617
rect 3541 19552 3549 19616
rect 3613 19552 3629 19616
rect 3693 19552 3709 19616
rect 3773 19552 3789 19616
rect 3853 19552 3861 19616
rect 3541 19551 3861 19552
rect 6138 19616 6458 19617
rect 6138 19552 6146 19616
rect 6210 19552 6226 19616
rect 6290 19552 6306 19616
rect 6370 19552 6386 19616
rect 6450 19552 6458 19616
rect 6138 19551 6458 19552
rect 9200 19546 10000 19576
rect 6686 19486 10000 19546
rect 6085 19410 6151 19413
rect 6686 19410 6746 19486
rect 9200 19456 10000 19486
rect 6085 19408 6746 19410
rect 6085 19352 6090 19408
rect 6146 19352 6746 19408
rect 6085 19350 6746 19352
rect 6085 19347 6151 19350
rect 5809 19274 5875 19277
rect 5809 19272 8034 19274
rect 5809 19216 5814 19272
rect 5870 19216 8034 19272
rect 5809 19214 8034 19216
rect 5809 19211 5875 19214
rect 2242 19072 2562 19073
rect 2242 19008 2250 19072
rect 2314 19008 2330 19072
rect 2394 19008 2410 19072
rect 2474 19008 2490 19072
rect 2554 19008 2562 19072
rect 2242 19007 2562 19008
rect 4840 19072 5160 19073
rect 4840 19008 4848 19072
rect 4912 19008 4928 19072
rect 4992 19008 5008 19072
rect 5072 19008 5088 19072
rect 5152 19008 5160 19072
rect 4840 19007 5160 19008
rect 7437 19072 7757 19073
rect 7437 19008 7445 19072
rect 7509 19008 7525 19072
rect 7589 19008 7605 19072
rect 7669 19008 7685 19072
rect 7749 19008 7757 19072
rect 7437 19007 7757 19008
rect 7974 19002 8034 19214
rect 9200 19002 10000 19032
rect 7974 18942 10000 19002
rect 9200 18912 10000 18942
rect 3541 18528 3861 18529
rect 3541 18464 3549 18528
rect 3613 18464 3629 18528
rect 3693 18464 3709 18528
rect 3773 18464 3789 18528
rect 3853 18464 3861 18528
rect 3541 18463 3861 18464
rect 6138 18528 6458 18529
rect 6138 18464 6146 18528
rect 6210 18464 6226 18528
rect 6290 18464 6306 18528
rect 6370 18464 6386 18528
rect 6450 18464 6458 18528
rect 6138 18463 6458 18464
rect 7189 18458 7255 18461
rect 9200 18458 10000 18488
rect 7189 18456 10000 18458
rect 7189 18400 7194 18456
rect 7250 18400 10000 18456
rect 7189 18398 10000 18400
rect 7189 18395 7255 18398
rect 9200 18368 10000 18398
rect 2242 17984 2562 17985
rect 2242 17920 2250 17984
rect 2314 17920 2330 17984
rect 2394 17920 2410 17984
rect 2474 17920 2490 17984
rect 2554 17920 2562 17984
rect 2242 17919 2562 17920
rect 4840 17984 5160 17985
rect 4840 17920 4848 17984
rect 4912 17920 4928 17984
rect 4992 17920 5008 17984
rect 5072 17920 5088 17984
rect 5152 17920 5160 17984
rect 4840 17919 5160 17920
rect 7437 17984 7757 17985
rect 7437 17920 7445 17984
rect 7509 17920 7525 17984
rect 7589 17920 7605 17984
rect 7669 17920 7685 17984
rect 7749 17920 7757 17984
rect 7437 17919 7757 17920
rect 7833 17914 7899 17917
rect 9200 17914 10000 17944
rect 7833 17912 10000 17914
rect 7833 17856 7838 17912
rect 7894 17856 10000 17912
rect 7833 17854 10000 17856
rect 7833 17851 7899 17854
rect 9200 17824 10000 17854
rect 4429 17642 4495 17645
rect 5257 17642 5323 17645
rect 4429 17640 5323 17642
rect 4429 17584 4434 17640
rect 4490 17584 5262 17640
rect 5318 17584 5323 17640
rect 4429 17582 5323 17584
rect 4429 17579 4495 17582
rect 5257 17579 5323 17582
rect 4061 17506 4127 17509
rect 5073 17506 5139 17509
rect 4061 17504 5139 17506
rect 4061 17448 4066 17504
rect 4122 17448 5078 17504
rect 5134 17448 5139 17504
rect 4061 17446 5139 17448
rect 4061 17443 4127 17446
rect 5073 17443 5139 17446
rect 3541 17440 3861 17441
rect 3541 17376 3549 17440
rect 3613 17376 3629 17440
rect 3693 17376 3709 17440
rect 3773 17376 3789 17440
rect 3853 17376 3861 17440
rect 3541 17375 3861 17376
rect 6138 17440 6458 17441
rect 6138 17376 6146 17440
rect 6210 17376 6226 17440
rect 6290 17376 6306 17440
rect 6370 17376 6386 17440
rect 6450 17376 6458 17440
rect 6138 17375 6458 17376
rect 6821 17370 6887 17373
rect 9200 17370 10000 17400
rect 6821 17368 10000 17370
rect 6821 17312 6826 17368
rect 6882 17312 10000 17368
rect 6821 17310 10000 17312
rect 6821 17307 6887 17310
rect 9200 17280 10000 17310
rect 2589 17098 2655 17101
rect 5349 17098 5415 17101
rect 2589 17096 5415 17098
rect 2589 17040 2594 17096
rect 2650 17040 5354 17096
rect 5410 17040 5415 17096
rect 2589 17038 5415 17040
rect 2589 17035 2655 17038
rect 5349 17035 5415 17038
rect 5809 17098 5875 17101
rect 5809 17096 8034 17098
rect 5809 17040 5814 17096
rect 5870 17040 8034 17096
rect 5809 17038 8034 17040
rect 5809 17035 5875 17038
rect 2242 16896 2562 16897
rect 2242 16832 2250 16896
rect 2314 16832 2330 16896
rect 2394 16832 2410 16896
rect 2474 16832 2490 16896
rect 2554 16832 2562 16896
rect 2242 16831 2562 16832
rect 4840 16896 5160 16897
rect 4840 16832 4848 16896
rect 4912 16832 4928 16896
rect 4992 16832 5008 16896
rect 5072 16832 5088 16896
rect 5152 16832 5160 16896
rect 4840 16831 5160 16832
rect 7437 16896 7757 16897
rect 7437 16832 7445 16896
rect 7509 16832 7525 16896
rect 7589 16832 7605 16896
rect 7669 16832 7685 16896
rect 7749 16832 7757 16896
rect 7437 16831 7757 16832
rect 7974 16826 8034 17038
rect 9200 16826 10000 16856
rect 7974 16766 10000 16826
rect 9200 16736 10000 16766
rect 3541 16352 3861 16353
rect 3541 16288 3549 16352
rect 3613 16288 3629 16352
rect 3693 16288 3709 16352
rect 3773 16288 3789 16352
rect 3853 16288 3861 16352
rect 3541 16287 3861 16288
rect 6138 16352 6458 16353
rect 6138 16288 6146 16352
rect 6210 16288 6226 16352
rect 6290 16288 6306 16352
rect 6370 16288 6386 16352
rect 6450 16288 6458 16352
rect 6138 16287 6458 16288
rect 6545 16282 6611 16285
rect 9200 16282 10000 16312
rect 6545 16280 10000 16282
rect 6545 16224 6550 16280
rect 6606 16224 10000 16280
rect 6545 16222 10000 16224
rect 6545 16219 6611 16222
rect 9200 16192 10000 16222
rect 2242 15808 2562 15809
rect 2242 15744 2250 15808
rect 2314 15744 2330 15808
rect 2394 15744 2410 15808
rect 2474 15744 2490 15808
rect 2554 15744 2562 15808
rect 2242 15743 2562 15744
rect 4840 15808 5160 15809
rect 4840 15744 4848 15808
rect 4912 15744 4928 15808
rect 4992 15744 5008 15808
rect 5072 15744 5088 15808
rect 5152 15744 5160 15808
rect 4840 15743 5160 15744
rect 7437 15808 7757 15809
rect 7437 15744 7445 15808
rect 7509 15744 7525 15808
rect 7589 15744 7605 15808
rect 7669 15744 7685 15808
rect 7749 15744 7757 15808
rect 7437 15743 7757 15744
rect 9200 15738 10000 15768
rect 7974 15678 10000 15738
rect 5717 15602 5783 15605
rect 7974 15602 8034 15678
rect 9200 15648 10000 15678
rect 5717 15600 8034 15602
rect 5717 15544 5722 15600
rect 5778 15544 8034 15600
rect 5717 15542 8034 15544
rect 5717 15539 5783 15542
rect 3541 15264 3861 15265
rect 3541 15200 3549 15264
rect 3613 15200 3629 15264
rect 3693 15200 3709 15264
rect 3773 15200 3789 15264
rect 3853 15200 3861 15264
rect 3541 15199 3861 15200
rect 6138 15264 6458 15265
rect 6138 15200 6146 15264
rect 6210 15200 6226 15264
rect 6290 15200 6306 15264
rect 6370 15200 6386 15264
rect 6450 15200 6458 15264
rect 6138 15199 6458 15200
rect 6637 15194 6703 15197
rect 9200 15194 10000 15224
rect 6637 15192 10000 15194
rect 6637 15136 6642 15192
rect 6698 15136 10000 15192
rect 6637 15134 10000 15136
rect 6637 15131 6703 15134
rect 9200 15104 10000 15134
rect 2242 14720 2562 14721
rect 2242 14656 2250 14720
rect 2314 14656 2330 14720
rect 2394 14656 2410 14720
rect 2474 14656 2490 14720
rect 2554 14656 2562 14720
rect 2242 14655 2562 14656
rect 4840 14720 5160 14721
rect 4840 14656 4848 14720
rect 4912 14656 4928 14720
rect 4992 14656 5008 14720
rect 5072 14656 5088 14720
rect 5152 14656 5160 14720
rect 4840 14655 5160 14656
rect 7437 14720 7757 14721
rect 7437 14656 7445 14720
rect 7509 14656 7525 14720
rect 7589 14656 7605 14720
rect 7669 14656 7685 14720
rect 7749 14656 7757 14720
rect 7437 14655 7757 14656
rect 9200 14650 10000 14680
rect 7974 14590 10000 14650
rect 5809 14514 5875 14517
rect 7974 14514 8034 14590
rect 9200 14560 10000 14590
rect 5809 14512 8034 14514
rect 5809 14456 5814 14512
rect 5870 14456 8034 14512
rect 5809 14454 8034 14456
rect 5809 14451 5875 14454
rect 3541 14176 3861 14177
rect 3541 14112 3549 14176
rect 3613 14112 3629 14176
rect 3693 14112 3709 14176
rect 3773 14112 3789 14176
rect 3853 14112 3861 14176
rect 3541 14111 3861 14112
rect 6138 14176 6458 14177
rect 6138 14112 6146 14176
rect 6210 14112 6226 14176
rect 6290 14112 6306 14176
rect 6370 14112 6386 14176
rect 6450 14112 6458 14176
rect 6138 14111 6458 14112
rect 9200 14106 10000 14136
rect 6686 14046 10000 14106
rect 5257 13970 5323 13973
rect 6686 13970 6746 14046
rect 9200 14016 10000 14046
rect 5257 13968 6746 13970
rect 5257 13912 5262 13968
rect 5318 13912 6746 13968
rect 5257 13910 6746 13912
rect 5257 13907 5323 13910
rect 2242 13632 2562 13633
rect 2242 13568 2250 13632
rect 2314 13568 2330 13632
rect 2394 13568 2410 13632
rect 2474 13568 2490 13632
rect 2554 13568 2562 13632
rect 2242 13567 2562 13568
rect 4840 13632 5160 13633
rect 4840 13568 4848 13632
rect 4912 13568 4928 13632
rect 4992 13568 5008 13632
rect 5072 13568 5088 13632
rect 5152 13568 5160 13632
rect 4840 13567 5160 13568
rect 7437 13632 7757 13633
rect 7437 13568 7445 13632
rect 7509 13568 7525 13632
rect 7589 13568 7605 13632
rect 7669 13568 7685 13632
rect 7749 13568 7757 13632
rect 7437 13567 7757 13568
rect 9200 13562 10000 13592
rect 7974 13502 10000 13562
rect 7189 13426 7255 13429
rect 7974 13426 8034 13502
rect 9200 13472 10000 13502
rect 7189 13424 8034 13426
rect 7189 13368 7194 13424
rect 7250 13368 8034 13424
rect 7189 13366 8034 13368
rect 7189 13363 7255 13366
rect 3541 13088 3861 13089
rect 3541 13024 3549 13088
rect 3613 13024 3629 13088
rect 3693 13024 3709 13088
rect 3773 13024 3789 13088
rect 3853 13024 3861 13088
rect 3541 13023 3861 13024
rect 6138 13088 6458 13089
rect 6138 13024 6146 13088
rect 6210 13024 6226 13088
rect 6290 13024 6306 13088
rect 6370 13024 6386 13088
rect 6450 13024 6458 13088
rect 6138 13023 6458 13024
rect 6637 13018 6703 13021
rect 9200 13018 10000 13048
rect 6637 13016 10000 13018
rect 6637 12960 6642 13016
rect 6698 12960 10000 13016
rect 6637 12958 10000 12960
rect 6637 12955 6703 12958
rect 9200 12928 10000 12958
rect 3049 12882 3115 12885
rect 7189 12882 7255 12885
rect 3049 12880 7255 12882
rect 3049 12824 3054 12880
rect 3110 12824 7194 12880
rect 7250 12824 7255 12880
rect 3049 12822 7255 12824
rect 3049 12819 3115 12822
rect 7189 12819 7255 12822
rect 6821 12746 6887 12749
rect 6821 12744 8034 12746
rect 6821 12688 6826 12744
rect 6882 12688 8034 12744
rect 6821 12686 8034 12688
rect 6821 12683 6887 12686
rect 2242 12544 2562 12545
rect 2242 12480 2250 12544
rect 2314 12480 2330 12544
rect 2394 12480 2410 12544
rect 2474 12480 2490 12544
rect 2554 12480 2562 12544
rect 2242 12479 2562 12480
rect 4840 12544 5160 12545
rect 4840 12480 4848 12544
rect 4912 12480 4928 12544
rect 4992 12480 5008 12544
rect 5072 12480 5088 12544
rect 5152 12480 5160 12544
rect 4840 12479 5160 12480
rect 7437 12544 7757 12545
rect 7437 12480 7445 12544
rect 7509 12480 7525 12544
rect 7589 12480 7605 12544
rect 7669 12480 7685 12544
rect 7749 12480 7757 12544
rect 7437 12479 7757 12480
rect 7974 12474 8034 12686
rect 9200 12474 10000 12504
rect 7974 12414 10000 12474
rect 9200 12384 10000 12414
rect 3541 12000 3861 12001
rect 3541 11936 3549 12000
rect 3613 11936 3629 12000
rect 3693 11936 3709 12000
rect 3773 11936 3789 12000
rect 3853 11936 3861 12000
rect 3541 11935 3861 11936
rect 6138 12000 6458 12001
rect 6138 11936 6146 12000
rect 6210 11936 6226 12000
rect 6290 11936 6306 12000
rect 6370 11936 6386 12000
rect 6450 11936 6458 12000
rect 6138 11935 6458 11936
rect 8201 11930 8267 11933
rect 9200 11930 10000 11960
rect 8201 11928 10000 11930
rect 8201 11872 8206 11928
rect 8262 11872 10000 11928
rect 8201 11870 10000 11872
rect 8201 11867 8267 11870
rect 9200 11840 10000 11870
rect 2242 11456 2562 11457
rect 2242 11392 2250 11456
rect 2314 11392 2330 11456
rect 2394 11392 2410 11456
rect 2474 11392 2490 11456
rect 2554 11392 2562 11456
rect 2242 11391 2562 11392
rect 4840 11456 5160 11457
rect 4840 11392 4848 11456
rect 4912 11392 4928 11456
rect 4992 11392 5008 11456
rect 5072 11392 5088 11456
rect 5152 11392 5160 11456
rect 4840 11391 5160 11392
rect 7437 11456 7757 11457
rect 7437 11392 7445 11456
rect 7509 11392 7525 11456
rect 7589 11392 7605 11456
rect 7669 11392 7685 11456
rect 7749 11392 7757 11456
rect 7437 11391 7757 11392
rect 7833 11386 7899 11389
rect 9200 11386 10000 11416
rect 7833 11384 10000 11386
rect 7833 11328 7838 11384
rect 7894 11328 10000 11384
rect 7833 11326 10000 11328
rect 7833 11323 7899 11326
rect 9200 11296 10000 11326
rect 3541 10912 3861 10913
rect 3541 10848 3549 10912
rect 3613 10848 3629 10912
rect 3693 10848 3709 10912
rect 3773 10848 3789 10912
rect 3853 10848 3861 10912
rect 3541 10847 3861 10848
rect 6138 10912 6458 10913
rect 6138 10848 6146 10912
rect 6210 10848 6226 10912
rect 6290 10848 6306 10912
rect 6370 10848 6386 10912
rect 6450 10848 6458 10912
rect 6138 10847 6458 10848
rect 7373 10842 7439 10845
rect 9200 10842 10000 10872
rect 7373 10840 10000 10842
rect 7373 10784 7378 10840
rect 7434 10784 10000 10840
rect 7373 10782 10000 10784
rect 7373 10779 7439 10782
rect 9200 10752 10000 10782
rect 2773 10706 2839 10709
rect 5809 10706 5875 10709
rect 2773 10704 5875 10706
rect 2773 10648 2778 10704
rect 2834 10648 5814 10704
rect 5870 10648 5875 10704
rect 2773 10646 5875 10648
rect 2773 10643 2839 10646
rect 5809 10643 5875 10646
rect 2681 10570 2747 10573
rect 6729 10570 6795 10573
rect 2681 10568 6795 10570
rect 2681 10512 2686 10568
rect 2742 10512 6734 10568
rect 6790 10512 6795 10568
rect 2681 10510 6795 10512
rect 2681 10507 2747 10510
rect 6729 10507 6795 10510
rect 2242 10368 2562 10369
rect 2242 10304 2250 10368
rect 2314 10304 2330 10368
rect 2394 10304 2410 10368
rect 2474 10304 2490 10368
rect 2554 10304 2562 10368
rect 2242 10303 2562 10304
rect 4840 10368 5160 10369
rect 4840 10304 4848 10368
rect 4912 10304 4928 10368
rect 4992 10304 5008 10368
rect 5072 10304 5088 10368
rect 5152 10304 5160 10368
rect 4840 10303 5160 10304
rect 7437 10368 7757 10369
rect 7437 10304 7445 10368
rect 7509 10304 7525 10368
rect 7589 10304 7605 10368
rect 7669 10304 7685 10368
rect 7749 10304 7757 10368
rect 7437 10303 7757 10304
rect 8109 10298 8175 10301
rect 9200 10298 10000 10328
rect 8109 10296 10000 10298
rect 8109 10240 8114 10296
rect 8170 10240 10000 10296
rect 8109 10238 10000 10240
rect 8109 10235 8175 10238
rect 9200 10208 10000 10238
rect 2589 10162 2655 10165
rect 5625 10162 5691 10165
rect 2589 10160 5691 10162
rect 2589 10104 2594 10160
rect 2650 10104 5630 10160
rect 5686 10104 5691 10160
rect 2589 10102 5691 10104
rect 2589 10099 2655 10102
rect 5625 10099 5691 10102
rect 1577 10026 1643 10029
rect 1577 10024 6010 10026
rect 1577 9968 1582 10024
rect 1638 9968 6010 10024
rect 1577 9966 6010 9968
rect 1577 9963 1643 9966
rect 3541 9824 3861 9825
rect 3541 9760 3549 9824
rect 3613 9760 3629 9824
rect 3693 9760 3709 9824
rect 3773 9760 3789 9824
rect 3853 9760 3861 9824
rect 3541 9759 3861 9760
rect 5950 9690 6010 9966
rect 8293 9890 8359 9893
rect 9200 9890 10000 9920
rect 8293 9888 10000 9890
rect 8293 9832 8298 9888
rect 8354 9832 10000 9888
rect 8293 9830 10000 9832
rect 8293 9827 8359 9830
rect 6138 9824 6458 9825
rect 6138 9760 6146 9824
rect 6210 9760 6226 9824
rect 6290 9760 6306 9824
rect 6370 9760 6386 9824
rect 6450 9760 6458 9824
rect 9200 9800 10000 9830
rect 6138 9759 6458 9760
rect 6177 9690 6243 9693
rect 5950 9688 6243 9690
rect 5950 9632 6182 9688
rect 6238 9632 6243 9688
rect 5950 9630 6243 9632
rect 6177 9627 6243 9630
rect 8109 9346 8175 9349
rect 9200 9346 10000 9376
rect 8109 9344 10000 9346
rect 8109 9288 8114 9344
rect 8170 9288 10000 9344
rect 8109 9286 10000 9288
rect 8109 9283 8175 9286
rect 2242 9280 2562 9281
rect 2242 9216 2250 9280
rect 2314 9216 2330 9280
rect 2394 9216 2410 9280
rect 2474 9216 2490 9280
rect 2554 9216 2562 9280
rect 2242 9215 2562 9216
rect 4840 9280 5160 9281
rect 4840 9216 4848 9280
rect 4912 9216 4928 9280
rect 4992 9216 5008 9280
rect 5072 9216 5088 9280
rect 5152 9216 5160 9280
rect 4840 9215 5160 9216
rect 7437 9280 7757 9281
rect 7437 9216 7445 9280
rect 7509 9216 7525 9280
rect 7589 9216 7605 9280
rect 7669 9216 7685 9280
rect 7749 9216 7757 9280
rect 9200 9256 10000 9286
rect 7437 9215 7757 9216
rect 6821 8802 6887 8805
rect 8201 8802 8267 8805
rect 9200 8802 10000 8832
rect 6821 8800 10000 8802
rect 6821 8744 6826 8800
rect 6882 8744 8206 8800
rect 8262 8744 10000 8800
rect 6821 8742 10000 8744
rect 6821 8739 6887 8742
rect 8201 8739 8267 8742
rect 3541 8736 3861 8737
rect 3541 8672 3549 8736
rect 3613 8672 3629 8736
rect 3693 8672 3709 8736
rect 3773 8672 3789 8736
rect 3853 8672 3861 8736
rect 3541 8671 3861 8672
rect 6138 8736 6458 8737
rect 6138 8672 6146 8736
rect 6210 8672 6226 8736
rect 6290 8672 6306 8736
rect 6370 8672 6386 8736
rect 6450 8672 6458 8736
rect 9200 8712 10000 8742
rect 6138 8671 6458 8672
rect 9200 8258 10000 8288
rect 7974 8198 10000 8258
rect 2242 8192 2562 8193
rect 2242 8128 2250 8192
rect 2314 8128 2330 8192
rect 2394 8128 2410 8192
rect 2474 8128 2490 8192
rect 2554 8128 2562 8192
rect 2242 8127 2562 8128
rect 4840 8192 5160 8193
rect 4840 8128 4848 8192
rect 4912 8128 4928 8192
rect 4992 8128 5008 8192
rect 5072 8128 5088 8192
rect 5152 8128 5160 8192
rect 4840 8127 5160 8128
rect 7437 8192 7757 8193
rect 7437 8128 7445 8192
rect 7509 8128 7525 8192
rect 7589 8128 7605 8192
rect 7669 8128 7685 8192
rect 7749 8128 7757 8192
rect 7437 8127 7757 8128
rect 6637 7986 6703 7989
rect 7974 7986 8034 8198
rect 9200 8168 10000 8198
rect 6637 7984 8034 7986
rect 6637 7928 6642 7984
rect 6698 7928 8034 7984
rect 6637 7926 8034 7928
rect 6637 7923 6703 7926
rect 7925 7714 7991 7717
rect 9200 7714 10000 7744
rect 7925 7712 10000 7714
rect 7925 7656 7930 7712
rect 7986 7656 10000 7712
rect 7925 7654 10000 7656
rect 7925 7651 7991 7654
rect 3541 7648 3861 7649
rect 3541 7584 3549 7648
rect 3613 7584 3629 7648
rect 3693 7584 3709 7648
rect 3773 7584 3789 7648
rect 3853 7584 3861 7648
rect 3541 7583 3861 7584
rect 6138 7648 6458 7649
rect 6138 7584 6146 7648
rect 6210 7584 6226 7648
rect 6290 7584 6306 7648
rect 6370 7584 6386 7648
rect 6450 7584 6458 7648
rect 9200 7624 10000 7654
rect 6138 7583 6458 7584
rect 1761 7306 1827 7309
rect 3785 7306 3851 7309
rect 1761 7304 7896 7306
rect 1761 7248 1766 7304
rect 1822 7248 3790 7304
rect 3846 7248 7896 7304
rect 1761 7246 7896 7248
rect 1761 7243 1827 7246
rect 3785 7243 3851 7246
rect 7836 7173 7896 7246
rect 7833 7170 7899 7173
rect 9200 7170 10000 7200
rect 7833 7168 10000 7170
rect 7833 7112 7838 7168
rect 7894 7112 10000 7168
rect 7833 7110 10000 7112
rect 7833 7107 7899 7110
rect 2242 7104 2562 7105
rect 2242 7040 2250 7104
rect 2314 7040 2330 7104
rect 2394 7040 2410 7104
rect 2474 7040 2490 7104
rect 2554 7040 2562 7104
rect 2242 7039 2562 7040
rect 4840 7104 5160 7105
rect 4840 7040 4848 7104
rect 4912 7040 4928 7104
rect 4992 7040 5008 7104
rect 5072 7040 5088 7104
rect 5152 7040 5160 7104
rect 4840 7039 5160 7040
rect 7437 7104 7757 7105
rect 7437 7040 7445 7104
rect 7509 7040 7525 7104
rect 7589 7040 7605 7104
rect 7669 7040 7685 7104
rect 7749 7040 7757 7104
rect 9200 7080 10000 7110
rect 7437 7039 7757 7040
rect 7925 6626 7991 6629
rect 9200 6626 10000 6656
rect 7925 6624 10000 6626
rect 7925 6568 7930 6624
rect 7986 6568 10000 6624
rect 7925 6566 10000 6568
rect 7925 6563 7991 6566
rect 3541 6560 3861 6561
rect 3541 6496 3549 6560
rect 3613 6496 3629 6560
rect 3693 6496 3709 6560
rect 3773 6496 3789 6560
rect 3853 6496 3861 6560
rect 3541 6495 3861 6496
rect 6138 6560 6458 6561
rect 6138 6496 6146 6560
rect 6210 6496 6226 6560
rect 6290 6496 6306 6560
rect 6370 6496 6386 6560
rect 6450 6496 6458 6560
rect 9200 6536 10000 6566
rect 6138 6495 6458 6496
rect 2589 6218 2655 6221
rect 5625 6218 5691 6221
rect 2589 6216 5691 6218
rect 2589 6160 2594 6216
rect 2650 6160 5630 6216
rect 5686 6160 5691 6216
rect 2589 6158 5691 6160
rect 2589 6155 2655 6158
rect 5625 6155 5691 6158
rect 8109 6082 8175 6085
rect 9200 6082 10000 6112
rect 8109 6080 10000 6082
rect 8109 6024 8114 6080
rect 8170 6024 10000 6080
rect 8109 6022 10000 6024
rect 8109 6019 8175 6022
rect 2242 6016 2562 6017
rect 2242 5952 2250 6016
rect 2314 5952 2330 6016
rect 2394 5952 2410 6016
rect 2474 5952 2490 6016
rect 2554 5952 2562 6016
rect 2242 5951 2562 5952
rect 4840 6016 5160 6017
rect 4840 5952 4848 6016
rect 4912 5952 4928 6016
rect 4992 5952 5008 6016
rect 5072 5952 5088 6016
rect 5152 5952 5160 6016
rect 4840 5951 5160 5952
rect 7437 6016 7757 6017
rect 7437 5952 7445 6016
rect 7509 5952 7525 6016
rect 7589 5952 7605 6016
rect 7669 5952 7685 6016
rect 7749 5952 7757 6016
rect 9200 5992 10000 6022
rect 7437 5951 7757 5952
rect 1577 5674 1643 5677
rect 5717 5674 5783 5677
rect 1577 5672 5783 5674
rect 1577 5616 1582 5672
rect 1638 5616 5722 5672
rect 5778 5616 5783 5672
rect 1577 5614 5783 5616
rect 1577 5611 1643 5614
rect 5717 5611 5783 5614
rect 8201 5538 8267 5541
rect 9200 5538 10000 5568
rect 8201 5536 10000 5538
rect 8201 5480 8206 5536
rect 8262 5480 10000 5536
rect 8201 5478 10000 5480
rect 8201 5475 8267 5478
rect 3541 5472 3861 5473
rect 3541 5408 3549 5472
rect 3613 5408 3629 5472
rect 3693 5408 3709 5472
rect 3773 5408 3789 5472
rect 3853 5408 3861 5472
rect 3541 5407 3861 5408
rect 6138 5472 6458 5473
rect 6138 5408 6146 5472
rect 6210 5408 6226 5472
rect 6290 5408 6306 5472
rect 6370 5408 6386 5472
rect 6450 5408 6458 5472
rect 9200 5448 10000 5478
rect 6138 5407 6458 5408
rect 1393 5130 1459 5133
rect 3417 5130 3483 5133
rect 1393 5128 3483 5130
rect 1393 5072 1398 5128
rect 1454 5072 3422 5128
rect 3478 5072 3483 5128
rect 1393 5070 3483 5072
rect 1393 5067 1459 5070
rect 3417 5067 3483 5070
rect 7925 4994 7991 4997
rect 9200 4994 10000 5024
rect 7925 4992 10000 4994
rect 7925 4936 7930 4992
rect 7986 4936 10000 4992
rect 7925 4934 10000 4936
rect 7925 4931 7991 4934
rect 2242 4928 2562 4929
rect 2242 4864 2250 4928
rect 2314 4864 2330 4928
rect 2394 4864 2410 4928
rect 2474 4864 2490 4928
rect 2554 4864 2562 4928
rect 2242 4863 2562 4864
rect 4840 4928 5160 4929
rect 4840 4864 4848 4928
rect 4912 4864 4928 4928
rect 4992 4864 5008 4928
rect 5072 4864 5088 4928
rect 5152 4864 5160 4928
rect 4840 4863 5160 4864
rect 7437 4928 7757 4929
rect 7437 4864 7445 4928
rect 7509 4864 7525 4928
rect 7589 4864 7605 4928
rect 7669 4864 7685 4928
rect 7749 4864 7757 4928
rect 9200 4904 10000 4934
rect 7437 4863 7757 4864
rect 8293 4450 8359 4453
rect 9200 4450 10000 4480
rect 8293 4448 10000 4450
rect 8293 4392 8298 4448
rect 8354 4392 10000 4448
rect 8293 4390 10000 4392
rect 8293 4387 8359 4390
rect 3541 4384 3861 4385
rect 3541 4320 3549 4384
rect 3613 4320 3629 4384
rect 3693 4320 3709 4384
rect 3773 4320 3789 4384
rect 3853 4320 3861 4384
rect 3541 4319 3861 4320
rect 6138 4384 6458 4385
rect 6138 4320 6146 4384
rect 6210 4320 6226 4384
rect 6290 4320 6306 4384
rect 6370 4320 6386 4384
rect 6450 4320 6458 4384
rect 9200 4360 10000 4390
rect 6138 4319 6458 4320
rect 6821 4042 6887 4045
rect 6821 4040 8034 4042
rect 6821 3984 6826 4040
rect 6882 3984 8034 4040
rect 6821 3982 8034 3984
rect 6821 3979 6887 3982
rect 7974 3906 8034 3982
rect 9200 3906 10000 3936
rect 7974 3846 10000 3906
rect 2242 3840 2562 3841
rect 2242 3776 2250 3840
rect 2314 3776 2330 3840
rect 2394 3776 2410 3840
rect 2474 3776 2490 3840
rect 2554 3776 2562 3840
rect 2242 3775 2562 3776
rect 4840 3840 5160 3841
rect 4840 3776 4848 3840
rect 4912 3776 4928 3840
rect 4992 3776 5008 3840
rect 5072 3776 5088 3840
rect 5152 3776 5160 3840
rect 4840 3775 5160 3776
rect 7437 3840 7757 3841
rect 7437 3776 7445 3840
rect 7509 3776 7525 3840
rect 7589 3776 7605 3840
rect 7669 3776 7685 3840
rect 7749 3776 7757 3840
rect 9200 3816 10000 3846
rect 7437 3775 7757 3776
rect 8201 3362 8267 3365
rect 9200 3362 10000 3392
rect 8201 3360 10000 3362
rect 8201 3304 8206 3360
rect 8262 3304 10000 3360
rect 8201 3302 10000 3304
rect 8201 3299 8267 3302
rect 3541 3296 3861 3297
rect 3541 3232 3549 3296
rect 3613 3232 3629 3296
rect 3693 3232 3709 3296
rect 3773 3232 3789 3296
rect 3853 3232 3861 3296
rect 3541 3231 3861 3232
rect 6138 3296 6458 3297
rect 6138 3232 6146 3296
rect 6210 3232 6226 3296
rect 6290 3232 6306 3296
rect 6370 3232 6386 3296
rect 6450 3232 6458 3296
rect 9200 3272 10000 3302
rect 6138 3231 6458 3232
rect 6637 2954 6703 2957
rect 6637 2952 8034 2954
rect 6637 2896 6642 2952
rect 6698 2896 8034 2952
rect 6637 2894 8034 2896
rect 6637 2891 6703 2894
rect 7974 2818 8034 2894
rect 9200 2818 10000 2848
rect 7974 2758 10000 2818
rect 2242 2752 2562 2753
rect 2242 2688 2250 2752
rect 2314 2688 2330 2752
rect 2394 2688 2410 2752
rect 2474 2688 2490 2752
rect 2554 2688 2562 2752
rect 2242 2687 2562 2688
rect 4840 2752 5160 2753
rect 4840 2688 4848 2752
rect 4912 2688 4928 2752
rect 4992 2688 5008 2752
rect 5072 2688 5088 2752
rect 5152 2688 5160 2752
rect 4840 2687 5160 2688
rect 7437 2752 7757 2753
rect 7437 2688 7445 2752
rect 7509 2688 7525 2752
rect 7589 2688 7605 2752
rect 7669 2688 7685 2752
rect 7749 2688 7757 2752
rect 9200 2728 10000 2758
rect 7437 2687 7757 2688
rect 8017 2274 8083 2277
rect 9200 2274 10000 2304
rect 8017 2272 10000 2274
rect 8017 2216 8022 2272
rect 8078 2216 10000 2272
rect 8017 2214 10000 2216
rect 8017 2211 8083 2214
rect 3541 2208 3861 2209
rect 3541 2144 3549 2208
rect 3613 2144 3629 2208
rect 3693 2144 3709 2208
rect 3773 2144 3789 2208
rect 3853 2144 3861 2208
rect 3541 2143 3861 2144
rect 6138 2208 6458 2209
rect 6138 2144 6146 2208
rect 6210 2144 6226 2208
rect 6290 2144 6306 2208
rect 6370 2144 6386 2208
rect 6450 2144 6458 2208
rect 9200 2184 10000 2214
rect 6138 2143 6458 2144
rect 6637 1730 6703 1733
rect 9200 1730 10000 1760
rect 6637 1728 10000 1730
rect 6637 1672 6642 1728
rect 6698 1672 10000 1728
rect 6637 1670 10000 1672
rect 6637 1667 6703 1670
rect 9200 1640 10000 1670
rect 5993 1186 6059 1189
rect 9200 1186 10000 1216
rect 5993 1184 10000 1186
rect 5993 1128 5998 1184
rect 6054 1128 10000 1184
rect 5993 1126 10000 1128
rect 5993 1123 6059 1126
rect 9200 1096 10000 1126
rect 6545 642 6611 645
rect 9200 642 10000 672
rect 6545 640 10000 642
rect 6545 584 6550 640
rect 6606 584 10000 640
rect 6545 582 10000 584
rect 6545 579 6611 582
rect 9200 552 10000 582
rect 6637 234 6703 237
rect 9200 234 10000 264
rect 6637 232 10000 234
rect 6637 176 6642 232
rect 6698 176 10000 232
rect 6637 174 10000 176
rect 6637 171 6703 174
rect 9200 144 10000 174
<< via3 >>
rect 2250 27772 2314 27776
rect 2250 27716 2254 27772
rect 2254 27716 2310 27772
rect 2310 27716 2314 27772
rect 2250 27712 2314 27716
rect 2330 27772 2394 27776
rect 2330 27716 2334 27772
rect 2334 27716 2390 27772
rect 2390 27716 2394 27772
rect 2330 27712 2394 27716
rect 2410 27772 2474 27776
rect 2410 27716 2414 27772
rect 2414 27716 2470 27772
rect 2470 27716 2474 27772
rect 2410 27712 2474 27716
rect 2490 27772 2554 27776
rect 2490 27716 2494 27772
rect 2494 27716 2550 27772
rect 2550 27716 2554 27772
rect 2490 27712 2554 27716
rect 4848 27772 4912 27776
rect 4848 27716 4852 27772
rect 4852 27716 4908 27772
rect 4908 27716 4912 27772
rect 4848 27712 4912 27716
rect 4928 27772 4992 27776
rect 4928 27716 4932 27772
rect 4932 27716 4988 27772
rect 4988 27716 4992 27772
rect 4928 27712 4992 27716
rect 5008 27772 5072 27776
rect 5008 27716 5012 27772
rect 5012 27716 5068 27772
rect 5068 27716 5072 27772
rect 5008 27712 5072 27716
rect 5088 27772 5152 27776
rect 5088 27716 5092 27772
rect 5092 27716 5148 27772
rect 5148 27716 5152 27772
rect 5088 27712 5152 27716
rect 7445 27772 7509 27776
rect 7445 27716 7449 27772
rect 7449 27716 7505 27772
rect 7505 27716 7509 27772
rect 7445 27712 7509 27716
rect 7525 27772 7589 27776
rect 7525 27716 7529 27772
rect 7529 27716 7585 27772
rect 7585 27716 7589 27772
rect 7525 27712 7589 27716
rect 7605 27772 7669 27776
rect 7605 27716 7609 27772
rect 7609 27716 7665 27772
rect 7665 27716 7669 27772
rect 7605 27712 7669 27716
rect 7685 27772 7749 27776
rect 7685 27716 7689 27772
rect 7689 27716 7745 27772
rect 7745 27716 7749 27772
rect 7685 27712 7749 27716
rect 3549 27228 3613 27232
rect 3549 27172 3553 27228
rect 3553 27172 3609 27228
rect 3609 27172 3613 27228
rect 3549 27168 3613 27172
rect 3629 27228 3693 27232
rect 3629 27172 3633 27228
rect 3633 27172 3689 27228
rect 3689 27172 3693 27228
rect 3629 27168 3693 27172
rect 3709 27228 3773 27232
rect 3709 27172 3713 27228
rect 3713 27172 3769 27228
rect 3769 27172 3773 27228
rect 3709 27168 3773 27172
rect 3789 27228 3853 27232
rect 3789 27172 3793 27228
rect 3793 27172 3849 27228
rect 3849 27172 3853 27228
rect 3789 27168 3853 27172
rect 6146 27228 6210 27232
rect 6146 27172 6150 27228
rect 6150 27172 6206 27228
rect 6206 27172 6210 27228
rect 6146 27168 6210 27172
rect 6226 27228 6290 27232
rect 6226 27172 6230 27228
rect 6230 27172 6286 27228
rect 6286 27172 6290 27228
rect 6226 27168 6290 27172
rect 6306 27228 6370 27232
rect 6306 27172 6310 27228
rect 6310 27172 6366 27228
rect 6366 27172 6370 27228
rect 6306 27168 6370 27172
rect 6386 27228 6450 27232
rect 6386 27172 6390 27228
rect 6390 27172 6446 27228
rect 6446 27172 6450 27228
rect 6386 27168 6450 27172
rect 2250 26684 2314 26688
rect 2250 26628 2254 26684
rect 2254 26628 2310 26684
rect 2310 26628 2314 26684
rect 2250 26624 2314 26628
rect 2330 26684 2394 26688
rect 2330 26628 2334 26684
rect 2334 26628 2390 26684
rect 2390 26628 2394 26684
rect 2330 26624 2394 26628
rect 2410 26684 2474 26688
rect 2410 26628 2414 26684
rect 2414 26628 2470 26684
rect 2470 26628 2474 26684
rect 2410 26624 2474 26628
rect 2490 26684 2554 26688
rect 2490 26628 2494 26684
rect 2494 26628 2550 26684
rect 2550 26628 2554 26684
rect 2490 26624 2554 26628
rect 4848 26684 4912 26688
rect 4848 26628 4852 26684
rect 4852 26628 4908 26684
rect 4908 26628 4912 26684
rect 4848 26624 4912 26628
rect 4928 26684 4992 26688
rect 4928 26628 4932 26684
rect 4932 26628 4988 26684
rect 4988 26628 4992 26684
rect 4928 26624 4992 26628
rect 5008 26684 5072 26688
rect 5008 26628 5012 26684
rect 5012 26628 5068 26684
rect 5068 26628 5072 26684
rect 5008 26624 5072 26628
rect 5088 26684 5152 26688
rect 5088 26628 5092 26684
rect 5092 26628 5148 26684
rect 5148 26628 5152 26684
rect 5088 26624 5152 26628
rect 7445 26684 7509 26688
rect 7445 26628 7449 26684
rect 7449 26628 7505 26684
rect 7505 26628 7509 26684
rect 7445 26624 7509 26628
rect 7525 26684 7589 26688
rect 7525 26628 7529 26684
rect 7529 26628 7585 26684
rect 7585 26628 7589 26684
rect 7525 26624 7589 26628
rect 7605 26684 7669 26688
rect 7605 26628 7609 26684
rect 7609 26628 7665 26684
rect 7665 26628 7669 26684
rect 7605 26624 7669 26628
rect 7685 26684 7749 26688
rect 7685 26628 7689 26684
rect 7689 26628 7745 26684
rect 7745 26628 7749 26684
rect 7685 26624 7749 26628
rect 3549 26140 3613 26144
rect 3549 26084 3553 26140
rect 3553 26084 3609 26140
rect 3609 26084 3613 26140
rect 3549 26080 3613 26084
rect 3629 26140 3693 26144
rect 3629 26084 3633 26140
rect 3633 26084 3689 26140
rect 3689 26084 3693 26140
rect 3629 26080 3693 26084
rect 3709 26140 3773 26144
rect 3709 26084 3713 26140
rect 3713 26084 3769 26140
rect 3769 26084 3773 26140
rect 3709 26080 3773 26084
rect 3789 26140 3853 26144
rect 3789 26084 3793 26140
rect 3793 26084 3849 26140
rect 3849 26084 3853 26140
rect 3789 26080 3853 26084
rect 6146 26140 6210 26144
rect 6146 26084 6150 26140
rect 6150 26084 6206 26140
rect 6206 26084 6210 26140
rect 6146 26080 6210 26084
rect 6226 26140 6290 26144
rect 6226 26084 6230 26140
rect 6230 26084 6286 26140
rect 6286 26084 6290 26140
rect 6226 26080 6290 26084
rect 6306 26140 6370 26144
rect 6306 26084 6310 26140
rect 6310 26084 6366 26140
rect 6366 26084 6370 26140
rect 6306 26080 6370 26084
rect 6386 26140 6450 26144
rect 6386 26084 6390 26140
rect 6390 26084 6446 26140
rect 6446 26084 6450 26140
rect 6386 26080 6450 26084
rect 2250 25596 2314 25600
rect 2250 25540 2254 25596
rect 2254 25540 2310 25596
rect 2310 25540 2314 25596
rect 2250 25536 2314 25540
rect 2330 25596 2394 25600
rect 2330 25540 2334 25596
rect 2334 25540 2390 25596
rect 2390 25540 2394 25596
rect 2330 25536 2394 25540
rect 2410 25596 2474 25600
rect 2410 25540 2414 25596
rect 2414 25540 2470 25596
rect 2470 25540 2474 25596
rect 2410 25536 2474 25540
rect 2490 25596 2554 25600
rect 2490 25540 2494 25596
rect 2494 25540 2550 25596
rect 2550 25540 2554 25596
rect 2490 25536 2554 25540
rect 4848 25596 4912 25600
rect 4848 25540 4852 25596
rect 4852 25540 4908 25596
rect 4908 25540 4912 25596
rect 4848 25536 4912 25540
rect 4928 25596 4992 25600
rect 4928 25540 4932 25596
rect 4932 25540 4988 25596
rect 4988 25540 4992 25596
rect 4928 25536 4992 25540
rect 5008 25596 5072 25600
rect 5008 25540 5012 25596
rect 5012 25540 5068 25596
rect 5068 25540 5072 25596
rect 5008 25536 5072 25540
rect 5088 25596 5152 25600
rect 5088 25540 5092 25596
rect 5092 25540 5148 25596
rect 5148 25540 5152 25596
rect 5088 25536 5152 25540
rect 7445 25596 7509 25600
rect 7445 25540 7449 25596
rect 7449 25540 7505 25596
rect 7505 25540 7509 25596
rect 7445 25536 7509 25540
rect 7525 25596 7589 25600
rect 7525 25540 7529 25596
rect 7529 25540 7585 25596
rect 7585 25540 7589 25596
rect 7525 25536 7589 25540
rect 7605 25596 7669 25600
rect 7605 25540 7609 25596
rect 7609 25540 7665 25596
rect 7665 25540 7669 25596
rect 7605 25536 7669 25540
rect 7685 25596 7749 25600
rect 7685 25540 7689 25596
rect 7689 25540 7745 25596
rect 7745 25540 7749 25596
rect 7685 25536 7749 25540
rect 3549 25052 3613 25056
rect 3549 24996 3553 25052
rect 3553 24996 3609 25052
rect 3609 24996 3613 25052
rect 3549 24992 3613 24996
rect 3629 25052 3693 25056
rect 3629 24996 3633 25052
rect 3633 24996 3689 25052
rect 3689 24996 3693 25052
rect 3629 24992 3693 24996
rect 3709 25052 3773 25056
rect 3709 24996 3713 25052
rect 3713 24996 3769 25052
rect 3769 24996 3773 25052
rect 3709 24992 3773 24996
rect 3789 25052 3853 25056
rect 3789 24996 3793 25052
rect 3793 24996 3849 25052
rect 3849 24996 3853 25052
rect 3789 24992 3853 24996
rect 6146 25052 6210 25056
rect 6146 24996 6150 25052
rect 6150 24996 6206 25052
rect 6206 24996 6210 25052
rect 6146 24992 6210 24996
rect 6226 25052 6290 25056
rect 6226 24996 6230 25052
rect 6230 24996 6286 25052
rect 6286 24996 6290 25052
rect 6226 24992 6290 24996
rect 6306 25052 6370 25056
rect 6306 24996 6310 25052
rect 6310 24996 6366 25052
rect 6366 24996 6370 25052
rect 6306 24992 6370 24996
rect 6386 25052 6450 25056
rect 6386 24996 6390 25052
rect 6390 24996 6446 25052
rect 6446 24996 6450 25052
rect 6386 24992 6450 24996
rect 2250 24508 2314 24512
rect 2250 24452 2254 24508
rect 2254 24452 2310 24508
rect 2310 24452 2314 24508
rect 2250 24448 2314 24452
rect 2330 24508 2394 24512
rect 2330 24452 2334 24508
rect 2334 24452 2390 24508
rect 2390 24452 2394 24508
rect 2330 24448 2394 24452
rect 2410 24508 2474 24512
rect 2410 24452 2414 24508
rect 2414 24452 2470 24508
rect 2470 24452 2474 24508
rect 2410 24448 2474 24452
rect 2490 24508 2554 24512
rect 2490 24452 2494 24508
rect 2494 24452 2550 24508
rect 2550 24452 2554 24508
rect 2490 24448 2554 24452
rect 4848 24508 4912 24512
rect 4848 24452 4852 24508
rect 4852 24452 4908 24508
rect 4908 24452 4912 24508
rect 4848 24448 4912 24452
rect 4928 24508 4992 24512
rect 4928 24452 4932 24508
rect 4932 24452 4988 24508
rect 4988 24452 4992 24508
rect 4928 24448 4992 24452
rect 5008 24508 5072 24512
rect 5008 24452 5012 24508
rect 5012 24452 5068 24508
rect 5068 24452 5072 24508
rect 5008 24448 5072 24452
rect 5088 24508 5152 24512
rect 5088 24452 5092 24508
rect 5092 24452 5148 24508
rect 5148 24452 5152 24508
rect 5088 24448 5152 24452
rect 7445 24508 7509 24512
rect 7445 24452 7449 24508
rect 7449 24452 7505 24508
rect 7505 24452 7509 24508
rect 7445 24448 7509 24452
rect 7525 24508 7589 24512
rect 7525 24452 7529 24508
rect 7529 24452 7585 24508
rect 7585 24452 7589 24508
rect 7525 24448 7589 24452
rect 7605 24508 7669 24512
rect 7605 24452 7609 24508
rect 7609 24452 7665 24508
rect 7665 24452 7669 24508
rect 7605 24448 7669 24452
rect 7685 24508 7749 24512
rect 7685 24452 7689 24508
rect 7689 24452 7745 24508
rect 7745 24452 7749 24508
rect 7685 24448 7749 24452
rect 3549 23964 3613 23968
rect 3549 23908 3553 23964
rect 3553 23908 3609 23964
rect 3609 23908 3613 23964
rect 3549 23904 3613 23908
rect 3629 23964 3693 23968
rect 3629 23908 3633 23964
rect 3633 23908 3689 23964
rect 3689 23908 3693 23964
rect 3629 23904 3693 23908
rect 3709 23964 3773 23968
rect 3709 23908 3713 23964
rect 3713 23908 3769 23964
rect 3769 23908 3773 23964
rect 3709 23904 3773 23908
rect 3789 23964 3853 23968
rect 3789 23908 3793 23964
rect 3793 23908 3849 23964
rect 3849 23908 3853 23964
rect 3789 23904 3853 23908
rect 6146 23964 6210 23968
rect 6146 23908 6150 23964
rect 6150 23908 6206 23964
rect 6206 23908 6210 23964
rect 6146 23904 6210 23908
rect 6226 23964 6290 23968
rect 6226 23908 6230 23964
rect 6230 23908 6286 23964
rect 6286 23908 6290 23964
rect 6226 23904 6290 23908
rect 6306 23964 6370 23968
rect 6306 23908 6310 23964
rect 6310 23908 6366 23964
rect 6366 23908 6370 23964
rect 6306 23904 6370 23908
rect 6386 23964 6450 23968
rect 6386 23908 6390 23964
rect 6390 23908 6446 23964
rect 6446 23908 6450 23964
rect 6386 23904 6450 23908
rect 2250 23420 2314 23424
rect 2250 23364 2254 23420
rect 2254 23364 2310 23420
rect 2310 23364 2314 23420
rect 2250 23360 2314 23364
rect 2330 23420 2394 23424
rect 2330 23364 2334 23420
rect 2334 23364 2390 23420
rect 2390 23364 2394 23420
rect 2330 23360 2394 23364
rect 2410 23420 2474 23424
rect 2410 23364 2414 23420
rect 2414 23364 2470 23420
rect 2470 23364 2474 23420
rect 2410 23360 2474 23364
rect 2490 23420 2554 23424
rect 2490 23364 2494 23420
rect 2494 23364 2550 23420
rect 2550 23364 2554 23420
rect 2490 23360 2554 23364
rect 4848 23420 4912 23424
rect 4848 23364 4852 23420
rect 4852 23364 4908 23420
rect 4908 23364 4912 23420
rect 4848 23360 4912 23364
rect 4928 23420 4992 23424
rect 4928 23364 4932 23420
rect 4932 23364 4988 23420
rect 4988 23364 4992 23420
rect 4928 23360 4992 23364
rect 5008 23420 5072 23424
rect 5008 23364 5012 23420
rect 5012 23364 5068 23420
rect 5068 23364 5072 23420
rect 5008 23360 5072 23364
rect 5088 23420 5152 23424
rect 5088 23364 5092 23420
rect 5092 23364 5148 23420
rect 5148 23364 5152 23420
rect 5088 23360 5152 23364
rect 7445 23420 7509 23424
rect 7445 23364 7449 23420
rect 7449 23364 7505 23420
rect 7505 23364 7509 23420
rect 7445 23360 7509 23364
rect 7525 23420 7589 23424
rect 7525 23364 7529 23420
rect 7529 23364 7585 23420
rect 7585 23364 7589 23420
rect 7525 23360 7589 23364
rect 7605 23420 7669 23424
rect 7605 23364 7609 23420
rect 7609 23364 7665 23420
rect 7665 23364 7669 23420
rect 7605 23360 7669 23364
rect 7685 23420 7749 23424
rect 7685 23364 7689 23420
rect 7689 23364 7745 23420
rect 7745 23364 7749 23420
rect 7685 23360 7749 23364
rect 3549 22876 3613 22880
rect 3549 22820 3553 22876
rect 3553 22820 3609 22876
rect 3609 22820 3613 22876
rect 3549 22816 3613 22820
rect 3629 22876 3693 22880
rect 3629 22820 3633 22876
rect 3633 22820 3689 22876
rect 3689 22820 3693 22876
rect 3629 22816 3693 22820
rect 3709 22876 3773 22880
rect 3709 22820 3713 22876
rect 3713 22820 3769 22876
rect 3769 22820 3773 22876
rect 3709 22816 3773 22820
rect 3789 22876 3853 22880
rect 3789 22820 3793 22876
rect 3793 22820 3849 22876
rect 3849 22820 3853 22876
rect 3789 22816 3853 22820
rect 6146 22876 6210 22880
rect 6146 22820 6150 22876
rect 6150 22820 6206 22876
rect 6206 22820 6210 22876
rect 6146 22816 6210 22820
rect 6226 22876 6290 22880
rect 6226 22820 6230 22876
rect 6230 22820 6286 22876
rect 6286 22820 6290 22876
rect 6226 22816 6290 22820
rect 6306 22876 6370 22880
rect 6306 22820 6310 22876
rect 6310 22820 6366 22876
rect 6366 22820 6370 22876
rect 6306 22816 6370 22820
rect 6386 22876 6450 22880
rect 6386 22820 6390 22876
rect 6390 22820 6446 22876
rect 6446 22820 6450 22876
rect 6386 22816 6450 22820
rect 2250 22332 2314 22336
rect 2250 22276 2254 22332
rect 2254 22276 2310 22332
rect 2310 22276 2314 22332
rect 2250 22272 2314 22276
rect 2330 22332 2394 22336
rect 2330 22276 2334 22332
rect 2334 22276 2390 22332
rect 2390 22276 2394 22332
rect 2330 22272 2394 22276
rect 2410 22332 2474 22336
rect 2410 22276 2414 22332
rect 2414 22276 2470 22332
rect 2470 22276 2474 22332
rect 2410 22272 2474 22276
rect 2490 22332 2554 22336
rect 2490 22276 2494 22332
rect 2494 22276 2550 22332
rect 2550 22276 2554 22332
rect 2490 22272 2554 22276
rect 4848 22332 4912 22336
rect 4848 22276 4852 22332
rect 4852 22276 4908 22332
rect 4908 22276 4912 22332
rect 4848 22272 4912 22276
rect 4928 22332 4992 22336
rect 4928 22276 4932 22332
rect 4932 22276 4988 22332
rect 4988 22276 4992 22332
rect 4928 22272 4992 22276
rect 5008 22332 5072 22336
rect 5008 22276 5012 22332
rect 5012 22276 5068 22332
rect 5068 22276 5072 22332
rect 5008 22272 5072 22276
rect 5088 22332 5152 22336
rect 5088 22276 5092 22332
rect 5092 22276 5148 22332
rect 5148 22276 5152 22332
rect 5088 22272 5152 22276
rect 7445 22332 7509 22336
rect 7445 22276 7449 22332
rect 7449 22276 7505 22332
rect 7505 22276 7509 22332
rect 7445 22272 7509 22276
rect 7525 22332 7589 22336
rect 7525 22276 7529 22332
rect 7529 22276 7585 22332
rect 7585 22276 7589 22332
rect 7525 22272 7589 22276
rect 7605 22332 7669 22336
rect 7605 22276 7609 22332
rect 7609 22276 7665 22332
rect 7665 22276 7669 22332
rect 7605 22272 7669 22276
rect 7685 22332 7749 22336
rect 7685 22276 7689 22332
rect 7689 22276 7745 22332
rect 7745 22276 7749 22332
rect 7685 22272 7749 22276
rect 3549 21788 3613 21792
rect 3549 21732 3553 21788
rect 3553 21732 3609 21788
rect 3609 21732 3613 21788
rect 3549 21728 3613 21732
rect 3629 21788 3693 21792
rect 3629 21732 3633 21788
rect 3633 21732 3689 21788
rect 3689 21732 3693 21788
rect 3629 21728 3693 21732
rect 3709 21788 3773 21792
rect 3709 21732 3713 21788
rect 3713 21732 3769 21788
rect 3769 21732 3773 21788
rect 3709 21728 3773 21732
rect 3789 21788 3853 21792
rect 3789 21732 3793 21788
rect 3793 21732 3849 21788
rect 3849 21732 3853 21788
rect 3789 21728 3853 21732
rect 6146 21788 6210 21792
rect 6146 21732 6150 21788
rect 6150 21732 6206 21788
rect 6206 21732 6210 21788
rect 6146 21728 6210 21732
rect 6226 21788 6290 21792
rect 6226 21732 6230 21788
rect 6230 21732 6286 21788
rect 6286 21732 6290 21788
rect 6226 21728 6290 21732
rect 6306 21788 6370 21792
rect 6306 21732 6310 21788
rect 6310 21732 6366 21788
rect 6366 21732 6370 21788
rect 6306 21728 6370 21732
rect 6386 21788 6450 21792
rect 6386 21732 6390 21788
rect 6390 21732 6446 21788
rect 6446 21732 6450 21788
rect 6386 21728 6450 21732
rect 2250 21244 2314 21248
rect 2250 21188 2254 21244
rect 2254 21188 2310 21244
rect 2310 21188 2314 21244
rect 2250 21184 2314 21188
rect 2330 21244 2394 21248
rect 2330 21188 2334 21244
rect 2334 21188 2390 21244
rect 2390 21188 2394 21244
rect 2330 21184 2394 21188
rect 2410 21244 2474 21248
rect 2410 21188 2414 21244
rect 2414 21188 2470 21244
rect 2470 21188 2474 21244
rect 2410 21184 2474 21188
rect 2490 21244 2554 21248
rect 2490 21188 2494 21244
rect 2494 21188 2550 21244
rect 2550 21188 2554 21244
rect 2490 21184 2554 21188
rect 4848 21244 4912 21248
rect 4848 21188 4852 21244
rect 4852 21188 4908 21244
rect 4908 21188 4912 21244
rect 4848 21184 4912 21188
rect 4928 21244 4992 21248
rect 4928 21188 4932 21244
rect 4932 21188 4988 21244
rect 4988 21188 4992 21244
rect 4928 21184 4992 21188
rect 5008 21244 5072 21248
rect 5008 21188 5012 21244
rect 5012 21188 5068 21244
rect 5068 21188 5072 21244
rect 5008 21184 5072 21188
rect 5088 21244 5152 21248
rect 5088 21188 5092 21244
rect 5092 21188 5148 21244
rect 5148 21188 5152 21244
rect 5088 21184 5152 21188
rect 7445 21244 7509 21248
rect 7445 21188 7449 21244
rect 7449 21188 7505 21244
rect 7505 21188 7509 21244
rect 7445 21184 7509 21188
rect 7525 21244 7589 21248
rect 7525 21188 7529 21244
rect 7529 21188 7585 21244
rect 7585 21188 7589 21244
rect 7525 21184 7589 21188
rect 7605 21244 7669 21248
rect 7605 21188 7609 21244
rect 7609 21188 7665 21244
rect 7665 21188 7669 21244
rect 7605 21184 7669 21188
rect 7685 21244 7749 21248
rect 7685 21188 7689 21244
rect 7689 21188 7745 21244
rect 7745 21188 7749 21244
rect 7685 21184 7749 21188
rect 3549 20700 3613 20704
rect 3549 20644 3553 20700
rect 3553 20644 3609 20700
rect 3609 20644 3613 20700
rect 3549 20640 3613 20644
rect 3629 20700 3693 20704
rect 3629 20644 3633 20700
rect 3633 20644 3689 20700
rect 3689 20644 3693 20700
rect 3629 20640 3693 20644
rect 3709 20700 3773 20704
rect 3709 20644 3713 20700
rect 3713 20644 3769 20700
rect 3769 20644 3773 20700
rect 3709 20640 3773 20644
rect 3789 20700 3853 20704
rect 3789 20644 3793 20700
rect 3793 20644 3849 20700
rect 3849 20644 3853 20700
rect 3789 20640 3853 20644
rect 6146 20700 6210 20704
rect 6146 20644 6150 20700
rect 6150 20644 6206 20700
rect 6206 20644 6210 20700
rect 6146 20640 6210 20644
rect 6226 20700 6290 20704
rect 6226 20644 6230 20700
rect 6230 20644 6286 20700
rect 6286 20644 6290 20700
rect 6226 20640 6290 20644
rect 6306 20700 6370 20704
rect 6306 20644 6310 20700
rect 6310 20644 6366 20700
rect 6366 20644 6370 20700
rect 6306 20640 6370 20644
rect 6386 20700 6450 20704
rect 6386 20644 6390 20700
rect 6390 20644 6446 20700
rect 6446 20644 6450 20700
rect 6386 20640 6450 20644
rect 2250 20156 2314 20160
rect 2250 20100 2254 20156
rect 2254 20100 2310 20156
rect 2310 20100 2314 20156
rect 2250 20096 2314 20100
rect 2330 20156 2394 20160
rect 2330 20100 2334 20156
rect 2334 20100 2390 20156
rect 2390 20100 2394 20156
rect 2330 20096 2394 20100
rect 2410 20156 2474 20160
rect 2410 20100 2414 20156
rect 2414 20100 2470 20156
rect 2470 20100 2474 20156
rect 2410 20096 2474 20100
rect 2490 20156 2554 20160
rect 2490 20100 2494 20156
rect 2494 20100 2550 20156
rect 2550 20100 2554 20156
rect 2490 20096 2554 20100
rect 4848 20156 4912 20160
rect 4848 20100 4852 20156
rect 4852 20100 4908 20156
rect 4908 20100 4912 20156
rect 4848 20096 4912 20100
rect 4928 20156 4992 20160
rect 4928 20100 4932 20156
rect 4932 20100 4988 20156
rect 4988 20100 4992 20156
rect 4928 20096 4992 20100
rect 5008 20156 5072 20160
rect 5008 20100 5012 20156
rect 5012 20100 5068 20156
rect 5068 20100 5072 20156
rect 5008 20096 5072 20100
rect 5088 20156 5152 20160
rect 5088 20100 5092 20156
rect 5092 20100 5148 20156
rect 5148 20100 5152 20156
rect 5088 20096 5152 20100
rect 7445 20156 7509 20160
rect 7445 20100 7449 20156
rect 7449 20100 7505 20156
rect 7505 20100 7509 20156
rect 7445 20096 7509 20100
rect 7525 20156 7589 20160
rect 7525 20100 7529 20156
rect 7529 20100 7585 20156
rect 7585 20100 7589 20156
rect 7525 20096 7589 20100
rect 7605 20156 7669 20160
rect 7605 20100 7609 20156
rect 7609 20100 7665 20156
rect 7665 20100 7669 20156
rect 7605 20096 7669 20100
rect 7685 20156 7749 20160
rect 7685 20100 7689 20156
rect 7689 20100 7745 20156
rect 7745 20100 7749 20156
rect 7685 20096 7749 20100
rect 3549 19612 3613 19616
rect 3549 19556 3553 19612
rect 3553 19556 3609 19612
rect 3609 19556 3613 19612
rect 3549 19552 3613 19556
rect 3629 19612 3693 19616
rect 3629 19556 3633 19612
rect 3633 19556 3689 19612
rect 3689 19556 3693 19612
rect 3629 19552 3693 19556
rect 3709 19612 3773 19616
rect 3709 19556 3713 19612
rect 3713 19556 3769 19612
rect 3769 19556 3773 19612
rect 3709 19552 3773 19556
rect 3789 19612 3853 19616
rect 3789 19556 3793 19612
rect 3793 19556 3849 19612
rect 3849 19556 3853 19612
rect 3789 19552 3853 19556
rect 6146 19612 6210 19616
rect 6146 19556 6150 19612
rect 6150 19556 6206 19612
rect 6206 19556 6210 19612
rect 6146 19552 6210 19556
rect 6226 19612 6290 19616
rect 6226 19556 6230 19612
rect 6230 19556 6286 19612
rect 6286 19556 6290 19612
rect 6226 19552 6290 19556
rect 6306 19612 6370 19616
rect 6306 19556 6310 19612
rect 6310 19556 6366 19612
rect 6366 19556 6370 19612
rect 6306 19552 6370 19556
rect 6386 19612 6450 19616
rect 6386 19556 6390 19612
rect 6390 19556 6446 19612
rect 6446 19556 6450 19612
rect 6386 19552 6450 19556
rect 2250 19068 2314 19072
rect 2250 19012 2254 19068
rect 2254 19012 2310 19068
rect 2310 19012 2314 19068
rect 2250 19008 2314 19012
rect 2330 19068 2394 19072
rect 2330 19012 2334 19068
rect 2334 19012 2390 19068
rect 2390 19012 2394 19068
rect 2330 19008 2394 19012
rect 2410 19068 2474 19072
rect 2410 19012 2414 19068
rect 2414 19012 2470 19068
rect 2470 19012 2474 19068
rect 2410 19008 2474 19012
rect 2490 19068 2554 19072
rect 2490 19012 2494 19068
rect 2494 19012 2550 19068
rect 2550 19012 2554 19068
rect 2490 19008 2554 19012
rect 4848 19068 4912 19072
rect 4848 19012 4852 19068
rect 4852 19012 4908 19068
rect 4908 19012 4912 19068
rect 4848 19008 4912 19012
rect 4928 19068 4992 19072
rect 4928 19012 4932 19068
rect 4932 19012 4988 19068
rect 4988 19012 4992 19068
rect 4928 19008 4992 19012
rect 5008 19068 5072 19072
rect 5008 19012 5012 19068
rect 5012 19012 5068 19068
rect 5068 19012 5072 19068
rect 5008 19008 5072 19012
rect 5088 19068 5152 19072
rect 5088 19012 5092 19068
rect 5092 19012 5148 19068
rect 5148 19012 5152 19068
rect 5088 19008 5152 19012
rect 7445 19068 7509 19072
rect 7445 19012 7449 19068
rect 7449 19012 7505 19068
rect 7505 19012 7509 19068
rect 7445 19008 7509 19012
rect 7525 19068 7589 19072
rect 7525 19012 7529 19068
rect 7529 19012 7585 19068
rect 7585 19012 7589 19068
rect 7525 19008 7589 19012
rect 7605 19068 7669 19072
rect 7605 19012 7609 19068
rect 7609 19012 7665 19068
rect 7665 19012 7669 19068
rect 7605 19008 7669 19012
rect 7685 19068 7749 19072
rect 7685 19012 7689 19068
rect 7689 19012 7745 19068
rect 7745 19012 7749 19068
rect 7685 19008 7749 19012
rect 3549 18524 3613 18528
rect 3549 18468 3553 18524
rect 3553 18468 3609 18524
rect 3609 18468 3613 18524
rect 3549 18464 3613 18468
rect 3629 18524 3693 18528
rect 3629 18468 3633 18524
rect 3633 18468 3689 18524
rect 3689 18468 3693 18524
rect 3629 18464 3693 18468
rect 3709 18524 3773 18528
rect 3709 18468 3713 18524
rect 3713 18468 3769 18524
rect 3769 18468 3773 18524
rect 3709 18464 3773 18468
rect 3789 18524 3853 18528
rect 3789 18468 3793 18524
rect 3793 18468 3849 18524
rect 3849 18468 3853 18524
rect 3789 18464 3853 18468
rect 6146 18524 6210 18528
rect 6146 18468 6150 18524
rect 6150 18468 6206 18524
rect 6206 18468 6210 18524
rect 6146 18464 6210 18468
rect 6226 18524 6290 18528
rect 6226 18468 6230 18524
rect 6230 18468 6286 18524
rect 6286 18468 6290 18524
rect 6226 18464 6290 18468
rect 6306 18524 6370 18528
rect 6306 18468 6310 18524
rect 6310 18468 6366 18524
rect 6366 18468 6370 18524
rect 6306 18464 6370 18468
rect 6386 18524 6450 18528
rect 6386 18468 6390 18524
rect 6390 18468 6446 18524
rect 6446 18468 6450 18524
rect 6386 18464 6450 18468
rect 2250 17980 2314 17984
rect 2250 17924 2254 17980
rect 2254 17924 2310 17980
rect 2310 17924 2314 17980
rect 2250 17920 2314 17924
rect 2330 17980 2394 17984
rect 2330 17924 2334 17980
rect 2334 17924 2390 17980
rect 2390 17924 2394 17980
rect 2330 17920 2394 17924
rect 2410 17980 2474 17984
rect 2410 17924 2414 17980
rect 2414 17924 2470 17980
rect 2470 17924 2474 17980
rect 2410 17920 2474 17924
rect 2490 17980 2554 17984
rect 2490 17924 2494 17980
rect 2494 17924 2550 17980
rect 2550 17924 2554 17980
rect 2490 17920 2554 17924
rect 4848 17980 4912 17984
rect 4848 17924 4852 17980
rect 4852 17924 4908 17980
rect 4908 17924 4912 17980
rect 4848 17920 4912 17924
rect 4928 17980 4992 17984
rect 4928 17924 4932 17980
rect 4932 17924 4988 17980
rect 4988 17924 4992 17980
rect 4928 17920 4992 17924
rect 5008 17980 5072 17984
rect 5008 17924 5012 17980
rect 5012 17924 5068 17980
rect 5068 17924 5072 17980
rect 5008 17920 5072 17924
rect 5088 17980 5152 17984
rect 5088 17924 5092 17980
rect 5092 17924 5148 17980
rect 5148 17924 5152 17980
rect 5088 17920 5152 17924
rect 7445 17980 7509 17984
rect 7445 17924 7449 17980
rect 7449 17924 7505 17980
rect 7505 17924 7509 17980
rect 7445 17920 7509 17924
rect 7525 17980 7589 17984
rect 7525 17924 7529 17980
rect 7529 17924 7585 17980
rect 7585 17924 7589 17980
rect 7525 17920 7589 17924
rect 7605 17980 7669 17984
rect 7605 17924 7609 17980
rect 7609 17924 7665 17980
rect 7665 17924 7669 17980
rect 7605 17920 7669 17924
rect 7685 17980 7749 17984
rect 7685 17924 7689 17980
rect 7689 17924 7745 17980
rect 7745 17924 7749 17980
rect 7685 17920 7749 17924
rect 3549 17436 3613 17440
rect 3549 17380 3553 17436
rect 3553 17380 3609 17436
rect 3609 17380 3613 17436
rect 3549 17376 3613 17380
rect 3629 17436 3693 17440
rect 3629 17380 3633 17436
rect 3633 17380 3689 17436
rect 3689 17380 3693 17436
rect 3629 17376 3693 17380
rect 3709 17436 3773 17440
rect 3709 17380 3713 17436
rect 3713 17380 3769 17436
rect 3769 17380 3773 17436
rect 3709 17376 3773 17380
rect 3789 17436 3853 17440
rect 3789 17380 3793 17436
rect 3793 17380 3849 17436
rect 3849 17380 3853 17436
rect 3789 17376 3853 17380
rect 6146 17436 6210 17440
rect 6146 17380 6150 17436
rect 6150 17380 6206 17436
rect 6206 17380 6210 17436
rect 6146 17376 6210 17380
rect 6226 17436 6290 17440
rect 6226 17380 6230 17436
rect 6230 17380 6286 17436
rect 6286 17380 6290 17436
rect 6226 17376 6290 17380
rect 6306 17436 6370 17440
rect 6306 17380 6310 17436
rect 6310 17380 6366 17436
rect 6366 17380 6370 17436
rect 6306 17376 6370 17380
rect 6386 17436 6450 17440
rect 6386 17380 6390 17436
rect 6390 17380 6446 17436
rect 6446 17380 6450 17436
rect 6386 17376 6450 17380
rect 2250 16892 2314 16896
rect 2250 16836 2254 16892
rect 2254 16836 2310 16892
rect 2310 16836 2314 16892
rect 2250 16832 2314 16836
rect 2330 16892 2394 16896
rect 2330 16836 2334 16892
rect 2334 16836 2390 16892
rect 2390 16836 2394 16892
rect 2330 16832 2394 16836
rect 2410 16892 2474 16896
rect 2410 16836 2414 16892
rect 2414 16836 2470 16892
rect 2470 16836 2474 16892
rect 2410 16832 2474 16836
rect 2490 16892 2554 16896
rect 2490 16836 2494 16892
rect 2494 16836 2550 16892
rect 2550 16836 2554 16892
rect 2490 16832 2554 16836
rect 4848 16892 4912 16896
rect 4848 16836 4852 16892
rect 4852 16836 4908 16892
rect 4908 16836 4912 16892
rect 4848 16832 4912 16836
rect 4928 16892 4992 16896
rect 4928 16836 4932 16892
rect 4932 16836 4988 16892
rect 4988 16836 4992 16892
rect 4928 16832 4992 16836
rect 5008 16892 5072 16896
rect 5008 16836 5012 16892
rect 5012 16836 5068 16892
rect 5068 16836 5072 16892
rect 5008 16832 5072 16836
rect 5088 16892 5152 16896
rect 5088 16836 5092 16892
rect 5092 16836 5148 16892
rect 5148 16836 5152 16892
rect 5088 16832 5152 16836
rect 7445 16892 7509 16896
rect 7445 16836 7449 16892
rect 7449 16836 7505 16892
rect 7505 16836 7509 16892
rect 7445 16832 7509 16836
rect 7525 16892 7589 16896
rect 7525 16836 7529 16892
rect 7529 16836 7585 16892
rect 7585 16836 7589 16892
rect 7525 16832 7589 16836
rect 7605 16892 7669 16896
rect 7605 16836 7609 16892
rect 7609 16836 7665 16892
rect 7665 16836 7669 16892
rect 7605 16832 7669 16836
rect 7685 16892 7749 16896
rect 7685 16836 7689 16892
rect 7689 16836 7745 16892
rect 7745 16836 7749 16892
rect 7685 16832 7749 16836
rect 3549 16348 3613 16352
rect 3549 16292 3553 16348
rect 3553 16292 3609 16348
rect 3609 16292 3613 16348
rect 3549 16288 3613 16292
rect 3629 16348 3693 16352
rect 3629 16292 3633 16348
rect 3633 16292 3689 16348
rect 3689 16292 3693 16348
rect 3629 16288 3693 16292
rect 3709 16348 3773 16352
rect 3709 16292 3713 16348
rect 3713 16292 3769 16348
rect 3769 16292 3773 16348
rect 3709 16288 3773 16292
rect 3789 16348 3853 16352
rect 3789 16292 3793 16348
rect 3793 16292 3849 16348
rect 3849 16292 3853 16348
rect 3789 16288 3853 16292
rect 6146 16348 6210 16352
rect 6146 16292 6150 16348
rect 6150 16292 6206 16348
rect 6206 16292 6210 16348
rect 6146 16288 6210 16292
rect 6226 16348 6290 16352
rect 6226 16292 6230 16348
rect 6230 16292 6286 16348
rect 6286 16292 6290 16348
rect 6226 16288 6290 16292
rect 6306 16348 6370 16352
rect 6306 16292 6310 16348
rect 6310 16292 6366 16348
rect 6366 16292 6370 16348
rect 6306 16288 6370 16292
rect 6386 16348 6450 16352
rect 6386 16292 6390 16348
rect 6390 16292 6446 16348
rect 6446 16292 6450 16348
rect 6386 16288 6450 16292
rect 2250 15804 2314 15808
rect 2250 15748 2254 15804
rect 2254 15748 2310 15804
rect 2310 15748 2314 15804
rect 2250 15744 2314 15748
rect 2330 15804 2394 15808
rect 2330 15748 2334 15804
rect 2334 15748 2390 15804
rect 2390 15748 2394 15804
rect 2330 15744 2394 15748
rect 2410 15804 2474 15808
rect 2410 15748 2414 15804
rect 2414 15748 2470 15804
rect 2470 15748 2474 15804
rect 2410 15744 2474 15748
rect 2490 15804 2554 15808
rect 2490 15748 2494 15804
rect 2494 15748 2550 15804
rect 2550 15748 2554 15804
rect 2490 15744 2554 15748
rect 4848 15804 4912 15808
rect 4848 15748 4852 15804
rect 4852 15748 4908 15804
rect 4908 15748 4912 15804
rect 4848 15744 4912 15748
rect 4928 15804 4992 15808
rect 4928 15748 4932 15804
rect 4932 15748 4988 15804
rect 4988 15748 4992 15804
rect 4928 15744 4992 15748
rect 5008 15804 5072 15808
rect 5008 15748 5012 15804
rect 5012 15748 5068 15804
rect 5068 15748 5072 15804
rect 5008 15744 5072 15748
rect 5088 15804 5152 15808
rect 5088 15748 5092 15804
rect 5092 15748 5148 15804
rect 5148 15748 5152 15804
rect 5088 15744 5152 15748
rect 7445 15804 7509 15808
rect 7445 15748 7449 15804
rect 7449 15748 7505 15804
rect 7505 15748 7509 15804
rect 7445 15744 7509 15748
rect 7525 15804 7589 15808
rect 7525 15748 7529 15804
rect 7529 15748 7585 15804
rect 7585 15748 7589 15804
rect 7525 15744 7589 15748
rect 7605 15804 7669 15808
rect 7605 15748 7609 15804
rect 7609 15748 7665 15804
rect 7665 15748 7669 15804
rect 7605 15744 7669 15748
rect 7685 15804 7749 15808
rect 7685 15748 7689 15804
rect 7689 15748 7745 15804
rect 7745 15748 7749 15804
rect 7685 15744 7749 15748
rect 3549 15260 3613 15264
rect 3549 15204 3553 15260
rect 3553 15204 3609 15260
rect 3609 15204 3613 15260
rect 3549 15200 3613 15204
rect 3629 15260 3693 15264
rect 3629 15204 3633 15260
rect 3633 15204 3689 15260
rect 3689 15204 3693 15260
rect 3629 15200 3693 15204
rect 3709 15260 3773 15264
rect 3709 15204 3713 15260
rect 3713 15204 3769 15260
rect 3769 15204 3773 15260
rect 3709 15200 3773 15204
rect 3789 15260 3853 15264
rect 3789 15204 3793 15260
rect 3793 15204 3849 15260
rect 3849 15204 3853 15260
rect 3789 15200 3853 15204
rect 6146 15260 6210 15264
rect 6146 15204 6150 15260
rect 6150 15204 6206 15260
rect 6206 15204 6210 15260
rect 6146 15200 6210 15204
rect 6226 15260 6290 15264
rect 6226 15204 6230 15260
rect 6230 15204 6286 15260
rect 6286 15204 6290 15260
rect 6226 15200 6290 15204
rect 6306 15260 6370 15264
rect 6306 15204 6310 15260
rect 6310 15204 6366 15260
rect 6366 15204 6370 15260
rect 6306 15200 6370 15204
rect 6386 15260 6450 15264
rect 6386 15204 6390 15260
rect 6390 15204 6446 15260
rect 6446 15204 6450 15260
rect 6386 15200 6450 15204
rect 2250 14716 2314 14720
rect 2250 14660 2254 14716
rect 2254 14660 2310 14716
rect 2310 14660 2314 14716
rect 2250 14656 2314 14660
rect 2330 14716 2394 14720
rect 2330 14660 2334 14716
rect 2334 14660 2390 14716
rect 2390 14660 2394 14716
rect 2330 14656 2394 14660
rect 2410 14716 2474 14720
rect 2410 14660 2414 14716
rect 2414 14660 2470 14716
rect 2470 14660 2474 14716
rect 2410 14656 2474 14660
rect 2490 14716 2554 14720
rect 2490 14660 2494 14716
rect 2494 14660 2550 14716
rect 2550 14660 2554 14716
rect 2490 14656 2554 14660
rect 4848 14716 4912 14720
rect 4848 14660 4852 14716
rect 4852 14660 4908 14716
rect 4908 14660 4912 14716
rect 4848 14656 4912 14660
rect 4928 14716 4992 14720
rect 4928 14660 4932 14716
rect 4932 14660 4988 14716
rect 4988 14660 4992 14716
rect 4928 14656 4992 14660
rect 5008 14716 5072 14720
rect 5008 14660 5012 14716
rect 5012 14660 5068 14716
rect 5068 14660 5072 14716
rect 5008 14656 5072 14660
rect 5088 14716 5152 14720
rect 5088 14660 5092 14716
rect 5092 14660 5148 14716
rect 5148 14660 5152 14716
rect 5088 14656 5152 14660
rect 7445 14716 7509 14720
rect 7445 14660 7449 14716
rect 7449 14660 7505 14716
rect 7505 14660 7509 14716
rect 7445 14656 7509 14660
rect 7525 14716 7589 14720
rect 7525 14660 7529 14716
rect 7529 14660 7585 14716
rect 7585 14660 7589 14716
rect 7525 14656 7589 14660
rect 7605 14716 7669 14720
rect 7605 14660 7609 14716
rect 7609 14660 7665 14716
rect 7665 14660 7669 14716
rect 7605 14656 7669 14660
rect 7685 14716 7749 14720
rect 7685 14660 7689 14716
rect 7689 14660 7745 14716
rect 7745 14660 7749 14716
rect 7685 14656 7749 14660
rect 3549 14172 3613 14176
rect 3549 14116 3553 14172
rect 3553 14116 3609 14172
rect 3609 14116 3613 14172
rect 3549 14112 3613 14116
rect 3629 14172 3693 14176
rect 3629 14116 3633 14172
rect 3633 14116 3689 14172
rect 3689 14116 3693 14172
rect 3629 14112 3693 14116
rect 3709 14172 3773 14176
rect 3709 14116 3713 14172
rect 3713 14116 3769 14172
rect 3769 14116 3773 14172
rect 3709 14112 3773 14116
rect 3789 14172 3853 14176
rect 3789 14116 3793 14172
rect 3793 14116 3849 14172
rect 3849 14116 3853 14172
rect 3789 14112 3853 14116
rect 6146 14172 6210 14176
rect 6146 14116 6150 14172
rect 6150 14116 6206 14172
rect 6206 14116 6210 14172
rect 6146 14112 6210 14116
rect 6226 14172 6290 14176
rect 6226 14116 6230 14172
rect 6230 14116 6286 14172
rect 6286 14116 6290 14172
rect 6226 14112 6290 14116
rect 6306 14172 6370 14176
rect 6306 14116 6310 14172
rect 6310 14116 6366 14172
rect 6366 14116 6370 14172
rect 6306 14112 6370 14116
rect 6386 14172 6450 14176
rect 6386 14116 6390 14172
rect 6390 14116 6446 14172
rect 6446 14116 6450 14172
rect 6386 14112 6450 14116
rect 2250 13628 2314 13632
rect 2250 13572 2254 13628
rect 2254 13572 2310 13628
rect 2310 13572 2314 13628
rect 2250 13568 2314 13572
rect 2330 13628 2394 13632
rect 2330 13572 2334 13628
rect 2334 13572 2390 13628
rect 2390 13572 2394 13628
rect 2330 13568 2394 13572
rect 2410 13628 2474 13632
rect 2410 13572 2414 13628
rect 2414 13572 2470 13628
rect 2470 13572 2474 13628
rect 2410 13568 2474 13572
rect 2490 13628 2554 13632
rect 2490 13572 2494 13628
rect 2494 13572 2550 13628
rect 2550 13572 2554 13628
rect 2490 13568 2554 13572
rect 4848 13628 4912 13632
rect 4848 13572 4852 13628
rect 4852 13572 4908 13628
rect 4908 13572 4912 13628
rect 4848 13568 4912 13572
rect 4928 13628 4992 13632
rect 4928 13572 4932 13628
rect 4932 13572 4988 13628
rect 4988 13572 4992 13628
rect 4928 13568 4992 13572
rect 5008 13628 5072 13632
rect 5008 13572 5012 13628
rect 5012 13572 5068 13628
rect 5068 13572 5072 13628
rect 5008 13568 5072 13572
rect 5088 13628 5152 13632
rect 5088 13572 5092 13628
rect 5092 13572 5148 13628
rect 5148 13572 5152 13628
rect 5088 13568 5152 13572
rect 7445 13628 7509 13632
rect 7445 13572 7449 13628
rect 7449 13572 7505 13628
rect 7505 13572 7509 13628
rect 7445 13568 7509 13572
rect 7525 13628 7589 13632
rect 7525 13572 7529 13628
rect 7529 13572 7585 13628
rect 7585 13572 7589 13628
rect 7525 13568 7589 13572
rect 7605 13628 7669 13632
rect 7605 13572 7609 13628
rect 7609 13572 7665 13628
rect 7665 13572 7669 13628
rect 7605 13568 7669 13572
rect 7685 13628 7749 13632
rect 7685 13572 7689 13628
rect 7689 13572 7745 13628
rect 7745 13572 7749 13628
rect 7685 13568 7749 13572
rect 3549 13084 3613 13088
rect 3549 13028 3553 13084
rect 3553 13028 3609 13084
rect 3609 13028 3613 13084
rect 3549 13024 3613 13028
rect 3629 13084 3693 13088
rect 3629 13028 3633 13084
rect 3633 13028 3689 13084
rect 3689 13028 3693 13084
rect 3629 13024 3693 13028
rect 3709 13084 3773 13088
rect 3709 13028 3713 13084
rect 3713 13028 3769 13084
rect 3769 13028 3773 13084
rect 3709 13024 3773 13028
rect 3789 13084 3853 13088
rect 3789 13028 3793 13084
rect 3793 13028 3849 13084
rect 3849 13028 3853 13084
rect 3789 13024 3853 13028
rect 6146 13084 6210 13088
rect 6146 13028 6150 13084
rect 6150 13028 6206 13084
rect 6206 13028 6210 13084
rect 6146 13024 6210 13028
rect 6226 13084 6290 13088
rect 6226 13028 6230 13084
rect 6230 13028 6286 13084
rect 6286 13028 6290 13084
rect 6226 13024 6290 13028
rect 6306 13084 6370 13088
rect 6306 13028 6310 13084
rect 6310 13028 6366 13084
rect 6366 13028 6370 13084
rect 6306 13024 6370 13028
rect 6386 13084 6450 13088
rect 6386 13028 6390 13084
rect 6390 13028 6446 13084
rect 6446 13028 6450 13084
rect 6386 13024 6450 13028
rect 2250 12540 2314 12544
rect 2250 12484 2254 12540
rect 2254 12484 2310 12540
rect 2310 12484 2314 12540
rect 2250 12480 2314 12484
rect 2330 12540 2394 12544
rect 2330 12484 2334 12540
rect 2334 12484 2390 12540
rect 2390 12484 2394 12540
rect 2330 12480 2394 12484
rect 2410 12540 2474 12544
rect 2410 12484 2414 12540
rect 2414 12484 2470 12540
rect 2470 12484 2474 12540
rect 2410 12480 2474 12484
rect 2490 12540 2554 12544
rect 2490 12484 2494 12540
rect 2494 12484 2550 12540
rect 2550 12484 2554 12540
rect 2490 12480 2554 12484
rect 4848 12540 4912 12544
rect 4848 12484 4852 12540
rect 4852 12484 4908 12540
rect 4908 12484 4912 12540
rect 4848 12480 4912 12484
rect 4928 12540 4992 12544
rect 4928 12484 4932 12540
rect 4932 12484 4988 12540
rect 4988 12484 4992 12540
rect 4928 12480 4992 12484
rect 5008 12540 5072 12544
rect 5008 12484 5012 12540
rect 5012 12484 5068 12540
rect 5068 12484 5072 12540
rect 5008 12480 5072 12484
rect 5088 12540 5152 12544
rect 5088 12484 5092 12540
rect 5092 12484 5148 12540
rect 5148 12484 5152 12540
rect 5088 12480 5152 12484
rect 7445 12540 7509 12544
rect 7445 12484 7449 12540
rect 7449 12484 7505 12540
rect 7505 12484 7509 12540
rect 7445 12480 7509 12484
rect 7525 12540 7589 12544
rect 7525 12484 7529 12540
rect 7529 12484 7585 12540
rect 7585 12484 7589 12540
rect 7525 12480 7589 12484
rect 7605 12540 7669 12544
rect 7605 12484 7609 12540
rect 7609 12484 7665 12540
rect 7665 12484 7669 12540
rect 7605 12480 7669 12484
rect 7685 12540 7749 12544
rect 7685 12484 7689 12540
rect 7689 12484 7745 12540
rect 7745 12484 7749 12540
rect 7685 12480 7749 12484
rect 3549 11996 3613 12000
rect 3549 11940 3553 11996
rect 3553 11940 3609 11996
rect 3609 11940 3613 11996
rect 3549 11936 3613 11940
rect 3629 11996 3693 12000
rect 3629 11940 3633 11996
rect 3633 11940 3689 11996
rect 3689 11940 3693 11996
rect 3629 11936 3693 11940
rect 3709 11996 3773 12000
rect 3709 11940 3713 11996
rect 3713 11940 3769 11996
rect 3769 11940 3773 11996
rect 3709 11936 3773 11940
rect 3789 11996 3853 12000
rect 3789 11940 3793 11996
rect 3793 11940 3849 11996
rect 3849 11940 3853 11996
rect 3789 11936 3853 11940
rect 6146 11996 6210 12000
rect 6146 11940 6150 11996
rect 6150 11940 6206 11996
rect 6206 11940 6210 11996
rect 6146 11936 6210 11940
rect 6226 11996 6290 12000
rect 6226 11940 6230 11996
rect 6230 11940 6286 11996
rect 6286 11940 6290 11996
rect 6226 11936 6290 11940
rect 6306 11996 6370 12000
rect 6306 11940 6310 11996
rect 6310 11940 6366 11996
rect 6366 11940 6370 11996
rect 6306 11936 6370 11940
rect 6386 11996 6450 12000
rect 6386 11940 6390 11996
rect 6390 11940 6446 11996
rect 6446 11940 6450 11996
rect 6386 11936 6450 11940
rect 2250 11452 2314 11456
rect 2250 11396 2254 11452
rect 2254 11396 2310 11452
rect 2310 11396 2314 11452
rect 2250 11392 2314 11396
rect 2330 11452 2394 11456
rect 2330 11396 2334 11452
rect 2334 11396 2390 11452
rect 2390 11396 2394 11452
rect 2330 11392 2394 11396
rect 2410 11452 2474 11456
rect 2410 11396 2414 11452
rect 2414 11396 2470 11452
rect 2470 11396 2474 11452
rect 2410 11392 2474 11396
rect 2490 11452 2554 11456
rect 2490 11396 2494 11452
rect 2494 11396 2550 11452
rect 2550 11396 2554 11452
rect 2490 11392 2554 11396
rect 4848 11452 4912 11456
rect 4848 11396 4852 11452
rect 4852 11396 4908 11452
rect 4908 11396 4912 11452
rect 4848 11392 4912 11396
rect 4928 11452 4992 11456
rect 4928 11396 4932 11452
rect 4932 11396 4988 11452
rect 4988 11396 4992 11452
rect 4928 11392 4992 11396
rect 5008 11452 5072 11456
rect 5008 11396 5012 11452
rect 5012 11396 5068 11452
rect 5068 11396 5072 11452
rect 5008 11392 5072 11396
rect 5088 11452 5152 11456
rect 5088 11396 5092 11452
rect 5092 11396 5148 11452
rect 5148 11396 5152 11452
rect 5088 11392 5152 11396
rect 7445 11452 7509 11456
rect 7445 11396 7449 11452
rect 7449 11396 7505 11452
rect 7505 11396 7509 11452
rect 7445 11392 7509 11396
rect 7525 11452 7589 11456
rect 7525 11396 7529 11452
rect 7529 11396 7585 11452
rect 7585 11396 7589 11452
rect 7525 11392 7589 11396
rect 7605 11452 7669 11456
rect 7605 11396 7609 11452
rect 7609 11396 7665 11452
rect 7665 11396 7669 11452
rect 7605 11392 7669 11396
rect 7685 11452 7749 11456
rect 7685 11396 7689 11452
rect 7689 11396 7745 11452
rect 7745 11396 7749 11452
rect 7685 11392 7749 11396
rect 3549 10908 3613 10912
rect 3549 10852 3553 10908
rect 3553 10852 3609 10908
rect 3609 10852 3613 10908
rect 3549 10848 3613 10852
rect 3629 10908 3693 10912
rect 3629 10852 3633 10908
rect 3633 10852 3689 10908
rect 3689 10852 3693 10908
rect 3629 10848 3693 10852
rect 3709 10908 3773 10912
rect 3709 10852 3713 10908
rect 3713 10852 3769 10908
rect 3769 10852 3773 10908
rect 3709 10848 3773 10852
rect 3789 10908 3853 10912
rect 3789 10852 3793 10908
rect 3793 10852 3849 10908
rect 3849 10852 3853 10908
rect 3789 10848 3853 10852
rect 6146 10908 6210 10912
rect 6146 10852 6150 10908
rect 6150 10852 6206 10908
rect 6206 10852 6210 10908
rect 6146 10848 6210 10852
rect 6226 10908 6290 10912
rect 6226 10852 6230 10908
rect 6230 10852 6286 10908
rect 6286 10852 6290 10908
rect 6226 10848 6290 10852
rect 6306 10908 6370 10912
rect 6306 10852 6310 10908
rect 6310 10852 6366 10908
rect 6366 10852 6370 10908
rect 6306 10848 6370 10852
rect 6386 10908 6450 10912
rect 6386 10852 6390 10908
rect 6390 10852 6446 10908
rect 6446 10852 6450 10908
rect 6386 10848 6450 10852
rect 2250 10364 2314 10368
rect 2250 10308 2254 10364
rect 2254 10308 2310 10364
rect 2310 10308 2314 10364
rect 2250 10304 2314 10308
rect 2330 10364 2394 10368
rect 2330 10308 2334 10364
rect 2334 10308 2390 10364
rect 2390 10308 2394 10364
rect 2330 10304 2394 10308
rect 2410 10364 2474 10368
rect 2410 10308 2414 10364
rect 2414 10308 2470 10364
rect 2470 10308 2474 10364
rect 2410 10304 2474 10308
rect 2490 10364 2554 10368
rect 2490 10308 2494 10364
rect 2494 10308 2550 10364
rect 2550 10308 2554 10364
rect 2490 10304 2554 10308
rect 4848 10364 4912 10368
rect 4848 10308 4852 10364
rect 4852 10308 4908 10364
rect 4908 10308 4912 10364
rect 4848 10304 4912 10308
rect 4928 10364 4992 10368
rect 4928 10308 4932 10364
rect 4932 10308 4988 10364
rect 4988 10308 4992 10364
rect 4928 10304 4992 10308
rect 5008 10364 5072 10368
rect 5008 10308 5012 10364
rect 5012 10308 5068 10364
rect 5068 10308 5072 10364
rect 5008 10304 5072 10308
rect 5088 10364 5152 10368
rect 5088 10308 5092 10364
rect 5092 10308 5148 10364
rect 5148 10308 5152 10364
rect 5088 10304 5152 10308
rect 7445 10364 7509 10368
rect 7445 10308 7449 10364
rect 7449 10308 7505 10364
rect 7505 10308 7509 10364
rect 7445 10304 7509 10308
rect 7525 10364 7589 10368
rect 7525 10308 7529 10364
rect 7529 10308 7585 10364
rect 7585 10308 7589 10364
rect 7525 10304 7589 10308
rect 7605 10364 7669 10368
rect 7605 10308 7609 10364
rect 7609 10308 7665 10364
rect 7665 10308 7669 10364
rect 7605 10304 7669 10308
rect 7685 10364 7749 10368
rect 7685 10308 7689 10364
rect 7689 10308 7745 10364
rect 7745 10308 7749 10364
rect 7685 10304 7749 10308
rect 3549 9820 3613 9824
rect 3549 9764 3553 9820
rect 3553 9764 3609 9820
rect 3609 9764 3613 9820
rect 3549 9760 3613 9764
rect 3629 9820 3693 9824
rect 3629 9764 3633 9820
rect 3633 9764 3689 9820
rect 3689 9764 3693 9820
rect 3629 9760 3693 9764
rect 3709 9820 3773 9824
rect 3709 9764 3713 9820
rect 3713 9764 3769 9820
rect 3769 9764 3773 9820
rect 3709 9760 3773 9764
rect 3789 9820 3853 9824
rect 3789 9764 3793 9820
rect 3793 9764 3849 9820
rect 3849 9764 3853 9820
rect 3789 9760 3853 9764
rect 6146 9820 6210 9824
rect 6146 9764 6150 9820
rect 6150 9764 6206 9820
rect 6206 9764 6210 9820
rect 6146 9760 6210 9764
rect 6226 9820 6290 9824
rect 6226 9764 6230 9820
rect 6230 9764 6286 9820
rect 6286 9764 6290 9820
rect 6226 9760 6290 9764
rect 6306 9820 6370 9824
rect 6306 9764 6310 9820
rect 6310 9764 6366 9820
rect 6366 9764 6370 9820
rect 6306 9760 6370 9764
rect 6386 9820 6450 9824
rect 6386 9764 6390 9820
rect 6390 9764 6446 9820
rect 6446 9764 6450 9820
rect 6386 9760 6450 9764
rect 2250 9276 2314 9280
rect 2250 9220 2254 9276
rect 2254 9220 2310 9276
rect 2310 9220 2314 9276
rect 2250 9216 2314 9220
rect 2330 9276 2394 9280
rect 2330 9220 2334 9276
rect 2334 9220 2390 9276
rect 2390 9220 2394 9276
rect 2330 9216 2394 9220
rect 2410 9276 2474 9280
rect 2410 9220 2414 9276
rect 2414 9220 2470 9276
rect 2470 9220 2474 9276
rect 2410 9216 2474 9220
rect 2490 9276 2554 9280
rect 2490 9220 2494 9276
rect 2494 9220 2550 9276
rect 2550 9220 2554 9276
rect 2490 9216 2554 9220
rect 4848 9276 4912 9280
rect 4848 9220 4852 9276
rect 4852 9220 4908 9276
rect 4908 9220 4912 9276
rect 4848 9216 4912 9220
rect 4928 9276 4992 9280
rect 4928 9220 4932 9276
rect 4932 9220 4988 9276
rect 4988 9220 4992 9276
rect 4928 9216 4992 9220
rect 5008 9276 5072 9280
rect 5008 9220 5012 9276
rect 5012 9220 5068 9276
rect 5068 9220 5072 9276
rect 5008 9216 5072 9220
rect 5088 9276 5152 9280
rect 5088 9220 5092 9276
rect 5092 9220 5148 9276
rect 5148 9220 5152 9276
rect 5088 9216 5152 9220
rect 7445 9276 7509 9280
rect 7445 9220 7449 9276
rect 7449 9220 7505 9276
rect 7505 9220 7509 9276
rect 7445 9216 7509 9220
rect 7525 9276 7589 9280
rect 7525 9220 7529 9276
rect 7529 9220 7585 9276
rect 7585 9220 7589 9276
rect 7525 9216 7589 9220
rect 7605 9276 7669 9280
rect 7605 9220 7609 9276
rect 7609 9220 7665 9276
rect 7665 9220 7669 9276
rect 7605 9216 7669 9220
rect 7685 9276 7749 9280
rect 7685 9220 7689 9276
rect 7689 9220 7745 9276
rect 7745 9220 7749 9276
rect 7685 9216 7749 9220
rect 3549 8732 3613 8736
rect 3549 8676 3553 8732
rect 3553 8676 3609 8732
rect 3609 8676 3613 8732
rect 3549 8672 3613 8676
rect 3629 8732 3693 8736
rect 3629 8676 3633 8732
rect 3633 8676 3689 8732
rect 3689 8676 3693 8732
rect 3629 8672 3693 8676
rect 3709 8732 3773 8736
rect 3709 8676 3713 8732
rect 3713 8676 3769 8732
rect 3769 8676 3773 8732
rect 3709 8672 3773 8676
rect 3789 8732 3853 8736
rect 3789 8676 3793 8732
rect 3793 8676 3849 8732
rect 3849 8676 3853 8732
rect 3789 8672 3853 8676
rect 6146 8732 6210 8736
rect 6146 8676 6150 8732
rect 6150 8676 6206 8732
rect 6206 8676 6210 8732
rect 6146 8672 6210 8676
rect 6226 8732 6290 8736
rect 6226 8676 6230 8732
rect 6230 8676 6286 8732
rect 6286 8676 6290 8732
rect 6226 8672 6290 8676
rect 6306 8732 6370 8736
rect 6306 8676 6310 8732
rect 6310 8676 6366 8732
rect 6366 8676 6370 8732
rect 6306 8672 6370 8676
rect 6386 8732 6450 8736
rect 6386 8676 6390 8732
rect 6390 8676 6446 8732
rect 6446 8676 6450 8732
rect 6386 8672 6450 8676
rect 2250 8188 2314 8192
rect 2250 8132 2254 8188
rect 2254 8132 2310 8188
rect 2310 8132 2314 8188
rect 2250 8128 2314 8132
rect 2330 8188 2394 8192
rect 2330 8132 2334 8188
rect 2334 8132 2390 8188
rect 2390 8132 2394 8188
rect 2330 8128 2394 8132
rect 2410 8188 2474 8192
rect 2410 8132 2414 8188
rect 2414 8132 2470 8188
rect 2470 8132 2474 8188
rect 2410 8128 2474 8132
rect 2490 8188 2554 8192
rect 2490 8132 2494 8188
rect 2494 8132 2550 8188
rect 2550 8132 2554 8188
rect 2490 8128 2554 8132
rect 4848 8188 4912 8192
rect 4848 8132 4852 8188
rect 4852 8132 4908 8188
rect 4908 8132 4912 8188
rect 4848 8128 4912 8132
rect 4928 8188 4992 8192
rect 4928 8132 4932 8188
rect 4932 8132 4988 8188
rect 4988 8132 4992 8188
rect 4928 8128 4992 8132
rect 5008 8188 5072 8192
rect 5008 8132 5012 8188
rect 5012 8132 5068 8188
rect 5068 8132 5072 8188
rect 5008 8128 5072 8132
rect 5088 8188 5152 8192
rect 5088 8132 5092 8188
rect 5092 8132 5148 8188
rect 5148 8132 5152 8188
rect 5088 8128 5152 8132
rect 7445 8188 7509 8192
rect 7445 8132 7449 8188
rect 7449 8132 7505 8188
rect 7505 8132 7509 8188
rect 7445 8128 7509 8132
rect 7525 8188 7589 8192
rect 7525 8132 7529 8188
rect 7529 8132 7585 8188
rect 7585 8132 7589 8188
rect 7525 8128 7589 8132
rect 7605 8188 7669 8192
rect 7605 8132 7609 8188
rect 7609 8132 7665 8188
rect 7665 8132 7669 8188
rect 7605 8128 7669 8132
rect 7685 8188 7749 8192
rect 7685 8132 7689 8188
rect 7689 8132 7745 8188
rect 7745 8132 7749 8188
rect 7685 8128 7749 8132
rect 3549 7644 3613 7648
rect 3549 7588 3553 7644
rect 3553 7588 3609 7644
rect 3609 7588 3613 7644
rect 3549 7584 3613 7588
rect 3629 7644 3693 7648
rect 3629 7588 3633 7644
rect 3633 7588 3689 7644
rect 3689 7588 3693 7644
rect 3629 7584 3693 7588
rect 3709 7644 3773 7648
rect 3709 7588 3713 7644
rect 3713 7588 3769 7644
rect 3769 7588 3773 7644
rect 3709 7584 3773 7588
rect 3789 7644 3853 7648
rect 3789 7588 3793 7644
rect 3793 7588 3849 7644
rect 3849 7588 3853 7644
rect 3789 7584 3853 7588
rect 6146 7644 6210 7648
rect 6146 7588 6150 7644
rect 6150 7588 6206 7644
rect 6206 7588 6210 7644
rect 6146 7584 6210 7588
rect 6226 7644 6290 7648
rect 6226 7588 6230 7644
rect 6230 7588 6286 7644
rect 6286 7588 6290 7644
rect 6226 7584 6290 7588
rect 6306 7644 6370 7648
rect 6306 7588 6310 7644
rect 6310 7588 6366 7644
rect 6366 7588 6370 7644
rect 6306 7584 6370 7588
rect 6386 7644 6450 7648
rect 6386 7588 6390 7644
rect 6390 7588 6446 7644
rect 6446 7588 6450 7644
rect 6386 7584 6450 7588
rect 2250 7100 2314 7104
rect 2250 7044 2254 7100
rect 2254 7044 2310 7100
rect 2310 7044 2314 7100
rect 2250 7040 2314 7044
rect 2330 7100 2394 7104
rect 2330 7044 2334 7100
rect 2334 7044 2390 7100
rect 2390 7044 2394 7100
rect 2330 7040 2394 7044
rect 2410 7100 2474 7104
rect 2410 7044 2414 7100
rect 2414 7044 2470 7100
rect 2470 7044 2474 7100
rect 2410 7040 2474 7044
rect 2490 7100 2554 7104
rect 2490 7044 2494 7100
rect 2494 7044 2550 7100
rect 2550 7044 2554 7100
rect 2490 7040 2554 7044
rect 4848 7100 4912 7104
rect 4848 7044 4852 7100
rect 4852 7044 4908 7100
rect 4908 7044 4912 7100
rect 4848 7040 4912 7044
rect 4928 7100 4992 7104
rect 4928 7044 4932 7100
rect 4932 7044 4988 7100
rect 4988 7044 4992 7100
rect 4928 7040 4992 7044
rect 5008 7100 5072 7104
rect 5008 7044 5012 7100
rect 5012 7044 5068 7100
rect 5068 7044 5072 7100
rect 5008 7040 5072 7044
rect 5088 7100 5152 7104
rect 5088 7044 5092 7100
rect 5092 7044 5148 7100
rect 5148 7044 5152 7100
rect 5088 7040 5152 7044
rect 7445 7100 7509 7104
rect 7445 7044 7449 7100
rect 7449 7044 7505 7100
rect 7505 7044 7509 7100
rect 7445 7040 7509 7044
rect 7525 7100 7589 7104
rect 7525 7044 7529 7100
rect 7529 7044 7585 7100
rect 7585 7044 7589 7100
rect 7525 7040 7589 7044
rect 7605 7100 7669 7104
rect 7605 7044 7609 7100
rect 7609 7044 7665 7100
rect 7665 7044 7669 7100
rect 7605 7040 7669 7044
rect 7685 7100 7749 7104
rect 7685 7044 7689 7100
rect 7689 7044 7745 7100
rect 7745 7044 7749 7100
rect 7685 7040 7749 7044
rect 3549 6556 3613 6560
rect 3549 6500 3553 6556
rect 3553 6500 3609 6556
rect 3609 6500 3613 6556
rect 3549 6496 3613 6500
rect 3629 6556 3693 6560
rect 3629 6500 3633 6556
rect 3633 6500 3689 6556
rect 3689 6500 3693 6556
rect 3629 6496 3693 6500
rect 3709 6556 3773 6560
rect 3709 6500 3713 6556
rect 3713 6500 3769 6556
rect 3769 6500 3773 6556
rect 3709 6496 3773 6500
rect 3789 6556 3853 6560
rect 3789 6500 3793 6556
rect 3793 6500 3849 6556
rect 3849 6500 3853 6556
rect 3789 6496 3853 6500
rect 6146 6556 6210 6560
rect 6146 6500 6150 6556
rect 6150 6500 6206 6556
rect 6206 6500 6210 6556
rect 6146 6496 6210 6500
rect 6226 6556 6290 6560
rect 6226 6500 6230 6556
rect 6230 6500 6286 6556
rect 6286 6500 6290 6556
rect 6226 6496 6290 6500
rect 6306 6556 6370 6560
rect 6306 6500 6310 6556
rect 6310 6500 6366 6556
rect 6366 6500 6370 6556
rect 6306 6496 6370 6500
rect 6386 6556 6450 6560
rect 6386 6500 6390 6556
rect 6390 6500 6446 6556
rect 6446 6500 6450 6556
rect 6386 6496 6450 6500
rect 2250 6012 2314 6016
rect 2250 5956 2254 6012
rect 2254 5956 2310 6012
rect 2310 5956 2314 6012
rect 2250 5952 2314 5956
rect 2330 6012 2394 6016
rect 2330 5956 2334 6012
rect 2334 5956 2390 6012
rect 2390 5956 2394 6012
rect 2330 5952 2394 5956
rect 2410 6012 2474 6016
rect 2410 5956 2414 6012
rect 2414 5956 2470 6012
rect 2470 5956 2474 6012
rect 2410 5952 2474 5956
rect 2490 6012 2554 6016
rect 2490 5956 2494 6012
rect 2494 5956 2550 6012
rect 2550 5956 2554 6012
rect 2490 5952 2554 5956
rect 4848 6012 4912 6016
rect 4848 5956 4852 6012
rect 4852 5956 4908 6012
rect 4908 5956 4912 6012
rect 4848 5952 4912 5956
rect 4928 6012 4992 6016
rect 4928 5956 4932 6012
rect 4932 5956 4988 6012
rect 4988 5956 4992 6012
rect 4928 5952 4992 5956
rect 5008 6012 5072 6016
rect 5008 5956 5012 6012
rect 5012 5956 5068 6012
rect 5068 5956 5072 6012
rect 5008 5952 5072 5956
rect 5088 6012 5152 6016
rect 5088 5956 5092 6012
rect 5092 5956 5148 6012
rect 5148 5956 5152 6012
rect 5088 5952 5152 5956
rect 7445 6012 7509 6016
rect 7445 5956 7449 6012
rect 7449 5956 7505 6012
rect 7505 5956 7509 6012
rect 7445 5952 7509 5956
rect 7525 6012 7589 6016
rect 7525 5956 7529 6012
rect 7529 5956 7585 6012
rect 7585 5956 7589 6012
rect 7525 5952 7589 5956
rect 7605 6012 7669 6016
rect 7605 5956 7609 6012
rect 7609 5956 7665 6012
rect 7665 5956 7669 6012
rect 7605 5952 7669 5956
rect 7685 6012 7749 6016
rect 7685 5956 7689 6012
rect 7689 5956 7745 6012
rect 7745 5956 7749 6012
rect 7685 5952 7749 5956
rect 3549 5468 3613 5472
rect 3549 5412 3553 5468
rect 3553 5412 3609 5468
rect 3609 5412 3613 5468
rect 3549 5408 3613 5412
rect 3629 5468 3693 5472
rect 3629 5412 3633 5468
rect 3633 5412 3689 5468
rect 3689 5412 3693 5468
rect 3629 5408 3693 5412
rect 3709 5468 3773 5472
rect 3709 5412 3713 5468
rect 3713 5412 3769 5468
rect 3769 5412 3773 5468
rect 3709 5408 3773 5412
rect 3789 5468 3853 5472
rect 3789 5412 3793 5468
rect 3793 5412 3849 5468
rect 3849 5412 3853 5468
rect 3789 5408 3853 5412
rect 6146 5468 6210 5472
rect 6146 5412 6150 5468
rect 6150 5412 6206 5468
rect 6206 5412 6210 5468
rect 6146 5408 6210 5412
rect 6226 5468 6290 5472
rect 6226 5412 6230 5468
rect 6230 5412 6286 5468
rect 6286 5412 6290 5468
rect 6226 5408 6290 5412
rect 6306 5468 6370 5472
rect 6306 5412 6310 5468
rect 6310 5412 6366 5468
rect 6366 5412 6370 5468
rect 6306 5408 6370 5412
rect 6386 5468 6450 5472
rect 6386 5412 6390 5468
rect 6390 5412 6446 5468
rect 6446 5412 6450 5468
rect 6386 5408 6450 5412
rect 2250 4924 2314 4928
rect 2250 4868 2254 4924
rect 2254 4868 2310 4924
rect 2310 4868 2314 4924
rect 2250 4864 2314 4868
rect 2330 4924 2394 4928
rect 2330 4868 2334 4924
rect 2334 4868 2390 4924
rect 2390 4868 2394 4924
rect 2330 4864 2394 4868
rect 2410 4924 2474 4928
rect 2410 4868 2414 4924
rect 2414 4868 2470 4924
rect 2470 4868 2474 4924
rect 2410 4864 2474 4868
rect 2490 4924 2554 4928
rect 2490 4868 2494 4924
rect 2494 4868 2550 4924
rect 2550 4868 2554 4924
rect 2490 4864 2554 4868
rect 4848 4924 4912 4928
rect 4848 4868 4852 4924
rect 4852 4868 4908 4924
rect 4908 4868 4912 4924
rect 4848 4864 4912 4868
rect 4928 4924 4992 4928
rect 4928 4868 4932 4924
rect 4932 4868 4988 4924
rect 4988 4868 4992 4924
rect 4928 4864 4992 4868
rect 5008 4924 5072 4928
rect 5008 4868 5012 4924
rect 5012 4868 5068 4924
rect 5068 4868 5072 4924
rect 5008 4864 5072 4868
rect 5088 4924 5152 4928
rect 5088 4868 5092 4924
rect 5092 4868 5148 4924
rect 5148 4868 5152 4924
rect 5088 4864 5152 4868
rect 7445 4924 7509 4928
rect 7445 4868 7449 4924
rect 7449 4868 7505 4924
rect 7505 4868 7509 4924
rect 7445 4864 7509 4868
rect 7525 4924 7589 4928
rect 7525 4868 7529 4924
rect 7529 4868 7585 4924
rect 7585 4868 7589 4924
rect 7525 4864 7589 4868
rect 7605 4924 7669 4928
rect 7605 4868 7609 4924
rect 7609 4868 7665 4924
rect 7665 4868 7669 4924
rect 7605 4864 7669 4868
rect 7685 4924 7749 4928
rect 7685 4868 7689 4924
rect 7689 4868 7745 4924
rect 7745 4868 7749 4924
rect 7685 4864 7749 4868
rect 3549 4380 3613 4384
rect 3549 4324 3553 4380
rect 3553 4324 3609 4380
rect 3609 4324 3613 4380
rect 3549 4320 3613 4324
rect 3629 4380 3693 4384
rect 3629 4324 3633 4380
rect 3633 4324 3689 4380
rect 3689 4324 3693 4380
rect 3629 4320 3693 4324
rect 3709 4380 3773 4384
rect 3709 4324 3713 4380
rect 3713 4324 3769 4380
rect 3769 4324 3773 4380
rect 3709 4320 3773 4324
rect 3789 4380 3853 4384
rect 3789 4324 3793 4380
rect 3793 4324 3849 4380
rect 3849 4324 3853 4380
rect 3789 4320 3853 4324
rect 6146 4380 6210 4384
rect 6146 4324 6150 4380
rect 6150 4324 6206 4380
rect 6206 4324 6210 4380
rect 6146 4320 6210 4324
rect 6226 4380 6290 4384
rect 6226 4324 6230 4380
rect 6230 4324 6286 4380
rect 6286 4324 6290 4380
rect 6226 4320 6290 4324
rect 6306 4380 6370 4384
rect 6306 4324 6310 4380
rect 6310 4324 6366 4380
rect 6366 4324 6370 4380
rect 6306 4320 6370 4324
rect 6386 4380 6450 4384
rect 6386 4324 6390 4380
rect 6390 4324 6446 4380
rect 6446 4324 6450 4380
rect 6386 4320 6450 4324
rect 2250 3836 2314 3840
rect 2250 3780 2254 3836
rect 2254 3780 2310 3836
rect 2310 3780 2314 3836
rect 2250 3776 2314 3780
rect 2330 3836 2394 3840
rect 2330 3780 2334 3836
rect 2334 3780 2390 3836
rect 2390 3780 2394 3836
rect 2330 3776 2394 3780
rect 2410 3836 2474 3840
rect 2410 3780 2414 3836
rect 2414 3780 2470 3836
rect 2470 3780 2474 3836
rect 2410 3776 2474 3780
rect 2490 3836 2554 3840
rect 2490 3780 2494 3836
rect 2494 3780 2550 3836
rect 2550 3780 2554 3836
rect 2490 3776 2554 3780
rect 4848 3836 4912 3840
rect 4848 3780 4852 3836
rect 4852 3780 4908 3836
rect 4908 3780 4912 3836
rect 4848 3776 4912 3780
rect 4928 3836 4992 3840
rect 4928 3780 4932 3836
rect 4932 3780 4988 3836
rect 4988 3780 4992 3836
rect 4928 3776 4992 3780
rect 5008 3836 5072 3840
rect 5008 3780 5012 3836
rect 5012 3780 5068 3836
rect 5068 3780 5072 3836
rect 5008 3776 5072 3780
rect 5088 3836 5152 3840
rect 5088 3780 5092 3836
rect 5092 3780 5148 3836
rect 5148 3780 5152 3836
rect 5088 3776 5152 3780
rect 7445 3836 7509 3840
rect 7445 3780 7449 3836
rect 7449 3780 7505 3836
rect 7505 3780 7509 3836
rect 7445 3776 7509 3780
rect 7525 3836 7589 3840
rect 7525 3780 7529 3836
rect 7529 3780 7585 3836
rect 7585 3780 7589 3836
rect 7525 3776 7589 3780
rect 7605 3836 7669 3840
rect 7605 3780 7609 3836
rect 7609 3780 7665 3836
rect 7665 3780 7669 3836
rect 7605 3776 7669 3780
rect 7685 3836 7749 3840
rect 7685 3780 7689 3836
rect 7689 3780 7745 3836
rect 7745 3780 7749 3836
rect 7685 3776 7749 3780
rect 3549 3292 3613 3296
rect 3549 3236 3553 3292
rect 3553 3236 3609 3292
rect 3609 3236 3613 3292
rect 3549 3232 3613 3236
rect 3629 3292 3693 3296
rect 3629 3236 3633 3292
rect 3633 3236 3689 3292
rect 3689 3236 3693 3292
rect 3629 3232 3693 3236
rect 3709 3292 3773 3296
rect 3709 3236 3713 3292
rect 3713 3236 3769 3292
rect 3769 3236 3773 3292
rect 3709 3232 3773 3236
rect 3789 3292 3853 3296
rect 3789 3236 3793 3292
rect 3793 3236 3849 3292
rect 3849 3236 3853 3292
rect 3789 3232 3853 3236
rect 6146 3292 6210 3296
rect 6146 3236 6150 3292
rect 6150 3236 6206 3292
rect 6206 3236 6210 3292
rect 6146 3232 6210 3236
rect 6226 3292 6290 3296
rect 6226 3236 6230 3292
rect 6230 3236 6286 3292
rect 6286 3236 6290 3292
rect 6226 3232 6290 3236
rect 6306 3292 6370 3296
rect 6306 3236 6310 3292
rect 6310 3236 6366 3292
rect 6366 3236 6370 3292
rect 6306 3232 6370 3236
rect 6386 3292 6450 3296
rect 6386 3236 6390 3292
rect 6390 3236 6446 3292
rect 6446 3236 6450 3292
rect 6386 3232 6450 3236
rect 2250 2748 2314 2752
rect 2250 2692 2254 2748
rect 2254 2692 2310 2748
rect 2310 2692 2314 2748
rect 2250 2688 2314 2692
rect 2330 2748 2394 2752
rect 2330 2692 2334 2748
rect 2334 2692 2390 2748
rect 2390 2692 2394 2748
rect 2330 2688 2394 2692
rect 2410 2748 2474 2752
rect 2410 2692 2414 2748
rect 2414 2692 2470 2748
rect 2470 2692 2474 2748
rect 2410 2688 2474 2692
rect 2490 2748 2554 2752
rect 2490 2692 2494 2748
rect 2494 2692 2550 2748
rect 2550 2692 2554 2748
rect 2490 2688 2554 2692
rect 4848 2748 4912 2752
rect 4848 2692 4852 2748
rect 4852 2692 4908 2748
rect 4908 2692 4912 2748
rect 4848 2688 4912 2692
rect 4928 2748 4992 2752
rect 4928 2692 4932 2748
rect 4932 2692 4988 2748
rect 4988 2692 4992 2748
rect 4928 2688 4992 2692
rect 5008 2748 5072 2752
rect 5008 2692 5012 2748
rect 5012 2692 5068 2748
rect 5068 2692 5072 2748
rect 5008 2688 5072 2692
rect 5088 2748 5152 2752
rect 5088 2692 5092 2748
rect 5092 2692 5148 2748
rect 5148 2692 5152 2748
rect 5088 2688 5152 2692
rect 7445 2748 7509 2752
rect 7445 2692 7449 2748
rect 7449 2692 7505 2748
rect 7505 2692 7509 2748
rect 7445 2688 7509 2692
rect 7525 2748 7589 2752
rect 7525 2692 7529 2748
rect 7529 2692 7585 2748
rect 7585 2692 7589 2748
rect 7525 2688 7589 2692
rect 7605 2748 7669 2752
rect 7605 2692 7609 2748
rect 7609 2692 7665 2748
rect 7665 2692 7669 2748
rect 7605 2688 7669 2692
rect 7685 2748 7749 2752
rect 7685 2692 7689 2748
rect 7689 2692 7745 2748
rect 7745 2692 7749 2748
rect 7685 2688 7749 2692
rect 3549 2204 3613 2208
rect 3549 2148 3553 2204
rect 3553 2148 3609 2204
rect 3609 2148 3613 2204
rect 3549 2144 3613 2148
rect 3629 2204 3693 2208
rect 3629 2148 3633 2204
rect 3633 2148 3689 2204
rect 3689 2148 3693 2204
rect 3629 2144 3693 2148
rect 3709 2204 3773 2208
rect 3709 2148 3713 2204
rect 3713 2148 3769 2204
rect 3769 2148 3773 2204
rect 3709 2144 3773 2148
rect 3789 2204 3853 2208
rect 3789 2148 3793 2204
rect 3793 2148 3849 2204
rect 3849 2148 3853 2204
rect 3789 2144 3853 2148
rect 6146 2204 6210 2208
rect 6146 2148 6150 2204
rect 6150 2148 6206 2204
rect 6206 2148 6210 2204
rect 6146 2144 6210 2148
rect 6226 2204 6290 2208
rect 6226 2148 6230 2204
rect 6230 2148 6286 2204
rect 6286 2148 6290 2204
rect 6226 2144 6290 2148
rect 6306 2204 6370 2208
rect 6306 2148 6310 2204
rect 6310 2148 6366 2204
rect 6366 2148 6370 2204
rect 6306 2144 6370 2148
rect 6386 2204 6450 2208
rect 6386 2148 6390 2204
rect 6390 2148 6446 2204
rect 6446 2148 6450 2204
rect 6386 2144 6450 2148
<< metal4 >>
rect 2242 27776 2563 27792
rect 2242 27712 2250 27776
rect 2314 27712 2330 27776
rect 2394 27712 2410 27776
rect 2474 27712 2490 27776
rect 2554 27712 2563 27776
rect 2242 26688 2563 27712
rect 2242 26624 2250 26688
rect 2314 26624 2330 26688
rect 2394 26624 2410 26688
rect 2474 26624 2490 26688
rect 2554 26624 2563 26688
rect 2242 25600 2563 26624
rect 2242 25536 2250 25600
rect 2314 25536 2330 25600
rect 2394 25536 2410 25600
rect 2474 25536 2490 25600
rect 2554 25536 2563 25600
rect 2242 24512 2563 25536
rect 2242 24448 2250 24512
rect 2314 24448 2330 24512
rect 2394 24448 2410 24512
rect 2474 24448 2490 24512
rect 2554 24448 2563 24512
rect 2242 23424 2563 24448
rect 2242 23360 2250 23424
rect 2314 23360 2330 23424
rect 2394 23360 2410 23424
rect 2474 23360 2490 23424
rect 2554 23360 2563 23424
rect 2242 22336 2563 23360
rect 2242 22272 2250 22336
rect 2314 22272 2330 22336
rect 2394 22272 2410 22336
rect 2474 22272 2490 22336
rect 2554 22272 2563 22336
rect 2242 21248 2563 22272
rect 2242 21184 2250 21248
rect 2314 21184 2330 21248
rect 2394 21184 2410 21248
rect 2474 21184 2490 21248
rect 2554 21184 2563 21248
rect 2242 20160 2563 21184
rect 2242 20096 2250 20160
rect 2314 20096 2330 20160
rect 2394 20096 2410 20160
rect 2474 20096 2490 20160
rect 2554 20096 2563 20160
rect 2242 19072 2563 20096
rect 2242 19008 2250 19072
rect 2314 19008 2330 19072
rect 2394 19008 2410 19072
rect 2474 19008 2490 19072
rect 2554 19008 2563 19072
rect 2242 17984 2563 19008
rect 2242 17920 2250 17984
rect 2314 17920 2330 17984
rect 2394 17920 2410 17984
rect 2474 17920 2490 17984
rect 2554 17920 2563 17984
rect 2242 16896 2563 17920
rect 2242 16832 2250 16896
rect 2314 16832 2330 16896
rect 2394 16832 2410 16896
rect 2474 16832 2490 16896
rect 2554 16832 2563 16896
rect 2242 15808 2563 16832
rect 2242 15744 2250 15808
rect 2314 15744 2330 15808
rect 2394 15744 2410 15808
rect 2474 15744 2490 15808
rect 2554 15744 2563 15808
rect 2242 14720 2563 15744
rect 2242 14656 2250 14720
rect 2314 14656 2330 14720
rect 2394 14656 2410 14720
rect 2474 14656 2490 14720
rect 2554 14656 2563 14720
rect 2242 13632 2563 14656
rect 2242 13568 2250 13632
rect 2314 13568 2330 13632
rect 2394 13568 2410 13632
rect 2474 13568 2490 13632
rect 2554 13568 2563 13632
rect 2242 12544 2563 13568
rect 2242 12480 2250 12544
rect 2314 12480 2330 12544
rect 2394 12480 2410 12544
rect 2474 12480 2490 12544
rect 2554 12480 2563 12544
rect 2242 11456 2563 12480
rect 2242 11392 2250 11456
rect 2314 11392 2330 11456
rect 2394 11392 2410 11456
rect 2474 11392 2490 11456
rect 2554 11392 2563 11456
rect 2242 10368 2563 11392
rect 2242 10304 2250 10368
rect 2314 10304 2330 10368
rect 2394 10304 2410 10368
rect 2474 10304 2490 10368
rect 2554 10304 2563 10368
rect 2242 9280 2563 10304
rect 2242 9216 2250 9280
rect 2314 9216 2330 9280
rect 2394 9216 2410 9280
rect 2474 9216 2490 9280
rect 2554 9216 2563 9280
rect 2242 8192 2563 9216
rect 2242 8128 2250 8192
rect 2314 8128 2330 8192
rect 2394 8128 2410 8192
rect 2474 8128 2490 8192
rect 2554 8128 2563 8192
rect 2242 7104 2563 8128
rect 2242 7040 2250 7104
rect 2314 7040 2330 7104
rect 2394 7040 2410 7104
rect 2474 7040 2490 7104
rect 2554 7040 2563 7104
rect 2242 6016 2563 7040
rect 2242 5952 2250 6016
rect 2314 5952 2330 6016
rect 2394 5952 2410 6016
rect 2474 5952 2490 6016
rect 2554 5952 2563 6016
rect 2242 4928 2563 5952
rect 2242 4864 2250 4928
rect 2314 4864 2330 4928
rect 2394 4864 2410 4928
rect 2474 4864 2490 4928
rect 2554 4864 2563 4928
rect 2242 3840 2563 4864
rect 2242 3776 2250 3840
rect 2314 3776 2330 3840
rect 2394 3776 2410 3840
rect 2474 3776 2490 3840
rect 2554 3776 2563 3840
rect 2242 2752 2563 3776
rect 2242 2688 2250 2752
rect 2314 2688 2330 2752
rect 2394 2688 2410 2752
rect 2474 2688 2490 2752
rect 2554 2688 2563 2752
rect 2242 2128 2563 2688
rect 3541 27232 3861 27792
rect 3541 27168 3549 27232
rect 3613 27168 3629 27232
rect 3693 27168 3709 27232
rect 3773 27168 3789 27232
rect 3853 27168 3861 27232
rect 3541 26144 3861 27168
rect 3541 26080 3549 26144
rect 3613 26080 3629 26144
rect 3693 26080 3709 26144
rect 3773 26080 3789 26144
rect 3853 26080 3861 26144
rect 3541 25056 3861 26080
rect 3541 24992 3549 25056
rect 3613 24992 3629 25056
rect 3693 24992 3709 25056
rect 3773 24992 3789 25056
rect 3853 24992 3861 25056
rect 3541 23968 3861 24992
rect 3541 23904 3549 23968
rect 3613 23904 3629 23968
rect 3693 23904 3709 23968
rect 3773 23904 3789 23968
rect 3853 23904 3861 23968
rect 3541 22880 3861 23904
rect 3541 22816 3549 22880
rect 3613 22816 3629 22880
rect 3693 22816 3709 22880
rect 3773 22816 3789 22880
rect 3853 22816 3861 22880
rect 3541 21792 3861 22816
rect 3541 21728 3549 21792
rect 3613 21728 3629 21792
rect 3693 21728 3709 21792
rect 3773 21728 3789 21792
rect 3853 21728 3861 21792
rect 3541 20704 3861 21728
rect 3541 20640 3549 20704
rect 3613 20640 3629 20704
rect 3693 20640 3709 20704
rect 3773 20640 3789 20704
rect 3853 20640 3861 20704
rect 3541 19616 3861 20640
rect 3541 19552 3549 19616
rect 3613 19552 3629 19616
rect 3693 19552 3709 19616
rect 3773 19552 3789 19616
rect 3853 19552 3861 19616
rect 3541 18528 3861 19552
rect 3541 18464 3549 18528
rect 3613 18464 3629 18528
rect 3693 18464 3709 18528
rect 3773 18464 3789 18528
rect 3853 18464 3861 18528
rect 3541 17440 3861 18464
rect 3541 17376 3549 17440
rect 3613 17376 3629 17440
rect 3693 17376 3709 17440
rect 3773 17376 3789 17440
rect 3853 17376 3861 17440
rect 3541 16352 3861 17376
rect 3541 16288 3549 16352
rect 3613 16288 3629 16352
rect 3693 16288 3709 16352
rect 3773 16288 3789 16352
rect 3853 16288 3861 16352
rect 3541 15264 3861 16288
rect 3541 15200 3549 15264
rect 3613 15200 3629 15264
rect 3693 15200 3709 15264
rect 3773 15200 3789 15264
rect 3853 15200 3861 15264
rect 3541 14176 3861 15200
rect 3541 14112 3549 14176
rect 3613 14112 3629 14176
rect 3693 14112 3709 14176
rect 3773 14112 3789 14176
rect 3853 14112 3861 14176
rect 3541 13088 3861 14112
rect 3541 13024 3549 13088
rect 3613 13024 3629 13088
rect 3693 13024 3709 13088
rect 3773 13024 3789 13088
rect 3853 13024 3861 13088
rect 3541 12000 3861 13024
rect 3541 11936 3549 12000
rect 3613 11936 3629 12000
rect 3693 11936 3709 12000
rect 3773 11936 3789 12000
rect 3853 11936 3861 12000
rect 3541 10912 3861 11936
rect 3541 10848 3549 10912
rect 3613 10848 3629 10912
rect 3693 10848 3709 10912
rect 3773 10848 3789 10912
rect 3853 10848 3861 10912
rect 3541 9824 3861 10848
rect 3541 9760 3549 9824
rect 3613 9760 3629 9824
rect 3693 9760 3709 9824
rect 3773 9760 3789 9824
rect 3853 9760 3861 9824
rect 3541 8736 3861 9760
rect 3541 8672 3549 8736
rect 3613 8672 3629 8736
rect 3693 8672 3709 8736
rect 3773 8672 3789 8736
rect 3853 8672 3861 8736
rect 3541 7648 3861 8672
rect 3541 7584 3549 7648
rect 3613 7584 3629 7648
rect 3693 7584 3709 7648
rect 3773 7584 3789 7648
rect 3853 7584 3861 7648
rect 3541 6560 3861 7584
rect 3541 6496 3549 6560
rect 3613 6496 3629 6560
rect 3693 6496 3709 6560
rect 3773 6496 3789 6560
rect 3853 6496 3861 6560
rect 3541 5472 3861 6496
rect 3541 5408 3549 5472
rect 3613 5408 3629 5472
rect 3693 5408 3709 5472
rect 3773 5408 3789 5472
rect 3853 5408 3861 5472
rect 3541 4384 3861 5408
rect 3541 4320 3549 4384
rect 3613 4320 3629 4384
rect 3693 4320 3709 4384
rect 3773 4320 3789 4384
rect 3853 4320 3861 4384
rect 3541 3296 3861 4320
rect 3541 3232 3549 3296
rect 3613 3232 3629 3296
rect 3693 3232 3709 3296
rect 3773 3232 3789 3296
rect 3853 3232 3861 3296
rect 3541 2208 3861 3232
rect 3541 2144 3549 2208
rect 3613 2144 3629 2208
rect 3693 2144 3709 2208
rect 3773 2144 3789 2208
rect 3853 2144 3861 2208
rect 3541 2128 3861 2144
rect 4840 27776 5160 27792
rect 4840 27712 4848 27776
rect 4912 27712 4928 27776
rect 4992 27712 5008 27776
rect 5072 27712 5088 27776
rect 5152 27712 5160 27776
rect 4840 26688 5160 27712
rect 4840 26624 4848 26688
rect 4912 26624 4928 26688
rect 4992 26624 5008 26688
rect 5072 26624 5088 26688
rect 5152 26624 5160 26688
rect 4840 25600 5160 26624
rect 4840 25536 4848 25600
rect 4912 25536 4928 25600
rect 4992 25536 5008 25600
rect 5072 25536 5088 25600
rect 5152 25536 5160 25600
rect 4840 24512 5160 25536
rect 4840 24448 4848 24512
rect 4912 24448 4928 24512
rect 4992 24448 5008 24512
rect 5072 24448 5088 24512
rect 5152 24448 5160 24512
rect 4840 23424 5160 24448
rect 4840 23360 4848 23424
rect 4912 23360 4928 23424
rect 4992 23360 5008 23424
rect 5072 23360 5088 23424
rect 5152 23360 5160 23424
rect 4840 22336 5160 23360
rect 4840 22272 4848 22336
rect 4912 22272 4928 22336
rect 4992 22272 5008 22336
rect 5072 22272 5088 22336
rect 5152 22272 5160 22336
rect 4840 21248 5160 22272
rect 4840 21184 4848 21248
rect 4912 21184 4928 21248
rect 4992 21184 5008 21248
rect 5072 21184 5088 21248
rect 5152 21184 5160 21248
rect 4840 20160 5160 21184
rect 4840 20096 4848 20160
rect 4912 20096 4928 20160
rect 4992 20096 5008 20160
rect 5072 20096 5088 20160
rect 5152 20096 5160 20160
rect 4840 19072 5160 20096
rect 4840 19008 4848 19072
rect 4912 19008 4928 19072
rect 4992 19008 5008 19072
rect 5072 19008 5088 19072
rect 5152 19008 5160 19072
rect 4840 17984 5160 19008
rect 4840 17920 4848 17984
rect 4912 17920 4928 17984
rect 4992 17920 5008 17984
rect 5072 17920 5088 17984
rect 5152 17920 5160 17984
rect 4840 16896 5160 17920
rect 4840 16832 4848 16896
rect 4912 16832 4928 16896
rect 4992 16832 5008 16896
rect 5072 16832 5088 16896
rect 5152 16832 5160 16896
rect 4840 15808 5160 16832
rect 4840 15744 4848 15808
rect 4912 15744 4928 15808
rect 4992 15744 5008 15808
rect 5072 15744 5088 15808
rect 5152 15744 5160 15808
rect 4840 14720 5160 15744
rect 4840 14656 4848 14720
rect 4912 14656 4928 14720
rect 4992 14656 5008 14720
rect 5072 14656 5088 14720
rect 5152 14656 5160 14720
rect 4840 13632 5160 14656
rect 4840 13568 4848 13632
rect 4912 13568 4928 13632
rect 4992 13568 5008 13632
rect 5072 13568 5088 13632
rect 5152 13568 5160 13632
rect 4840 12544 5160 13568
rect 4840 12480 4848 12544
rect 4912 12480 4928 12544
rect 4992 12480 5008 12544
rect 5072 12480 5088 12544
rect 5152 12480 5160 12544
rect 4840 11456 5160 12480
rect 4840 11392 4848 11456
rect 4912 11392 4928 11456
rect 4992 11392 5008 11456
rect 5072 11392 5088 11456
rect 5152 11392 5160 11456
rect 4840 10368 5160 11392
rect 4840 10304 4848 10368
rect 4912 10304 4928 10368
rect 4992 10304 5008 10368
rect 5072 10304 5088 10368
rect 5152 10304 5160 10368
rect 4840 9280 5160 10304
rect 4840 9216 4848 9280
rect 4912 9216 4928 9280
rect 4992 9216 5008 9280
rect 5072 9216 5088 9280
rect 5152 9216 5160 9280
rect 4840 8192 5160 9216
rect 4840 8128 4848 8192
rect 4912 8128 4928 8192
rect 4992 8128 5008 8192
rect 5072 8128 5088 8192
rect 5152 8128 5160 8192
rect 4840 7104 5160 8128
rect 4840 7040 4848 7104
rect 4912 7040 4928 7104
rect 4992 7040 5008 7104
rect 5072 7040 5088 7104
rect 5152 7040 5160 7104
rect 4840 6016 5160 7040
rect 4840 5952 4848 6016
rect 4912 5952 4928 6016
rect 4992 5952 5008 6016
rect 5072 5952 5088 6016
rect 5152 5952 5160 6016
rect 4840 4928 5160 5952
rect 4840 4864 4848 4928
rect 4912 4864 4928 4928
rect 4992 4864 5008 4928
rect 5072 4864 5088 4928
rect 5152 4864 5160 4928
rect 4840 3840 5160 4864
rect 4840 3776 4848 3840
rect 4912 3776 4928 3840
rect 4992 3776 5008 3840
rect 5072 3776 5088 3840
rect 5152 3776 5160 3840
rect 4840 2752 5160 3776
rect 4840 2688 4848 2752
rect 4912 2688 4928 2752
rect 4992 2688 5008 2752
rect 5072 2688 5088 2752
rect 5152 2688 5160 2752
rect 4840 2128 5160 2688
rect 6138 27232 6458 27792
rect 6138 27168 6146 27232
rect 6210 27168 6226 27232
rect 6290 27168 6306 27232
rect 6370 27168 6386 27232
rect 6450 27168 6458 27232
rect 6138 26144 6458 27168
rect 6138 26080 6146 26144
rect 6210 26080 6226 26144
rect 6290 26080 6306 26144
rect 6370 26080 6386 26144
rect 6450 26080 6458 26144
rect 6138 25056 6458 26080
rect 6138 24992 6146 25056
rect 6210 24992 6226 25056
rect 6290 24992 6306 25056
rect 6370 24992 6386 25056
rect 6450 24992 6458 25056
rect 6138 23968 6458 24992
rect 6138 23904 6146 23968
rect 6210 23904 6226 23968
rect 6290 23904 6306 23968
rect 6370 23904 6386 23968
rect 6450 23904 6458 23968
rect 6138 22880 6458 23904
rect 6138 22816 6146 22880
rect 6210 22816 6226 22880
rect 6290 22816 6306 22880
rect 6370 22816 6386 22880
rect 6450 22816 6458 22880
rect 6138 21792 6458 22816
rect 6138 21728 6146 21792
rect 6210 21728 6226 21792
rect 6290 21728 6306 21792
rect 6370 21728 6386 21792
rect 6450 21728 6458 21792
rect 6138 20704 6458 21728
rect 6138 20640 6146 20704
rect 6210 20640 6226 20704
rect 6290 20640 6306 20704
rect 6370 20640 6386 20704
rect 6450 20640 6458 20704
rect 6138 19616 6458 20640
rect 6138 19552 6146 19616
rect 6210 19552 6226 19616
rect 6290 19552 6306 19616
rect 6370 19552 6386 19616
rect 6450 19552 6458 19616
rect 6138 18528 6458 19552
rect 6138 18464 6146 18528
rect 6210 18464 6226 18528
rect 6290 18464 6306 18528
rect 6370 18464 6386 18528
rect 6450 18464 6458 18528
rect 6138 17440 6458 18464
rect 6138 17376 6146 17440
rect 6210 17376 6226 17440
rect 6290 17376 6306 17440
rect 6370 17376 6386 17440
rect 6450 17376 6458 17440
rect 6138 16352 6458 17376
rect 6138 16288 6146 16352
rect 6210 16288 6226 16352
rect 6290 16288 6306 16352
rect 6370 16288 6386 16352
rect 6450 16288 6458 16352
rect 6138 15264 6458 16288
rect 6138 15200 6146 15264
rect 6210 15200 6226 15264
rect 6290 15200 6306 15264
rect 6370 15200 6386 15264
rect 6450 15200 6458 15264
rect 6138 14176 6458 15200
rect 6138 14112 6146 14176
rect 6210 14112 6226 14176
rect 6290 14112 6306 14176
rect 6370 14112 6386 14176
rect 6450 14112 6458 14176
rect 6138 13088 6458 14112
rect 6138 13024 6146 13088
rect 6210 13024 6226 13088
rect 6290 13024 6306 13088
rect 6370 13024 6386 13088
rect 6450 13024 6458 13088
rect 6138 12000 6458 13024
rect 6138 11936 6146 12000
rect 6210 11936 6226 12000
rect 6290 11936 6306 12000
rect 6370 11936 6386 12000
rect 6450 11936 6458 12000
rect 6138 10912 6458 11936
rect 6138 10848 6146 10912
rect 6210 10848 6226 10912
rect 6290 10848 6306 10912
rect 6370 10848 6386 10912
rect 6450 10848 6458 10912
rect 6138 9824 6458 10848
rect 6138 9760 6146 9824
rect 6210 9760 6226 9824
rect 6290 9760 6306 9824
rect 6370 9760 6386 9824
rect 6450 9760 6458 9824
rect 6138 8736 6458 9760
rect 6138 8672 6146 8736
rect 6210 8672 6226 8736
rect 6290 8672 6306 8736
rect 6370 8672 6386 8736
rect 6450 8672 6458 8736
rect 6138 7648 6458 8672
rect 6138 7584 6146 7648
rect 6210 7584 6226 7648
rect 6290 7584 6306 7648
rect 6370 7584 6386 7648
rect 6450 7584 6458 7648
rect 6138 6560 6458 7584
rect 6138 6496 6146 6560
rect 6210 6496 6226 6560
rect 6290 6496 6306 6560
rect 6370 6496 6386 6560
rect 6450 6496 6458 6560
rect 6138 5472 6458 6496
rect 6138 5408 6146 5472
rect 6210 5408 6226 5472
rect 6290 5408 6306 5472
rect 6370 5408 6386 5472
rect 6450 5408 6458 5472
rect 6138 4384 6458 5408
rect 6138 4320 6146 4384
rect 6210 4320 6226 4384
rect 6290 4320 6306 4384
rect 6370 4320 6386 4384
rect 6450 4320 6458 4384
rect 6138 3296 6458 4320
rect 6138 3232 6146 3296
rect 6210 3232 6226 3296
rect 6290 3232 6306 3296
rect 6370 3232 6386 3296
rect 6450 3232 6458 3296
rect 6138 2208 6458 3232
rect 6138 2144 6146 2208
rect 6210 2144 6226 2208
rect 6290 2144 6306 2208
rect 6370 2144 6386 2208
rect 6450 2144 6458 2208
rect 6138 2128 6458 2144
rect 7437 27776 7757 27792
rect 7437 27712 7445 27776
rect 7509 27712 7525 27776
rect 7589 27712 7605 27776
rect 7669 27712 7685 27776
rect 7749 27712 7757 27776
rect 7437 26688 7757 27712
rect 7437 26624 7445 26688
rect 7509 26624 7525 26688
rect 7589 26624 7605 26688
rect 7669 26624 7685 26688
rect 7749 26624 7757 26688
rect 7437 25600 7757 26624
rect 7437 25536 7445 25600
rect 7509 25536 7525 25600
rect 7589 25536 7605 25600
rect 7669 25536 7685 25600
rect 7749 25536 7757 25600
rect 7437 24512 7757 25536
rect 7437 24448 7445 24512
rect 7509 24448 7525 24512
rect 7589 24448 7605 24512
rect 7669 24448 7685 24512
rect 7749 24448 7757 24512
rect 7437 23424 7757 24448
rect 7437 23360 7445 23424
rect 7509 23360 7525 23424
rect 7589 23360 7605 23424
rect 7669 23360 7685 23424
rect 7749 23360 7757 23424
rect 7437 22336 7757 23360
rect 7437 22272 7445 22336
rect 7509 22272 7525 22336
rect 7589 22272 7605 22336
rect 7669 22272 7685 22336
rect 7749 22272 7757 22336
rect 7437 21248 7757 22272
rect 7437 21184 7445 21248
rect 7509 21184 7525 21248
rect 7589 21184 7605 21248
rect 7669 21184 7685 21248
rect 7749 21184 7757 21248
rect 7437 20160 7757 21184
rect 7437 20096 7445 20160
rect 7509 20096 7525 20160
rect 7589 20096 7605 20160
rect 7669 20096 7685 20160
rect 7749 20096 7757 20160
rect 7437 19072 7757 20096
rect 7437 19008 7445 19072
rect 7509 19008 7525 19072
rect 7589 19008 7605 19072
rect 7669 19008 7685 19072
rect 7749 19008 7757 19072
rect 7437 17984 7757 19008
rect 7437 17920 7445 17984
rect 7509 17920 7525 17984
rect 7589 17920 7605 17984
rect 7669 17920 7685 17984
rect 7749 17920 7757 17984
rect 7437 16896 7757 17920
rect 7437 16832 7445 16896
rect 7509 16832 7525 16896
rect 7589 16832 7605 16896
rect 7669 16832 7685 16896
rect 7749 16832 7757 16896
rect 7437 15808 7757 16832
rect 7437 15744 7445 15808
rect 7509 15744 7525 15808
rect 7589 15744 7605 15808
rect 7669 15744 7685 15808
rect 7749 15744 7757 15808
rect 7437 14720 7757 15744
rect 7437 14656 7445 14720
rect 7509 14656 7525 14720
rect 7589 14656 7605 14720
rect 7669 14656 7685 14720
rect 7749 14656 7757 14720
rect 7437 13632 7757 14656
rect 7437 13568 7445 13632
rect 7509 13568 7525 13632
rect 7589 13568 7605 13632
rect 7669 13568 7685 13632
rect 7749 13568 7757 13632
rect 7437 12544 7757 13568
rect 7437 12480 7445 12544
rect 7509 12480 7525 12544
rect 7589 12480 7605 12544
rect 7669 12480 7685 12544
rect 7749 12480 7757 12544
rect 7437 11456 7757 12480
rect 7437 11392 7445 11456
rect 7509 11392 7525 11456
rect 7589 11392 7605 11456
rect 7669 11392 7685 11456
rect 7749 11392 7757 11456
rect 7437 10368 7757 11392
rect 7437 10304 7445 10368
rect 7509 10304 7525 10368
rect 7589 10304 7605 10368
rect 7669 10304 7685 10368
rect 7749 10304 7757 10368
rect 7437 9280 7757 10304
rect 7437 9216 7445 9280
rect 7509 9216 7525 9280
rect 7589 9216 7605 9280
rect 7669 9216 7685 9280
rect 7749 9216 7757 9280
rect 7437 8192 7757 9216
rect 7437 8128 7445 8192
rect 7509 8128 7525 8192
rect 7589 8128 7605 8192
rect 7669 8128 7685 8192
rect 7749 8128 7757 8192
rect 7437 7104 7757 8128
rect 7437 7040 7445 7104
rect 7509 7040 7525 7104
rect 7589 7040 7605 7104
rect 7669 7040 7685 7104
rect 7749 7040 7757 7104
rect 7437 6016 7757 7040
rect 7437 5952 7445 6016
rect 7509 5952 7525 6016
rect 7589 5952 7605 6016
rect 7669 5952 7685 6016
rect 7749 5952 7757 6016
rect 7437 4928 7757 5952
rect 7437 4864 7445 4928
rect 7509 4864 7525 4928
rect 7589 4864 7605 4928
rect 7669 4864 7685 4928
rect 7749 4864 7757 4928
rect 7437 3840 7757 4864
rect 7437 3776 7445 3840
rect 7509 3776 7525 3840
rect 7589 3776 7605 3840
rect 7669 3776 7685 3840
rect 7749 3776 7757 3840
rect 7437 2752 7757 3776
rect 7437 2688 7445 2752
rect 7509 2688 7525 2752
rect 7589 2688 7605 2752
rect 7669 2688 7685 2752
rect 7749 2688 7757 2752
rect 7437 2128 7757 2688
use sky130_fd_sc_hd__clkbuf_2  ring.x6.x1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635107566
transform -1 0 2208 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_1  ring.x5.x3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635107566
transform -1 0 1932 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635107566
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1635107566
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_7 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635107566
transform 1 0 1748 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635107566
transform 1 0 1380 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9
timestamp 1635107566
transform 1 0 1932 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3
timestamp 1635107566
transform 1 0 1380 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ring.x38
timestamp 1635107566
transform 1 0 2944 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ring.x2.x5 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635107566
transform -1 0 2576 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_12
timestamp 1635107566
transform 1 0 2208 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16
timestamp 1635107566
transform 1 0 2576 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_2  ring.x27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635107566
transform 1 0 2576 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24
timestamp 1635107566
transform 1 0 3312 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_37
timestamp 1635107566
transform 1 0 4508 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635107566
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__mux4_2  ring.x30 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635107566
transform 1 0 3772 0 1 2176
box -38 -48 1694 592
use sky130_fd_sc_hd__clkbuf_8  ring.x35 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635107566
transform 1 0 4876 0 -1 3264
box -38 -48 1050 592
use sky130_fd_sc_hd__decap_4  FILLER_1_52
timestamp 1635107566
transform 1 0 5888 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635107566
transform 1 0 5428 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_2  ring.x6.x6 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635107566
transform -1 0 7176 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1635107566
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1635107566
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_59
timestamp 1635107566
transform 1 0 6532 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635107566
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55
timestamp 1635107566
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x2.x2_TE_B $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635107566
transform 1 0 6348 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__einvn_4  ring.x5.x2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635107566
transform -1 0 7912 0 -1 3264
box -38 -48 1050 592
use sky130_fd_sc_hd__decap_4  FILLER_0_66
timestamp 1635107566
transform 1 0 7176 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_77
timestamp 1635107566
transform 1 0 8188 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_74 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635107566
transform 1 0 7912 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_80
timestamp 1635107566
transform 1 0 8464 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1635107566
transform -1 0 8832 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1635107566
transform -1 0 8832 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ring.x5.x4
timestamp 1635107566
transform -1 0 8188 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1635107566
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_2  ring.x28
timestamp 1635107566
transform -1 0 3312 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_4  FILLER_2_24
timestamp 1635107566
transform 1 0 3312 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_29
timestamp 1635107566
transform 1 0 3772 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_33
timestamp 1635107566
transform 1 0 4140 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1635107566
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__einvn_8  ring.x2.x7 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635107566
transform -1 0 5888 0 1 3264
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_6  FILLER_2_52
timestamp 1635107566
transform 1 0 5888 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_58
timestamp 1635107566
transform 1 0 6440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__einvn_8  ring.x5.x7
timestamp 1635107566
transform -1 0 8188 0 1 3264
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_4  FILLER_2_77
timestamp 1635107566
transform 1 0 8188 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1635107566
transform -1 0 8832 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3
timestamp 1635107566
transform 1 0 1380 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_7
timestamp 1635107566
transform 1 0 1748 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1635107566
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  ring.x2.x3
timestamp 1635107566
transform -1 0 1748 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_2  ring.x29
timestamp 1635107566
transform 1 0 2116 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_4  FILLER_3_32
timestamp 1635107566
transform 1 0 4048 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__einvn_4  ring.x2.x2
timestamp 1635107566
transform -1 0 5428 0 -1 4352
box -38 -48 1050 592
use sky130_fd_sc_hd__decap_8  FILLER_3_47
timestamp 1635107566
transform 1 0 5428 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1635107566
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1635107566
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__einvn_8  ring.x4.x7
timestamp 1635107566
transform -1 0 8004 0 -1 4352
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_6  FILLER_3_75
timestamp 1635107566
transform 1 0 8004 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1635107566
transform -1 0 8832 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_16
timestamp 1635107566
transform 1 0 2576 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_3
timestamp 1635107566
transform 1 0 1380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_8
timestamp 1635107566
transform 1 0 1840 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1635107566
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ring.x3.x1
timestamp 1635107566
transform -1 0 3312 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_1  ring.x4.x3
timestamp 1635107566
transform -1 0 1840 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ring.x5.x1
timestamp 1635107566
transform -1 0 2576 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_24
timestamp 1635107566
transform 1 0 3312 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_36
timestamp 1635107566
transform 1 0 4416 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1635107566
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__einvp_2  ring.x2.x4
timestamp 1635107566
transform -1 0 5428 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ring.x2.x6
timestamp 1635107566
transform -1 0 4416 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_4_47
timestamp 1635107566
transform 1 0 5428 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_51
timestamp 1635107566
transform 1 0 5796 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_63
timestamp 1635107566
transform 1 0 6900 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__einvn_4  ring.x4.x2
timestamp 1635107566
transform -1 0 6900 0 1 4352
box -38 -48 1050 592
use sky130_fd_sc_hd__decap_6  FILLER_4_74
timestamp 1635107566
transform 1 0 7912 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_80
timestamp 1635107566
transform 1 0 8464 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1635107566
transform -1 0 8832 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ring.x4.x6
timestamp 1635107566
transform -1 0 7912 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1635107566
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_2  ring.x31
timestamp 1635107566
transform 1 0 1380 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_4  FILLER_5_24
timestamp 1635107566
transform 1 0 3312 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_2  ring.x32
timestamp 1635107566
transform 1 0 3680 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_6  FILLER_5_49
timestamp 1635107566
transform 1 0 5612 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1635107566
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_64
timestamp 1635107566
transform 1 0 6992 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1635107566
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__einvp_2  ring.x4.x4
timestamp 1635107566
transform -1 0 6992 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_5_75
timestamp 1635107566
transform 1 0 8004 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1635107566
transform -1 0 8832 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ring.x5.x6
timestamp 1635107566
transform -1 0 8004 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  ring.x6.x5
timestamp 1635107566
transform -1 0 1656 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  ring.x6.x3
timestamp 1635107566
transform -1 0 2300 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ring.x5.x5
timestamp 1635107566
transform -1 0 1932 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1635107566
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1635107566
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_6
timestamp 1635107566
transform 1 0 1656 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_9
timestamp 1635107566
transform 1 0 1932 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_6_3
timestamp 1635107566
transform 1 0 1380 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ring.x4.x5
timestamp 1635107566
transform -1 0 2576 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ring.x4.x1
timestamp 1635107566
transform -1 0 3312 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_13
timestamp 1635107566
transform 1 0 2300 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_16
timestamp 1635107566
transform 1 0 2576 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_2  ring.x33
timestamp 1635107566
transform -1 0 4600 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_4  FILLER_6_24
timestamp 1635107566
transform 1 0 3312 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_29
timestamp 1635107566
transform 1 0 3772 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_33
timestamp 1635107566
transform 1 0 4140 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_41
timestamp 1635107566
transform 1 0 4876 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_38
timestamp 1635107566
transform 1 0 4600 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1635107566
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__einvp_2  ring.x1.x4
timestamp 1635107566
transform -1 0 5612 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ring.x6.x4
timestamp 1635107566
transform -1 0 4876 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x1.x4_TE
timestamp 1635107566
transform 1 0 6624 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_56
timestamp 1635107566
transform 1 0 6256 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_62
timestamp 1635107566
transform 1 0 6808 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_49
timestamp 1635107566
transform 1 0 5612 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1635107566
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_57
timestamp 1635107566
transform 1 0 6348 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1635107566
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__einvn_4  ring.x3.x2
timestamp 1635107566
transform -1 0 6256 0 1 5440
box -38 -48 1050 592
use sky130_fd_sc_hd__einvn_8  ring.x6.x7
timestamp 1635107566
transform -1 0 8188 0 -1 6528
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_4  FILLER_6_77
timestamp 1635107566
transform 1 0 8188 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_77
timestamp 1635107566
transform 1 0 8188 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1635107566
transform -1 0 8832 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1635107566
transform -1 0 8832 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__einvn_4  ring.x6.x2
timestamp 1635107566
transform -1 0 8188 0 1 5440
box -38 -48 1050 592
use sky130_fd_sc_hd__decap_4  FILLER_8_13
timestamp 1635107566
transform 1 0 2300 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_6
timestamp 1635107566
transform 1 0 1656 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1635107566
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ring.x1.x5
timestamp 1635107566
transform -1 0 2300 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  ring.x3.x3
timestamp 1635107566
transform -1 0 1656 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ring.x3.x6
timestamp 1635107566
transform 1 0 2668 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_8_24
timestamp 1635107566
transform 1 0 3312 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_29
timestamp 1635107566
transform 1 0 3772 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1635107566
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__einvn_8  ring.x1.x7
timestamp 1635107566
transform -1 0 5612 0 1 6528
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_4  FILLER_8_49
timestamp 1635107566
transform 1 0 5612 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__einvn_8  ring.x3.x7
timestamp 1635107566
transform -1 0 7636 0 1 6528
box -38 -48 1694 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x1.x7_TE_B
timestamp 1635107566
transform -1 0 8188 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_71
timestamp 1635107566
transform 1 0 7636 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_77
timestamp 1635107566
transform 1 0 8188 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1635107566
transform -1 0 8832 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_11
timestamp 1635107566
transform 1 0 2116 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_19
timestamp 1635107566
transform 1 0 2852 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_3
timestamp 1635107566
transform 1 0 1380 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_7
timestamp 1635107566
transform 1 0 1748 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1635107566
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ring.x7.x1
timestamp 1635107566
transform -1 0 2852 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_1  ring.x7.x3
timestamp 1635107566
transform -1 0 2116 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_30
timestamp 1635107566
transform 1 0 3864 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__einvn_4  ring.x1.x2
timestamp 1635107566
transform -1 0 5244 0 -1 7616
box -38 -48 1050 592
use sky130_fd_sc_hd__einvp_2  ring.x7.x6
timestamp 1635107566
transform -1 0 3864 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_9_45
timestamp 1635107566
transform 1 0 5244 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_52
timestamp 1635107566
transform 1 0 5888 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1635107566
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_1  ring.x1.x3
timestamp 1635107566
transform 1 0 5612 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__einvn_8  ring.x7.x7
timestamp 1635107566
transform -1 0 8004 0 -1 7616
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_6  FILLER_9_75
timestamp 1635107566
transform 1 0 8004 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1635107566
transform -1 0 8832 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x2.x4_TE
timestamp 1635107566
transform -1 0 2024 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_10
timestamp 1635107566
transform 1 0 2024 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_17
timestamp 1635107566
transform 1 0 2668 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_3
timestamp 1635107566
transform 1 0 1380 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_7
timestamp 1635107566
transform 1 0 1748 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1635107566
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ring.x3.x5
timestamp 1635107566
transform -1 0 3312 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ring.x7.x5
timestamp 1635107566
transform -1 0 2668 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x1.x2_TE_B
timestamp 1635107566
transform 1 0 3772 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_24
timestamp 1635107566
transform 1 0 3312 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_31
timestamp 1635107566
transform 1 0 3956 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_42
timestamp 1635107566
transform 1 0 4968 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1635107566
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__einvp_2  ring.x1.x6
timestamp 1635107566
transform -1 0 4968 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_10_48
timestamp 1635107566
transform 1 0 5520 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_56
timestamp 1635107566
transform 1 0 6256 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_60
timestamp 1635107566
transform 1 0 6624 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__einvp_2  ring.x3.x4
timestamp 1635107566
transform -1 0 6256 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_4  ring.x7.x2
timestamp 1635107566
transform -1 0 7728 0 1 7616
box -38 -48 1050 592
use sky130_fd_sc_hd__decap_8  FILLER_10_72
timestamp 1635107566
transform 1 0 7728 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_80
timestamp 1635107566
transform 1 0 8464 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1635107566
transform -1 0 8832 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x1.x6_TE
timestamp 1635107566
transform -1 0 2668 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x2.x6_TE
timestamp 1635107566
transform -1 0 2116 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x3.x4_TE
timestamp 1635107566
transform -1 0 1564 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_11
timestamp 1635107566
transform 1 0 2116 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_17
timestamp 1635107566
transform 1 0 2668 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_5
timestamp 1635107566
transform 1 0 1564 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1635107566
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ring.x8.x1
timestamp 1635107566
transform -1 0 3404 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_25
timestamp 1635107566
transform 1 0 3404 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_40
timestamp 1635107566
transform 1 0 4784 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_8  ring.x26
timestamp 1635107566
transform 1 0 3772 0 -1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__fill_1  FILLER_11_44
timestamp 1635107566
transform 1 0 5152 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_52
timestamp 1635107566
transform 1 0 5888 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_61
timestamp 1635107566
transform 1 0 6716 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_65
timestamp 1635107566
transform 1 0 7084 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1635107566
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  ring.x2.x1
timestamp 1635107566
transform -1 0 6716 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_2  ring.x7.x4
timestamp 1635107566
transform -1 0 5888 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_11_77
timestamp 1635107566
transform 1 0 8188 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1635107566
transform -1 0 8832 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__einvn_4  ring.x9.x2
timestamp 1635107566
transform -1 0 8188 0 -1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x2.x7_TE_B
timestamp 1635107566
transform -1 0 2668 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x3.x2_TE_B
timestamp 1635107566
transform -1 0 2116 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x3.x7_TE_B
timestamp 1635107566
transform -1 0 1564 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_11
timestamp 1635107566
transform 1 0 2116 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_17
timestamp 1635107566
transform 1 0 2668 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_5
timestamp 1635107566
transform 1 0 1564 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1635107566
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ring.x8.x5
timestamp 1635107566
transform -1 0 3312 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_24
timestamp 1635107566
transform 1 0 3312 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_12_29
timestamp 1635107566
transform 1 0 3772 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_36
timestamp 1635107566
transform 1 0 4416 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1635107566
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  ring.x1.x1
timestamp 1635107566
transform -1 0 5152 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  ring.x36
timestamp 1635107566
transform -1 0 4416 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_44
timestamp 1635107566
transform 1 0 5152 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_55
timestamp 1635107566
transform 1 0 6164 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_2  ring.x8.x6
timestamp 1635107566
transform -1 0 6164 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ring.x9.x7
timestamp 1635107566
transform 1 0 6532 0 1 8704
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_4  FILLER_12_77
timestamp 1635107566
transform 1 0 8188 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1635107566
transform -1 0 8832 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1635107566
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1635107566
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_3
timestamp 1635107566
transform 1 0 1380 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x4.x2_TE_B
timestamp 1635107566
transform -1 0 1564 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_5
timestamp 1635107566
transform 1 0 1564 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_7
timestamp 1635107566
transform 1 0 1748 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x38_A
timestamp 1635107566
transform -1 0 2116 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x30_S0
timestamp 1635107566
transform -1 0 2024 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  ring.x9.x5
timestamp 1635107566
transform -1 0 2668 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_11
timestamp 1635107566
transform 1 0 2116 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_10
timestamp 1635107566
transform 1 0 2024 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_17
timestamp 1635107566
transform 1 0 2668 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_17
timestamp 1635107566
transform 1 0 2668 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x30_S1
timestamp 1635107566
transform -1 0 2668 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__clkinv_1  ring.x9.x3
timestamp 1635107566
transform -1 0 3312 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ring.x9.x1
timestamp 1635107566
transform -1 0 3404 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  ring.x37
timestamp 1635107566
transform 1 0 3956 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  ring.x34 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635107566
transform 1 0 3772 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1635107566
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_29
timestamp 1635107566
transform 1 0 3772 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_24
timestamp 1635107566
transform 1 0 3312 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_25
timestamp 1635107566
transform 1 0 3404 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_4  ring.x47 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635107566
transform -1 0 5520 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_14_35
timestamp 1635107566
transform 1 0 4324 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_38
timestamp 1635107566
transform 1 0 4600 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_4  ring.x21
timestamp 1635107566
transform -1 0 5796 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1635107566
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1635107566
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_48
timestamp 1635107566
transform 1 0 5520 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_63
timestamp 1635107566
transform 1 0 6900 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1635107566
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__einvn_4  ring.x8.x2
timestamp 1635107566
transform -1 0 6900 0 1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__einvn_8  ring.x8.x7
timestamp 1635107566
transform -1 0 8004 0 -1 9792
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_6  FILLER_13_75
timestamp 1635107566
transform 1 0 8004 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_14_74
timestamp 1635107566
transform 1 0 7912 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_80
timestamp 1635107566
transform 1 0 8464 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1635107566
transform -1 0 8832 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1635107566
transform -1 0 8832 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ring.x8.x4
timestamp 1635107566
transform -1 0 7912 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x34_S
timestamp 1635107566
transform -1 0 2944 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x39.x6_TE
timestamp 1635107566
transform -1 0 2392 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x4.x4_TE
timestamp 1635107566
transform -1 0 1840 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_14
timestamp 1635107566
transform 1 0 2392 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_20
timestamp 1635107566
transform 1 0 2944 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_15_3
timestamp 1635107566
transform 1 0 1380 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_8
timestamp 1635107566
transform 1 0 1840 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1635107566
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x3.x6_TE
timestamp 1635107566
transform -1 0 3496 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_26
timestamp 1635107566
transform 1 0 3496 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_33
timestamp 1635107566
transform 1 0 4140 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_41
timestamp 1635107566
transform 1 0 4876 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  ring.x13.x1
timestamp 1635107566
transform -1 0 4876 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_1  ring.x8.x3
timestamp 1635107566
transform -1 0 4140 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_52
timestamp 1635107566
transform 1 0 5888 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_64
timestamp 1635107566
transform 1 0 6992 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1635107566
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__einvp_2  ring.x39.x6
timestamp 1635107566
transform -1 0 6992 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ring.x9.x6
timestamp 1635107566
transform -1 0 5888 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_15_77
timestamp 1635107566
transform 1 0 8188 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1635107566
transform -1 0 8832 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ring.x9.x4
timestamp 1635107566
transform -1 0 8188 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x39.x4_TE
timestamp 1635107566
transform 1 0 2576 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x4.x6_TE
timestamp 1635107566
transform -1 0 2208 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x40.x4_TE
timestamp 1635107566
transform -1 0 1656 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_12
timestamp 1635107566
transform 1 0 2208 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_18
timestamp 1635107566
transform 1 0 2760 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_3
timestamp 1635107566
transform 1 0 1380 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_6
timestamp 1635107566
transform 1 0 1656 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1635107566
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x11.x2_TE_B
timestamp 1635107566
transform -1 0 3956 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x11.x4_TE
timestamp 1635107566
transform 1 0 3128 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_24
timestamp 1635107566
transform 1 0 3312 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_31
timestamp 1635107566
transform 1 0 3956 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_42
timestamp 1635107566
transform 1 0 4968 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1635107566
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__einvp_2  ring.x40.x4
timestamp 1635107566
transform -1 0 4968 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_16_46
timestamp 1635107566
transform 1 0 5336 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_54
timestamp 1635107566
transform 1 0 6072 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_2  ring.x11.x4
timestamp 1635107566
transform -1 0 7452 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ring.x39.x4
timestamp 1635107566
transform -1 0 6072 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_16_69
timestamp 1635107566
transform 1 0 7452 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_77
timestamp 1635107566
transform 1 0 8188 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1635107566
transform -1 0 8832 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ring.x10.x1
timestamp 1635107566
transform -1 0 8188 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x11.x7_TE_B
timestamp 1635107566
transform -1 0 2852 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x4.x7_TE_B
timestamp 1635107566
transform -1 0 2300 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x40.x7_TE_B
timestamp 1635107566
transform 1 0 1564 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_13
timestamp 1635107566
transform 1 0 2300 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_19
timestamp 1635107566
transform 1 0 2852 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_3
timestamp 1635107566
transform 1 0 1380 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_7
timestamp 1635107566
transform 1 0 1748 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1635107566
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_26
timestamp 1635107566
transform 1 0 3496 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_1  ring.x39.x3
timestamp 1635107566
transform -1 0 3496 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__einvn_8  ring.x40.x7
timestamp 1635107566
transform -1 0 5520 0 -1 11968
box -38 -48 1694 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x10.x2_TE_B
timestamp 1635107566
transform 1 0 6348 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_48
timestamp 1635107566
transform 1 0 5520 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_59
timestamp 1635107566
transform 1 0 6532 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1635107566
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__einvn_4  ring.x11.x2
timestamp 1635107566
transform -1 0 7912 0 -1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__decap_6  FILLER_17_74
timestamp 1635107566
transform 1 0 7912 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_80
timestamp 1635107566
transform 1 0 8464 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1635107566
transform -1 0 8832 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x39.x7_TE_B
timestamp 1635107566
transform -1 0 2024 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_10
timestamp 1635107566
transform 1 0 2024 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_17
timestamp 1635107566
transform 1 0 2668 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_3
timestamp 1635107566
transform 1 0 1380 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_7
timestamp 1635107566
transform 1 0 1748 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1635107566
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ring.x11.x5
timestamp 1635107566
transform -1 0 3312 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ring.x39.x5
timestamp 1635107566
transform -1 0 2668 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_24
timestamp 1635107566
transform 1 0 3312 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_32
timestamp 1635107566
transform 1 0 4048 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1635107566
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_1  ring.x11.x3
timestamp 1635107566
transform -1 0 4048 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__einvn_8  ring.x39.x7
timestamp 1635107566
transform -1 0 6072 0 1 11968
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_4  FILLER_18_54
timestamp 1635107566
transform 1 0 6072 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__einvn_8  ring.x11.x7
timestamp 1635107566
transform -1 0 8096 0 1 11968
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_4  FILLER_18_76
timestamp 1635107566
transform 1 0 8096 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_80
timestamp 1635107566
transform 1 0 8464 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1635107566
transform -1 0 8832 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1635107566
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1635107566
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_3
timestamp 1635107566
transform 1 0 1380 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_3
timestamp 1635107566
transform 1 0 1380 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x5.x4_TE
timestamp 1635107566
transform -1 0 1656 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_6
timestamp 1635107566
transform 1 0 1656 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_8
timestamp 1635107566
transform 1 0 1840 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x40.x2_TE_B
timestamp 1635107566
transform -1 0 1840 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  ring.x40.x5
timestamp 1635107566
transform -1 0 2484 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_12
timestamp 1635107566
transform 1 0 2208 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x40.x6_TE
timestamp 1635107566
transform 1 0 2024 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__clkinv_1  ring.x40.x3
timestamp 1635107566
transform -1 0 3128 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_18
timestamp 1635107566
transform 1 0 2760 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_15
timestamp 1635107566
transform 1 0 2484 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x11.x6_TE
timestamp 1635107566
transform -1 0 2760 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  ring.x40.x1
timestamp 1635107566
transform -1 0 3864 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ring.x10.x5
timestamp 1635107566
transform -1 0 4048 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1635107566
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_32
timestamp 1635107566
transform 1 0 4048 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_24
timestamp 1635107566
transform 1 0 3312 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_30
timestamp 1635107566
transform 1 0 3864 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_22
timestamp 1635107566
transform 1 0 3128 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x10.x6_TE
timestamp 1635107566
transform -1 0 3312 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_2  ring.x40.x6
timestamp 1635107566
transform -1 0 5060 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_20_43
timestamp 1635107566
transform 1 0 5060 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__einvn_4  ring.x40.x2
timestamp 1635107566
transform -1 0 5244 0 -1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__decap_4  FILLER_19_45
timestamp 1635107566
transform 1 0 5244 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_52
timestamp 1635107566
transform 1 0 5888 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_57
timestamp 1635107566
transform 1 0 6348 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_58
timestamp 1635107566
transform 1 0 6440 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1635107566
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_1  ring.x10.x3
timestamp 1635107566
transform -1 0 5888 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ring.x11.x6
timestamp 1635107566
transform -1 0 7176 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_4  ring.x39.x2
timestamp 1635107566
transform -1 0 6440 0 1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__decap_4  FILLER_19_66
timestamp 1635107566
transform 1 0 7176 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_77
timestamp 1635107566
transform 1 0 8188 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_77
timestamp 1635107566
transform 1 0 8188 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1635107566
transform -1 0 8832 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1635107566
transform -1 0 8832 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__einvn_4  ring.x10.x2
timestamp 1635107566
transform -1 0 8188 0 1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__einvp_2  ring.x10.x6
timestamp 1635107566
transform -1 0 8188 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x39.x2_TE_B
timestamp 1635107566
transform -1 0 3220 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x5.x2_TE_B
timestamp 1635107566
transform -1 0 2668 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x5.x7_TE_B
timestamp 1635107566
transform -1 0 2116 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x6.x4_TE
timestamp 1635107566
transform -1 0 1564 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_11
timestamp 1635107566
transform 1 0 2116 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_17
timestamp 1635107566
transform 1 0 2668 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_5
timestamp 1635107566
transform 1 0 1564 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1635107566
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x10.x7_TE_B
timestamp 1635107566
transform -1 0 3772 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_23
timestamp 1635107566
transform 1 0 3220 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_29
timestamp 1635107566
transform 1 0 3772 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_36
timestamp 1635107566
transform 1 0 4416 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  ring.x12.x1
timestamp 1635107566
transform -1 0 5152 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_1  ring.x12.x3
timestamp 1635107566
transform -1 0 4416 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_44
timestamp 1635107566
transform 1 0 5152 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_52
timestamp 1635107566
transform 1 0 5888 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_57
timestamp 1635107566
transform 1 0 6348 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1635107566
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__einvn_8  ring.x10.x7
timestamp 1635107566
transform -1 0 8188 0 -1 14144
box -38 -48 1694 592
use sky130_fd_sc_hd__clkbuf_2  ring.x11.x1
timestamp 1635107566
transform -1 0 5888 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_77
timestamp 1635107566
transform 1 0 8188 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1635107566
transform -1 0 8832 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x5.x6_TE
timestamp 1635107566
transform -1 0 2760 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x6.x2_TE_B
timestamp 1635107566
transform -1 0 2208 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x6.x7_TE_B
timestamp 1635107566
transform -1 0 1656 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_12
timestamp 1635107566
transform 1 0 2208 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_18
timestamp 1635107566
transform 1 0 2760 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_3
timestamp 1635107566
transform 1 0 1380 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_6
timestamp 1635107566
transform 1 0 1656 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1635107566
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x10.x4_TE
timestamp 1635107566
transform -1 0 3956 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x12.x2_TE_B
timestamp 1635107566
transform -1 0 3312 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_24
timestamp 1635107566
transform 1 0 3312 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_31
timestamp 1635107566
transform 1 0 3956 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_39
timestamp 1635107566
transform 1 0 4692 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1635107566
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__einvp_2  ring.x12.x6
timestamp 1635107566
transform -1 0 5704 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  ring.x39.x1
timestamp 1635107566
transform -1 0 4692 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_50
timestamp 1635107566
transform 1 0 5704 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_65
timestamp 1635107566
transform 1 0 7084 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__einvn_4  ring.x12.x2
timestamp 1635107566
transform -1 0 7084 0 1 14144
box -38 -48 1050 592
use sky130_fd_sc_hd__fill_1  FILLER_22_69
timestamp 1635107566
transform 1 0 7452 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_77
timestamp 1635107566
transform 1 0 8188 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1635107566
transform -1 0 8832 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ring.x10.x4
timestamp 1635107566
transform -1 0 8188 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x12.x7_TE_B
timestamp 1635107566
transform -1 0 3128 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x6.x6_TE
timestamp 1635107566
transform -1 0 2576 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x7.x2_TE_B
timestamp 1635107566
transform 1 0 1840 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_10
timestamp 1635107566
transform 1 0 2024 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_16
timestamp 1635107566
transform 1 0 2576 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_3
timestamp 1635107566
transform 1 0 1380 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_7
timestamp 1635107566
transform 1 0 1748 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1635107566
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x12.x6_TE
timestamp 1635107566
transform -1 0 3680 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_22
timestamp 1635107566
transform 1 0 3128 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_28
timestamp 1635107566
transform 1 0 3680 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_35
timestamp 1635107566
transform 1 0 4324 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ring.x12.x5
timestamp 1635107566
transform -1 0 4324 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__einvn_4  ring.x13.x2
timestamp 1635107566
transform -1 0 5704 0 -1 15232
box -38 -48 1050 592
use sky130_fd_sc_hd__decap_6  FILLER_23_50
timestamp 1635107566
transform 1 0 5704 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1635107566
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__einvn_8  ring.x12.x7
timestamp 1635107566
transform -1 0 8004 0 -1 15232
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_6  FILLER_23_75
timestamp 1635107566
transform 1 0 8004 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1635107566
transform -1 0 8832 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x13.x7_TE_B
timestamp 1635107566
transform -1 0 2760 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x7.x4_TE
timestamp 1635107566
transform 1 0 2024 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x7.x6_TE
timestamp 1635107566
transform -1 0 1656 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_12
timestamp 1635107566
transform 1 0 2208 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_18
timestamp 1635107566
transform 1 0 2760 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_3
timestamp 1635107566
transform 1 0 1380 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_6
timestamp 1635107566
transform 1 0 1656 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1635107566
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x12.x4_TE
timestamp 1635107566
transform -1 0 3956 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x13.x2_TE_B
timestamp 1635107566
transform -1 0 3312 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_24
timestamp 1635107566
transform 1 0 3312 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_31
timestamp 1635107566
transform 1 0 3956 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1635107566
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__einvn_8  ring.x13.x7
timestamp 1635107566
transform -1 0 5980 0 1 15232
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_4  FILLER_24_53
timestamp 1635107566
transform 1 0 5980 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_64
timestamp 1635107566
transform 1 0 6992 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_2  ring.x12.x4
timestamp 1635107566
transform -1 0 6992 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_24_75
timestamp 1635107566
transform 1 0 8004 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1635107566
transform -1 0 8832 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ring.x17.x4
timestamp 1635107566
transform -1 0 8004 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x17.x4_TE
timestamp 1635107566
transform 1 0 2576 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x18.x2_TE_B
timestamp 1635107566
transform -1 0 2208 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x7.x7_TE_B
timestamp 1635107566
transform -1 0 1656 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_12
timestamp 1635107566
transform 1 0 2208 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_18
timestamp 1635107566
transform 1 0 2760 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_3
timestamp 1635107566
transform 1 0 1380 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_6
timestamp 1635107566
transform 1 0 1656 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1635107566
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x13.x4_TE
timestamp 1635107566
transform 1 0 3128 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_24
timestamp 1635107566
transform 1 0 3312 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_31
timestamp 1635107566
transform 1 0 3956 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_38
timestamp 1635107566
transform 1 0 4600 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_1  ring.x13.x3
timestamp 1635107566
transform -1 0 4600 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ring.x13.x4
timestamp 1635107566
transform -1 0 5612 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  ring.x13.x5
timestamp 1635107566
transform -1 0 3956 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_25_49
timestamp 1635107566
transform 1 0 5612 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1635107566
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_61
timestamp 1635107566
transform 1 0 6716 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_65
timestamp 1635107566
transform 1 0 7084 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1635107566
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  ring.x14.x1
timestamp 1635107566
transform -1 0 6716 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_77
timestamp 1635107566
transform 1 0 8188 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1635107566
transform -1 0 8832 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__einvn_4  ring.x18.x2
timestamp 1635107566
transform -1 0 8188 0 -1 16320
box -38 -48 1050 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1635107566
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1635107566
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_3
timestamp 1635107566
transform 1 0 1380 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x8.x2_TE_B
timestamp 1635107566
transform -1 0 1564 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_7
timestamp 1635107566
transform 1 0 1748 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_5
timestamp 1635107566
transform 1 0 1564 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x8.x4_TE
timestamp 1635107566
transform 1 0 1564 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x17.x7_TE_B
timestamp 1635107566
transform -1 0 2116 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_13
timestamp 1635107566
transform 1 0 2300 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_11
timestamp 1635107566
transform 1 0 2116 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x17.x2_TE_B
timestamp 1635107566
transform -1 0 2300 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__clkinv_1  ring.x18.x3
timestamp 1635107566
transform -1 0 2944 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_17
timestamp 1635107566
transform 1 0 2668 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x17.x6_TE
timestamp 1635107566
transform -1 0 2668 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  ring.x18.x5
timestamp 1635107566
transform -1 0 3312 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_20
timestamp 1635107566
transform 1 0 2944 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ring.x17.x5
timestamp 1635107566
transform -1 0 3588 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1635107566
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_27
timestamp 1635107566
transform 1 0 3588 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_29
timestamp 1635107566
transform 1 0 3772 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_24
timestamp 1635107566
transform 1 0 3312 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_1  ring.x17.x3
timestamp 1635107566
transform -1 0 4508 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ring.x15.x5
timestamp 1635107566
transform -1 0 4232 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_34
timestamp 1635107566
transform 1 0 4232 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_37
timestamp 1635107566
transform 1 0 4508 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_33
timestamp 1635107566
transform 1 0 4140 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  ring.x14.x5
timestamp 1635107566
transform -1 0 4876 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ring.x13.x6
timestamp 1635107566
transform -1 0 5520 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_27_41
timestamp 1635107566
transform 1 0 4876 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_48
timestamp 1635107566
transform 1 0 5520 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_54
timestamp 1635107566
transform 1 0 6072 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_52
timestamp 1635107566
transform 1 0 5888 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1635107566
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__einvn_4  ring.x17.x2
timestamp 1635107566
transform -1 0 7360 0 -1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__einvp_2  ring.x17.x6
timestamp 1635107566
transform -1 0 5888 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ring.x17.x7
timestamp 1635107566
transform 1 0 6164 0 1 16320
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_8  FILLER_26_73
timestamp 1635107566
transform 1 0 7820 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_68
timestamp 1635107566
transform 1 0 7360 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_76
timestamp 1635107566
transform 1 0 8096 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_80
timestamp 1635107566
transform 1 0 8464 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1635107566
transform -1 0 8832 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1635107566
transform -1 0 8832 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ring.x18.x1
timestamp 1635107566
transform -1 0 8096 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x15.x2_TE_B
timestamp 1635107566
transform 1 0 2576 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x18.x7_TE_B
timestamp 1635107566
transform 1 0 2024 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x8.x6_TE
timestamp 1635107566
transform -1 0 1656 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_12
timestamp 1635107566
transform 1 0 2208 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_18
timestamp 1635107566
transform 1 0 2760 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_3
timestamp 1635107566
transform 1 0 1380 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_6
timestamp 1635107566
transform 1 0 1656 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1635107566
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x14.x6_TE
timestamp 1635107566
transform -1 0 3312 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_24
timestamp 1635107566
transform 1 0 3312 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_29
timestamp 1635107566
transform 1 0 3772 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_40
timestamp 1635107566
transform 1 0 4784 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1635107566
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__einvp_2  ring.x14.x6
timestamp 1635107566
transform 1 0 4140 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_28_55
timestamp 1635107566
transform 1 0 6164 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__einvn_4  ring.x15.x2
timestamp 1635107566
transform -1 0 6164 0 1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__einvn_8  ring.x18.x7
timestamp 1635107566
transform -1 0 8188 0 1 17408
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_4  FILLER_28_77
timestamp 1635107566
transform 1 0 8188 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1635107566
transform -1 0 8832 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x15.x6_TE
timestamp 1635107566
transform -1 0 2668 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x18.x4_TE
timestamp 1635107566
transform -1 0 2116 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x8.x7_TE_B
timestamp 1635107566
transform -1 0 1564 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_11
timestamp 1635107566
transform 1 0 2116 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_17
timestamp 1635107566
transform 1 0 2668 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_5
timestamp 1635107566
transform 1 0 1564 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1635107566
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  ring.x15.x3
timestamp 1635107566
transform -1 0 3312 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_24
timestamp 1635107566
transform 1 0 3312 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_31
timestamp 1635107566
transform 1 0 3956 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__einvn_4  ring.x14.x2
timestamp 1635107566
transform -1 0 5336 0 -1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ring.x14.x3
timestamp 1635107566
transform -1 0 3956 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x13.x6_TE
timestamp 1635107566
transform -1 0 5888 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_46
timestamp 1635107566
transform 1 0 5336 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_52
timestamp 1635107566
transform 1 0 5888 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_64
timestamp 1635107566
transform 1 0 6992 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1635107566
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__einvp_2  ring.x15.x6
timestamp 1635107566
transform -1 0 6992 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_29_77
timestamp 1635107566
transform 1 0 8188 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1635107566
transform -1 0 8832 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ring.x18.x4
timestamp 1635107566
transform -1 0 8188 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x16.x4_TE
timestamp 1635107566
transform 1 0 2576 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x18.x6_TE
timestamp 1635107566
transform -1 0 2208 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x9.x2_TE_B
timestamp 1635107566
transform -1 0 1656 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_12
timestamp 1635107566
transform 1 0 2208 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_18
timestamp 1635107566
transform 1 0 2760 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_3
timestamp 1635107566
transform 1 0 1380 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_6
timestamp 1635107566
transform 1 0 1656 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1635107566
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x14.x7_TE_B
timestamp 1635107566
transform -1 0 3312 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_24
timestamp 1635107566
transform 1 0 3312 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_29
timestamp 1635107566
transform 1 0 3772 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1635107566
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__einvn_8  ring.x14.x7
timestamp 1635107566
transform -1 0 5796 0 1 18496
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_6  FILLER_30_51
timestamp 1635107566
transform 1 0 5796 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_57
timestamp 1635107566
transform 1 0 6348 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_65
timestamp 1635107566
transform 1 0 7084 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_2  ring.x16.x4
timestamp 1635107566
transform -1 0 7084 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_30_69
timestamp 1635107566
transform 1 0 7452 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_77
timestamp 1635107566
transform 1 0 8188 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1635107566
transform -1 0 8832 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ring.x18.x6
timestamp 1635107566
transform -1 0 8188 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x15.x4_TE
timestamp 1635107566
transform -1 0 3036 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x19.x4_TE
timestamp 1635107566
transform -1 0 2484 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x9.x4_TE
timestamp 1635107566
transform 1 0 1748 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_15
timestamp 1635107566
transform 1 0 2484 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_21
timestamp 1635107566
transform 1 0 3036 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_3
timestamp 1635107566
transform 1 0 1380 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_9
timestamp 1635107566
transform 1 0 1932 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1635107566
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x14.x4_TE
timestamp 1635107566
transform 1 0 3404 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_27
timestamp 1635107566
transform 1 0 3588 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_35
timestamp 1635107566
transform 1 0 4324 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_2  ring.x14.x4
timestamp 1635107566
transform -1 0 5336 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  ring.x15.x1
timestamp 1635107566
transform -1 0 4324 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x14.x2_TE_B
timestamp 1635107566
transform -1 0 5888 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_46
timestamp 1635107566
transform 1 0 5336 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_52
timestamp 1635107566
transform 1 0 5888 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_64
timestamp 1635107566
transform 1 0 6992 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1635107566
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__einvp_2  ring.x15.x4
timestamp 1635107566
transform -1 0 6992 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_31_77
timestamp 1635107566
transform 1 0 8188 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1635107566
transform -1 0 8832 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ring.x19.x4
timestamp 1635107566
transform -1 0 8188 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x19.x2_TE_B
timestamp 1635107566
transform -1 0 2760 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x9.x6_TE
timestamp 1635107566
transform -1 0 2208 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x9.x7_TE_B
timestamp 1635107566
transform -1 0 1656 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_12
timestamp 1635107566
transform 1 0 2208 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_18
timestamp 1635107566
transform 1 0 2760 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_3
timestamp 1635107566
transform 1 0 1380 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_6
timestamp 1635107566
transform 1 0 1656 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1635107566
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x15.x7_TE_B
timestamp 1635107566
transform -1 0 3312 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_24
timestamp 1635107566
transform 1 0 3312 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_29
timestamp 1635107566
transform 1 0 3772 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_37
timestamp 1635107566
transform 1 0 4508 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1635107566
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__einvn_8  ring.x15.x7
timestamp 1635107566
transform 1 0 4876 0 1 19584
box -38 -48 1694 592
use sky130_fd_sc_hd__clkbuf_2  ring.x17.x1
timestamp 1635107566
transform -1 0 4508 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_59
timestamp 1635107566
transform 1 0 6532 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_65
timestamp 1635107566
transform 1 0 7084 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_77
timestamp 1635107566
transform 1 0 8188 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1635107566
transform -1 0 8832 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__einvn_4  ring.x19.x2
timestamp 1635107566
transform -1 0 8188 0 1 19584
box -38 -48 1050 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1635107566
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1635107566
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_33_3
timestamp 1635107566
transform 1 0 1380 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  ring.x19.x5
timestamp 1635107566
transform -1 0 3220 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_18
timestamp 1635107566
transform 1 0 2760 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_15
timestamp 1635107566
transform 1 0 2484 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_16
timestamp 1635107566
transform 1 0 2576 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_33_11
timestamp 1635107566
transform 1 0 2116 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x19.x7_TE_B
timestamp 1635107566
transform 1 0 2576 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x16.x7_TE_B
timestamp 1635107566
transform -1 0 2576 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635107566
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__clkinv_1  ring.x19.x3
timestamp 1635107566
transform -1 0 3864 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1635107566
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_29
timestamp 1635107566
transform 1 0 3772 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_24
timestamp 1635107566
transform 1 0 3312 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_30
timestamp 1635107566
transform 1 0 3864 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_23
timestamp 1635107566
transform 1 0 3220 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x16.x2_TE_B
timestamp 1635107566
transform -1 0 3312 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  ring.x19.x1
timestamp 1635107566
transform -1 0 5152 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ring.x16.x5
timestamp 1635107566
transform -1 0 4416 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  ring.x16.x3
timestamp 1635107566
transform -1 0 4508 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_36
timestamp 1635107566
transform 1 0 4416 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_37
timestamp 1635107566
transform 1 0 4508 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__einvn_4  ring.x16.x2
timestamp 1635107566
transform -1 0 5888 0 -1 20672
box -38 -48 1050 592
use sky130_fd_sc_hd__decap_4  FILLER_33_52
timestamp 1635107566
transform 1 0 5888 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_44
timestamp 1635107566
transform 1 0 5152 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_55
timestamp 1635107566
transform 1 0 6164 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1635107566
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__einvp_2  ring.x16.x6
timestamp 1635107566
transform -1 0 6164 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ring.x16.x7
timestamp 1635107566
transform -1 0 8004 0 -1 20672
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_8  ring.x19.x7
timestamp 1635107566
transform 1 0 6532 0 1 20672
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_6  FILLER_33_75
timestamp 1635107566
transform 1 0 8004 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_77
timestamp 1635107566
transform 1 0 8188 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1635107566
transform -1 0 8832 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1635107566
transform -1 0 8832 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x42.x2_TE_B
timestamp 1635107566
transform -1 0 2760 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_15
timestamp 1635107566
transform 1 0 2484 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_18
timestamp 1635107566
transform 1 0 2760 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_3
timestamp 1635107566
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1635107566
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x16.x6_TE
timestamp 1635107566
transform -1 0 3864 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x19.x6_TE
timestamp 1635107566
transform 1 0 3128 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_24
timestamp 1635107566
transform 1 0 3312 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_30
timestamp 1635107566
transform 1 0 3864 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_37
timestamp 1635107566
transform 1 0 4508 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__einvn_4  ring.x42.x2
timestamp 1635107566
transform -1 0 5888 0 -1 21760
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_1  ring.x42.x5
timestamp 1635107566
transform -1 0 4508 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_52
timestamp 1635107566
transform 1 0 5888 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_61
timestamp 1635107566
transform 1 0 6716 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1635107566
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  ring.x16.x1
timestamp 1635107566
transform 1 0 6348 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_69
timestamp 1635107566
transform 1 0 7452 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_77
timestamp 1635107566
transform 1 0 8188 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1635107566
transform -1 0 8832 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ring.x19.x6
timestamp 1635107566
transform -1 0 8188 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x42.x7_TE_B
timestamp 1635107566
transform 1 0 2576 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_36_15
timestamp 1635107566
transform 1 0 2484 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_18
timestamp 1635107566
transform 1 0 2760 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_3
timestamp 1635107566
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1635107566
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x20.x2_TE_B
timestamp 1635107566
transform -1 0 3312 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_24
timestamp 1635107566
transform 1 0 3312 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_32
timestamp 1635107566
transform 1 0 4048 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1635107566
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_1  ring.x42.x3
timestamp 1635107566
transform -1 0 4048 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__einvn_8  ring.x42.x7
timestamp 1635107566
transform -1 0 6072 0 1 21760
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_8  FILLER_36_54
timestamp 1635107566
transform 1 0 6072 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__einvn_4  ring.x20.x2
timestamp 1635107566
transform -1 0 7820 0 1 21760
box -38 -48 1050 592
use sky130_fd_sc_hd__decap_8  FILLER_36_73
timestamp 1635107566
transform 1 0 7820 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1635107566
transform -1 0 8832 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x20.x7_TE_B
timestamp 1635107566
transform -1 0 3128 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x42.x4_TE
timestamp 1635107566
transform -1 0 2576 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_11
timestamp 1635107566
transform 1 0 2116 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_16
timestamp 1635107566
transform 1 0 2576 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_3
timestamp 1635107566
transform 1 0 1380 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1635107566
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_22
timestamp 1635107566
transform 1 0 3128 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_29
timestamp 1635107566
transform 1 0 3772 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_37
timestamp 1635107566
transform 1 0 4508 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ring.x20.x5
timestamp 1635107566
transform -1 0 3772 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ring.x42.x1
timestamp 1635107566
transform 1 0 4140 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_2  ring.x42.x4
timestamp 1635107566
transform -1 0 5520 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_37_48
timestamp 1635107566
transform 1 0 5520 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_57
timestamp 1635107566
transform 1 0 6348 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1635107566
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__einvn_8  ring.x20.x7
timestamp 1635107566
transform -1 0 8188 0 -1 22848
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_4  FILLER_37_77
timestamp 1635107566
transform 1 0 8188 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1635107566
transform -1 0 8832 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x42.x6_TE
timestamp 1635107566
transform -1 0 2760 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_15
timestamp 1635107566
transform 1 0 2484 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_18
timestamp 1635107566
transform 1 0 2760 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_3
timestamp 1635107566
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1635107566
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x20.x4_TE
timestamp 1635107566
transform -1 0 3956 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x20.x6_TE
timestamp 1635107566
transform -1 0 3312 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_24
timestamp 1635107566
transform 1 0 3312 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_31
timestamp 1635107566
transform 1 0 3956 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_38
timestamp 1635107566
transform 1 0 4600 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1635107566
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_1  ring.x20.x3
timestamp 1635107566
transform -1 0 4600 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ring.x42.x6
timestamp 1635107566
transform -1 0 5612 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_38_49
timestamp 1635107566
transform 1 0 5612 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_53
timestamp 1635107566
transform 1 0 5980 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_61
timestamp 1635107566
transform 1 0 6716 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_2  ring.x20.x4
timestamp 1635107566
transform -1 0 7728 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ring.x20.x6
timestamp 1635107566
transform -1 0 6716 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_38_72
timestamp 1635107566
transform 1 0 7728 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_80
timestamp 1635107566
transform 1 0 8464 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1635107566
transform -1 0 8832 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1635107566
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1635107566
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_40_9
timestamp 1635107566
transform 1 0 1932 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_3
timestamp 1635107566
transform 1 0 1380 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x24.x7_TE_B
timestamp 1635107566
transform -1 0 2208 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_18
timestamp 1635107566
transform 1 0 2760 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_12
timestamp 1635107566
transform 1 0 2208 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_21
timestamp 1635107566
transform 1 0 3036 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_15
timestamp 1635107566
transform 1 0 2484 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x24.x6_TE
timestamp 1635107566
transform -1 0 2760 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x24.x4_TE
timestamp 1635107566
transform -1 0 3036 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_3
timestamp 1635107566
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1635107566
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_40_29
timestamp 1635107566
transform 1 0 3772 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_24
timestamp 1635107566
transform 1 0 3312 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_27
timestamp 1635107566
transform 1 0 3588 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x22.x6_TE
timestamp 1635107566
transform -1 0 3312 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x22.x2_TE_B
timestamp 1635107566
transform -1 0 3588 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_2  ring.x24.x6
timestamp 1635107566
transform -1 0 5152 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  ring.x24.x5
timestamp 1635107566
transform -1 0 4232 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  ring.x24.x3
timestamp 1635107566
transform -1 0 4140 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_33
timestamp 1635107566
transform 1 0 4140 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_34
timestamp 1635107566
transform 1 0 4232 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ring.x22.x5
timestamp 1635107566
transform -1 0 4876 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_41
timestamp 1635107566
transform 1 0 4876 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_52
timestamp 1635107566
transform 1 0 5888 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_57
timestamp 1635107566
transform 1 0 6348 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_62
timestamp 1635107566
transform 1 0 6808 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_44
timestamp 1635107566
transform 1 0 5152 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1635107566
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  ring.x22.x1
timestamp 1635107566
transform -1 0 6808 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_2  ring.x24.x4
timestamp 1635107566
transform -1 0 5888 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ring.x24.x7
timestamp 1635107566
transform -1 0 7176 0 1 23936
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_4  FILLER_39_77
timestamp 1635107566
transform 1 0 8188 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_66
timestamp 1635107566
transform 1 0 7176 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_77
timestamp 1635107566
transform 1 0 8188 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1635107566
transform -1 0 8832 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1635107566
transform -1 0 8832 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__einvn_4  ring.x22.x2
timestamp 1635107566
transform -1 0 8188 0 -1 23936
box -38 -48 1050 592
use sky130_fd_sc_hd__einvp_2  ring.x22.x6
timestamp 1635107566
transform -1 0 8188 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x24.x2_TE_B
timestamp 1635107566
transform 1 0 2852 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x41.x4_TE
timestamp 1635107566
transform -1 0 2484 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x41.x7_TE_B
timestamp 1635107566
transform -1 0 1932 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_15
timestamp 1635107566
transform 1 0 2484 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_21
timestamp 1635107566
transform 1 0 3036 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_3
timestamp 1635107566
transform 1 0 1380 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_9
timestamp 1635107566
transform 1 0 1932 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1635107566
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_28
timestamp 1635107566
transform 1 0 3680 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ring.x41.x5
timestamp 1635107566
transform -1 0 3680 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__einvn_8  ring.x41.x7
timestamp 1635107566
transform -1 0 5704 0 -1 25024
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_6  FILLER_41_50
timestamp 1635107566
transform 1 0 5704 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1635107566
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__einvn_4  ring.x24.x2
timestamp 1635107566
transform -1 0 7360 0 -1 25024
box -38 -48 1050 592
use sky130_fd_sc_hd__decap_4  FILLER_41_68
timestamp 1635107566
transform 1 0 7360 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_72
timestamp 1635107566
transform 1 0 7728 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_77
timestamp 1635107566
transform 1 0 8188 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1635107566
transform -1 0 8832 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ring.x20.x1
timestamp 1635107566
transform -1 0 8188 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x22.x7_TE_B
timestamp 1635107566
transform -1 0 2668 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x25.x4_TE
timestamp 1635107566
transform 1 0 1932 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_11
timestamp 1635107566
transform 1 0 2116 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_17
timestamp 1635107566
transform 1 0 2668 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_3
timestamp 1635107566
transform 1 0 1380 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1635107566
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  ring.x41.x3
timestamp 1635107566
transform -1 0 3312 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_24
timestamp 1635107566
transform 1 0 3312 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_29
timestamp 1635107566
transform 1 0 3772 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_40
timestamp 1635107566
transform 1 0 4784 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1635107566
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__einvp_2  ring.x41.x4
timestamp 1635107566
transform -1 0 4784 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_42_51
timestamp 1635107566
transform 1 0 5796 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__einvn_8  ring.x22.x7
timestamp 1635107566
transform -1 0 8188 0 1 25024
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_2  ring.x25.x4
timestamp 1635107566
transform -1 0 5796 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_42_77
timestamp 1635107566
transform 1 0 8188 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1635107566
transform -1 0 8832 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x23.x2_TE_B
timestamp 1635107566
transform -1 0 2392 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x25.x7_TE_B
timestamp 1635107566
transform -1 0 1840 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_14
timestamp 1635107566
transform 1 0 2392 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_43_3
timestamp 1635107566
transform 1 0 1380 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_8
timestamp 1635107566
transform 1 0 1840 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1635107566
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ring.x41.x1
timestamp 1635107566
transform 1 0 2760 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_22
timestamp 1635107566
transform 1 0 3128 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_30
timestamp 1635107566
transform 1 0 3864 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  ring.x25.x1
timestamp 1635107566
transform 1 0 3496 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__einvn_8  ring.x25.x7
timestamp 1635107566
transform 1 0 4232 0 -1 26112
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_4  FILLER_43_52
timestamp 1635107566
transform 1 0 5888 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_60
timestamp 1635107566
transform 1 0 6624 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1635107566
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_1  ring.x22.x3
timestamp 1635107566
transform -1 0 6624 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__einvn_4  ring.x23.x2
timestamp 1635107566
transform -1 0 8004 0 -1 26112
box -38 -48 1050 592
use sky130_fd_sc_hd__decap_6  FILLER_43_75
timestamp 1635107566
transform 1 0 8004 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1635107566
transform -1 0 8832 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x23.x7_TE_B
timestamp 1635107566
transform -1 0 2668 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x25.x6_TE
timestamp 1635107566
transform -1 0 2116 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_11
timestamp 1635107566
transform 1 0 2116 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_17
timestamp 1635107566
transform 1 0 2668 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_3
timestamp 1635107566
transform 1 0 1380 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1635107566
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ring.x23.x5
timestamp 1635107566
transform -1 0 3312 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_24
timestamp 1635107566
transform 1 0 3312 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_29
timestamp 1635107566
transform 1 0 3772 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_38
timestamp 1635107566
transform 1 0 4600 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1635107566
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__einvn_4  ring.x25.x2
timestamp 1635107566
transform -1 0 5980 0 1 26112
box -38 -48 1050 592
use sky130_fd_sc_hd__einvp_2  ring.x25.x6
timestamp 1635107566
transform -1 0 4600 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_44_53
timestamp 1635107566
transform 1 0 5980 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__einvn_8  ring.x23.x7
timestamp 1635107566
transform -1 0 8004 0 1 26112
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_6  FILLER_44_75
timestamp 1635107566
transform 1 0 8004 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1635107566
transform -1 0 8832 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x25.x2_TE_B
timestamp 1635107566
transform 1 0 2484 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x41.x2_TE_B
timestamp 1635107566
transform -1 0 2116 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_11
timestamp 1635107566
transform 1 0 2116 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_17
timestamp 1635107566
transform 1 0 2668 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_3
timestamp 1635107566
transform 1 0 1380 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1635107566
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  ring.x25.x3
timestamp 1635107566
transform -1 0 3312 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_24
timestamp 1635107566
transform 1 0 3312 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_31
timestamp 1635107566
transform 1 0 3956 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_1  ring.x23.x3
timestamp 1635107566
transform -1 0 3956 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__einvn_4  ring.x41.x2
timestamp 1635107566
transform -1 0 5336 0 -1 27200
box -38 -48 1050 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x22.x4_TE
timestamp 1635107566
transform 1 0 5704 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_46
timestamp 1635107566
transform 1 0 5336 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_52
timestamp 1635107566
transform 1 0 5888 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_57
timestamp 1635107566
transform 1 0 6348 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1635107566
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__einvp_2  ring.x23.x4
timestamp 1635107566
transform -1 0 7176 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_45_66
timestamp 1635107566
transform 1 0 7176 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_77
timestamp 1635107566
transform 1 0 8188 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1635107566
transform -1 0 8832 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ring.x22.x4
timestamp 1635107566
transform -1 0 8188 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x23.x6_TE
timestamp 1635107566
transform -1 0 2760 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x41.x6_TE
timestamp 1635107566
transform 1 0 2024 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_12
timestamp 1635107566
transform 1 0 2208 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_18
timestamp 1635107566
transform 1 0 2760 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_3
timestamp 1635107566
transform 1 0 1380 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_9
timestamp 1635107566
transform 1 0 1932 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1635107566
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ring.x23.x4_TE
timestamp 1635107566
transform -1 0 3312 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_24
timestamp 1635107566
transform 1 0 3312 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_32
timestamp 1635107566
transform 1 0 4048 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_43
timestamp 1635107566
transform 1 0 5060 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1635107566
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  ring.x25.x5
timestamp 1635107566
transform -1 0 4048 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ring.x41.x6
timestamp 1635107566
transform -1 0 5060 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_46_47
timestamp 1635107566
transform 1 0 5428 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_52
timestamp 1635107566
transform 1 0 5888 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_57
timestamp 1635107566
transform 1 0 6348 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_63
timestamp 1635107566
transform 1 0 6900 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1635107566
transform 1 0 6256 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  ring.x23.x1
timestamp 1635107566
transform -1 0 6900 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  ring.x24.x1
timestamp 1635107566
transform -1 0 5888 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_74
timestamp 1635107566
transform 1 0 7912 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_80
timestamp 1635107566
transform 1 0 8464 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1635107566
transform -1 0 8832 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ring.x23.x6
timestamp 1635107566
transform -1 0 7912 0 1 27200
box -38 -48 682 592
<< labels >>
rlabel metal2 s 6918 0 6974 800 6 clk_out
port 0 nsew signal tristate
rlabel metal2 s 938 0 994 800 6 clkmux[0]
port 1 nsew signal input
rlabel metal2 s 2870 0 2926 800 6 clkmux[1]
port 2 nsew signal input
rlabel metal2 s 4894 0 4950 800 6 clkmux[2]
port 3 nsew signal input
rlabel metal2 s 8942 0 8998 800 6 start
port 4 nsew signal input
rlabel metal3 s 9200 144 10000 264 6 trim_a[0]
port 5 nsew signal input
rlabel metal3 s 9200 5448 10000 5568 6 trim_a[10]
port 6 nsew signal input
rlabel metal3 s 9200 5992 10000 6112 6 trim_a[11]
port 7 nsew signal input
rlabel metal3 s 9200 6536 10000 6656 6 trim_a[12]
port 8 nsew signal input
rlabel metal3 s 9200 7080 10000 7200 6 trim_a[13]
port 9 nsew signal input
rlabel metal3 s 9200 7624 10000 7744 6 trim_a[14]
port 10 nsew signal input
rlabel metal3 s 9200 8168 10000 8288 6 trim_a[15]
port 11 nsew signal input
rlabel metal3 s 9200 8712 10000 8832 6 trim_a[16]
port 12 nsew signal input
rlabel metal3 s 9200 9256 10000 9376 6 trim_a[17]
port 13 nsew signal input
rlabel metal3 s 9200 9800 10000 9920 6 trim_a[18]
port 14 nsew signal input
rlabel metal3 s 9200 10208 10000 10328 6 trim_a[19]
port 15 nsew signal input
rlabel metal3 s 9200 552 10000 672 6 trim_a[1]
port 16 nsew signal input
rlabel metal3 s 9200 10752 10000 10872 6 trim_a[20]
port 17 nsew signal input
rlabel metal3 s 9200 11296 10000 11416 6 trim_a[21]
port 18 nsew signal input
rlabel metal3 s 9200 11840 10000 11960 6 trim_a[22]
port 19 nsew signal input
rlabel metal3 s 9200 12384 10000 12504 6 trim_a[23]
port 20 nsew signal input
rlabel metal3 s 9200 12928 10000 13048 6 trim_a[24]
port 21 nsew signal input
rlabel metal3 s 9200 13472 10000 13592 6 trim_a[25]
port 22 nsew signal input
rlabel metal3 s 9200 14016 10000 14136 6 trim_a[26]
port 23 nsew signal input
rlabel metal3 s 9200 14560 10000 14680 6 trim_a[27]
port 24 nsew signal input
rlabel metal3 s 9200 1096 10000 1216 6 trim_a[2]
port 25 nsew signal input
rlabel metal3 s 9200 1640 10000 1760 6 trim_a[3]
port 26 nsew signal input
rlabel metal3 s 9200 2184 10000 2304 6 trim_a[4]
port 27 nsew signal input
rlabel metal3 s 9200 2728 10000 2848 6 trim_a[5]
port 28 nsew signal input
rlabel metal3 s 9200 3272 10000 3392 6 trim_a[6]
port 29 nsew signal input
rlabel metal3 s 9200 3816 10000 3936 6 trim_a[7]
port 30 nsew signal input
rlabel metal3 s 9200 4360 10000 4480 6 trim_a[8]
port 31 nsew signal input
rlabel metal3 s 9200 4904 10000 5024 6 trim_a[9]
port 32 nsew signal input
rlabel metal3 s 9200 15104 10000 15224 6 trim_b[0]
port 33 nsew signal input
rlabel metal3 s 9200 20408 10000 20528 6 trim_b[10]
port 34 nsew signal input
rlabel metal3 s 9200 20952 10000 21072 6 trim_b[11]
port 35 nsew signal input
rlabel metal3 s 9200 21496 10000 21616 6 trim_b[12]
port 36 nsew signal input
rlabel metal3 s 9200 22040 10000 22160 6 trim_b[13]
port 37 nsew signal input
rlabel metal3 s 9200 22584 10000 22704 6 trim_b[14]
port 38 nsew signal input
rlabel metal3 s 9200 23128 10000 23248 6 trim_b[15]
port 39 nsew signal input
rlabel metal3 s 9200 23672 10000 23792 6 trim_b[16]
port 40 nsew signal input
rlabel metal3 s 9200 24216 10000 24336 6 trim_b[17]
port 41 nsew signal input
rlabel metal3 s 9200 24760 10000 24880 6 trim_b[18]
port 42 nsew signal input
rlabel metal3 s 9200 25304 10000 25424 6 trim_b[19]
port 43 nsew signal input
rlabel metal3 s 9200 15648 10000 15768 6 trim_b[1]
port 44 nsew signal input
rlabel metal3 s 9200 25848 10000 25968 6 trim_b[20]
port 45 nsew signal input
rlabel metal3 s 9200 26392 10000 26512 6 trim_b[21]
port 46 nsew signal input
rlabel metal3 s 9200 26936 10000 27056 6 trim_b[22]
port 47 nsew signal input
rlabel metal3 s 9200 27480 10000 27600 6 trim_b[23]
port 48 nsew signal input
rlabel metal3 s 9200 28024 10000 28144 6 trim_b[24]
port 49 nsew signal input
rlabel metal3 s 9200 28568 10000 28688 6 trim_b[25]
port 50 nsew signal input
rlabel metal3 s 9200 29112 10000 29232 6 trim_b[26]
port 51 nsew signal input
rlabel metal3 s 9200 29656 10000 29776 6 trim_b[27]
port 52 nsew signal input
rlabel metal3 s 9200 16192 10000 16312 6 trim_b[2]
port 53 nsew signal input
rlabel metal3 s 9200 16736 10000 16856 6 trim_b[3]
port 54 nsew signal input
rlabel metal3 s 9200 17280 10000 17400 6 trim_b[4]
port 55 nsew signal input
rlabel metal3 s 9200 17824 10000 17944 6 trim_b[5]
port 56 nsew signal input
rlabel metal3 s 9200 18368 10000 18488 6 trim_b[6]
port 57 nsew signal input
rlabel metal3 s 9200 18912 10000 19032 6 trim_b[7]
port 58 nsew signal input
rlabel metal3 s 9200 19456 10000 19576 6 trim_b[8]
port 59 nsew signal input
rlabel metal3 s 9200 20000 10000 20120 6 trim_b[9]
port 60 nsew signal input
rlabel metal4 s 2243 2128 2563 27792 6 vccd1
port 61 nsew power input
rlabel metal4 s 4840 2128 5160 27792 6 vccd1
port 61 nsew power input
rlabel metal4 s 7437 2128 7757 27792 6 vccd1
port 61 nsew power input
rlabel metal4 s 3541 2128 3861 27792 6 vssd1
port 62 nsew ground input
rlabel metal4 s 6138 2128 6458 27792 6 vssd1
port 62 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 10000 30000
<< end >>
