magic
tech sky130A
magscale 1 2
timestamp 1641029093
<< metal1 >>
rect 331214 702992 331220 703044
rect 331272 703032 331278 703044
rect 332502 703032 332508 703044
rect 331272 703004 332508 703032
rect 331272 702992 331278 703004
rect 332502 702992 332508 703004
rect 332560 702992 332566 703044
rect 170306 700884 170312 700936
rect 170364 700924 170370 700936
rect 171042 700924 171048 700936
rect 170364 700896 171048 700924
rect 170364 700884 170370 700896
rect 171042 700884 171048 700896
rect 171100 700884 171106 700936
rect 252462 700612 252468 700664
rect 252520 700652 252526 700664
rect 283834 700652 283840 700664
rect 252520 700624 283840 700652
rect 252520 700612 252526 700624
rect 283834 700612 283840 700624
rect 283892 700612 283898 700664
rect 246942 700544 246948 700596
rect 247000 700584 247006 700596
rect 413646 700584 413652 700596
rect 247000 700556 413652 700584
rect 247000 700544 247006 700556
rect 413646 700544 413652 700556
rect 413704 700544 413710 700596
rect 72970 700476 72976 700528
rect 73028 700516 73034 700528
rect 258074 700516 258080 700528
rect 73028 700488 258080 700516
rect 73028 700476 73034 700488
rect 258074 700476 258080 700488
rect 258132 700476 258138 700528
rect 40494 700408 40500 700460
rect 40552 700448 40558 700460
rect 41322 700448 41328 700460
rect 40552 700420 41328 700448
rect 40552 700408 40558 700420
rect 41322 700408 41328 700420
rect 41380 700408 41386 700460
rect 235166 700408 235172 700460
rect 235224 700448 235230 700460
rect 242158 700448 242164 700460
rect 235224 700420 242164 700448
rect 235224 700408 235230 700420
rect 242158 700408 242164 700420
rect 242216 700408 242222 700460
rect 244182 700408 244188 700460
rect 244240 700448 244246 700460
rect 478506 700448 478512 700460
rect 244240 700420 478512 700448
rect 244240 700408 244246 700420
rect 478506 700408 478512 700420
rect 478564 700408 478570 700460
rect 24302 700340 24308 700392
rect 24360 700380 24366 700392
rect 260098 700380 260104 700392
rect 24360 700352 260104 700380
rect 24360 700340 24366 700352
rect 260098 700340 260104 700352
rect 260156 700340 260162 700392
rect 479518 700340 479524 700392
rect 479576 700380 479582 700392
rect 527174 700380 527180 700392
rect 479576 700352 527180 700380
rect 479576 700340 479582 700352
rect 527174 700340 527180 700352
rect 527232 700340 527238 700392
rect 218974 700272 218980 700324
rect 219032 700312 219038 700324
rect 222838 700312 222844 700324
rect 219032 700284 222844 700312
rect 219032 700272 219038 700284
rect 222838 700272 222844 700284
rect 222896 700272 222902 700324
rect 241422 700272 241428 700324
rect 241480 700312 241486 700324
rect 543458 700312 543464 700324
rect 241480 700284 543464 700312
rect 241480 700272 241486 700284
rect 543458 700272 543464 700284
rect 543516 700272 543522 700324
rect 105446 699660 105452 699712
rect 105504 699700 105510 699712
rect 106182 699700 106188 699712
rect 105504 699672 106188 699700
rect 105504 699660 105510 699672
rect 106182 699660 106188 699672
rect 106240 699660 106246 699712
rect 154114 699660 154120 699712
rect 154172 699700 154178 699712
rect 155218 699700 155224 699712
rect 154172 699672 155224 699700
rect 154172 699660 154178 699672
rect 155218 699660 155224 699672
rect 155276 699660 155282 699712
rect 347038 699660 347044 699712
rect 347096 699700 347102 699712
rect 348786 699700 348792 699712
rect 347096 699672 348792 699700
rect 347096 699660 347102 699672
rect 348786 699660 348792 699672
rect 348844 699660 348850 699712
rect 359458 699660 359464 699712
rect 359516 699700 359522 699712
rect 364978 699700 364984 699712
rect 359516 699672 364984 699700
rect 359516 699660 359522 699672
rect 364978 699660 364984 699672
rect 365036 699660 365042 699712
rect 396718 699660 396724 699712
rect 396776 699700 396782 699712
rect 397454 699700 397460 699712
rect 396776 699672 397460 699700
rect 396776 699660 396782 699672
rect 397454 699660 397460 699672
rect 397512 699660 397518 699712
rect 249058 698912 249064 698964
rect 249116 698952 249122 698964
rect 462314 698952 462320 698964
rect 249116 698924 462320 698952
rect 249116 698912 249122 698924
rect 462314 698912 462320 698924
rect 462372 698912 462378 698964
rect 266354 697552 266360 697604
rect 266412 697592 266418 697604
rect 267642 697592 267648 697604
rect 266412 697564 267648 697592
rect 266412 697552 266418 697564
rect 267642 697552 267648 697564
rect 267700 697552 267706 697604
rect 238662 696940 238668 696992
rect 238720 696980 238726 696992
rect 580166 696980 580172 696992
rect 238720 696952 580172 696980
rect 238720 696940 238726 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 3418 683204 3424 683256
rect 3476 683244 3482 683256
rect 262214 683244 262220 683256
rect 3476 683216 262220 683244
rect 3476 683204 3482 683216
rect 262214 683204 262220 683216
rect 262272 683204 262278 683256
rect 238570 683136 238576 683188
rect 238628 683176 238634 683188
rect 580166 683176 580172 683188
rect 238628 683148 580172 683176
rect 238628 683136 238634 683148
rect 580166 683136 580172 683148
rect 580224 683136 580230 683188
rect 237282 670692 237288 670744
rect 237340 670732 237346 670744
rect 580166 670732 580172 670744
rect 237340 670704 580172 670732
rect 237340 670692 237346 670704
rect 580166 670692 580172 670704
rect 580224 670692 580230 670744
rect 3510 656888 3516 656940
rect 3568 656928 3574 656940
rect 263686 656928 263692 656940
rect 3568 656900 263692 656928
rect 3568 656888 3574 656900
rect 263686 656888 263692 656900
rect 263744 656888 263750 656940
rect 235902 643084 235908 643136
rect 235960 643124 235966 643136
rect 580166 643124 580172 643136
rect 235960 643096 580172 643124
rect 235960 643084 235966 643096
rect 580166 643084 580172 643096
rect 580224 643084 580230 643136
rect 3510 632068 3516 632120
rect 3568 632108 3574 632120
rect 264974 632108 264980 632120
rect 3568 632080 264980 632108
rect 3568 632068 3574 632080
rect 264974 632068 264980 632080
rect 265032 632068 265038 632120
rect 237190 630640 237196 630692
rect 237248 630680 237254 630692
rect 580166 630680 580172 630692
rect 237248 630652 580172 630680
rect 237248 630640 237254 630652
rect 580166 630640 580172 630652
rect 580224 630640 580230 630692
rect 3510 618264 3516 618316
rect 3568 618304 3574 618316
rect 217318 618304 217324 618316
rect 3568 618276 217324 618304
rect 3568 618264 3574 618276
rect 217318 618264 217324 618276
rect 217376 618264 217382 618316
rect 234522 616836 234528 616888
rect 234580 616876 234586 616888
rect 580166 616876 580172 616888
rect 234580 616848 580172 616876
rect 234580 616836 234586 616848
rect 580166 616836 580172 616848
rect 580224 616836 580230 616888
rect 250990 607860 250996 607912
rect 251048 607900 251054 607912
rect 266354 607900 266360 607912
rect 251048 607872 266360 607900
rect 251048 607860 251054 607872
rect 266354 607860 266360 607872
rect 266412 607860 266418 607912
rect 3510 605820 3516 605872
rect 3568 605860 3574 605872
rect 266354 605860 266360 605872
rect 3568 605832 266360 605860
rect 3568 605820 3574 605832
rect 266354 605820 266360 605832
rect 266412 605820 266418 605872
rect 233142 590656 233148 590708
rect 233200 590696 233206 590708
rect 579798 590696 579804 590708
rect 233200 590668 579804 590696
rect 233200 590656 233206 590668
rect 579798 590656 579804 590668
rect 579856 590656 579862 590708
rect 3326 579640 3332 579692
rect 3384 579680 3390 579692
rect 267734 579680 267740 579692
rect 3384 579652 267740 579680
rect 3384 579640 3390 579652
rect 267734 579640 267740 579652
rect 267792 579640 267798 579692
rect 234430 576852 234436 576904
rect 234488 576892 234494 576904
rect 580166 576892 580172 576904
rect 234488 576864 580172 576892
rect 234488 576852 234494 576864
rect 580166 576852 580172 576864
rect 580224 576852 580230 576904
rect 3234 565836 3240 565888
rect 3292 565876 3298 565888
rect 215938 565876 215944 565888
rect 3292 565848 215944 565876
rect 3292 565836 3298 565848
rect 215938 565836 215944 565848
rect 215996 565836 216002 565888
rect 231762 563048 231768 563100
rect 231820 563088 231826 563100
rect 579798 563088 579804 563100
rect 231820 563060 579804 563088
rect 231820 563048 231826 563060
rect 579798 563048 579804 563060
rect 579856 563048 579862 563100
rect 3326 553392 3332 553444
rect 3384 553432 3390 553444
rect 267826 553432 267832 553444
rect 3384 553404 267832 553432
rect 3384 553392 3390 553404
rect 267826 553392 267832 553404
rect 267884 553392 267890 553444
rect 230382 536800 230388 536852
rect 230440 536840 230446 536852
rect 580166 536840 580172 536852
rect 230440 536812 580172 536840
rect 230440 536800 230446 536812
rect 580166 536800 580172 536812
rect 580224 536800 580230 536852
rect 2958 527144 2964 527196
rect 3016 527184 3022 527196
rect 270494 527184 270500 527196
rect 3016 527156 270500 527184
rect 3016 527144 3022 527156
rect 270494 527144 270500 527156
rect 270552 527144 270558 527196
rect 231670 524424 231676 524476
rect 231728 524464 231734 524476
rect 580166 524464 580172 524476
rect 231728 524436 580172 524464
rect 231728 524424 231734 524436
rect 580166 524424 580172 524436
rect 580224 524424 580230 524476
rect 3510 514768 3516 514820
rect 3568 514808 3574 514820
rect 269758 514808 269764 514820
rect 3568 514780 269764 514808
rect 3568 514768 3574 514780
rect 269758 514768 269764 514780
rect 269816 514768 269822 514820
rect 229002 510620 229008 510672
rect 229060 510660 229066 510672
rect 580166 510660 580172 510672
rect 229060 510632 580172 510660
rect 229060 510620 229066 510632
rect 580166 510620 580172 510632
rect 580224 510620 580230 510672
rect 3050 500964 3056 501016
rect 3108 501004 3114 501016
rect 270586 501004 270592 501016
rect 3108 500976 270592 501004
rect 3108 500964 3114 500976
rect 270586 500964 270592 500976
rect 270644 500964 270650 501016
rect 227622 484372 227628 484424
rect 227680 484412 227686 484424
rect 580166 484412 580172 484424
rect 227680 484384 580172 484412
rect 227680 484372 227686 484384
rect 580166 484372 580172 484384
rect 580224 484372 580230 484424
rect 3050 474716 3056 474768
rect 3108 474756 3114 474768
rect 273254 474756 273260 474768
rect 3108 474728 273260 474756
rect 3108 474716 3114 474728
rect 273254 474716 273260 474728
rect 273312 474716 273318 474768
rect 228910 470568 228916 470620
rect 228968 470608 228974 470620
rect 579982 470608 579988 470620
rect 228968 470580 579988 470608
rect 228968 470568 228974 470580
rect 579982 470568 579988 470580
rect 580040 470568 580046 470620
rect 3510 462340 3516 462392
rect 3568 462380 3574 462392
rect 214558 462380 214564 462392
rect 3568 462352 214564 462380
rect 3568 462340 3574 462352
rect 214558 462340 214564 462352
rect 214616 462340 214622 462392
rect 227530 456764 227536 456816
rect 227588 456804 227594 456816
rect 580166 456804 580172 456816
rect 227588 456776 580172 456804
rect 227588 456764 227594 456776
rect 580166 456764 580172 456776
rect 580224 456764 580230 456816
rect 3142 448536 3148 448588
rect 3200 448576 3206 448588
rect 273346 448576 273352 448588
rect 3200 448548 273352 448576
rect 3200 448536 3206 448548
rect 273346 448536 273352 448548
rect 273404 448536 273410 448588
rect 224862 430584 224868 430636
rect 224920 430624 224926 430636
rect 580166 430624 580172 430636
rect 224920 430596 580172 430624
rect 224920 430584 224926 430596
rect 580166 430584 580172 430596
rect 580224 430584 580230 430636
rect 3510 422288 3516 422340
rect 3568 422328 3574 422340
rect 276014 422328 276020 422340
rect 3568 422300 276020 422328
rect 3568 422288 3574 422300
rect 276014 422288 276020 422300
rect 276072 422288 276078 422340
rect 226242 418140 226248 418192
rect 226300 418180 226306 418192
rect 580166 418180 580172 418192
rect 226300 418152 580172 418180
rect 226300 418140 226306 418152
rect 580166 418140 580172 418152
rect 580224 418140 580230 418192
rect 2866 409844 2872 409896
rect 2924 409884 2930 409896
rect 213178 409884 213184 409896
rect 2924 409856 213184 409884
rect 2924 409844 2930 409856
rect 213178 409844 213184 409856
rect 213236 409844 213242 409896
rect 224770 404336 224776 404388
rect 224828 404376 224834 404388
rect 580166 404376 580172 404388
rect 224828 404348 580172 404376
rect 224828 404336 224834 404348
rect 580166 404336 580172 404348
rect 580224 404336 580230 404388
rect 3510 397468 3516 397520
rect 3568 397508 3574 397520
rect 276106 397508 276112 397520
rect 3568 397480 276112 397508
rect 3568 397468 3574 397480
rect 276106 397468 276112 397480
rect 276164 397468 276170 397520
rect 3510 371220 3516 371272
rect 3568 371260 3574 371272
rect 277394 371260 277400 371272
rect 3568 371232 277400 371260
rect 3568 371220 3574 371232
rect 277394 371220 277400 371232
rect 277452 371220 277458 371272
rect 371602 368908 371608 368960
rect 371660 368948 371666 368960
rect 374178 368948 374184 368960
rect 371660 368920 374184 368948
rect 371660 368908 371666 368920
rect 374178 368908 374184 368920
rect 374236 368908 374242 368960
rect 445202 368500 445208 368552
rect 445260 368540 445266 368552
rect 454034 368540 454040 368552
rect 445260 368512 454040 368540
rect 445260 368500 445266 368512
rect 454034 368500 454040 368512
rect 454092 368500 454098 368552
rect 371602 367140 371608 367192
rect 371660 367180 371666 367192
rect 378134 367180 378140 367192
rect 371660 367152 378140 367180
rect 371660 367140 371666 367152
rect 378134 367140 378140 367152
rect 378192 367140 378198 367192
rect 371694 367072 371700 367124
rect 371752 367112 371758 367124
rect 383654 367112 383660 367124
rect 371752 367084 383660 367112
rect 371752 367072 371758 367084
rect 383654 367072 383660 367084
rect 383712 367072 383718 367124
rect 445662 367072 445668 367124
rect 445720 367112 445726 367124
rect 449894 367112 449900 367124
rect 445720 367084 449900 367112
rect 445720 367072 445726 367084
rect 449894 367072 449900 367084
rect 449952 367072 449958 367124
rect 371602 365848 371608 365900
rect 371660 365888 371666 365900
rect 376938 365888 376944 365900
rect 371660 365860 376944 365888
rect 371660 365848 371666 365860
rect 376938 365848 376944 365860
rect 376996 365848 377002 365900
rect 371234 365780 371240 365832
rect 371292 365820 371298 365832
rect 382274 365820 382280 365832
rect 371292 365792 382280 365820
rect 371292 365780 371298 365792
rect 382274 365780 382280 365792
rect 382332 365780 382338 365832
rect 371510 365712 371516 365764
rect 371568 365752 371574 365764
rect 385034 365752 385040 365764
rect 371568 365724 385040 365752
rect 371568 365712 371574 365724
rect 385034 365712 385040 365724
rect 385092 365712 385098 365764
rect 445294 365712 445300 365764
rect 445352 365752 445358 365764
rect 456794 365752 456800 365764
rect 445352 365724 456800 365752
rect 445352 365712 445358 365724
rect 456794 365712 456800 365724
rect 456852 365712 456858 365764
rect 371234 364624 371240 364676
rect 371292 364664 371298 364676
rect 375558 364664 375564 364676
rect 371292 364636 375564 364664
rect 371292 364624 371298 364636
rect 375558 364624 375564 364636
rect 375616 364624 375622 364676
rect 371602 364352 371608 364404
rect 371660 364392 371666 364404
rect 382366 364392 382372 364404
rect 371660 364364 382372 364392
rect 371660 364352 371666 364364
rect 382366 364352 382372 364364
rect 382424 364352 382430 364404
rect 445662 364352 445668 364404
rect 445720 364392 445726 364404
rect 452746 364392 452752 364404
rect 445720 364364 452752 364392
rect 445720 364352 445726 364364
rect 452746 364352 452752 364364
rect 452804 364352 452810 364404
rect 371602 363060 371608 363112
rect 371660 363100 371666 363112
rect 378318 363100 378324 363112
rect 371660 363072 378324 363100
rect 371660 363060 371666 363072
rect 378318 363060 378324 363072
rect 378376 363060 378382 363112
rect 371694 362924 371700 362976
rect 371752 362964 371758 362976
rect 374270 362964 374276 362976
rect 371752 362936 374276 362964
rect 371752 362924 371758 362936
rect 374270 362924 374276 362936
rect 374328 362924 374334 362976
rect 444926 362924 444932 362976
rect 444984 362964 444990 362976
rect 448606 362964 448612 362976
rect 444984 362936 448612 362964
rect 444984 362924 444990 362936
rect 448606 362924 448612 362936
rect 448664 362924 448670 362976
rect 371602 361632 371608 361684
rect 371660 361672 371666 361684
rect 377030 361672 377036 361684
rect 371660 361644 377036 361672
rect 371660 361632 371666 361644
rect 377030 361632 377036 361644
rect 377088 361632 377094 361684
rect 371694 361564 371700 361616
rect 371752 361604 371758 361616
rect 380986 361604 380992 361616
rect 371752 361576 380992 361604
rect 371752 361564 371758 361576
rect 380986 361564 380992 361576
rect 381044 361564 381050 361616
rect 445202 361564 445208 361616
rect 445260 361604 445266 361616
rect 454126 361604 454132 361616
rect 445260 361576 454132 361604
rect 445260 361564 445266 361576
rect 454126 361564 454132 361576
rect 454184 361564 454190 361616
rect 371602 361496 371608 361548
rect 371660 361536 371666 361548
rect 375374 361536 375380 361548
rect 371660 361508 375380 361536
rect 371660 361496 371666 361508
rect 375374 361496 375380 361508
rect 375432 361496 375438 361548
rect 445110 360748 445116 360800
rect 445168 360788 445174 360800
rect 449986 360788 449992 360800
rect 445168 360760 449992 360788
rect 445168 360748 445174 360760
rect 449986 360748 449992 360760
rect 450044 360748 450050 360800
rect 371602 360408 371608 360460
rect 371660 360448 371666 360460
rect 374454 360448 374460 360460
rect 371660 360420 374460 360448
rect 371660 360408 371666 360420
rect 374454 360408 374460 360420
rect 374512 360408 374518 360460
rect 371418 360340 371424 360392
rect 371476 360380 371482 360392
rect 378226 360380 378232 360392
rect 371476 360352 378232 360380
rect 371476 360340 371482 360352
rect 378226 360340 378232 360352
rect 378284 360340 378290 360392
rect 444558 360272 444564 360324
rect 444616 360312 444622 360324
rect 452654 360312 452660 360324
rect 444616 360284 452660 360312
rect 444616 360272 444622 360284
rect 452654 360272 452660 360284
rect 452712 360272 452718 360324
rect 371878 359524 371884 359576
rect 371936 359564 371942 359576
rect 379514 359564 379520 359576
rect 371936 359536 379520 359564
rect 371936 359524 371942 359536
rect 379514 359524 379520 359536
rect 379572 359524 379578 359576
rect 372062 359456 372068 359508
rect 372120 359496 372126 359508
rect 372890 359496 372896 359508
rect 372120 359468 372896 359496
rect 372120 359456 372126 359468
rect 372890 359456 372896 359468
rect 372948 359456 372954 359508
rect 371694 357484 371700 357536
rect 371752 357524 371758 357536
rect 376754 357524 376760 357536
rect 371752 357496 376760 357524
rect 371752 357484 371758 357496
rect 376754 357484 376760 357496
rect 376812 357484 376818 357536
rect 3142 357416 3148 357468
rect 3200 357456 3206 357468
rect 253198 357456 253204 357468
rect 3200 357428 253204 357456
rect 3200 357416 3206 357428
rect 253198 357416 253204 357428
rect 253256 357416 253262 357468
rect 371602 357416 371608 357468
rect 371660 357456 371666 357468
rect 382550 357456 382556 357468
rect 371660 357428 382556 357456
rect 371660 357416 371666 357428
rect 382550 357416 382556 357428
rect 382608 357416 382614 357468
rect 444558 357416 444564 357468
rect 444616 357456 444622 357468
rect 448514 357456 448520 357468
rect 444616 357428 448520 357456
rect 444616 357416 444622 357428
rect 448514 357416 448520 357428
rect 448572 357416 448578 357468
rect 371602 356192 371608 356244
rect 371660 356232 371666 356244
rect 375650 356232 375656 356244
rect 371660 356204 375656 356232
rect 371660 356192 371666 356204
rect 375650 356192 375656 356204
rect 375708 356192 375714 356244
rect 444374 356192 444380 356244
rect 444432 356232 444438 356244
rect 447134 356232 447140 356244
rect 444432 356204 447140 356232
rect 444432 356192 444438 356204
rect 447134 356192 447140 356204
rect 447192 356192 447198 356244
rect 371234 356124 371240 356176
rect 371292 356164 371298 356176
rect 381078 356164 381084 356176
rect 371292 356136 381084 356164
rect 371292 356124 371298 356136
rect 381078 356124 381084 356136
rect 381136 356124 381142 356176
rect 371510 356056 371516 356108
rect 371568 356096 371574 356108
rect 385218 356096 385224 356108
rect 371568 356068 385224 356096
rect 371568 356056 371574 356068
rect 385218 356056 385224 356068
rect 385276 356056 385282 356108
rect 444742 355036 444748 355088
rect 444800 355076 444806 355088
rect 450078 355076 450084 355088
rect 444800 355048 450084 355076
rect 444800 355036 444806 355048
rect 450078 355036 450084 355048
rect 450136 355036 450142 355088
rect 371510 354764 371516 354816
rect 371568 354804 371574 354816
rect 376846 354804 376852 354816
rect 371568 354776 376852 354804
rect 371568 354764 371574 354776
rect 376846 354764 376852 354776
rect 376904 354764 376910 354816
rect 371602 354696 371608 354748
rect 371660 354736 371666 354748
rect 380894 354736 380900 354748
rect 371660 354708 380900 354736
rect 371660 354696 371666 354708
rect 380894 354696 380900 354708
rect 380952 354696 380958 354748
rect 371970 353948 371976 354000
rect 372028 353988 372034 354000
rect 383746 353988 383752 354000
rect 372028 353960 383752 353988
rect 372028 353948 372034 353960
rect 383746 353948 383752 353960
rect 383804 353948 383810 354000
rect 371326 353336 371332 353388
rect 371384 353376 371390 353388
rect 375466 353376 375472 353388
rect 371384 353348 375472 353376
rect 371384 353336 371390 353348
rect 375466 353336 375472 353348
rect 375524 353336 375530 353388
rect 371694 353268 371700 353320
rect 371752 353308 371758 353320
rect 374086 353308 374092 353320
rect 371752 353280 374092 353308
rect 371752 353268 371758 353280
rect 374086 353268 374092 353280
rect 374144 353268 374150 353320
rect 372154 352588 372160 352640
rect 372212 352628 372218 352640
rect 378410 352628 378416 352640
rect 372212 352600 378416 352628
rect 372212 352588 372218 352600
rect 378410 352588 378416 352600
rect 378468 352588 378474 352640
rect 372338 352520 372344 352572
rect 372396 352560 372402 352572
rect 379606 352560 379612 352572
rect 372396 352532 379612 352560
rect 372396 352520 372402 352532
rect 379606 352520 379612 352532
rect 379664 352520 379670 352572
rect 444742 352452 444748 352504
rect 444800 352492 444806 352504
rect 448698 352492 448704 352504
rect 444800 352464 448704 352492
rect 444800 352452 444806 352464
rect 448698 352452 448704 352464
rect 448756 352452 448762 352504
rect 444466 351976 444472 352028
rect 444524 352016 444530 352028
rect 447226 352016 447232 352028
rect 444524 351988 447232 352016
rect 444524 351976 444530 351988
rect 447226 351976 447232 351988
rect 447284 351976 447290 352028
rect 371602 349256 371608 349308
rect 371660 349296 371666 349308
rect 373994 349296 374000 349308
rect 371660 349268 374000 349296
rect 371660 349256 371666 349268
rect 373994 349256 374000 349268
rect 374052 349256 374058 349308
rect 371602 348168 371608 348220
rect 371660 348208 371666 348220
rect 374362 348208 374368 348220
rect 371660 348180 374368 348208
rect 371660 348168 371666 348180
rect 374362 348168 374368 348180
rect 374420 348168 374426 348220
rect 445662 347760 445668 347812
rect 445720 347800 445726 347812
rect 454218 347800 454224 347812
rect 445720 347772 454224 347800
rect 445720 347760 445726 347772
rect 454218 347760 454224 347772
rect 454276 347760 454282 347812
rect 444650 346400 444656 346452
rect 444708 346440 444714 346452
rect 447502 346440 447508 346452
rect 444708 346412 447508 346440
rect 444708 346400 444714 346412
rect 447502 346400 447508 346412
rect 447560 346400 447566 346452
rect 445294 345108 445300 345160
rect 445352 345148 445358 345160
rect 452838 345148 452844 345160
rect 445352 345120 452844 345148
rect 445352 345108 445358 345120
rect 452838 345108 452844 345120
rect 452896 345108 452902 345160
rect 3326 345040 3332 345092
rect 3384 345080 3390 345092
rect 278774 345080 278780 345092
rect 3384 345052 278780 345080
rect 3384 345040 3390 345052
rect 278774 345040 278780 345052
rect 278832 345040 278838 345092
rect 445662 345040 445668 345092
rect 445720 345080 445726 345092
rect 456886 345080 456892 345092
rect 445720 345052 456892 345080
rect 445720 345040 445726 345052
rect 456886 345040 456892 345052
rect 456944 345040 456950 345092
rect 445662 343680 445668 343732
rect 445720 343720 445726 343732
rect 451274 343720 451280 343732
rect 445720 343692 451280 343720
rect 445720 343680 445726 343692
rect 451274 343680 451280 343692
rect 451332 343680 451338 343732
rect 445018 342252 445024 342304
rect 445076 342292 445082 342304
rect 458174 342292 458180 342304
rect 445076 342264 458180 342292
rect 445076 342252 445082 342264
rect 458174 342252 458180 342264
rect 458232 342252 458238 342304
rect 444558 341232 444564 341284
rect 444616 341272 444622 341284
rect 447410 341272 447416 341284
rect 444616 341244 447416 341272
rect 444616 341232 444622 341244
rect 447410 341232 447416 341244
rect 447468 341232 447474 341284
rect 369946 340552 369952 340604
rect 370004 340592 370010 340604
rect 370130 340592 370136 340604
rect 370004 340564 370136 340592
rect 370004 340552 370010 340564
rect 370130 340552 370136 340564
rect 370188 340552 370194 340604
rect 444558 340144 444564 340196
rect 444616 340184 444622 340196
rect 446030 340184 446036 340196
rect 444616 340156 446036 340184
rect 444616 340144 444622 340156
rect 446030 340144 446036 340156
rect 446088 340144 446094 340196
rect 300762 337424 300768 337476
rect 300820 337464 300826 337476
rect 438946 337464 438952 337476
rect 300820 337436 438952 337464
rect 300820 337424 300826 337436
rect 438946 337424 438952 337436
rect 439004 337424 439010 337476
rect 198550 337356 198556 337408
rect 198608 337396 198614 337408
rect 366910 337396 366916 337408
rect 198608 337368 366916 337396
rect 198608 337356 198614 337368
rect 366910 337356 366916 337368
rect 366968 337356 366974 337408
rect 441246 336744 441252 336796
rect 441304 336784 441310 336796
rect 441614 336784 441620 336796
rect 441304 336756 441620 336784
rect 441304 336744 441310 336756
rect 441614 336744 441620 336756
rect 441672 336744 441678 336796
rect 369026 335316 369032 335368
rect 369084 335356 369090 335368
rect 369302 335356 369308 335368
rect 369084 335328 369308 335356
rect 369084 335316 369090 335328
rect 369302 335316 369308 335328
rect 369360 335316 369366 335368
rect 137922 326340 137928 326392
rect 137980 326380 137986 326392
rect 255314 326380 255320 326392
rect 137980 326352 255320 326380
rect 137980 326340 137986 326352
rect 255314 326340 255320 326352
rect 255372 326340 255378 326392
rect 220722 324300 220728 324352
rect 220780 324340 220786 324352
rect 580166 324340 580172 324352
rect 220780 324312 580172 324340
rect 220780 324300 220786 324312
rect 580166 324300 580172 324312
rect 580224 324300 580230 324352
rect 3326 318792 3332 318844
rect 3384 318832 3390 318844
rect 280890 318832 280896 318844
rect 3384 318804 280896 318832
rect 3384 318792 3390 318804
rect 280890 318792 280896 318804
rect 280948 318792 280954 318844
rect 220630 311856 220636 311908
rect 220688 311896 220694 311908
rect 580166 311896 580172 311908
rect 220688 311868 580172 311896
rect 220688 311856 220694 311868
rect 580166 311856 580172 311868
rect 580224 311856 580230 311908
rect 245470 309748 245476 309800
rect 245528 309788 245534 309800
rect 396718 309788 396724 309800
rect 245528 309760 396724 309788
rect 245528 309748 245534 309760
rect 396718 309748 396724 309760
rect 396776 309748 396782 309800
rect 3418 308388 3424 308440
rect 3476 308428 3482 308440
rect 263226 308428 263232 308440
rect 3476 308400 263232 308428
rect 3476 308388 3482 308400
rect 263226 308388 263232 308400
rect 263284 308388 263290 308440
rect 253198 307504 253204 307556
rect 253256 307544 253262 307556
rect 280338 307544 280344 307556
rect 253256 307516 280344 307544
rect 253256 307504 253262 307516
rect 280338 307504 280344 307516
rect 280396 307504 280402 307556
rect 217318 307436 217324 307488
rect 217376 307476 217382 307488
rect 267274 307476 267280 307488
rect 217376 307448 267280 307476
rect 217376 307436 217382 307448
rect 267274 307436 267280 307448
rect 267332 307436 267338 307488
rect 215938 307368 215944 307420
rect 215996 307408 216002 307420
rect 269942 307408 269948 307420
rect 215996 307380 269948 307408
rect 215996 307368 216002 307380
rect 269942 307368 269948 307380
rect 270000 307368 270006 307420
rect 213178 307300 213184 307352
rect 213236 307340 213242 307352
rect 277762 307340 277768 307352
rect 213236 307312 277768 307340
rect 213236 307300 213242 307312
rect 277762 307300 277768 307312
rect 277820 307300 277826 307352
rect 249426 307232 249432 307284
rect 249484 307272 249490 307284
rect 347038 307272 347044 307284
rect 249484 307244 347044 307272
rect 249484 307232 249490 307244
rect 347038 307232 347044 307244
rect 347096 307232 347102 307284
rect 89622 307164 89628 307216
rect 89680 307204 89686 307216
rect 256234 307204 256240 307216
rect 89680 307176 256240 307204
rect 89680 307164 89686 307176
rect 256234 307164 256240 307176
rect 256292 307164 256298 307216
rect 8202 307096 8208 307148
rect 8260 307136 8266 307148
rect 258074 307136 258080 307148
rect 8260 307108 258080 307136
rect 8260 307096 8266 307108
rect 258074 307096 258080 307108
rect 258132 307096 258138 307148
rect 222930 307028 222936 307080
rect 222988 307068 222994 307080
rect 582466 307068 582472 307080
rect 222988 307040 582472 307068
rect 222988 307028 222994 307040
rect 582466 307028 582472 307040
rect 582524 307028 582530 307080
rect 222838 306076 222844 306128
rect 222896 306116 222902 306128
rect 254302 306116 254308 306128
rect 222896 306088 254308 306116
rect 222896 306076 222902 306088
rect 254302 306076 254308 306088
rect 254360 306076 254366 306128
rect 214558 306008 214564 306060
rect 214616 306048 214622 306060
rect 275094 306048 275100 306060
rect 214616 306020 275100 306048
rect 214616 306008 214622 306020
rect 275094 306008 275100 306020
rect 275152 306008 275158 306060
rect 248414 305940 248420 305992
rect 248472 305980 248478 305992
rect 331214 305980 331220 305992
rect 248472 305952 331220 305980
rect 248472 305940 248478 305952
rect 331214 305940 331220 305952
rect 331272 305940 331278 305992
rect 155218 305872 155224 305924
rect 155276 305912 155282 305924
rect 256878 305912 256884 305924
rect 155276 305884 256884 305912
rect 155276 305872 155282 305884
rect 256878 305872 256884 305884
rect 256936 305872 256942 305924
rect 41322 305804 41328 305856
rect 41380 305844 41386 305856
rect 260374 305844 260380 305856
rect 41380 305816 260380 305844
rect 41380 305804 41386 305816
rect 260374 305804 260380 305816
rect 260432 305804 260438 305856
rect 240318 305736 240324 305788
rect 240376 305776 240382 305788
rect 479518 305776 479524 305788
rect 240376 305748 479524 305776
rect 240376 305736 240382 305748
rect 479518 305736 479524 305748
rect 479576 305736 479582 305788
rect 222102 305668 222108 305720
rect 222160 305708 222166 305720
rect 582374 305708 582380 305720
rect 222160 305680 582380 305708
rect 222160 305668 222166 305680
rect 582374 305668 582380 305680
rect 582432 305668 582438 305720
rect 221182 305600 221188 305652
rect 221240 305640 221246 305652
rect 582558 305640 582564 305652
rect 221240 305612 582564 305640
rect 221240 305600 221246 305612
rect 582558 305600 582564 305612
rect 582616 305600 582622 305652
rect 3234 304988 3240 305040
rect 3292 305028 3298 305040
rect 282822 305028 282828 305040
rect 3292 305000 282828 305028
rect 3292 304988 3298 305000
rect 282822 304988 282828 305000
rect 282880 304988 282886 305040
rect 242158 304784 242164 304836
rect 242216 304824 242222 304836
rect 252554 304824 252560 304836
rect 242216 304796 252560 304824
rect 242216 304784 242222 304796
rect 252554 304784 252560 304796
rect 252612 304784 252618 304836
rect 249886 304716 249892 304768
rect 249944 304756 249950 304768
rect 299474 304756 299480 304768
rect 249944 304728 299480 304756
rect 249944 304716 249950 304728
rect 299474 304716 299480 304728
rect 299532 304716 299538 304768
rect 202782 304648 202788 304700
rect 202840 304688 202846 304700
rect 251818 304688 251824 304700
rect 202840 304660 251824 304688
rect 202840 304648 202846 304660
rect 251818 304648 251824 304660
rect 251876 304648 251882 304700
rect 171042 304580 171048 304632
rect 171100 304620 171106 304632
rect 255130 304620 255136 304632
rect 171100 304592 255136 304620
rect 171100 304580 171106 304592
rect 255130 304580 255136 304592
rect 255188 304580 255194 304632
rect 247310 304512 247316 304564
rect 247368 304552 247374 304564
rect 359458 304552 359464 304564
rect 247368 304524 359464 304552
rect 247368 304512 247374 304524
rect 359458 304512 359464 304524
rect 359516 304512 359522 304564
rect 106182 304444 106188 304496
rect 106240 304484 106246 304496
rect 257706 304484 257712 304496
rect 106240 304456 257712 304484
rect 106240 304444 106246 304456
rect 257706 304444 257712 304456
rect 257764 304444 257770 304496
rect 244734 304376 244740 304428
rect 244792 304416 244798 304428
rect 429194 304416 429200 304428
rect 244792 304388 429200 304416
rect 244792 304376 244798 304388
rect 429194 304376 429200 304388
rect 429252 304376 429258 304428
rect 242066 304308 242072 304360
rect 242124 304348 242130 304360
rect 494054 304348 494060 304360
rect 242124 304320 494060 304348
rect 242124 304308 242130 304320
rect 494054 304308 494060 304320
rect 494112 304308 494118 304360
rect 239490 304240 239496 304292
rect 239548 304280 239554 304292
rect 558914 304280 558920 304292
rect 239548 304252 558920 304280
rect 239548 304240 239554 304252
rect 558914 304240 558920 304252
rect 558972 304240 558978 304292
rect 128998 303696 129004 303748
rect 129056 303736 129062 303748
rect 297726 303736 297732 303748
rect 129056 303708 297732 303736
rect 129056 303696 129062 303708
rect 297726 303696 297732 303708
rect 297784 303696 297790 303748
rect 202046 303628 202052 303680
rect 202104 303668 202110 303680
rect 582466 303668 582472 303680
rect 202104 303640 582472 303668
rect 202104 303628 202110 303640
rect 582466 303628 582472 303640
rect 582524 303628 582530 303680
rect 242986 303492 242992 303544
rect 243044 303532 243050 303544
rect 249058 303532 249064 303544
rect 243044 303504 249064 303532
rect 243044 303492 243050 303504
rect 249058 303492 249064 303504
rect 249116 303492 249122 303544
rect 256234 303288 256240 303340
rect 256292 303328 256298 303340
rect 259454 303328 259460 303340
rect 256292 303300 259460 303328
rect 256292 303288 256298 303300
rect 259454 303288 259460 303300
rect 259512 303288 259518 303340
rect 209866 303084 209872 303136
rect 209924 303124 209930 303136
rect 548518 303124 548524 303136
rect 209924 303096 548524 303124
rect 209924 303084 209930 303096
rect 548518 303084 548524 303096
rect 548576 303084 548582 303136
rect 258074 303016 258080 303068
rect 258132 303056 258138 303068
rect 261202 303056 261208 303068
rect 258132 303028 261208 303056
rect 258132 303016 258138 303028
rect 261202 303016 261208 303028
rect 261260 303016 261266 303068
rect 237742 302948 237748 303000
rect 237800 302988 237806 303000
rect 238662 302988 238668 303000
rect 237800 302960 238668 302988
rect 237800 302948 237806 302960
rect 238662 302948 238668 302960
rect 238720 302948 238726 303000
rect 251634 302948 251640 303000
rect 251692 302988 251698 303000
rect 252462 302988 252468 303000
rect 251692 302960 252468 302988
rect 251692 302948 251698 302960
rect 252462 302948 252468 302960
rect 252520 302948 252526 303000
rect 260098 302948 260104 303000
rect 260156 302988 260162 303000
rect 262122 302988 262128 303000
rect 260156 302960 262128 302988
rect 260156 302948 260162 302960
rect 262122 302948 262128 302960
rect 262180 302948 262186 303000
rect 263226 302948 263232 303000
rect 263284 302988 263290 303000
rect 264698 302988 264704 303000
rect 263284 302960 264704 302988
rect 263284 302948 263290 302960
rect 264698 302948 264704 302960
rect 264756 302948 264762 303000
rect 269758 302948 269764 303000
rect 269816 302988 269822 303000
rect 272518 302988 272524 303000
rect 269816 302960 272524 302988
rect 269816 302948 269822 302960
rect 272518 302948 272524 302960
rect 272576 302948 272582 303000
rect 211614 302880 211620 302932
rect 211672 302920 211678 302932
rect 311158 302920 311164 302932
rect 211672 302892 311164 302920
rect 211672 302880 211678 302892
rect 311158 302880 311164 302892
rect 311216 302880 311222 302932
rect 209038 302812 209044 302864
rect 209096 302852 209102 302864
rect 309778 302852 309784 302864
rect 209096 302824 309784 302852
rect 209096 302812 209102 302824
rect 309778 302812 309784 302824
rect 309836 302812 309842 302864
rect 180058 302744 180064 302796
rect 180116 302784 180122 302796
rect 285582 302784 285588 302796
rect 180116 302756 285588 302784
rect 180116 302744 180122 302756
rect 285582 302744 285588 302756
rect 285640 302744 285646 302796
rect 299474 302744 299480 302796
rect 299532 302784 299538 302796
rect 300762 302784 300768 302796
rect 299532 302756 300768 302784
rect 299532 302744 299538 302756
rect 300762 302744 300768 302756
rect 300820 302744 300826 302796
rect 212534 302676 212540 302728
rect 212592 302716 212598 302728
rect 318058 302716 318064 302728
rect 212592 302688 318064 302716
rect 212592 302676 212598 302688
rect 318058 302676 318064 302688
rect 318116 302676 318122 302728
rect 204714 302608 204720 302660
rect 204772 302648 204778 302660
rect 313918 302648 313924 302660
rect 204772 302620 313924 302648
rect 204772 302608 204778 302620
rect 313918 302608 313924 302620
rect 313976 302608 313982 302660
rect 207290 302540 207296 302592
rect 207348 302580 207354 302592
rect 316678 302580 316684 302592
rect 207348 302552 316684 302580
rect 207348 302540 207354 302552
rect 316678 302540 316684 302552
rect 316736 302540 316742 302592
rect 166258 302472 166264 302524
rect 166316 302512 166322 302524
rect 288158 302512 288164 302524
rect 166316 302484 288164 302512
rect 166316 302472 166322 302484
rect 288158 302472 288164 302484
rect 288216 302472 288222 302524
rect 148318 302404 148324 302456
rect 148376 302444 148382 302456
rect 290826 302444 290832 302456
rect 148376 302416 290832 302444
rect 148376 302404 148382 302416
rect 290826 302404 290832 302416
rect 290884 302404 290890 302456
rect 215110 302336 215116 302388
rect 215168 302376 215174 302388
rect 443638 302376 443644 302388
rect 215168 302348 443644 302376
rect 215168 302336 215174 302348
rect 443638 302336 443644 302348
rect 443696 302336 443702 302388
rect 14458 302268 14464 302320
rect 14516 302308 14522 302320
rect 293402 302308 293408 302320
rect 14516 302280 293408 302308
rect 14516 302268 14522 302280
rect 293402 302268 293408 302280
rect 293460 302268 293466 302320
rect 251818 302200 251824 302252
rect 251876 302240 251882 302252
rect 253382 302240 253388 302252
rect 251876 302212 253388 302240
rect 251876 302200 251882 302212
rect 253382 302200 253388 302212
rect 253440 302200 253446 302252
rect 285674 302200 285680 302252
rect 285732 302240 285738 302252
rect 289906 302240 289912 302252
rect 285732 302212 289912 302240
rect 285732 302200 285738 302212
rect 289906 302200 289912 302212
rect 289964 302200 289970 302252
rect 223850 302064 223856 302116
rect 223908 302104 223914 302116
rect 224770 302104 224776 302116
rect 223908 302076 224776 302104
rect 223908 302064 223914 302076
rect 224770 302064 224776 302076
rect 224828 302064 224834 302116
rect 228174 302064 228180 302116
rect 228232 302104 228238 302116
rect 228910 302104 228916 302116
rect 228232 302076 228916 302104
rect 228232 302064 228238 302076
rect 228910 302064 228916 302076
rect 228968 302064 228974 302116
rect 230750 302064 230756 302116
rect 230808 302104 230814 302116
rect 231670 302104 231676 302116
rect 230808 302076 231676 302104
rect 230808 302064 230814 302076
rect 231670 302064 231676 302076
rect 231728 302064 231734 302116
rect 233418 302064 233424 302116
rect 233476 302104 233482 302116
rect 234430 302104 234436 302116
rect 233476 302076 234436 302104
rect 233476 302064 233482 302076
rect 234430 302064 234436 302076
rect 234488 302064 234494 302116
rect 235166 302064 235172 302116
rect 235224 302104 235230 302116
rect 235902 302104 235908 302116
rect 235224 302076 235908 302104
rect 235224 302064 235230 302076
rect 235902 302064 235908 302076
rect 235960 302064 235966 302116
rect 235994 302064 236000 302116
rect 236052 302104 236058 302116
rect 237190 302104 237196 302116
rect 236052 302076 237196 302104
rect 236052 302064 236058 302076
rect 237190 302064 237196 302076
rect 237248 302064 237254 302116
rect 216030 301588 216036 301640
rect 216088 301628 216094 301640
rect 301498 301628 301504 301640
rect 216088 301600 301504 301628
rect 216088 301588 216094 301600
rect 301498 301588 301504 301600
rect 301556 301588 301562 301640
rect 199378 301520 199384 301572
rect 199436 301560 199442 301572
rect 286410 301560 286416 301572
rect 199436 301532 286416 301560
rect 199436 301520 199442 301532
rect 286410 301520 286416 301532
rect 286468 301520 286474 301572
rect 206462 301452 206468 301504
rect 206520 301492 206526 301504
rect 307018 301492 307024 301504
rect 206520 301464 307024 301492
rect 206520 301452 206526 301464
rect 307018 301452 307024 301464
rect 307076 301452 307082 301504
rect 174538 301384 174544 301436
rect 174596 301424 174602 301436
rect 284662 301424 284668 301436
rect 174596 301396 284668 301424
rect 174596 301384 174602 301396
rect 284662 301384 284668 301396
rect 284720 301384 284726 301436
rect 152458 301316 152464 301368
rect 152516 301356 152522 301368
rect 292482 301356 292488 301368
rect 152516 301328 292488 301356
rect 152516 301316 152522 301328
rect 292482 301316 292488 301328
rect 292540 301316 292546 301368
rect 156598 301248 156604 301300
rect 156656 301288 156662 301300
rect 296898 301288 296904 301300
rect 156656 301260 296904 301288
rect 156656 301248 156662 301260
rect 296898 301248 296904 301260
rect 296956 301248 296962 301300
rect 144178 301180 144184 301232
rect 144236 301220 144242 301232
rect 298646 301220 298652 301232
rect 144236 301192 298652 301220
rect 144236 301180 144242 301192
rect 298646 301180 298652 301192
rect 298704 301180 298710 301232
rect 90358 301112 90364 301164
rect 90416 301152 90422 301164
rect 283834 301152 283840 301164
rect 90416 301124 283840 301152
rect 90416 301112 90422 301124
rect 283834 301112 283840 301124
rect 283892 301112 283898 301164
rect 210786 301044 210792 301096
rect 210844 301084 210850 301096
rect 582926 301084 582932 301096
rect 210844 301056 582932 301084
rect 210844 301044 210850 301056
rect 582926 301044 582932 301056
rect 582984 301044 582990 301096
rect 202966 300976 202972 301028
rect 203024 301016 203030 301028
rect 582650 301016 582656 301028
rect 203024 300988 582656 301016
rect 203024 300976 203030 300988
rect 582650 300976 582656 300988
rect 582708 300976 582714 301028
rect 200390 300908 200396 300960
rect 200448 300948 200454 300960
rect 582374 300948 582380 300960
rect 200448 300920 582380 300948
rect 200448 300908 200454 300920
rect 582374 300908 582380 300920
rect 582432 300908 582438 300960
rect 201218 300840 201224 300892
rect 201276 300880 201282 300892
rect 583110 300880 583116 300892
rect 201276 300852 583116 300880
rect 201276 300840 201282 300852
rect 583110 300840 583116 300852
rect 583168 300840 583174 300892
rect 213362 300296 213368 300348
rect 213420 300336 213426 300348
rect 219342 300336 219348 300348
rect 213420 300308 219348 300336
rect 213420 300296 213426 300308
rect 219342 300296 219348 300308
rect 219400 300296 219406 300348
rect 219434 300296 219440 300348
rect 219492 300336 219498 300348
rect 220722 300336 220728 300348
rect 219492 300308 220728 300336
rect 219492 300296 219498 300308
rect 220722 300296 220728 300308
rect 220780 300296 220786 300348
rect 226426 300296 226432 300348
rect 226484 300336 226490 300348
rect 227530 300336 227536 300348
rect 226484 300308 227536 300336
rect 226484 300296 226490 300308
rect 227530 300296 227536 300308
rect 227588 300296 227594 300348
rect 196618 300228 196624 300280
rect 196676 300268 196682 300280
rect 282086 300268 282092 300280
rect 196676 300240 282092 300268
rect 196676 300228 196682 300240
rect 282086 300228 282092 300240
rect 282144 300228 282150 300280
rect 203794 300160 203800 300212
rect 203852 300200 203858 300212
rect 305638 300200 305644 300212
rect 203852 300172 305644 300200
rect 203852 300160 203858 300172
rect 305638 300160 305644 300172
rect 305696 300160 305702 300212
rect 159358 300092 159364 300144
rect 159416 300132 159422 300144
rect 291654 300132 291660 300144
rect 159416 300104 291660 300132
rect 159416 300092 159422 300104
rect 291654 300092 291660 300104
rect 291712 300092 291718 300144
rect 155218 300024 155224 300076
rect 155276 300064 155282 300076
rect 287146 300064 287152 300076
rect 155276 300036 287152 300064
rect 155276 300024 155282 300036
rect 287146 300024 287152 300036
rect 287204 300024 287210 300076
rect 157978 299956 157984 300008
rect 158036 299996 158042 300008
rect 293954 299996 293960 300008
rect 158036 299968 293960 299996
rect 158036 299956 158042 299968
rect 293954 299956 293960 299968
rect 294012 299956 294018 300008
rect 151078 299888 151084 299940
rect 151136 299928 151142 299940
rect 294782 299928 294788 299940
rect 151136 299900 294788 299928
rect 151136 299888 151142 299900
rect 294782 299888 294788 299900
rect 294840 299888 294846 299940
rect 146938 299820 146944 299872
rect 146996 299860 147002 299872
rect 295702 299860 295708 299872
rect 146996 299832 295708 299860
rect 146996 299820 147002 299832
rect 295702 299820 295708 299832
rect 295760 299820 295766 299872
rect 88978 299752 88984 299804
rect 89036 299792 89042 299804
rect 288710 299792 288716 299804
rect 89036 299764 288716 299792
rect 89036 299752 89042 299764
rect 288710 299752 288716 299764
rect 288768 299752 288774 299804
rect 218882 299684 218888 299736
rect 218940 299724 218946 299736
rect 579890 299724 579896 299736
rect 218940 299696 579896 299724
rect 218940 299684 218946 299696
rect 579890 299684 579896 299696
rect 579948 299684 579954 299736
rect 219342 299616 219348 299668
rect 219400 299656 219406 299668
rect 583018 299656 583024 299668
rect 219400 299628 583024 299656
rect 219400 299616 219406 299628
rect 583018 299616 583024 299628
rect 583076 299616 583082 299668
rect 208302 299548 208308 299600
rect 208360 299588 208366 299600
rect 582834 299588 582840 299600
rect 208360 299560 582840 299588
rect 208360 299548 208366 299560
rect 582834 299548 582840 299560
rect 582892 299548 582898 299600
rect 205634 299480 205640 299532
rect 205692 299520 205698 299532
rect 582558 299520 582564 299532
rect 205692 299492 582564 299520
rect 205692 299480 205698 299492
rect 582558 299480 582564 299492
rect 582616 299480 582622 299532
rect 216766 299412 216772 299464
rect 216824 299452 216830 299464
rect 216824 299424 231854 299452
rect 216824 299412 216830 299424
rect 214650 299344 214656 299396
rect 214708 299384 214714 299396
rect 214708 299356 217916 299384
rect 214708 299344 214714 299356
rect 216766 299316 216772 299328
rect 216646 299288 216772 299316
rect 216646 299044 216674 299288
rect 216766 299276 216772 299288
rect 216824 299276 216830 299328
rect 217410 299276 217416 299328
rect 217468 299276 217474 299328
rect 217686 299276 217692 299328
rect 217744 299276 217750 299328
rect 212506 299016 216674 299044
rect 3418 298800 3424 298852
rect 3476 298840 3482 298852
rect 3476 298812 200114 298840
rect 3476 298800 3482 298812
rect 200086 298772 200114 298812
rect 212506 298772 212534 299016
rect 200086 298744 212534 298772
rect 208366 298676 209774 298704
rect 208366 298432 208394 298676
rect 200086 298404 208394 298432
rect 199838 298256 199844 298308
rect 199896 298296 199902 298308
rect 200086 298296 200114 298404
rect 199896 298268 200114 298296
rect 199896 298256 199902 298268
rect 209746 298024 209774 298676
rect 217428 298024 217456 299276
rect 217704 298160 217732 299276
rect 217888 298636 217916 299356
rect 217962 299344 217968 299396
rect 218020 299344 218026 299396
rect 217980 299248 218008 299344
rect 218054 299276 218060 299328
rect 218112 299316 218118 299328
rect 218112 299288 224954 299316
rect 218112 299276 218118 299288
rect 217980 299220 222194 299248
rect 222166 298636 222194 299220
rect 224926 298908 224954 299288
rect 231826 299180 231854 299424
rect 285674 299316 285680 299328
rect 277366 299288 285680 299316
rect 231826 299152 237374 299180
rect 224926 298880 231854 298908
rect 231826 298772 231854 298880
rect 237346 298840 237374 299152
rect 277366 298840 277394 299288
rect 285674 299276 285680 299288
rect 285732 299276 285738 299328
rect 237346 298812 277394 298840
rect 580258 298772 580264 298784
rect 231826 298744 580264 298772
rect 580258 298732 580264 298744
rect 580316 298732 580322 298784
rect 223546 298676 226334 298704
rect 223546 298636 223574 298676
rect 217888 298608 220952 298636
rect 222166 298608 223574 298636
rect 226306 298636 226334 298676
rect 226306 298608 235994 298636
rect 220924 298500 220952 298608
rect 235966 298568 235994 298608
rect 235966 298540 237374 298568
rect 237346 298500 237374 298540
rect 238726 298540 240134 298568
rect 238726 298500 238754 298540
rect 220924 298472 223252 298500
rect 237346 298472 238754 298500
rect 240106 298500 240134 298540
rect 240106 298472 241514 298500
rect 223224 298296 223252 298472
rect 224926 298404 238754 298432
rect 224926 298364 224954 298404
rect 223546 298336 224954 298364
rect 223546 298296 223574 298336
rect 223224 298268 223574 298296
rect 238726 298296 238754 298404
rect 241486 298296 241514 298472
rect 302786 298324 302792 298376
rect 302844 298364 302850 298376
rect 323578 298364 323584 298376
rect 302844 298336 323584 298364
rect 302844 298324 302850 298336
rect 323578 298324 323584 298336
rect 323636 298324 323642 298376
rect 359458 298296 359464 298308
rect 238726 298268 240134 298296
rect 241486 298268 359464 298296
rect 240106 298228 240134 298268
rect 359458 298256 359464 298268
rect 359516 298256 359522 298308
rect 312538 298228 312544 298240
rect 240106 298200 312544 298228
rect 312538 298188 312544 298200
rect 312596 298188 312602 298240
rect 442258 298160 442264 298172
rect 217704 298132 222194 298160
rect 222166 298092 222194 298132
rect 223546 298132 442264 298160
rect 223546 298092 223574 298132
rect 442258 298120 442264 298132
rect 442316 298120 442322 298172
rect 222166 298064 223574 298092
rect 209746 297996 217456 298024
rect 436094 297644 436100 297696
rect 436152 297684 436158 297696
rect 442994 297684 443000 297696
rect 436152 297656 443000 297684
rect 436152 297644 436158 297656
rect 442994 297644 443000 297656
rect 443052 297644 443058 297696
rect 434714 297576 434720 297628
rect 434772 297616 434778 297628
rect 441706 297616 441712 297628
rect 434772 297588 441712 297616
rect 434772 297576 434778 297588
rect 441706 297576 441712 297588
rect 441764 297576 441770 297628
rect 373258 297440 373264 297492
rect 373316 297480 373322 297492
rect 379514 297480 379520 297492
rect 373316 297452 379520 297480
rect 373316 297440 373322 297452
rect 379514 297440 379520 297452
rect 379572 297440 379578 297492
rect 374178 297372 374184 297424
rect 374236 297412 374242 297424
rect 385126 297412 385132 297424
rect 374236 297384 385132 297412
rect 374236 297372 374242 297384
rect 385126 297372 385132 297384
rect 385184 297372 385190 297424
rect 450170 297372 450176 297424
rect 450228 297412 450234 297424
rect 454034 297412 454040 297424
rect 450228 297384 454040 297412
rect 450228 297372 450234 297384
rect 454034 297372 454040 297384
rect 454092 297372 454098 297424
rect 445662 297032 445668 297084
rect 445720 297072 445726 297084
rect 450170 297072 450176 297084
rect 445720 297044 450176 297072
rect 445720 297032 445726 297044
rect 450170 297032 450176 297044
rect 450228 297032 450234 297084
rect 302970 296760 302976 296812
rect 303028 296800 303034 296812
rect 369486 296800 369492 296812
rect 303028 296772 369492 296800
rect 303028 296760 303034 296772
rect 369486 296760 369492 296772
rect 369544 296800 369550 296812
rect 373258 296800 373264 296812
rect 369544 296772 373264 296800
rect 369544 296760 369550 296772
rect 373258 296760 373264 296772
rect 373316 296760 373322 296812
rect 302878 296692 302884 296744
rect 302936 296732 302942 296744
rect 369394 296732 369400 296744
rect 302936 296704 369400 296732
rect 302936 296692 302942 296704
rect 369394 296692 369400 296704
rect 369452 296732 369458 296744
rect 374178 296732 374184 296744
rect 369452 296704 374184 296732
rect 369452 296692 369458 296704
rect 374178 296692 374184 296704
rect 374236 296692 374242 296744
rect 370130 296080 370136 296132
rect 370188 296120 370194 296132
rect 378134 296120 378140 296132
rect 370188 296092 378140 296120
rect 370188 296080 370194 296092
rect 378134 296080 378140 296092
rect 378192 296080 378198 296132
rect 372890 296012 372896 296064
rect 372948 296052 372954 296064
rect 379514 296052 379520 296064
rect 372948 296024 379520 296052
rect 372948 296012 372954 296024
rect 379514 296012 379520 296024
rect 379572 296012 379578 296064
rect 369394 295944 369400 295996
rect 369452 295944 369458 295996
rect 383654 295984 383660 295996
rect 373966 295956 383660 295984
rect 327718 295876 327724 295928
rect 327776 295916 327782 295928
rect 369412 295916 369440 295944
rect 327776 295888 369440 295916
rect 327776 295876 327782 295888
rect 352558 295808 352564 295860
rect 352616 295848 352622 295860
rect 369394 295848 369400 295860
rect 352616 295820 369400 295848
rect 352616 295808 352622 295820
rect 369394 295808 369400 295820
rect 369452 295848 369458 295860
rect 373966 295848 373994 295956
rect 383654 295944 383660 295956
rect 383712 295944 383718 295996
rect 445754 295944 445760 295996
rect 445812 295984 445818 295996
rect 458266 295984 458272 295996
rect 445812 295956 458272 295984
rect 445812 295944 445818 295956
rect 458266 295944 458272 295956
rect 458324 295944 458330 295996
rect 369452 295820 373994 295848
rect 369452 295808 369458 295820
rect 302786 295332 302792 295384
rect 302844 295372 302850 295384
rect 322198 295372 322204 295384
rect 302844 295344 322204 295372
rect 302844 295332 302850 295344
rect 322198 295332 322204 295344
rect 322256 295332 322262 295384
rect 371234 295264 371240 295316
rect 371292 295304 371298 295316
rect 376938 295304 376944 295316
rect 371292 295276 376944 295304
rect 371292 295264 371298 295276
rect 376938 295264 376944 295276
rect 376996 295304 377002 295316
rect 385402 295304 385408 295316
rect 376996 295276 385408 295304
rect 376996 295264 377002 295276
rect 385402 295264 385408 295276
rect 385460 295264 385466 295316
rect 445662 295264 445668 295316
rect 445720 295304 445726 295316
rect 449894 295304 449900 295316
rect 445720 295276 449900 295304
rect 445720 295264 445726 295276
rect 449894 295264 449900 295276
rect 449952 295264 449958 295316
rect 449894 294652 449900 294704
rect 449952 294692 449958 294704
rect 454034 294692 454040 294704
rect 449952 294664 454040 294692
rect 449952 294652 449958 294664
rect 454034 294652 454040 294664
rect 454092 294652 454098 294704
rect 371694 294584 371700 294636
rect 371752 294624 371758 294636
rect 382274 294624 382280 294636
rect 371752 294596 382280 294624
rect 371752 294584 371758 294596
rect 382274 294584 382280 294596
rect 382332 294584 382338 294636
rect 445662 294584 445668 294636
rect 445720 294624 445726 294636
rect 448790 294624 448796 294636
rect 445720 294596 448796 294624
rect 445720 294584 445726 294596
rect 448790 294584 448796 294596
rect 448848 294624 448854 294636
rect 456794 294624 456800 294636
rect 448848 294596 456800 294624
rect 448848 294584 448854 294596
rect 456794 294584 456800 294596
rect 456852 294584 456858 294636
rect 170398 293972 170404 294024
rect 170456 294012 170462 294024
rect 197906 294012 197912 294024
rect 170456 293984 197912 294012
rect 170456 293972 170462 293984
rect 197906 293972 197912 293984
rect 197964 293972 197970 294024
rect 371694 293972 371700 294024
rect 371752 294012 371758 294024
rect 376938 294012 376944 294024
rect 371752 293984 376944 294012
rect 371752 293972 371758 293984
rect 376938 293972 376944 293984
rect 376996 294012 377002 294024
rect 385034 294012 385040 294024
rect 376996 293984 385040 294012
rect 376996 293972 377002 293984
rect 385034 293972 385040 293984
rect 385092 293972 385098 294024
rect 3050 293904 3056 293956
rect 3108 293944 3114 293956
rect 196618 293944 196624 293956
rect 3108 293916 196624 293944
rect 3108 293904 3114 293916
rect 196618 293904 196624 293916
rect 196676 293904 196682 293956
rect 373350 293904 373356 293956
rect 373408 293944 373414 293956
rect 375558 293944 375564 293956
rect 373408 293916 375564 293944
rect 373408 293904 373414 293916
rect 375558 293904 375564 293916
rect 375616 293904 375622 293956
rect 372154 293428 372160 293480
rect 372212 293468 372218 293480
rect 373350 293468 373356 293480
rect 372212 293440 373356 293468
rect 372212 293428 372218 293440
rect 373350 293428 373356 293440
rect 373408 293428 373414 293480
rect 371694 293224 371700 293276
rect 371752 293264 371758 293276
rect 376018 293264 376024 293276
rect 371752 293236 376024 293264
rect 371752 293224 371758 293236
rect 376018 293224 376024 293236
rect 376076 293264 376082 293276
rect 382366 293264 382372 293276
rect 376076 293236 382372 293264
rect 376076 293224 376082 293236
rect 382366 293224 382372 293236
rect 382424 293224 382430 293276
rect 445662 293224 445668 293276
rect 445720 293264 445726 293276
rect 452746 293264 452752 293276
rect 445720 293236 452752 293264
rect 445720 293224 445726 293236
rect 452746 293224 452752 293236
rect 452804 293264 452810 293276
rect 456794 293264 456800 293276
rect 452804 293236 456800 293264
rect 452804 293224 452810 293236
rect 456794 293224 456800 293236
rect 456852 293224 456858 293276
rect 371234 292408 371240 292460
rect 371292 292448 371298 292460
rect 378318 292448 378324 292460
rect 371292 292420 378324 292448
rect 371292 292408 371298 292420
rect 378318 292408 378324 292420
rect 378376 292408 378382 292460
rect 371694 292340 371700 292392
rect 371752 292380 371758 292392
rect 374178 292380 374184 292392
rect 371752 292352 374184 292380
rect 371752 292340 371758 292352
rect 374178 292340 374184 292352
rect 374236 292340 374242 292392
rect 378318 292000 378324 292052
rect 378376 292040 378382 292052
rect 382366 292040 382372 292052
rect 378376 292012 382372 292040
rect 378376 292000 378382 292012
rect 382366 292000 382372 292012
rect 382424 292000 382430 292052
rect 372154 291932 372160 291984
rect 372212 291972 372218 291984
rect 372706 291972 372712 291984
rect 372212 291944 372712 291972
rect 372212 291932 372218 291944
rect 372706 291932 372712 291944
rect 372764 291972 372770 291984
rect 378502 291972 378508 291984
rect 372764 291944 378508 291972
rect 372764 291932 372770 291944
rect 378502 291932 378508 291944
rect 378560 291932 378566 291984
rect 302234 291456 302240 291508
rect 302292 291496 302298 291508
rect 304258 291496 304264 291508
rect 302292 291468 304264 291496
rect 302292 291456 302298 291468
rect 304258 291456 304264 291468
rect 304316 291456 304322 291508
rect 175918 291184 175924 291236
rect 175976 291224 175982 291236
rect 197538 291224 197544 291236
rect 175976 291196 197544 291224
rect 175976 291184 175982 291196
rect 197538 291184 197544 291196
rect 197596 291184 197602 291236
rect 445662 291184 445668 291236
rect 445720 291224 445726 291236
rect 448606 291224 448612 291236
rect 445720 291196 448612 291224
rect 445720 291184 445726 291196
rect 448606 291184 448612 291196
rect 448664 291224 448670 291236
rect 452746 291224 452752 291236
rect 448664 291196 452752 291224
rect 448664 291184 448670 291196
rect 452746 291184 452752 291196
rect 452804 291184 452810 291236
rect 371234 290504 371240 290556
rect 371292 290544 371298 290556
rect 377030 290544 377036 290556
rect 371292 290516 377036 290544
rect 371292 290504 371298 290516
rect 377030 290504 377036 290516
rect 377088 290504 377094 290556
rect 371694 290436 371700 290488
rect 371752 290476 371758 290488
rect 380986 290476 380992 290488
rect 371752 290448 380992 290476
rect 371752 290436 371758 290448
rect 380986 290436 380992 290448
rect 381044 290436 381050 290488
rect 445754 290436 445760 290488
rect 445812 290476 445818 290488
rect 454126 290476 454132 290488
rect 445812 290448 454132 290476
rect 445812 290436 445818 290448
rect 454126 290436 454132 290448
rect 454184 290436 454190 290488
rect 371694 289552 371700 289604
rect 371752 289592 371758 289604
rect 375374 289592 375380 289604
rect 371752 289564 375380 289592
rect 371752 289552 371758 289564
rect 375374 289552 375380 289564
rect 375432 289592 375438 289604
rect 375558 289592 375564 289604
rect 375432 289564 375564 289592
rect 375432 289552 375438 289564
rect 375558 289552 375564 289564
rect 375616 289552 375622 289604
rect 445662 289144 445668 289196
rect 445720 289184 445726 289196
rect 449986 289184 449992 289196
rect 445720 289156 449992 289184
rect 445720 289144 445726 289156
rect 449986 289144 449992 289156
rect 450044 289184 450050 289196
rect 454126 289184 454132 289196
rect 450044 289156 454132 289184
rect 450044 289144 450050 289156
rect 454126 289144 454132 289156
rect 454184 289144 454190 289196
rect 371694 289076 371700 289128
rect 371752 289116 371758 289128
rect 378226 289116 378232 289128
rect 371752 289088 378232 289116
rect 371752 289076 371758 289088
rect 378226 289076 378232 289088
rect 378284 289076 378290 289128
rect 371694 288464 371700 288516
rect 371752 288504 371758 288516
rect 374454 288504 374460 288516
rect 371752 288476 374460 288504
rect 371752 288464 371758 288476
rect 374454 288464 374460 288476
rect 374512 288464 374518 288516
rect 302694 288396 302700 288448
rect 302752 288436 302758 288448
rect 320818 288436 320824 288448
rect 302752 288408 320824 288436
rect 302752 288396 302758 288408
rect 320818 288396 320824 288408
rect 320876 288396 320882 288448
rect 371694 288328 371700 288380
rect 371752 288368 371758 288380
rect 379606 288368 379612 288380
rect 371752 288340 379612 288368
rect 371752 288328 371758 288340
rect 379606 288328 379612 288340
rect 379664 288328 379670 288380
rect 371694 287648 371700 287700
rect 371752 287688 371758 287700
rect 378410 287688 378416 287700
rect 371752 287660 378416 287688
rect 371752 287648 371758 287660
rect 378410 287648 378416 287660
rect 378468 287648 378474 287700
rect 449986 287376 449992 287428
rect 450044 287416 450050 287428
rect 452654 287416 452660 287428
rect 450044 287388 452660 287416
rect 450044 287376 450050 287388
rect 452654 287376 452660 287388
rect 452712 287376 452718 287428
rect 445478 287240 445484 287292
rect 445536 287280 445542 287292
rect 445846 287280 445852 287292
rect 445536 287252 445852 287280
rect 445536 287240 445542 287252
rect 445846 287240 445852 287252
rect 445904 287280 445910 287292
rect 452654 287280 452660 287292
rect 445904 287252 452660 287280
rect 445904 287240 445910 287252
rect 452654 287240 452660 287252
rect 452712 287240 452718 287292
rect 445662 287104 445668 287156
rect 445720 287144 445726 287156
rect 449986 287144 449992 287156
rect 445720 287116 449992 287144
rect 445720 287104 445726 287116
rect 449986 287104 449992 287116
rect 450044 287104 450050 287156
rect 176010 287036 176016 287088
rect 176068 287076 176074 287088
rect 197538 287076 197544 287088
rect 176068 287048 197544 287076
rect 176068 287036 176074 287048
rect 197538 287036 197544 287048
rect 197596 287036 197602 287088
rect 379606 287036 379612 287088
rect 379664 287076 379670 287088
rect 385310 287076 385316 287088
rect 379664 287048 385316 287076
rect 379664 287036 379670 287048
rect 385310 287036 385316 287048
rect 385368 287036 385374 287088
rect 371694 286968 371700 287020
rect 371752 287008 371758 287020
rect 376754 287008 376760 287020
rect 371752 286980 376760 287008
rect 371752 286968 371758 286980
rect 376754 286968 376760 286980
rect 376812 286968 376818 287020
rect 371970 286628 371976 286680
rect 372028 286668 372034 286680
rect 372154 286668 372160 286680
rect 372028 286640 372160 286668
rect 372028 286628 372034 286640
rect 372154 286628 372160 286640
rect 372212 286628 372218 286680
rect 371602 286492 371608 286544
rect 371660 286532 371666 286544
rect 371970 286532 371976 286544
rect 371660 286504 371976 286532
rect 371660 286492 371666 286504
rect 371970 286492 371976 286504
rect 372028 286492 372034 286544
rect 371602 286356 371608 286408
rect 371660 286396 371666 286408
rect 374638 286396 374644 286408
rect 371660 286368 374644 286396
rect 371660 286356 371666 286368
rect 374638 286356 374644 286368
rect 374696 286396 374702 286408
rect 382550 286396 382556 286408
rect 374696 286368 382556 286396
rect 374696 286356 374702 286368
rect 382550 286356 382556 286368
rect 382608 286356 382614 286408
rect 371234 286288 371240 286340
rect 371292 286328 371298 286340
rect 383746 286328 383752 286340
rect 371292 286300 383752 286328
rect 371292 286288 371298 286300
rect 383746 286288 383752 286300
rect 383804 286288 383810 286340
rect 445662 285948 445668 286000
rect 445720 285988 445726 286000
rect 448514 285988 448520 286000
rect 445720 285960 448520 285988
rect 445720 285948 445726 285960
rect 448514 285948 448520 285960
rect 448572 285948 448578 286000
rect 302786 285676 302792 285728
rect 302844 285716 302850 285728
rect 324958 285716 324964 285728
rect 302844 285688 324964 285716
rect 302844 285676 302850 285688
rect 324958 285676 324964 285688
rect 325016 285676 325022 285728
rect 376754 285676 376760 285728
rect 376812 285716 376818 285728
rect 381262 285716 381268 285728
rect 376812 285688 381268 285716
rect 376812 285676 376818 285688
rect 381262 285676 381268 285688
rect 381320 285676 381326 285728
rect 371694 285608 371700 285660
rect 371752 285648 371758 285660
rect 381078 285648 381084 285660
rect 371752 285620 381084 285648
rect 371752 285608 371758 285620
rect 381078 285608 381084 285620
rect 381136 285608 381142 285660
rect 371602 285472 371608 285524
rect 371660 285512 371666 285524
rect 375374 285512 375380 285524
rect 371660 285484 375380 285512
rect 371660 285472 371666 285484
rect 375374 285472 375380 285484
rect 375432 285512 375438 285524
rect 375650 285512 375656 285524
rect 375432 285484 375656 285512
rect 375432 285472 375438 285484
rect 375650 285472 375656 285484
rect 375708 285472 375714 285524
rect 445386 284792 445392 284844
rect 445444 284832 445450 284844
rect 447134 284832 447140 284844
rect 445444 284804 447140 284832
rect 445444 284792 445450 284804
rect 447134 284792 447140 284804
rect 447192 284792 447198 284844
rect 381078 284384 381084 284436
rect 381136 284424 381142 284436
rect 382274 284424 382280 284436
rect 381136 284396 382280 284424
rect 381136 284384 381142 284396
rect 382274 284384 382280 284396
rect 382332 284384 382338 284436
rect 371602 284316 371608 284368
rect 371660 284356 371666 284368
rect 377398 284356 377404 284368
rect 371660 284328 377404 284356
rect 371660 284316 371666 284328
rect 377398 284316 377404 284328
rect 377456 284356 377462 284368
rect 385218 284356 385224 284368
rect 377456 284328 385224 284356
rect 377456 284316 377462 284328
rect 385218 284316 385224 284328
rect 385276 284316 385282 284368
rect 447134 284316 447140 284368
rect 447192 284356 447198 284368
rect 447318 284356 447324 284368
rect 447192 284328 447324 284356
rect 447192 284316 447198 284328
rect 447318 284316 447324 284328
rect 447376 284316 447382 284368
rect 371694 283636 371700 283688
rect 371752 283676 371758 283688
rect 376754 283676 376760 283688
rect 371752 283648 376760 283676
rect 371752 283636 371758 283648
rect 376754 283636 376760 283648
rect 376812 283636 376818 283688
rect 371602 283568 371608 283620
rect 371660 283608 371666 283620
rect 380894 283608 380900 283620
rect 371660 283580 380900 283608
rect 371660 283568 371666 283580
rect 380894 283568 380900 283580
rect 380952 283568 380958 283620
rect 445662 283568 445668 283620
rect 445720 283608 445726 283620
rect 450078 283608 450084 283620
rect 445720 283580 450084 283608
rect 445720 283568 445726 283580
rect 450078 283568 450084 283580
rect 450136 283568 450142 283620
rect 178678 282888 178684 282940
rect 178736 282928 178742 282940
rect 197354 282928 197360 282940
rect 178736 282900 197360 282928
rect 178736 282888 178742 282900
rect 197354 282888 197360 282900
rect 197412 282888 197418 282940
rect 380894 282888 380900 282940
rect 380952 282928 380958 282940
rect 381170 282928 381176 282940
rect 380952 282900 381176 282928
rect 380952 282888 380958 282900
rect 381170 282888 381176 282900
rect 381228 282888 381234 282940
rect 371602 282684 371608 282736
rect 371660 282724 371666 282736
rect 375466 282724 375472 282736
rect 371660 282696 375472 282724
rect 371660 282684 371666 282696
rect 375466 282684 375472 282696
rect 375524 282684 375530 282736
rect 371602 282140 371608 282192
rect 371660 282180 371666 282192
rect 374086 282180 374092 282192
rect 371660 282152 374092 282180
rect 371660 282140 371666 282152
rect 374086 282140 374092 282152
rect 374144 282180 374150 282192
rect 374270 282180 374276 282192
rect 374144 282152 374276 282180
rect 374144 282140 374150 282152
rect 374270 282140 374276 282152
rect 374328 282140 374334 282192
rect 181438 281528 181444 281580
rect 181496 281568 181502 281580
rect 197354 281568 197360 281580
rect 181496 281540 197360 281568
rect 181496 281528 181502 281540
rect 197354 281528 197360 281540
rect 197412 281528 197418 281580
rect 302510 281528 302516 281580
rect 302568 281568 302574 281580
rect 353938 281568 353944 281580
rect 302568 281540 353944 281568
rect 302568 281528 302574 281540
rect 353938 281528 353944 281540
rect 353996 281528 354002 281580
rect 445662 281324 445668 281376
rect 445720 281364 445726 281376
rect 448698 281364 448704 281376
rect 445720 281336 448704 281364
rect 445720 281324 445726 281336
rect 448698 281324 448704 281336
rect 448756 281324 448762 281376
rect 445018 280236 445024 280288
rect 445076 280276 445082 280288
rect 447226 280276 447232 280288
rect 445076 280248 447232 280276
rect 445076 280236 445082 280248
rect 447226 280236 447232 280248
rect 447284 280236 447290 280288
rect 444374 279624 444380 279676
rect 444432 279664 444438 279676
rect 444650 279664 444656 279676
rect 444432 279636 444656 279664
rect 444432 279624 444438 279636
rect 444650 279624 444656 279636
rect 444708 279624 444714 279676
rect 371970 278944 371976 278996
rect 372028 278984 372034 278996
rect 374086 278984 374092 278996
rect 372028 278956 374092 278984
rect 372028 278944 372034 278956
rect 374086 278944 374092 278956
rect 374144 278944 374150 278996
rect 173158 278740 173164 278792
rect 173216 278780 173222 278792
rect 197722 278780 197728 278792
rect 173216 278752 197728 278780
rect 173216 278740 173222 278752
rect 197722 278740 197728 278752
rect 197780 278740 197786 278792
rect 302786 278740 302792 278792
rect 302844 278780 302850 278792
rect 356698 278780 356704 278792
rect 302844 278752 356704 278780
rect 302844 278740 302850 278752
rect 356698 278740 356704 278752
rect 356756 278740 356762 278792
rect 369118 278604 369124 278656
rect 369176 278644 369182 278656
rect 369394 278644 369400 278656
rect 369176 278616 369400 278644
rect 369176 278604 369182 278616
rect 369394 278604 369400 278616
rect 369452 278604 369458 278656
rect 371694 277312 371700 277364
rect 371752 277352 371758 277364
rect 373994 277352 374000 277364
rect 371752 277324 374000 277352
rect 371752 277312 371758 277324
rect 373994 277312 374000 277324
rect 374052 277312 374058 277364
rect 445662 276632 445668 276684
rect 445720 276672 445726 276684
rect 454218 276672 454224 276684
rect 445720 276644 454224 276672
rect 445720 276632 445726 276644
rect 454218 276632 454224 276644
rect 454276 276632 454282 276684
rect 371694 276088 371700 276140
rect 371752 276128 371758 276140
rect 374362 276128 374368 276140
rect 371752 276100 374368 276128
rect 371752 276088 371758 276100
rect 374362 276088 374368 276100
rect 374420 276128 374426 276140
rect 375098 276128 375104 276140
rect 374420 276100 375104 276128
rect 374420 276088 374426 276100
rect 375098 276088 375104 276100
rect 375156 276088 375162 276140
rect 169662 276020 169668 276072
rect 169720 276060 169726 276072
rect 197354 276060 197360 276072
rect 169720 276032 197360 276060
rect 169720 276020 169726 276032
rect 197354 276020 197360 276032
rect 197412 276020 197418 276072
rect 302786 276020 302792 276072
rect 302844 276060 302850 276072
rect 360194 276060 360200 276072
rect 302844 276032 360200 276060
rect 302844 276020 302850 276032
rect 360194 276020 360200 276032
rect 360252 276060 360258 276072
rect 360654 276060 360660 276072
rect 360252 276032 360660 276060
rect 360252 276020 360258 276032
rect 360654 276020 360660 276032
rect 360712 276020 360718 276072
rect 373994 276020 374000 276072
rect 374052 276060 374058 276072
rect 374546 276060 374552 276072
rect 374052 276032 374552 276060
rect 374052 276020 374058 276032
rect 374546 276020 374552 276032
rect 374604 276020 374610 276072
rect 445662 275952 445668 276004
rect 445720 275992 445726 276004
rect 447502 275992 447508 276004
rect 445720 275964 447508 275992
rect 445720 275952 445726 275964
rect 447502 275952 447508 275964
rect 447560 275952 447566 276004
rect 369210 275340 369216 275392
rect 369268 275380 369274 275392
rect 369394 275380 369400 275392
rect 369268 275352 369400 275380
rect 369268 275340 369274 275352
rect 369394 275340 369400 275352
rect 369452 275340 369458 275392
rect 447502 275272 447508 275324
rect 447560 275312 447566 275324
rect 458358 275312 458364 275324
rect 447560 275284 458364 275312
rect 447560 275272 447566 275284
rect 458358 275272 458364 275284
rect 458416 275272 458422 275324
rect 372614 274728 372620 274780
rect 372672 274768 372678 274780
rect 373074 274768 373080 274780
rect 372672 274740 373080 274768
rect 372672 274728 372678 274740
rect 373074 274728 373080 274740
rect 373132 274728 373138 274780
rect 196618 274660 196624 274712
rect 196676 274700 196682 274712
rect 198642 274700 198648 274712
rect 196676 274672 198648 274700
rect 196676 274660 196682 274672
rect 198642 274660 198648 274672
rect 198700 274660 198706 274712
rect 370314 274660 370320 274712
rect 370372 274700 370378 274712
rect 372890 274700 372896 274712
rect 370372 274672 372896 274700
rect 370372 274660 370378 274672
rect 372890 274660 372896 274672
rect 372948 274660 372954 274712
rect 445662 274592 445668 274644
rect 445720 274632 445726 274644
rect 446398 274632 446404 274644
rect 445720 274604 446404 274632
rect 445720 274592 445726 274604
rect 446398 274592 446404 274604
rect 446456 274632 446462 274644
rect 452838 274632 452844 274644
rect 446456 274604 452844 274632
rect 446456 274592 446462 274604
rect 452838 274592 452844 274604
rect 452896 274592 452902 274644
rect 445018 273912 445024 273964
rect 445076 273952 445082 273964
rect 453298 273952 453304 273964
rect 445076 273924 453304 273952
rect 445076 273912 445082 273924
rect 453298 273912 453304 273924
rect 453356 273952 453362 273964
rect 456886 273952 456892 273964
rect 453356 273924 456892 273952
rect 453356 273912 453362 273924
rect 456886 273912 456892 273924
rect 456944 273912 456950 273964
rect 442258 273164 442264 273216
rect 442316 273204 442322 273216
rect 579890 273204 579896 273216
rect 442316 273176 579896 273204
rect 442316 273164 442322 273176
rect 579890 273164 579896 273176
rect 579948 273164 579954 273216
rect 445662 272484 445668 272536
rect 445720 272524 445726 272536
rect 451274 272524 451280 272536
rect 445720 272496 451280 272524
rect 445720 272484 445726 272496
rect 451274 272484 451280 272496
rect 451332 272524 451338 272536
rect 456886 272524 456892 272536
rect 451332 272496 456892 272524
rect 451332 272484 451338 272496
rect 456886 272484 456892 272496
rect 456944 272484 456950 272536
rect 177298 271872 177304 271924
rect 177356 271912 177362 271924
rect 197538 271912 197544 271924
rect 177356 271884 197544 271912
rect 177356 271872 177362 271884
rect 197538 271872 197544 271884
rect 197596 271872 197602 271924
rect 195238 270512 195244 270564
rect 195296 270552 195302 270564
rect 197722 270552 197728 270564
rect 195296 270524 197728 270552
rect 195296 270512 195302 270524
rect 197722 270512 197728 270524
rect 197780 270512 197786 270564
rect 445662 270512 445668 270564
rect 445720 270552 445726 270564
rect 451366 270552 451372 270564
rect 445720 270524 451372 270552
rect 445720 270512 445726 270524
rect 451366 270512 451372 270524
rect 451424 270552 451430 270564
rect 458174 270552 458180 270564
rect 451424 270524 458180 270552
rect 451424 270512 451430 270524
rect 458174 270512 458180 270524
rect 458232 270512 458238 270564
rect 447226 270444 447232 270496
rect 447284 270484 447290 270496
rect 447410 270484 447416 270496
rect 447284 270456 447416 270484
rect 447284 270444 447290 270456
rect 447410 270444 447416 270456
rect 447468 270444 447474 270496
rect 445386 269764 445392 269816
rect 445444 269804 445450 269816
rect 447226 269804 447232 269816
rect 445444 269776 447232 269804
rect 445444 269764 445450 269776
rect 447226 269764 447232 269776
rect 447284 269764 447290 269816
rect 369026 268744 369032 268796
rect 369084 268784 369090 268796
rect 369084 268756 369164 268784
rect 369084 268744 369090 268756
rect 369136 268456 369164 268756
rect 444558 268676 444564 268728
rect 444616 268716 444622 268728
rect 446030 268716 446036 268728
rect 444616 268688 446036 268716
rect 444616 268676 444622 268688
rect 446030 268676 446036 268688
rect 446088 268676 446094 268728
rect 369118 268404 369124 268456
rect 369176 268404 369182 268456
rect 303246 268336 303252 268388
rect 303304 268376 303310 268388
rect 327718 268376 327724 268388
rect 303304 268348 327724 268376
rect 303304 268336 303310 268348
rect 327718 268336 327724 268348
rect 327776 268336 327782 268388
rect 192478 268132 192484 268184
rect 192536 268172 192542 268184
rect 197814 268172 197820 268184
rect 192536 268144 197820 268172
rect 192536 268132 192542 268144
rect 197814 268132 197820 268144
rect 197872 268132 197878 268184
rect 3510 267656 3516 267708
rect 3568 267696 3574 267708
rect 90358 267696 90364 267708
rect 3568 267668 90364 267696
rect 3568 267656 3574 267668
rect 90358 267656 90364 267668
rect 90416 267656 90422 267708
rect 323578 267656 323584 267708
rect 323636 267696 323642 267708
rect 438854 267696 438860 267708
rect 323636 267668 438860 267696
rect 323636 267656 323642 267668
rect 438854 267656 438860 267668
rect 438912 267656 438918 267708
rect 191098 266432 191104 266484
rect 191156 266472 191162 266484
rect 197354 266472 197360 266484
rect 191156 266444 197360 266472
rect 191156 266432 191162 266444
rect 197354 266432 197360 266444
rect 197412 266432 197418 266484
rect 359458 266296 359464 266348
rect 359516 266336 359522 266348
rect 366910 266336 366916 266348
rect 359516 266308 366916 266336
rect 359516 266296 359522 266308
rect 366910 266296 366916 266308
rect 366968 266296 366974 266348
rect 435174 266336 435180 266348
rect 369826 266308 435180 266336
rect 362862 266228 362868 266280
rect 362920 266268 362926 266280
rect 369826 266268 369854 266308
rect 435174 266296 435180 266308
rect 435232 266336 435238 266348
rect 441614 266336 441620 266348
rect 435232 266308 441620 266336
rect 435232 266296 435238 266308
rect 441614 266296 441620 266308
rect 441672 266296 441678 266348
rect 437382 266268 437388 266280
rect 362920 266240 369854 266268
rect 373966 266240 437388 266268
rect 362920 266228 362926 266240
rect 324958 266160 324964 266212
rect 325016 266200 325022 266212
rect 325016 266172 354674 266200
rect 325016 266160 325022 266172
rect 354646 266132 354674 266172
rect 364886 266160 364892 266212
rect 364944 266200 364950 266212
rect 373966 266200 373994 266240
rect 437382 266228 437388 266240
rect 437440 266268 437446 266280
rect 442994 266268 443000 266280
rect 437440 266240 443000 266268
rect 437440 266228 437446 266240
rect 442994 266228 443000 266240
rect 443052 266228 443058 266280
rect 364944 266172 373994 266200
rect 364944 266160 364950 266172
rect 368474 266132 368480 266144
rect 354646 266104 368480 266132
rect 368474 266092 368480 266104
rect 368532 266092 368538 266144
rect 360194 265684 360200 265736
rect 360252 265724 360258 265736
rect 360930 265724 360936 265736
rect 360252 265696 360936 265724
rect 360252 265684 360258 265696
rect 360930 265684 360936 265696
rect 360988 265724 360994 265736
rect 431954 265724 431960 265736
rect 360988 265696 431960 265724
rect 360988 265684 360994 265696
rect 431954 265684 431960 265696
rect 432012 265724 432018 265736
rect 432598 265724 432604 265736
rect 432012 265696 432604 265724
rect 432012 265684 432018 265696
rect 432598 265684 432604 265696
rect 432656 265684 432662 265736
rect 368474 265616 368480 265668
rect 368532 265656 368538 265668
rect 369302 265656 369308 265668
rect 368532 265628 369308 265656
rect 368532 265616 368538 265628
rect 369302 265616 369308 265628
rect 369360 265656 369366 265668
rect 440878 265656 440884 265668
rect 369360 265628 440884 265656
rect 369360 265616 369366 265628
rect 440878 265616 440884 265628
rect 440936 265616 440942 265668
rect 302786 264868 302792 264920
rect 302844 264908 302850 264920
rect 352558 264908 352564 264920
rect 302844 264880 352564 264908
rect 302844 264868 302850 264880
rect 352558 264868 352564 264880
rect 352616 264868 352622 264920
rect 188430 263576 188436 263628
rect 188488 263616 188494 263628
rect 197354 263616 197360 263628
rect 188488 263588 197360 263616
rect 188488 263576 188494 263588
rect 197354 263576 197360 263588
rect 197412 263576 197418 263628
rect 187050 262216 187056 262268
rect 187108 262256 187114 262268
rect 197354 262256 197360 262268
rect 187108 262228 197360 262256
rect 187108 262216 187114 262228
rect 197354 262216 197360 262228
rect 197412 262216 197418 262268
rect 302786 262148 302792 262200
rect 302844 262188 302850 262200
rect 370130 262188 370136 262200
rect 302844 262160 370136 262188
rect 302844 262148 302850 262160
rect 370130 262148 370136 262160
rect 370188 262148 370194 262200
rect 184290 259428 184296 259480
rect 184348 259468 184354 259480
rect 197722 259468 197728 259480
rect 184348 259440 197728 259468
rect 184348 259428 184354 259440
rect 197722 259428 197728 259440
rect 197780 259428 197786 259480
rect 182818 256708 182824 256760
rect 182876 256748 182882 256760
rect 197538 256748 197544 256760
rect 182876 256720 197544 256748
rect 182876 256708 182882 256720
rect 197538 256708 197544 256720
rect 197596 256708 197602 256760
rect 302786 256708 302792 256760
rect 302844 256748 302850 256760
rect 370498 256748 370504 256760
rect 302844 256720 370504 256748
rect 302844 256708 302850 256720
rect 370498 256708 370504 256720
rect 370556 256708 370562 256760
rect 181530 255280 181536 255332
rect 181588 255320 181594 255332
rect 197906 255320 197912 255332
rect 181588 255292 197912 255320
rect 181588 255280 181594 255292
rect 197906 255280 197912 255292
rect 197964 255280 197970 255332
rect 3142 255212 3148 255264
rect 3200 255252 3206 255264
rect 180058 255252 180064 255264
rect 3200 255224 180064 255252
rect 3200 255212 3206 255224
rect 180058 255212 180064 255224
rect 180116 255212 180122 255264
rect 302326 253920 302332 253972
rect 302384 253960 302390 253972
rect 359458 253960 359464 253972
rect 302384 253932 359464 253960
rect 302384 253920 302390 253932
rect 359458 253920 359464 253932
rect 359516 253920 359522 253972
rect 180058 252560 180064 252612
rect 180116 252600 180122 252612
rect 197538 252600 197544 252612
rect 180116 252572 197544 252600
rect 180116 252560 180122 252572
rect 197538 252560 197544 252572
rect 197596 252560 197602 252612
rect 178770 251200 178776 251252
rect 178828 251240 178834 251252
rect 197354 251240 197360 251252
rect 178828 251212 197360 251240
rect 178828 251200 178834 251212
rect 197354 251200 197360 251212
rect 197412 251200 197418 251252
rect 370222 249704 370228 249756
rect 370280 249744 370286 249756
rect 373350 249744 373356 249756
rect 370280 249716 373356 249744
rect 370280 249704 370286 249716
rect 373350 249704 373356 249716
rect 373408 249704 373414 249756
rect 171778 248412 171784 248464
rect 171836 248452 171842 248464
rect 197630 248452 197636 248464
rect 171836 248424 197636 248452
rect 171836 248412 171842 248424
rect 197630 248412 197636 248424
rect 197688 248412 197694 248464
rect 302786 248412 302792 248464
rect 302844 248452 302850 248464
rect 370222 248452 370228 248464
rect 302844 248424 370228 248452
rect 302844 248412 302850 248424
rect 370222 248412 370228 248424
rect 370280 248412 370286 248464
rect 301498 245556 301504 245608
rect 301556 245596 301562 245608
rect 580166 245596 580172 245608
rect 301556 245568 580172 245596
rect 301556 245556 301562 245568
rect 580166 245556 580172 245568
rect 580224 245556 580230 245608
rect 173250 244264 173256 244316
rect 173308 244304 173314 244316
rect 197354 244304 197360 244316
rect 173308 244276 197360 244304
rect 173308 244264 173314 244276
rect 197354 244264 197360 244276
rect 197412 244264 197418 244316
rect 191190 241476 191196 241528
rect 191248 241516 191254 241528
rect 197906 241516 197912 241528
rect 191248 241488 197912 241516
rect 191248 241476 191254 241488
rect 197906 241476 197912 241488
rect 197964 241476 197970 241528
rect 3510 241408 3516 241460
rect 3568 241448 3574 241460
rect 174538 241448 174544 241460
rect 3568 241420 174544 241448
rect 3568 241408 3574 241420
rect 174538 241408 174544 241420
rect 174596 241408 174602 241460
rect 180150 240116 180156 240168
rect 180208 240156 180214 240168
rect 197722 240156 197728 240168
rect 180208 240128 197728 240156
rect 180208 240116 180214 240128
rect 197722 240116 197728 240128
rect 197780 240116 197786 240168
rect 302970 239368 302976 239420
rect 303028 239408 303034 239420
rect 370314 239408 370320 239420
rect 303028 239380 370320 239408
rect 303028 239368 303034 239380
rect 370314 239368 370320 239380
rect 370372 239368 370378 239420
rect 192570 237396 192576 237448
rect 192628 237436 192634 237448
rect 197538 237436 197544 237448
rect 192628 237408 197544 237436
rect 192628 237396 192634 237408
rect 197538 237396 197544 237408
rect 197596 237396 197602 237448
rect 195330 236104 195336 236156
rect 195388 236144 195394 236156
rect 197722 236144 197728 236156
rect 195388 236116 197728 236144
rect 195388 236104 195394 236116
rect 197722 236104 197728 236116
rect 197780 236104 197786 236156
rect 193858 233792 193864 233844
rect 193916 233832 193922 233844
rect 197722 233832 197728 233844
rect 193916 233804 197728 233832
rect 193916 233792 193922 233804
rect 197722 233792 197728 233804
rect 197780 233792 197786 233844
rect 312538 233180 312544 233232
rect 312596 233220 312602 233232
rect 579982 233220 579988 233232
rect 312596 233192 579988 233220
rect 312596 233180 312602 233192
rect 579982 233180 579988 233192
rect 580040 233180 580046 233232
rect 196710 231888 196716 231940
rect 196768 231928 196774 231940
rect 198366 231928 198372 231940
rect 196768 231900 198372 231928
rect 196768 231888 196774 231900
rect 198366 231888 198372 231900
rect 198424 231888 198430 231940
rect 303062 231072 303068 231124
rect 303120 231112 303126 231124
rect 369578 231112 369584 231124
rect 303120 231084 369584 231112
rect 303120 231072 303126 231084
rect 369578 231072 369584 231084
rect 369636 231112 369642 231124
rect 374178 231112 374184 231124
rect 369636 231084 374184 231112
rect 369636 231072 369642 231084
rect 374178 231072 374184 231084
rect 374236 231072 374242 231124
rect 303154 229712 303160 229764
rect 303212 229752 303218 229764
rect 372798 229752 372804 229764
rect 303212 229724 372804 229752
rect 303212 229712 303218 229724
rect 372798 229712 372804 229724
rect 372856 229712 372862 229764
rect 177390 229100 177396 229152
rect 177448 229140 177454 229152
rect 197630 229140 197636 229152
rect 177448 229112 197636 229140
rect 177448 229100 177454 229112
rect 197630 229100 197636 229112
rect 197688 229100 197694 229152
rect 311158 228352 311164 228404
rect 311216 228392 311222 228404
rect 580258 228392 580264 228404
rect 311216 228364 580264 228392
rect 311216 228352 311222 228364
rect 580258 228352 580264 228364
rect 580316 228352 580322 228404
rect 186958 227740 186964 227792
rect 187016 227780 187022 227792
rect 197354 227780 197360 227792
rect 187016 227752 197360 227780
rect 187016 227740 187022 227752
rect 197354 227740 197360 227752
rect 197412 227740 197418 227792
rect 303246 226992 303252 227044
rect 303304 227032 303310 227044
rect 372614 227032 372620 227044
rect 303304 227004 372620 227032
rect 303304 226992 303310 227004
rect 372614 226992 372620 227004
rect 372672 226992 372678 227044
rect 440878 226244 440884 226296
rect 440936 226284 440942 226296
rect 442994 226284 443000 226296
rect 440936 226256 443000 226284
rect 440936 226244 440942 226256
rect 442994 226244 443000 226256
rect 443052 226244 443058 226296
rect 437382 226176 437388 226228
rect 437440 226216 437446 226228
rect 441706 226216 441712 226228
rect 437440 226188 441712 226216
rect 437440 226176 437446 226188
rect 441706 226176 441712 226188
rect 441764 226176 441770 226228
rect 371602 225700 371608 225752
rect 371660 225740 371666 225752
rect 372338 225740 372344 225752
rect 371660 225712 372344 225740
rect 371660 225700 371666 225712
rect 372338 225700 372344 225712
rect 372396 225700 372402 225752
rect 372982 225700 372988 225752
rect 373040 225740 373046 225752
rect 373534 225740 373540 225752
rect 373040 225712 373540 225740
rect 373040 225700 373046 225712
rect 373534 225700 373540 225712
rect 373592 225740 373598 225752
rect 378410 225740 378416 225752
rect 373592 225712 378416 225740
rect 373592 225700 373598 225712
rect 378410 225700 378416 225712
rect 378468 225700 378474 225752
rect 372246 225632 372252 225684
rect 372304 225672 372310 225684
rect 373258 225672 373264 225684
rect 372304 225644 373264 225672
rect 372304 225632 372310 225644
rect 373258 225632 373264 225644
rect 373316 225672 373322 225684
rect 381078 225672 381084 225684
rect 373316 225644 381084 225672
rect 373316 225632 373322 225644
rect 381078 225632 381084 225644
rect 381136 225632 381142 225684
rect 302878 225564 302884 225616
rect 302936 225604 302942 225616
rect 369854 225604 369860 225616
rect 302936 225576 369860 225604
rect 302936 225564 302942 225576
rect 369854 225564 369860 225576
rect 369912 225564 369918 225616
rect 371602 225564 371608 225616
rect 371660 225604 371666 225616
rect 385126 225604 385132 225616
rect 371660 225576 385132 225604
rect 371660 225564 371666 225576
rect 385126 225564 385132 225576
rect 385184 225564 385190 225616
rect 359642 225292 359648 225344
rect 359700 225332 359706 225344
rect 372982 225332 372988 225344
rect 359700 225304 372988 225332
rect 359700 225292 359706 225304
rect 372982 225292 372988 225304
rect 373040 225292 373046 225344
rect 372798 225224 372804 225276
rect 372856 225264 372862 225276
rect 373166 225264 373172 225276
rect 372856 225236 373172 225264
rect 372856 225224 372862 225236
rect 373166 225224 373172 225236
rect 373224 225224 373230 225276
rect 359366 225156 359372 225208
rect 359424 225196 359430 225208
rect 374362 225196 374368 225208
rect 359424 225168 374368 225196
rect 359424 225156 359430 225168
rect 374362 225156 374368 225168
rect 374420 225196 374426 225208
rect 378318 225196 378324 225208
rect 374420 225168 378324 225196
rect 374420 225156 374426 225168
rect 378318 225156 378324 225168
rect 378376 225156 378382 225208
rect 359550 225088 359556 225140
rect 359608 225128 359614 225140
rect 383746 225128 383752 225140
rect 359608 225100 383752 225128
rect 359608 225088 359614 225100
rect 383746 225088 383752 225100
rect 383804 225088 383810 225140
rect 371234 225020 371240 225072
rect 371292 225060 371298 225072
rect 372798 225060 372804 225072
rect 371292 225032 372804 225060
rect 371292 225020 371298 225032
rect 372798 225020 372804 225032
rect 372856 225060 372862 225072
rect 441798 225060 441804 225072
rect 372856 225032 441804 225060
rect 372856 225020 372862 225032
rect 441798 225020 441804 225032
rect 441856 225060 441862 225072
rect 441856 225032 449940 225060
rect 441856 225020 441862 225032
rect 449912 225004 449940 225032
rect 184198 224952 184204 225004
rect 184256 224992 184262 225004
rect 197354 224992 197360 225004
rect 184256 224964 197360 224992
rect 184256 224952 184262 224964
rect 197354 224952 197360 224964
rect 197412 224952 197418 225004
rect 372522 224952 372528 225004
rect 372580 224992 372586 225004
rect 372982 224992 372988 225004
rect 372580 224964 372988 224992
rect 372580 224952 372586 224964
rect 372982 224952 372988 224964
rect 373040 224992 373046 225004
rect 444558 224992 444564 225004
rect 373040 224964 444564 224992
rect 373040 224952 373046 224964
rect 444558 224952 444564 224964
rect 444616 224952 444622 225004
rect 449894 224952 449900 225004
rect 449952 224992 449958 225004
rect 450170 224992 450176 225004
rect 449952 224964 450176 224992
rect 449952 224952 449958 224964
rect 450170 224952 450176 224964
rect 450228 224952 450234 225004
rect 359458 224408 359464 224460
rect 359516 224448 359522 224460
rect 369394 224448 369400 224460
rect 359516 224420 369400 224448
rect 359516 224408 359522 224420
rect 369394 224408 369400 224420
rect 369452 224408 369458 224460
rect 302786 224340 302792 224392
rect 302844 224380 302850 224392
rect 369946 224380 369952 224392
rect 302844 224352 369952 224380
rect 302844 224340 302850 224352
rect 369946 224340 369952 224352
rect 370004 224340 370010 224392
rect 302694 224272 302700 224324
rect 302752 224312 302758 224324
rect 370222 224312 370228 224324
rect 302752 224284 370228 224312
rect 302752 224272 302758 224284
rect 370222 224272 370228 224284
rect 370280 224272 370286 224324
rect 371326 224272 371332 224324
rect 371384 224312 371390 224324
rect 379514 224312 379520 224324
rect 371384 224284 379520 224312
rect 371384 224272 371390 224284
rect 379514 224272 379520 224284
rect 379572 224272 379578 224324
rect 302970 224204 302976 224256
rect 303028 224244 303034 224256
rect 370406 224244 370412 224256
rect 303028 224216 370412 224244
rect 303028 224204 303034 224216
rect 370406 224204 370412 224216
rect 370464 224204 370470 224256
rect 371602 224204 371608 224256
rect 371660 224244 371666 224256
rect 383654 224244 383660 224256
rect 371660 224216 383660 224244
rect 371660 224204 371666 224216
rect 383654 224204 383660 224216
rect 383712 224204 383718 224256
rect 441798 224244 441804 224256
rect 431926 224216 441804 224244
rect 359734 223932 359740 223984
rect 359792 223972 359798 223984
rect 385310 223972 385316 223984
rect 359792 223944 385316 223972
rect 359792 223932 359798 223944
rect 385310 223932 385316 223944
rect 385368 223932 385374 223984
rect 359458 223864 359464 223916
rect 359516 223904 359522 223916
rect 374454 223904 374460 223916
rect 359516 223876 374460 223904
rect 359516 223864 359522 223876
rect 374454 223864 374460 223876
rect 374512 223864 374518 223916
rect 431926 223904 431954 224216
rect 441798 224204 441804 224216
rect 441856 224244 441862 224256
rect 458266 224244 458272 224256
rect 441856 224216 458272 224244
rect 441856 224204 441862 224216
rect 458266 224204 458272 224216
rect 458324 224204 458330 224256
rect 383626 223876 431954 223904
rect 373994 223796 374000 223848
rect 374052 223836 374058 223848
rect 383626 223836 383654 223876
rect 374052 223808 383654 223836
rect 374052 223796 374058 223808
rect 302786 223524 302792 223576
rect 302844 223564 302850 223576
rect 359366 223564 359372 223576
rect 302844 223536 359372 223564
rect 302844 223524 302850 223536
rect 359366 223524 359372 223536
rect 359424 223524 359430 223576
rect 378318 223524 378324 223576
rect 378376 223564 378382 223576
rect 382458 223564 382464 223576
rect 378376 223536 382464 223564
rect 378376 223524 378382 223536
rect 382458 223524 382464 223536
rect 382516 223524 382522 223576
rect 444558 223524 444564 223576
rect 444616 223564 444622 223576
rect 454034 223564 454040 223576
rect 444616 223536 454040 223564
rect 444616 223524 444622 223536
rect 454034 223524 454040 223536
rect 454092 223524 454098 223576
rect 371602 222844 371608 222896
rect 371660 222884 371666 222896
rect 374914 222884 374920 222896
rect 371660 222856 374920 222884
rect 371660 222844 371666 222856
rect 374914 222844 374920 222856
rect 374972 222884 374978 222896
rect 378134 222884 378140 222896
rect 374972 222856 378140 222884
rect 374972 222844 374978 222856
rect 378134 222844 378140 222856
rect 378192 222844 378198 222896
rect 371234 222368 371240 222420
rect 371292 222408 371298 222420
rect 375650 222408 375656 222420
rect 371292 222380 375656 222408
rect 371292 222368 371298 222380
rect 375650 222368 375656 222380
rect 375708 222408 375714 222420
rect 376938 222408 376944 222420
rect 375708 222380 376944 222408
rect 375708 222368 375714 222380
rect 376938 222368 376944 222380
rect 376996 222368 377002 222420
rect 371602 222300 371608 222352
rect 371660 222340 371666 222352
rect 372338 222340 372344 222352
rect 371660 222312 372344 222340
rect 371660 222300 371666 222312
rect 372338 222300 372344 222312
rect 372396 222340 372402 222352
rect 373994 222340 374000 222352
rect 372396 222312 374000 222340
rect 372396 222300 372402 222312
rect 373994 222300 374000 222312
rect 374052 222300 374058 222352
rect 371326 222232 371332 222284
rect 371384 222272 371390 222284
rect 378318 222272 378324 222284
rect 371384 222244 378324 222272
rect 371384 222232 371390 222244
rect 378318 222232 378324 222244
rect 378376 222232 378382 222284
rect 188338 222164 188344 222216
rect 188396 222204 188402 222216
rect 197354 222204 197360 222216
rect 188396 222176 197360 222204
rect 188396 222164 188402 222176
rect 197354 222164 197360 222176
rect 197412 222164 197418 222216
rect 445662 222096 445668 222148
rect 445720 222136 445726 222148
rect 448606 222136 448612 222148
rect 445720 222108 448612 222136
rect 445720 222096 445726 222108
rect 448606 222096 448612 222108
rect 448664 222136 448670 222148
rect 448790 222136 448796 222148
rect 448664 222108 448796 222136
rect 448664 222096 448670 222108
rect 448790 222096 448796 222108
rect 448848 222096 448854 222148
rect 370130 221416 370136 221468
rect 370188 221456 370194 221468
rect 385034 221456 385040 221468
rect 370188 221428 385040 221456
rect 370188 221416 370194 221428
rect 385034 221416 385040 221428
rect 385092 221416 385098 221468
rect 371234 220872 371240 220924
rect 371292 220912 371298 220924
rect 382458 220912 382464 220924
rect 371292 220884 382464 220912
rect 371292 220872 371298 220884
rect 382458 220872 382464 220884
rect 382516 220912 382522 220924
rect 385402 220912 385408 220924
rect 382516 220884 385408 220912
rect 382516 220872 382522 220884
rect 385402 220872 385408 220884
rect 385460 220872 385466 220924
rect 302786 220736 302792 220788
rect 302844 220776 302850 220788
rect 359458 220776 359464 220788
rect 302844 220748 359464 220776
rect 302844 220736 302850 220748
rect 359458 220736 359464 220748
rect 359516 220736 359522 220788
rect 369854 220736 369860 220788
rect 369912 220776 369918 220788
rect 376018 220776 376024 220788
rect 369912 220748 376024 220776
rect 369912 220736 369918 220748
rect 376018 220736 376024 220748
rect 376076 220776 376082 220788
rect 380894 220776 380900 220788
rect 376076 220748 380900 220776
rect 376076 220736 376082 220748
rect 380894 220736 380900 220748
rect 380952 220736 380958 220788
rect 456794 220736 456800 220788
rect 456852 220776 456858 220788
rect 456978 220776 456984 220788
rect 456852 220748 456984 220776
rect 456852 220736 456858 220748
rect 456978 220736 456984 220748
rect 457036 220736 457042 220788
rect 371234 220668 371240 220720
rect 371292 220708 371298 220720
rect 372798 220708 372804 220720
rect 371292 220680 372804 220708
rect 371292 220668 371298 220680
rect 372798 220668 372804 220680
rect 372856 220668 372862 220720
rect 373166 220668 373172 220720
rect 373224 220708 373230 220720
rect 382366 220708 382372 220720
rect 373224 220680 382372 220708
rect 373224 220668 373230 220680
rect 382366 220668 382372 220680
rect 382424 220668 382430 220720
rect 372062 220600 372068 220652
rect 372120 220640 372126 220652
rect 373184 220640 373212 220668
rect 372120 220612 373212 220640
rect 372120 220600 372126 220612
rect 445110 220056 445116 220108
rect 445168 220096 445174 220108
rect 456978 220096 456984 220108
rect 445168 220068 456984 220096
rect 445168 220056 445174 220068
rect 456978 220056 456984 220068
rect 457036 220056 457042 220108
rect 445662 219580 445668 219632
rect 445720 219620 445726 219632
rect 452746 219620 452752 219632
rect 445720 219592 452752 219620
rect 445720 219580 445726 219592
rect 452746 219580 452752 219592
rect 452804 219580 452810 219632
rect 372614 219376 372620 219428
rect 372672 219416 372678 219428
rect 380986 219416 380992 219428
rect 372672 219388 380992 219416
rect 372672 219376 372678 219388
rect 380986 219376 380992 219388
rect 381044 219376 381050 219428
rect 443638 219376 443644 219428
rect 443696 219416 443702 219428
rect 579890 219416 579896 219428
rect 443696 219388 579896 219416
rect 443696 219376 443702 219388
rect 579890 219376 579896 219388
rect 579948 219376 579954 219428
rect 370406 218696 370412 218748
rect 370464 218736 370470 218748
rect 378502 218736 378508 218748
rect 370464 218708 378508 218736
rect 370464 218696 370470 218708
rect 378502 218696 378508 218708
rect 378560 218696 378566 218748
rect 378226 218220 378232 218272
rect 378284 218260 378290 218272
rect 378502 218260 378508 218272
rect 378284 218232 378508 218260
rect 378284 218220 378290 218232
rect 378502 218220 378508 218232
rect 378560 218220 378566 218272
rect 371050 218084 371056 218136
rect 371108 218124 371114 218136
rect 375926 218124 375932 218136
rect 371108 218096 375932 218124
rect 371108 218084 371114 218096
rect 375926 218084 375932 218096
rect 375984 218124 375990 218136
rect 377030 218124 377036 218136
rect 375984 218096 377036 218124
rect 375984 218084 375990 218096
rect 377030 218084 377036 218096
rect 377088 218084 377094 218136
rect 174538 218016 174544 218068
rect 174596 218056 174602 218068
rect 197538 218056 197544 218068
rect 174596 218028 197544 218056
rect 174596 218016 174602 218028
rect 197538 218016 197544 218028
rect 197596 218016 197602 218068
rect 445754 218016 445760 218068
rect 445812 218056 445818 218068
rect 446122 218056 446128 218068
rect 445812 218028 446128 218056
rect 445812 218016 445818 218028
rect 446122 218016 446128 218028
rect 446180 218016 446186 218068
rect 302510 217948 302516 218000
rect 302568 217988 302574 218000
rect 359734 217988 359740 218000
rect 302568 217960 359740 217988
rect 302568 217948 302574 217960
rect 359734 217948 359740 217960
rect 359792 217948 359798 218000
rect 370222 217948 370228 218000
rect 370280 217988 370286 218000
rect 375558 217988 375564 218000
rect 370280 217960 375564 217988
rect 370280 217948 370286 217960
rect 375558 217948 375564 217960
rect 375616 217948 375622 218000
rect 445662 217268 445668 217320
rect 445720 217308 445726 217320
rect 454126 217308 454132 217320
rect 445720 217280 454132 217308
rect 445720 217268 445726 217280
rect 454126 217268 454132 217280
rect 454184 217268 454190 217320
rect 371602 217132 371608 217184
rect 371660 217172 371666 217184
rect 372246 217172 372252 217184
rect 371660 217144 372252 217172
rect 371660 217132 371666 217144
rect 372246 217132 372252 217144
rect 372304 217132 372310 217184
rect 371602 216996 371608 217048
rect 371660 217036 371666 217048
rect 374362 217036 374368 217048
rect 371660 217008 374368 217036
rect 371660 216996 371666 217008
rect 374362 216996 374368 217008
rect 374420 216996 374426 217048
rect 174630 216656 174636 216708
rect 174688 216696 174694 216708
rect 197354 216696 197360 216708
rect 174688 216668 197360 216696
rect 174688 216656 174694 216668
rect 197354 216656 197360 216668
rect 197412 216656 197418 216708
rect 375558 216656 375564 216708
rect 375616 216696 375622 216708
rect 376938 216696 376944 216708
rect 375616 216668 376944 216696
rect 375616 216656 375622 216668
rect 376938 216656 376944 216668
rect 376996 216656 377002 216708
rect 445662 216112 445668 216164
rect 445720 216152 445726 216164
rect 449986 216152 449992 216164
rect 445720 216124 449992 216152
rect 445720 216112 445726 216124
rect 449986 216112 449992 216124
rect 450044 216112 450050 216164
rect 371326 215976 371332 216028
rect 371384 216016 371390 216028
rect 374454 216016 374460 216028
rect 371384 215988 374460 216016
rect 371384 215976 371390 215988
rect 374454 215976 374460 215988
rect 374512 216016 374518 216028
rect 378134 216016 378140 216028
rect 374512 215988 378140 216016
rect 374512 215976 374518 215988
rect 378134 215976 378140 215988
rect 378192 215976 378198 216028
rect 371602 215908 371608 215960
rect 371660 215948 371666 215960
rect 375558 215948 375564 215960
rect 371660 215920 375564 215948
rect 371660 215908 371666 215920
rect 375558 215908 375564 215920
rect 375616 215948 375622 215960
rect 385218 215948 385224 215960
rect 375616 215920 385224 215948
rect 375616 215908 375622 215920
rect 385218 215908 385224 215920
rect 385276 215908 385282 215960
rect 372338 215432 372344 215484
rect 372396 215472 372402 215484
rect 373534 215472 373540 215484
rect 372396 215444 373540 215472
rect 372396 215432 372402 215444
rect 373534 215432 373540 215444
rect 373592 215472 373598 215484
rect 375006 215472 375012 215484
rect 373592 215444 375012 215472
rect 373592 215432 373598 215444
rect 375006 215432 375012 215444
rect 375064 215432 375070 215484
rect 449986 215296 449992 215348
rect 450044 215336 450050 215348
rect 450170 215336 450176 215348
rect 450044 215308 450176 215336
rect 450044 215296 450050 215308
rect 450170 215296 450176 215308
rect 450228 215296 450234 215348
rect 3326 215228 3332 215280
rect 3384 215268 3390 215280
rect 199378 215268 199384 215280
rect 3384 215240 199384 215268
rect 3384 215228 3390 215240
rect 199378 215228 199384 215240
rect 199436 215228 199442 215280
rect 302786 215228 302792 215280
rect 302844 215268 302850 215280
rect 359642 215268 359648 215280
rect 302844 215240 359648 215268
rect 302844 215228 302850 215240
rect 359642 215228 359648 215240
rect 359700 215228 359706 215280
rect 371602 215228 371608 215280
rect 371660 215268 371666 215280
rect 371660 215240 373994 215268
rect 371660 215228 371666 215240
rect 373966 215200 373994 215240
rect 383746 215200 383752 215212
rect 373966 215172 383752 215200
rect 383746 215160 383752 215172
rect 383804 215200 383810 215212
rect 385218 215200 385224 215212
rect 383804 215172 385224 215200
rect 383804 215160 383810 215172
rect 385218 215160 385224 215172
rect 385276 215160 385282 215212
rect 378410 214344 378416 214396
rect 378468 214384 378474 214396
rect 381262 214384 381268 214396
rect 378468 214356 381268 214384
rect 378468 214344 378474 214356
rect 381262 214344 381268 214356
rect 381320 214344 381326 214396
rect 445662 214004 445668 214056
rect 445720 214044 445726 214056
rect 452654 214044 452660 214056
rect 445720 214016 452660 214044
rect 445720 214004 445726 214016
rect 452654 214004 452660 214016
rect 452712 214044 452718 214056
rect 452838 214044 452844 214056
rect 452712 214016 452844 214044
rect 452712 214004 452718 214016
rect 452838 214004 452844 214016
rect 452896 214004 452902 214056
rect 174722 213936 174728 213988
rect 174780 213976 174786 213988
rect 197538 213976 197544 213988
rect 174780 213948 197544 213976
rect 174780 213936 174786 213948
rect 197538 213936 197544 213948
rect 197596 213936 197602 213988
rect 371602 213936 371608 213988
rect 371660 213976 371666 213988
rect 378410 213976 378416 213988
rect 371660 213948 378416 213976
rect 371660 213936 371666 213948
rect 378410 213936 378416 213948
rect 378468 213936 378474 213988
rect 445662 213868 445668 213920
rect 445720 213908 445726 213920
rect 448514 213908 448520 213920
rect 445720 213880 448520 213908
rect 445720 213868 445726 213880
rect 448514 213868 448520 213880
rect 448572 213868 448578 213920
rect 372062 213732 372068 213784
rect 372120 213772 372126 213784
rect 377398 213772 377404 213784
rect 372120 213744 377404 213772
rect 372120 213732 372126 213744
rect 377398 213732 377404 213744
rect 377456 213772 377462 213784
rect 382550 213772 382556 213784
rect 377456 213744 382556 213772
rect 377456 213732 377462 213744
rect 382550 213732 382556 213744
rect 382608 213732 382614 213784
rect 371326 213256 371332 213308
rect 371384 213296 371390 213308
rect 374638 213296 374644 213308
rect 371384 213268 374644 213296
rect 371384 213256 371390 213268
rect 374638 213256 374644 213268
rect 374696 213296 374702 213308
rect 377030 213296 377036 213308
rect 374696 213268 377036 213296
rect 374696 213256 374702 213268
rect 377030 213256 377036 213268
rect 377088 213256 377094 213308
rect 371602 213188 371608 213240
rect 371660 213228 371666 213240
rect 375374 213228 375380 213240
rect 371660 213200 375380 213228
rect 371660 213188 371666 213200
rect 375374 213188 375380 213200
rect 375432 213228 375438 213240
rect 383746 213228 383752 213240
rect 375432 213200 383752 213228
rect 375432 213188 375438 213200
rect 383746 213188 383752 213200
rect 383804 213188 383810 213240
rect 371326 213120 371332 213172
rect 371384 213160 371390 213172
rect 372246 213160 372252 213172
rect 371384 213132 372252 213160
rect 371384 213120 371390 213132
rect 372246 213120 372252 213132
rect 372304 213120 372310 213172
rect 445294 212780 445300 212832
rect 445352 212820 445358 212832
rect 447318 212820 447324 212832
rect 445352 212792 447324 212820
rect 445352 212780 445358 212792
rect 447318 212780 447324 212792
rect 447376 212780 447382 212832
rect 170490 212508 170496 212560
rect 170548 212548 170554 212560
rect 197354 212548 197360 212560
rect 170548 212520 197360 212548
rect 170548 212508 170554 212520
rect 197354 212508 197360 212520
rect 197412 212508 197418 212560
rect 376846 212440 376852 212492
rect 376904 212480 376910 212492
rect 381170 212480 381176 212492
rect 376904 212452 381176 212480
rect 376904 212440 376910 212452
rect 381170 212440 381176 212452
rect 381228 212440 381234 212492
rect 372246 211760 372252 211812
rect 372304 211800 372310 211812
rect 373166 211800 373172 211812
rect 372304 211772 373172 211800
rect 372304 211760 372310 211772
rect 373166 211760 373172 211772
rect 373224 211800 373230 211812
rect 382274 211800 382280 211812
rect 373224 211772 382280 211800
rect 373224 211760 373230 211772
rect 382274 211760 382280 211772
rect 382332 211760 382338 211812
rect 445662 211556 445668 211608
rect 445720 211596 445726 211608
rect 450078 211596 450084 211608
rect 445720 211568 450084 211596
rect 445720 211556 445726 211568
rect 450078 211556 450084 211568
rect 450136 211556 450142 211608
rect 371602 211216 371608 211268
rect 371660 211256 371666 211268
rect 376754 211256 376760 211268
rect 371660 211228 376760 211256
rect 371660 211216 371666 211228
rect 376754 211216 376760 211228
rect 376812 211216 376818 211268
rect 370406 211148 370412 211200
rect 370464 211188 370470 211200
rect 376846 211188 376852 211200
rect 370464 211160 376852 211188
rect 370464 211148 370470 211160
rect 376846 211148 376852 211160
rect 376904 211148 376910 211200
rect 302786 211080 302792 211132
rect 302844 211120 302850 211132
rect 359550 211120 359556 211132
rect 302844 211092 359556 211120
rect 302844 211080 302850 211092
rect 359550 211080 359556 211092
rect 359608 211080 359614 211132
rect 374730 211080 374736 211132
rect 374788 211120 374794 211132
rect 375466 211120 375472 211132
rect 374788 211092 375472 211120
rect 374788 211080 374794 211092
rect 375466 211080 375472 211092
rect 375524 211080 375530 211132
rect 445846 211080 445852 211132
rect 445904 211120 445910 211132
rect 446030 211120 446036 211132
rect 445904 211092 446036 211120
rect 445904 211080 445910 211092
rect 446030 211080 446036 211092
rect 446088 211080 446094 211132
rect 371602 210604 371608 210656
rect 371660 210644 371666 210656
rect 374730 210644 374736 210656
rect 371660 210616 374736 210644
rect 371660 210604 371666 210616
rect 374730 210604 374736 210616
rect 374788 210604 374794 210656
rect 444558 210468 444564 210520
rect 444616 210508 444622 210520
rect 446030 210508 446036 210520
rect 444616 210480 446036 210508
rect 444616 210468 444622 210480
rect 446030 210468 446036 210480
rect 446088 210468 446094 210520
rect 372706 210060 372712 210112
rect 372764 210100 372770 210112
rect 374270 210100 374276 210112
rect 372764 210072 374276 210100
rect 372764 210060 372770 210072
rect 374270 210060 374276 210072
rect 374328 210060 374334 210112
rect 182910 209788 182916 209840
rect 182968 209828 182974 209840
rect 197354 209828 197360 209840
rect 182968 209800 197360 209828
rect 182968 209788 182974 209800
rect 197354 209788 197360 209800
rect 197412 209788 197418 209840
rect 375834 209788 375840 209840
rect 375892 209828 375898 209840
rect 376754 209828 376760 209840
rect 375892 209800 376760 209828
rect 375892 209788 375898 209800
rect 376754 209788 376760 209800
rect 376812 209788 376818 209840
rect 445662 209176 445668 209228
rect 445720 209216 445726 209228
rect 448698 209216 448704 209228
rect 445720 209188 448704 209216
rect 445720 209176 445726 209188
rect 448698 209176 448704 209188
rect 448756 209176 448762 209228
rect 160002 209040 160008 209092
rect 160060 209080 160066 209092
rect 198090 209080 198096 209092
rect 160060 209052 198096 209080
rect 160060 209040 160066 209052
rect 198090 209040 198096 209052
rect 198148 209040 198154 209092
rect 369670 208700 369676 208752
rect 369728 208740 369734 208752
rect 372982 208740 372988 208752
rect 369728 208712 372988 208740
rect 369728 208700 369734 208712
rect 372982 208700 372988 208712
rect 373040 208700 373046 208752
rect 445110 208156 445116 208208
rect 445168 208196 445174 208208
rect 447134 208196 447140 208208
rect 445168 208168 447140 208196
rect 445168 208156 445174 208168
rect 447134 208156 447140 208168
rect 447192 208156 447198 208208
rect 302326 207000 302332 207052
rect 302384 207040 302390 207052
rect 359458 207040 359464 207052
rect 302384 207012 359464 207040
rect 302384 207000 302390 207012
rect 359458 207000 359464 207012
rect 359516 207000 359522 207052
rect 369762 206932 369768 206984
rect 369820 206972 369826 206984
rect 374086 206972 374092 206984
rect 369820 206944 374092 206972
rect 369820 206932 369826 206944
rect 374086 206932 374092 206944
rect 374144 206932 374150 206984
rect 369302 206456 369308 206508
rect 369360 206456 369366 206508
rect 369210 206252 369216 206304
rect 369268 206292 369274 206304
rect 369320 206292 369348 206456
rect 369268 206264 369348 206292
rect 369268 206252 369274 206264
rect 369118 206116 369124 206168
rect 369176 206156 369182 206168
rect 369394 206156 369400 206168
rect 369176 206128 369400 206156
rect 369176 206116 369182 206128
rect 369394 206116 369400 206128
rect 369452 206116 369458 206168
rect 371602 205776 371608 205828
rect 371660 205816 371666 205828
rect 372614 205816 372620 205828
rect 371660 205788 372620 205816
rect 371660 205776 371666 205788
rect 372614 205776 372620 205788
rect 372672 205816 372678 205828
rect 373258 205816 373264 205828
rect 372672 205788 373264 205816
rect 372672 205776 372678 205788
rect 373258 205776 373264 205788
rect 373316 205776 373322 205828
rect 181622 205640 181628 205692
rect 181680 205680 181686 205692
rect 197354 205680 197360 205692
rect 181680 205652 197360 205680
rect 181680 205640 181686 205652
rect 197354 205640 197360 205652
rect 197412 205640 197418 205692
rect 445294 205572 445300 205624
rect 445352 205612 445358 205624
rect 454218 205612 454224 205624
rect 445352 205584 454224 205612
rect 445352 205572 445358 205584
rect 454218 205572 454224 205584
rect 454276 205612 454282 205624
rect 458174 205612 458180 205624
rect 454276 205584 458180 205612
rect 454276 205572 454282 205584
rect 458174 205572 458180 205584
rect 458232 205572 458238 205624
rect 371602 205300 371608 205352
rect 371660 205340 371666 205352
rect 374546 205340 374552 205352
rect 371660 205312 374552 205340
rect 371660 205300 371666 205312
rect 374546 205300 374552 205312
rect 374604 205300 374610 205352
rect 371602 204756 371608 204808
rect 371660 204796 371666 204808
rect 372890 204796 372896 204808
rect 371660 204768 372896 204796
rect 371660 204756 371666 204768
rect 372890 204756 372896 204768
rect 372948 204756 372954 204808
rect 302694 204280 302700 204332
rect 302752 204320 302758 204332
rect 359550 204320 359556 204332
rect 302752 204292 359556 204320
rect 302752 204280 302758 204292
rect 359550 204280 359556 204292
rect 359608 204280 359614 204332
rect 371602 204212 371608 204264
rect 371660 204252 371666 204264
rect 373994 204252 374000 204264
rect 371660 204224 374000 204252
rect 371660 204212 371666 204224
rect 373994 204212 374000 204224
rect 374052 204252 374058 204264
rect 375098 204252 375104 204264
rect 374052 204224 375104 204252
rect 374052 204212 374058 204224
rect 375098 204212 375104 204224
rect 375156 204212 375162 204264
rect 454218 204212 454224 204264
rect 454276 204252 454282 204264
rect 458358 204252 458364 204264
rect 454276 204224 458364 204252
rect 454276 204212 454282 204224
rect 458358 204212 458364 204224
rect 458416 204212 458422 204264
rect 369578 204008 369584 204060
rect 369636 204008 369642 204060
rect 369596 203856 369624 204008
rect 369578 203804 369584 203856
rect 369636 203804 369642 203856
rect 445018 202852 445024 202904
rect 445076 202892 445082 202904
rect 454218 202892 454224 202904
rect 445076 202864 454224 202892
rect 445076 202852 445082 202864
rect 454218 202852 454224 202864
rect 454276 202852 454282 202904
rect 3050 202784 3056 202836
rect 3108 202824 3114 202836
rect 166258 202824 166264 202836
rect 3108 202796 166264 202824
rect 3108 202784 3114 202796
rect 166258 202784 166264 202796
rect 166316 202784 166322 202836
rect 372062 202784 372068 202836
rect 372120 202824 372126 202836
rect 373074 202824 373080 202836
rect 372120 202796 373080 202824
rect 372120 202784 372126 202796
rect 373074 202784 373080 202796
rect 373132 202824 373138 202836
rect 373350 202824 373356 202836
rect 373132 202796 373356 202824
rect 373132 202784 373138 202796
rect 373350 202784 373356 202796
rect 373408 202784 373414 202836
rect 371234 202444 371240 202496
rect 371292 202484 371298 202496
rect 374638 202484 374644 202496
rect 371292 202456 374644 202484
rect 371292 202444 371298 202456
rect 374638 202444 374644 202456
rect 374696 202444 374702 202496
rect 370038 201560 370044 201612
rect 370096 201600 370102 201612
rect 373994 201600 374000 201612
rect 370096 201572 374000 201600
rect 370096 201560 370102 201572
rect 373994 201560 374000 201572
rect 374052 201560 374058 201612
rect 180242 201492 180248 201544
rect 180300 201532 180306 201544
rect 197354 201532 197360 201544
rect 180300 201504 197360 201532
rect 180300 201492 180306 201504
rect 197354 201492 197360 201504
rect 197412 201492 197418 201544
rect 302786 201492 302792 201544
rect 302844 201532 302850 201544
rect 360102 201532 360108 201544
rect 302844 201504 360108 201532
rect 302844 201492 302850 201504
rect 360102 201492 360108 201504
rect 360160 201492 360166 201544
rect 445662 201492 445668 201544
rect 445720 201532 445726 201544
rect 446398 201532 446404 201544
rect 445720 201504 446404 201532
rect 445720 201492 445726 201504
rect 446398 201492 446404 201504
rect 446456 201532 446462 201544
rect 451274 201532 451280 201544
rect 446456 201504 451280 201532
rect 446456 201492 446462 201504
rect 451274 201492 451280 201504
rect 451332 201492 451338 201544
rect 445662 200744 445668 200796
rect 445720 200784 445726 200796
rect 453298 200784 453304 200796
rect 445720 200756 453304 200784
rect 445720 200744 445726 200756
rect 453298 200744 453304 200756
rect 453356 200784 453362 200796
rect 456794 200784 456800 200796
rect 453356 200756 456800 200784
rect 453356 200744 453362 200756
rect 456794 200744 456800 200756
rect 456852 200744 456858 200796
rect 445662 199384 445668 199436
rect 445720 199424 445726 199436
rect 452654 199424 452660 199436
rect 445720 199396 452660 199424
rect 445720 199384 445726 199396
rect 452654 199384 452660 199396
rect 452712 199424 452718 199436
rect 456886 199424 456892 199436
rect 452712 199396 456892 199424
rect 452712 199384 452718 199396
rect 456886 199384 456892 199396
rect 456944 199384 456950 199436
rect 445662 198772 445668 198824
rect 445720 198812 445726 198824
rect 451366 198812 451372 198824
rect 445720 198784 451372 198812
rect 445720 198772 445726 198784
rect 451366 198772 451372 198784
rect 451424 198772 451430 198824
rect 193950 198704 193956 198756
rect 194008 198744 194014 198756
rect 198274 198744 198280 198756
rect 194008 198716 198280 198744
rect 194008 198704 194014 198716
rect 198274 198704 198280 198716
rect 198332 198704 198338 198756
rect 445386 197616 445392 197668
rect 445444 197656 445450 197668
rect 447226 197656 447232 197668
rect 445444 197628 447232 197656
rect 445444 197616 445450 197628
rect 447226 197616 447232 197628
rect 447284 197616 447290 197668
rect 173342 197344 173348 197396
rect 173400 197384 173406 197396
rect 197354 197384 197360 197396
rect 173400 197356 197360 197384
rect 173400 197344 173406 197356
rect 197354 197344 197360 197356
rect 197412 197344 197418 197396
rect 302786 197344 302792 197396
rect 302844 197384 302850 197396
rect 302844 197356 359504 197384
rect 302844 197344 302850 197356
rect 359476 197180 359504 197356
rect 441338 197276 441344 197328
rect 441396 197316 441402 197328
rect 442994 197316 443000 197328
rect 441396 197288 443000 197316
rect 441396 197276 441402 197288
rect 442994 197276 443000 197288
rect 443052 197276 443058 197328
rect 360102 197208 360108 197260
rect 360160 197248 360166 197260
rect 383746 197248 383752 197260
rect 360160 197220 383752 197248
rect 360160 197208 360166 197220
rect 383746 197208 383752 197220
rect 383804 197208 383810 197260
rect 382550 197180 382556 197192
rect 359476 197152 382556 197180
rect 382550 197140 382556 197152
rect 382608 197140 382614 197192
rect 359458 197072 359464 197124
rect 359516 197112 359522 197124
rect 378410 197112 378416 197124
rect 359516 197084 378416 197112
rect 359516 197072 359522 197084
rect 378410 197072 378416 197084
rect 378468 197072 378474 197124
rect 359550 197004 359556 197056
rect 359608 197044 359614 197056
rect 377030 197044 377036 197056
rect 359608 197016 377036 197044
rect 359608 197004 359614 197016
rect 377030 197004 377036 197016
rect 377088 197004 377094 197056
rect 382274 196732 382280 196784
rect 382332 196772 382338 196784
rect 382550 196772 382556 196784
rect 382332 196744 382556 196772
rect 382332 196732 382338 196744
rect 382550 196732 382556 196744
rect 382608 196732 382614 196784
rect 302878 195984 302884 196036
rect 302936 196024 302942 196036
rect 369486 196024 369492 196036
rect 302936 195996 369492 196024
rect 302936 195984 302942 195996
rect 369486 195984 369492 195996
rect 369544 195984 369550 196036
rect 302326 195916 302332 195968
rect 302384 195956 302390 195968
rect 302384 195928 354674 195956
rect 302384 195916 302390 195928
rect 354646 195888 354674 195928
rect 371234 195916 371240 195968
rect 371292 195956 371298 195968
rect 374086 195956 374092 195968
rect 371292 195928 374092 195956
rect 371292 195916 371298 195928
rect 374086 195916 374092 195928
rect 374144 195916 374150 195968
rect 373166 195888 373172 195900
rect 354646 195860 373172 195888
rect 373166 195848 373172 195860
rect 373224 195848 373230 195900
rect 302970 195236 302976 195288
rect 303028 195276 303034 195288
rect 372614 195276 372620 195288
rect 303028 195248 372620 195276
rect 303028 195236 303034 195248
rect 372614 195236 372620 195248
rect 372672 195276 372678 195288
rect 374178 195276 374184 195288
rect 372672 195248 374184 195276
rect 372672 195236 372678 195248
rect 374178 195236 374184 195248
rect 374236 195236 374242 195288
rect 173434 194556 173440 194608
rect 173492 194596 173498 194608
rect 197630 194596 197636 194608
rect 173492 194568 197636 194596
rect 173492 194556 173498 194568
rect 197630 194556 197636 194568
rect 197688 194556 197694 194608
rect 304258 194488 304264 194540
rect 304316 194528 304322 194540
rect 366910 194528 366916 194540
rect 304316 194500 366916 194528
rect 304316 194488 304322 194500
rect 366910 194488 366916 194500
rect 366968 194488 366974 194540
rect 436002 194488 436008 194540
rect 436060 194528 436066 194540
rect 441614 194528 441620 194540
rect 436060 194500 441620 194528
rect 436060 194488 436066 194500
rect 441614 194488 441620 194500
rect 441672 194488 441678 194540
rect 437198 194420 437204 194472
rect 437256 194460 437262 194472
rect 441706 194460 441712 194472
rect 437256 194432 441712 194460
rect 437256 194420 437262 194432
rect 441706 194420 441712 194432
rect 441764 194460 441770 194472
rect 443178 194460 443184 194472
rect 441764 194432 443184 194460
rect 441764 194420 441770 194432
rect 443178 194420 443184 194432
rect 443236 194420 443242 194472
rect 301498 193808 301504 193860
rect 301556 193848 301562 193860
rect 438946 193848 438952 193860
rect 301556 193820 438952 193848
rect 301556 193808 301562 193820
rect 438946 193808 438952 193820
rect 439004 193808 439010 193860
rect 435174 193672 435180 193724
rect 435232 193712 435238 193724
rect 436002 193712 436008 193724
rect 435232 193684 436008 193712
rect 435232 193672 435238 193684
rect 436002 193672 436008 193684
rect 436060 193672 436066 193724
rect 176102 193196 176108 193248
rect 176160 193236 176166 193248
rect 197354 193236 197360 193248
rect 176160 193208 197360 193236
rect 176160 193196 176166 193208
rect 197354 193196 197360 193208
rect 197412 193196 197418 193248
rect 171870 193128 171876 193180
rect 171928 193168 171934 193180
rect 173250 193168 173256 193180
rect 171928 193140 173256 193168
rect 171928 193128 171934 193140
rect 173250 193128 173256 193140
rect 173308 193128 173314 193180
rect 302786 193128 302792 193180
rect 302844 193168 302850 193180
rect 370406 193168 370412 193180
rect 302844 193140 370412 193168
rect 302844 193128 302850 193140
rect 370406 193128 370412 193140
rect 370464 193128 370470 193180
rect 191282 191632 191288 191684
rect 191340 191672 191346 191684
rect 198182 191672 198188 191684
rect 191340 191644 198188 191672
rect 191340 191632 191346 191644
rect 198182 191632 198188 191644
rect 198240 191632 198246 191684
rect 172422 190136 172428 190188
rect 172480 190176 172486 190188
rect 178678 190176 178684 190188
rect 172480 190148 178684 190176
rect 172480 190136 172486 190148
rect 178678 190136 178684 190148
rect 178736 190136 178742 190188
rect 183002 189048 183008 189100
rect 183060 189088 183066 189100
rect 197354 189088 197360 189100
rect 183060 189060 197360 189088
rect 183060 189048 183066 189060
rect 197354 189048 197360 189060
rect 197412 189048 197418 189100
rect 3510 188980 3516 189032
rect 3568 189020 3574 189032
rect 155218 189020 155224 189032
rect 3568 188992 155224 189020
rect 3568 188980 3574 188992
rect 155218 188980 155224 188992
rect 155276 188980 155282 189032
rect 172054 188980 172060 189032
rect 172112 189020 172118 189032
rect 181438 189020 181444 189032
rect 172112 188992 181444 189020
rect 172112 188980 172118 188992
rect 181438 188980 181444 188992
rect 181496 188980 181502 189032
rect 302786 188980 302792 189032
rect 302844 189020 302850 189032
rect 375834 189020 375840 189032
rect 302844 188992 375840 189020
rect 302844 188980 302850 188992
rect 375834 188980 375840 188992
rect 375892 188980 375898 189032
rect 172146 187620 172152 187672
rect 172204 187660 172210 187672
rect 173158 187660 173164 187672
rect 172204 187632 173164 187660
rect 172204 187620 172210 187632
rect 173158 187620 173164 187632
rect 173216 187620 173222 187672
rect 178678 186328 178684 186380
rect 178736 186368 178742 186380
rect 197354 186368 197360 186380
rect 178736 186340 197360 186368
rect 178736 186328 178742 186340
rect 197354 186328 197360 186340
rect 197412 186328 197418 186380
rect 302694 186260 302700 186312
rect 302752 186300 302758 186312
rect 374730 186300 374736 186312
rect 302752 186272 374736 186300
rect 302752 186260 302758 186272
rect 374730 186260 374736 186272
rect 374788 186300 374794 186312
rect 375282 186300 375288 186312
rect 374788 186272 375288 186300
rect 374788 186260 374794 186272
rect 375282 186260 375288 186272
rect 375340 186260 375346 186312
rect 171962 185512 171968 185564
rect 172020 185552 172026 185564
rect 180150 185552 180156 185564
rect 172020 185524 180156 185552
rect 172020 185512 172026 185524
rect 180150 185512 180156 185524
rect 180208 185512 180214 185564
rect 195422 185172 195428 185224
rect 195480 185212 195486 185224
rect 198090 185212 198096 185224
rect 195480 185184 198096 185212
rect 195480 185172 195486 185184
rect 198090 185172 198096 185184
rect 198148 185172 198154 185224
rect 172422 184832 172428 184884
rect 172480 184872 172486 184884
rect 196618 184872 196624 184884
rect 172480 184844 196624 184872
rect 172480 184832 172486 184844
rect 196618 184832 196624 184844
rect 196676 184832 196682 184884
rect 171686 184764 171692 184816
rect 171744 184804 171750 184816
rect 177298 184804 177304 184816
rect 171744 184776 177304 184804
rect 171744 184764 171750 184776
rect 177298 184764 177304 184776
rect 177356 184764 177362 184816
rect 196802 184152 196808 184204
rect 196860 184192 196866 184204
rect 198366 184192 198372 184204
rect 196860 184164 198372 184192
rect 196860 184152 196866 184164
rect 198366 184152 198372 184164
rect 198424 184152 198430 184204
rect 172422 183472 172428 183524
rect 172480 183512 172486 183524
rect 195238 183512 195244 183524
rect 172480 183484 195244 183512
rect 172480 183472 172486 183484
rect 195238 183472 195244 183484
rect 195296 183472 195302 183524
rect 181438 182792 181444 182844
rect 181496 182832 181502 182844
rect 197354 182832 197360 182844
rect 181496 182804 197360 182832
rect 181496 182792 181502 182804
rect 197354 182792 197360 182804
rect 197412 182792 197418 182844
rect 172054 182112 172060 182164
rect 172112 182152 172118 182164
rect 192478 182152 192484 182164
rect 172112 182124 192484 182152
rect 172112 182112 172118 182124
rect 192478 182112 192484 182124
rect 192536 182112 192542 182164
rect 436002 181636 436008 181688
rect 436060 181676 436066 181688
rect 441706 181676 441712 181688
rect 436060 181648 441712 181676
rect 436060 181636 436066 181648
rect 441706 181636 441712 181648
rect 441764 181636 441770 181688
rect 172422 180752 172428 180804
rect 172480 180792 172486 180804
rect 191098 180792 191104 180804
rect 172480 180764 191104 180792
rect 172480 180752 172486 180764
rect 191098 180752 191104 180764
rect 191156 180752 191162 180804
rect 302786 180072 302792 180124
rect 302844 180112 302850 180124
rect 370314 180112 370320 180124
rect 302844 180084 370320 180112
rect 302844 180072 302850 180084
rect 370314 180072 370320 180084
rect 370372 180072 370378 180124
rect 192478 179392 192484 179444
rect 192536 179432 192542 179444
rect 198366 179432 198372 179444
rect 192536 179404 198372 179432
rect 192536 179392 192542 179404
rect 198366 179392 198372 179404
rect 198424 179392 198430 179444
rect 172422 179324 172428 179376
rect 172480 179364 172486 179376
rect 188430 179364 188436 179376
rect 172480 179336 188436 179364
rect 172480 179324 172486 179336
rect 188430 179324 188436 179336
rect 188488 179324 188494 179376
rect 318058 179324 318064 179376
rect 318116 179364 318122 179376
rect 580166 179364 580172 179376
rect 318116 179336 580172 179364
rect 318116 179324 318122 179336
rect 580166 179324 580172 179336
rect 580224 179324 580230 179376
rect 188522 178032 188528 178084
rect 188580 178072 188586 178084
rect 197354 178072 197360 178084
rect 188580 178044 197360 178072
rect 188580 178032 188586 178044
rect 197354 178032 197360 178044
rect 197412 178032 197418 178084
rect 172422 177964 172428 178016
rect 172480 178004 172486 178016
rect 187050 178004 187056 178016
rect 172480 177976 187056 178004
rect 172480 177964 172486 177976
rect 187050 177964 187056 177976
rect 187108 177964 187114 178016
rect 172330 177896 172336 177948
rect 172388 177936 172394 177948
rect 184290 177936 184296 177948
rect 172388 177908 184296 177936
rect 172388 177896 172394 177908
rect 184290 177896 184296 177908
rect 184348 177896 184354 177948
rect 172238 176604 172244 176656
rect 172296 176644 172302 176656
rect 182818 176644 182824 176656
rect 172296 176616 182824 176644
rect 172296 176604 172302 176616
rect 182818 176604 182824 176616
rect 182876 176604 182882 176656
rect 302786 175924 302792 175976
rect 302844 175964 302850 175976
rect 370130 175964 370136 175976
rect 302844 175936 370136 175964
rect 302844 175924 302850 175936
rect 370130 175924 370136 175936
rect 370188 175964 370194 175976
rect 370774 175964 370780 175976
rect 370188 175936 370780 175964
rect 370188 175924 370194 175936
rect 370774 175924 370780 175936
rect 370832 175924 370838 175976
rect 177298 175244 177304 175296
rect 177356 175284 177362 175296
rect 197630 175284 197636 175296
rect 177356 175256 197636 175284
rect 177356 175244 177362 175256
rect 197630 175244 197636 175256
rect 197688 175244 197694 175296
rect 172422 175176 172428 175228
rect 172480 175216 172486 175228
rect 181530 175216 181536 175228
rect 172480 175188 181536 175216
rect 172480 175176 172486 175188
rect 181530 175176 181536 175188
rect 181588 175176 181594 175228
rect 370590 175176 370596 175228
rect 370648 175216 370654 175228
rect 375742 175216 375748 175228
rect 370648 175188 375748 175216
rect 370648 175176 370654 175188
rect 375742 175176 375748 175188
rect 375800 175216 375806 175228
rect 448606 175216 448612 175228
rect 375800 175188 448612 175216
rect 375800 175176 375806 175188
rect 448606 175176 448612 175188
rect 448664 175176 448670 175228
rect 184290 173884 184296 173936
rect 184348 173924 184354 173936
rect 197354 173924 197360 173936
rect 184348 173896 197360 173924
rect 184348 173884 184354 173896
rect 197354 173884 197360 173896
rect 197412 173884 197418 173936
rect 172422 173612 172428 173664
rect 172480 173652 172486 173664
rect 180058 173652 180064 173664
rect 172480 173624 180064 173652
rect 172480 173612 172486 173624
rect 180058 173612 180064 173624
rect 180116 173612 180122 173664
rect 180150 173136 180156 173188
rect 180208 173176 180214 173188
rect 198090 173176 198096 173188
rect 180208 173148 198096 173176
rect 180208 173136 180214 173148
rect 198090 173136 198096 173148
rect 198148 173136 198154 173188
rect 374546 172456 374552 172508
rect 374604 172496 374610 172508
rect 450170 172496 450176 172508
rect 374604 172468 450176 172496
rect 374604 172456 374610 172468
rect 450170 172456 450176 172468
rect 450228 172456 450234 172508
rect 172422 172388 172428 172440
rect 172480 172428 172486 172440
rect 178770 172428 178776 172440
rect 172480 172400 178776 172428
rect 172480 172388 172486 172400
rect 178770 172388 178776 172400
rect 178828 172388 178834 172440
rect 369670 171096 369676 171148
rect 369728 171136 369734 171148
rect 374546 171136 374552 171148
rect 369728 171108 374552 171136
rect 369728 171096 369734 171108
rect 374546 171096 374552 171108
rect 374604 171096 374610 171148
rect 172238 171028 172244 171080
rect 172296 171068 172302 171080
rect 197998 171068 198004 171080
rect 172296 171040 198004 171068
rect 172296 171028 172302 171040
rect 197998 171028 198004 171040
rect 198056 171028 198062 171080
rect 302786 170348 302792 170400
rect 302844 170388 302850 170400
rect 370590 170388 370596 170400
rect 302844 170360 370596 170388
rect 302844 170348 302850 170360
rect 370590 170348 370596 170360
rect 370648 170348 370654 170400
rect 172238 168988 172244 169040
rect 172296 169028 172302 169040
rect 193858 169028 193864 169040
rect 172296 169000 193864 169028
rect 172296 168988 172302 169000
rect 193858 168988 193864 169000
rect 193916 168988 193922 169040
rect 446122 168416 446128 168428
rect 371252 168388 446128 168416
rect 172422 168308 172428 168360
rect 172480 168348 172486 168360
rect 191190 168348 191196 168360
rect 172480 168320 191196 168348
rect 172480 168308 172486 168320
rect 191190 168308 191196 168320
rect 191248 168308 191254 168360
rect 370038 168308 370044 168360
rect 370096 168348 370102 168360
rect 371252 168348 371280 168388
rect 446122 168376 446128 168388
rect 446180 168376 446186 168428
rect 370096 168320 371280 168348
rect 370096 168308 370102 168320
rect 369118 167900 369124 167952
rect 369176 167940 369182 167952
rect 370038 167940 370044 167952
rect 369176 167912 370044 167940
rect 369176 167900 369182 167912
rect 370038 167900 370044 167912
rect 370096 167900 370102 167952
rect 449986 167056 449992 167068
rect 371252 167028 449992 167056
rect 369302 166948 369308 167000
rect 369360 166988 369366 167000
rect 370498 166988 370504 167000
rect 369360 166960 370504 166988
rect 369360 166948 369366 166960
rect 370498 166948 370504 166960
rect 370556 166988 370562 167000
rect 371252 166988 371280 167028
rect 449986 167016 449992 167028
rect 450044 167016 450050 167068
rect 370556 166960 371280 166988
rect 370556 166948 370562 166960
rect 178770 166336 178776 166388
rect 178828 166376 178834 166388
rect 197722 166376 197728 166388
rect 178828 166348 197728 166376
rect 178828 166336 178834 166348
rect 197722 166336 197728 166348
rect 197780 166336 197786 166388
rect 171778 166268 171784 166320
rect 171836 166308 171842 166320
rect 192478 166308 192484 166320
rect 171836 166280 192484 166308
rect 171836 166268 171842 166280
rect 192478 166268 192484 166280
rect 192536 166268 192542 166320
rect 172054 165520 172060 165572
rect 172112 165560 172118 165572
rect 192570 165560 192576 165572
rect 172112 165532 192576 165560
rect 172112 165520 172118 165532
rect 192570 165520 192576 165532
rect 192628 165520 192634 165572
rect 192478 164500 192484 164552
rect 192536 164540 192542 164552
rect 197538 164540 197544 164552
rect 192536 164512 197544 164540
rect 192536 164500 192542 164512
rect 197538 164500 197544 164512
rect 197596 164500 197602 164552
rect 448698 164268 448704 164280
rect 370516 164240 448704 164268
rect 370516 164212 370544 164240
rect 448698 164228 448704 164240
rect 448756 164228 448762 164280
rect 3234 164160 3240 164212
rect 3292 164200 3298 164212
rect 88978 164200 88984 164212
rect 3292 164172 88984 164200
rect 3292 164160 3298 164172
rect 88978 164160 88984 164172
rect 89036 164160 89042 164212
rect 172422 164160 172428 164212
rect 172480 164200 172486 164212
rect 195330 164200 195336 164212
rect 172480 164172 195336 164200
rect 172480 164160 172486 164172
rect 195330 164160 195336 164172
rect 195388 164160 195394 164212
rect 370222 164160 370228 164212
rect 370280 164200 370286 164212
rect 370498 164200 370504 164212
rect 370280 164172 370504 164200
rect 370280 164160 370286 164172
rect 370498 164160 370504 164172
rect 370556 164160 370562 164212
rect 370590 164160 370596 164212
rect 370648 164200 370654 164212
rect 372890 164200 372896 164212
rect 370648 164172 372896 164200
rect 370648 164160 370654 164172
rect 372890 164160 372896 164172
rect 372948 164200 372954 164212
rect 452838 164200 452844 164212
rect 372948 164172 452844 164200
rect 372948 164160 372954 164172
rect 452838 164160 452844 164172
rect 452896 164160 452902 164212
rect 172146 162800 172152 162852
rect 172204 162840 172210 162852
rect 172204 162812 180794 162840
rect 172204 162800 172210 162812
rect 180766 162772 180794 162812
rect 196618 162800 196624 162852
rect 196676 162840 196682 162852
rect 198182 162840 198188 162852
rect 196676 162812 198188 162840
rect 196676 162800 196682 162812
rect 198182 162800 198188 162812
rect 198240 162800 198246 162852
rect 196710 162772 196716 162784
rect 180766 162744 196716 162772
rect 196710 162732 196716 162744
rect 196768 162732 196774 162784
rect 373258 162120 373264 162172
rect 373316 162160 373322 162172
rect 454126 162160 454132 162172
rect 373316 162132 454132 162160
rect 373316 162120 373322 162132
rect 454126 162120 454132 162132
rect 454184 162120 454190 162172
rect 303062 161372 303068 161424
rect 303120 161412 303126 161424
rect 369762 161412 369768 161424
rect 303120 161384 369768 161412
rect 303120 161372 303126 161384
rect 369762 161372 369768 161384
rect 369820 161412 369826 161424
rect 370222 161412 370228 161424
rect 369820 161384 370228 161412
rect 369820 161372 369826 161384
rect 370222 161372 370228 161384
rect 370280 161372 370286 161424
rect 172422 161168 172428 161220
rect 172480 161208 172486 161220
rect 177390 161208 177396 161220
rect 172480 161180 177396 161208
rect 172480 161168 172486 161180
rect 177390 161168 177396 161180
rect 177448 161168 177454 161220
rect 169202 160760 169208 160812
rect 169260 160800 169266 160812
rect 175918 160800 175924 160812
rect 169260 160772 175924 160800
rect 169260 160760 169266 160772
rect 175918 160760 175924 160772
rect 175976 160760 175982 160812
rect 198734 160732 198740 160744
rect 171106 160704 198740 160732
rect 165154 160488 165160 160540
rect 165212 160528 165218 160540
rect 171106 160528 171134 160704
rect 198734 160692 198740 160704
rect 198792 160692 198798 160744
rect 372614 160692 372620 160744
rect 372672 160732 372678 160744
rect 373350 160732 373356 160744
rect 372672 160704 373356 160732
rect 372672 160692 372678 160704
rect 373350 160692 373356 160704
rect 373408 160732 373414 160744
rect 445938 160732 445944 160744
rect 373408 160704 445944 160732
rect 373408 160692 373414 160704
rect 445938 160692 445944 160704
rect 445996 160692 446002 160744
rect 165212 160500 171134 160528
rect 165212 160488 165218 160500
rect 177482 160080 177488 160132
rect 177540 160120 177546 160132
rect 197538 160120 197544 160132
rect 177540 160092 197544 160120
rect 177540 160080 177546 160092
rect 197538 160080 197544 160092
rect 197596 160080 197602 160132
rect 192570 158788 192576 158840
rect 192628 158828 192634 158840
rect 197354 158828 197360 158840
rect 192628 158800 197360 158828
rect 192628 158788 192634 158800
rect 197354 158788 197360 158800
rect 197412 158788 197418 158840
rect 162854 158652 162860 158704
rect 162912 158692 162918 158704
rect 176010 158692 176016 158704
rect 162912 158664 176016 158692
rect 162912 158652 162918 158664
rect 176010 158652 176016 158664
rect 176068 158652 176074 158704
rect 369394 158652 369400 158704
rect 369452 158692 369458 158704
rect 373902 158692 373908 158704
rect 369452 158664 373908 158692
rect 369452 158652 369458 158664
rect 373902 158652 373908 158664
rect 373960 158692 373966 158704
rect 448514 158692 448520 158704
rect 373960 158664 448520 158692
rect 373960 158652 373966 158664
rect 448514 158652 448520 158664
rect 448572 158652 448578 158704
rect 166902 157972 166908 158024
rect 166960 158012 166966 158024
rect 195238 158012 195244 158024
rect 166960 157984 195244 158012
rect 166960 157972 166966 157984
rect 195238 157972 195244 157984
rect 195296 157972 195302 158024
rect 372062 156680 372068 156732
rect 372120 156720 372126 156732
rect 444466 156720 444472 156732
rect 372120 156692 444472 156720
rect 372120 156680 372126 156692
rect 444466 156680 444472 156692
rect 444524 156680 444530 156732
rect 171962 156612 171968 156664
rect 172020 156652 172026 156664
rect 188522 156652 188528 156664
rect 172020 156624 188528 156652
rect 172020 156612 172026 156624
rect 188522 156612 188528 156624
rect 188580 156612 188586 156664
rect 309778 156612 309784 156664
rect 309836 156652 309842 156664
rect 579614 156652 579620 156664
rect 309836 156624 579620 156652
rect 309836 156612 309842 156624
rect 579614 156612 579620 156624
rect 579672 156612 579678 156664
rect 191098 155932 191104 155984
rect 191156 155972 191162 155984
rect 197814 155972 197820 155984
rect 191156 155944 197820 155972
rect 191156 155932 191162 155944
rect 197814 155932 197820 155944
rect 197872 155932 197878 155984
rect 302878 155864 302884 155916
rect 302936 155904 302942 155916
rect 369578 155904 369584 155916
rect 302936 155876 369584 155904
rect 302936 155864 302942 155876
rect 369578 155864 369584 155876
rect 369636 155904 369642 155916
rect 370866 155904 370872 155916
rect 369636 155876 370872 155904
rect 369636 155864 369642 155876
rect 370866 155864 370872 155876
rect 370924 155864 370930 155916
rect 444558 155864 444564 155916
rect 444616 155904 444622 155916
rect 447318 155904 447324 155916
rect 444616 155876 447324 155904
rect 444616 155864 444622 155876
rect 447318 155864 447324 155876
rect 447376 155864 447382 155916
rect 182818 154572 182824 154624
rect 182876 154612 182882 154624
rect 197354 154612 197360 154624
rect 182876 154584 197360 154612
rect 182876 154572 182882 154584
rect 197354 154572 197360 154584
rect 197412 154572 197418 154624
rect 374638 154572 374644 154624
rect 374696 154612 374702 154624
rect 444558 154612 444564 154624
rect 374696 154584 444564 154612
rect 374696 154572 374702 154584
rect 444558 154572 444564 154584
rect 444616 154572 444622 154624
rect 171594 154504 171600 154556
rect 171652 154544 171658 154556
rect 174538 154544 174544 154556
rect 171652 154516 174544 154544
rect 171652 154504 171658 154516
rect 174538 154504 174544 154516
rect 174596 154504 174602 154556
rect 371970 154504 371976 154556
rect 372028 154544 372034 154556
rect 385126 154544 385132 154556
rect 372028 154516 385132 154544
rect 372028 154504 372034 154516
rect 385126 154504 385132 154516
rect 385184 154504 385190 154556
rect 371418 154436 371424 154488
rect 371476 154476 371482 154488
rect 381078 154476 381084 154488
rect 371476 154448 381084 154476
rect 371476 154436 371482 154448
rect 381078 154436 381084 154448
rect 381136 154436 381142 154488
rect 444926 154028 444932 154080
rect 444984 154068 444990 154080
rect 449894 154068 449900 154080
rect 444984 154040 449900 154068
rect 444984 154028 444990 154040
rect 449894 154028 449900 154040
rect 449952 154028 449958 154080
rect 171686 153756 171692 153808
rect 171744 153796 171750 153808
rect 174630 153796 174636 153808
rect 171744 153768 174636 153796
rect 171744 153756 171750 153768
rect 174630 153756 174636 153768
rect 174688 153756 174694 153808
rect 444374 153388 444380 153400
rect 431926 153360 444380 153388
rect 370866 153280 370872 153332
rect 370924 153320 370930 153332
rect 431926 153320 431954 153360
rect 444374 153348 444380 153360
rect 444432 153388 444438 153400
rect 452746 153388 452752 153400
rect 444432 153360 452752 153388
rect 444432 153348 444438 153360
rect 452746 153348 452752 153360
rect 452804 153348 452810 153400
rect 370924 153292 431954 153320
rect 370924 153280 370930 153292
rect 370222 153212 370228 153264
rect 370280 153252 370286 153264
rect 441798 153252 441804 153264
rect 370280 153224 441804 153252
rect 370280 153212 370286 153224
rect 441798 153212 441804 153224
rect 441856 153252 441862 153264
rect 445294 153252 445300 153264
rect 441856 153224 445300 153252
rect 441856 153212 441862 153224
rect 445294 153212 445300 153224
rect 445352 153212 445358 153264
rect 171594 153144 171600 153196
rect 171652 153184 171658 153196
rect 174722 153184 174728 153196
rect 171652 153156 174728 153184
rect 171652 153144 171658 153156
rect 174722 153144 174728 153156
rect 174780 153144 174786 153196
rect 302510 153144 302516 153196
rect 302568 153184 302574 153196
rect 302568 153156 368152 153184
rect 302568 153144 302574 153156
rect 302602 153076 302608 153128
rect 302660 153116 302666 153128
rect 302660 153088 367968 153116
rect 302660 153076 302666 153088
rect 302786 153008 302792 153060
rect 302844 153048 302850 153060
rect 302844 153020 354674 153048
rect 302844 153008 302850 153020
rect 354646 152844 354674 153020
rect 367940 152912 367968 153088
rect 368124 153048 368152 153156
rect 369302 153144 369308 153196
rect 369360 153184 369366 153196
rect 369578 153184 369584 153196
rect 369360 153156 369584 153184
rect 369360 153144 369366 153156
rect 369578 153144 369584 153156
rect 369636 153144 369642 153196
rect 370130 153144 370136 153196
rect 370188 153184 370194 153196
rect 370590 153184 370596 153196
rect 370188 153156 370596 153184
rect 370188 153144 370194 153156
rect 370590 153144 370596 153156
rect 370648 153144 370654 153196
rect 371878 153144 371884 153196
rect 371936 153184 371942 153196
rect 383654 153184 383660 153196
rect 371936 153156 383660 153184
rect 371936 153144 371942 153156
rect 383654 153144 383660 153156
rect 383712 153144 383718 153196
rect 445662 153144 445668 153196
rect 445720 153184 445726 153196
rect 458266 153184 458272 153196
rect 445720 153156 458272 153184
rect 445720 153144 445726 153156
rect 458266 153144 458272 153156
rect 458324 153144 458330 153196
rect 371418 153076 371424 153128
rect 371476 153116 371482 153128
rect 379514 153116 379520 153128
rect 371476 153088 379520 153116
rect 371476 153076 371482 153088
rect 379514 153076 379520 153088
rect 379572 153076 379578 153128
rect 370038 153048 370044 153060
rect 368124 153020 370044 153048
rect 370038 153008 370044 153020
rect 370096 153008 370102 153060
rect 369670 152912 369676 152924
rect 367940 152884 369676 152912
rect 369670 152872 369676 152884
rect 369728 152872 369734 152924
rect 369302 152844 369308 152856
rect 354646 152816 369308 152844
rect 369302 152804 369308 152816
rect 369360 152804 369366 152856
rect 359458 152124 359464 152176
rect 359516 152164 359522 152176
rect 369118 152164 369124 152176
rect 359516 152136 369124 152164
rect 359516 152124 359522 152136
rect 369118 152124 369124 152136
rect 369176 152164 369182 152176
rect 372614 152164 372620 152176
rect 369176 152136 372620 152164
rect 369176 152124 369182 152136
rect 372614 152124 372620 152136
rect 372672 152124 372678 152176
rect 358906 152056 358912 152108
rect 358964 152096 358970 152108
rect 369210 152096 369216 152108
rect 358964 152068 369216 152096
rect 358964 152056 358970 152068
rect 369210 152056 369216 152068
rect 369268 152096 369274 152108
rect 374638 152096 374644 152108
rect 369268 152068 374644 152096
rect 369268 152056 369274 152068
rect 374638 152056 374644 152068
rect 374696 152056 374702 152108
rect 360102 151988 360108 152040
rect 360160 152028 360166 152040
rect 369394 152028 369400 152040
rect 360160 152000 369400 152028
rect 360160 151988 360166 152000
rect 369394 151988 369400 152000
rect 369452 151988 369458 152040
rect 359550 151920 359556 151972
rect 359608 151960 359614 151972
rect 369578 151960 369584 151972
rect 359608 151932 369584 151960
rect 359608 151920 359614 151932
rect 369578 151920 369584 151932
rect 369636 151920 369642 151972
rect 370130 151892 370136 151904
rect 360120 151864 370136 151892
rect 175918 151784 175924 151836
rect 175976 151824 175982 151836
rect 197354 151824 197360 151836
rect 175976 151796 197360 151824
rect 175976 151784 175982 151796
rect 197354 151784 197360 151796
rect 197412 151784 197418 151836
rect 172238 151716 172244 151768
rect 172296 151756 172302 151768
rect 191282 151756 191288 151768
rect 172296 151728 191288 151756
rect 172296 151716 172302 151728
rect 191282 151716 191288 151728
rect 191340 151716 191346 151768
rect 302694 151716 302700 151768
rect 302752 151756 302758 151768
rect 360120 151756 360148 151864
rect 370130 151852 370136 151864
rect 370188 151852 370194 151904
rect 302752 151728 360148 151756
rect 302752 151716 302758 151728
rect 371418 151716 371424 151768
rect 371476 151756 371482 151768
rect 374914 151756 374920 151768
rect 371476 151728 374920 151756
rect 371476 151716 371482 151728
rect 374914 151716 374920 151728
rect 374972 151716 374978 151768
rect 444926 151716 444932 151768
rect 444984 151756 444990 151768
rect 454034 151756 454040 151768
rect 444984 151728 454040 151756
rect 444984 151716 444990 151728
rect 454034 151716 454040 151728
rect 454092 151716 454098 151768
rect 172422 151648 172428 151700
rect 172480 151688 172486 151700
rect 182910 151688 182916 151700
rect 172480 151660 182916 151688
rect 172480 151648 172486 151660
rect 182910 151648 182916 151660
rect 182968 151648 182974 151700
rect 171686 151580 171692 151632
rect 171744 151620 171750 151632
rect 181622 151620 181628 151632
rect 171744 151592 181628 151620
rect 171744 151580 171750 151592
rect 181622 151580 181628 151592
rect 181680 151580 181686 151632
rect 371970 151580 371976 151632
rect 372028 151620 372034 151632
rect 378318 151620 378324 151632
rect 372028 151592 378324 151620
rect 372028 151580 372034 151592
rect 378318 151580 378324 151592
rect 378376 151580 378382 151632
rect 371418 150900 371424 150952
rect 371476 150940 371482 150952
rect 375650 150940 375656 150952
rect 371476 150912 375656 150940
rect 371476 150900 371482 150912
rect 375650 150900 375656 150912
rect 375708 150900 375714 150952
rect 3510 150356 3516 150408
rect 3568 150396 3574 150408
rect 148318 150396 148324 150408
rect 3568 150368 148324 150396
rect 3568 150356 3574 150368
rect 148318 150356 148324 150368
rect 148376 150356 148382 150408
rect 172422 150356 172428 150408
rect 172480 150396 172486 150408
rect 193950 150396 193956 150408
rect 172480 150368 193956 150396
rect 172480 150356 172486 150368
rect 193950 150356 193956 150368
rect 194008 150356 194014 150408
rect 371970 150356 371976 150408
rect 372028 150396 372034 150408
rect 385034 150396 385040 150408
rect 372028 150368 385040 150396
rect 372028 150356 372034 150368
rect 385034 150356 385040 150368
rect 385092 150356 385098 150408
rect 371418 150288 371424 150340
rect 371476 150328 371482 150340
rect 382458 150328 382464 150340
rect 371476 150300 382464 150328
rect 371476 150288 371482 150300
rect 382458 150288 382464 150300
rect 382516 150288 382522 150340
rect 444926 150152 444932 150204
rect 444984 150192 444990 150204
rect 448606 150192 448612 150204
rect 444984 150164 448612 150192
rect 444984 150152 444990 150164
rect 448606 150152 448612 150164
rect 448664 150152 448670 150204
rect 171502 149744 171508 149796
rect 171560 149784 171566 149796
rect 180242 149784 180248 149796
rect 171560 149756 180248 149784
rect 171560 149744 171566 149756
rect 180242 149744 180248 149756
rect 180300 149744 180306 149796
rect 174538 149064 174544 149116
rect 174596 149104 174602 149116
rect 197354 149104 197360 149116
rect 174596 149076 197360 149104
rect 174596 149064 174602 149076
rect 197354 149064 197360 149076
rect 197412 149064 197418 149116
rect 302326 148996 302332 149048
rect 302384 149036 302390 149048
rect 360102 149036 360108 149048
rect 302384 149008 360108 149036
rect 302384 148996 302390 149008
rect 360102 148996 360108 149008
rect 360160 148996 360166 149048
rect 371970 148996 371976 149048
rect 372028 149036 372034 149048
rect 382366 149036 382372 149048
rect 372028 149008 382372 149036
rect 372028 148996 372034 149008
rect 382366 148996 382372 149008
rect 382424 148996 382430 149048
rect 445294 148996 445300 149048
rect 445352 149036 445358 149048
rect 456978 149036 456984 149048
rect 445352 149008 456984 149036
rect 445352 148996 445358 149008
rect 456978 148996 456984 149008
rect 457036 148996 457042 149048
rect 371418 148928 371424 148980
rect 371476 148968 371482 148980
rect 380894 148968 380900 148980
rect 371476 148940 380900 148968
rect 371476 148928 371482 148940
rect 380894 148928 380900 148940
rect 380952 148928 380958 148980
rect 172422 148860 172428 148912
rect 172480 148900 172486 148912
rect 195422 148900 195428 148912
rect 172480 148872 195428 148900
rect 172480 148860 172486 148872
rect 195422 148860 195428 148872
rect 195480 148860 195486 148912
rect 171686 148316 171692 148368
rect 171744 148356 171750 148368
rect 173342 148356 173348 148368
rect 171744 148328 173348 148356
rect 171744 148316 171750 148328
rect 173342 148316 173348 148328
rect 173400 148316 173406 148368
rect 198090 148356 198096 148368
rect 180766 148328 198096 148356
rect 173158 148248 173164 148300
rect 173216 148288 173222 148300
rect 180766 148288 180794 148328
rect 198090 148316 198096 148328
rect 198148 148316 198154 148368
rect 173216 148260 180794 148288
rect 173216 148248 173222 148260
rect 171502 147976 171508 148028
rect 171560 148016 171566 148028
rect 173434 148016 173440 148028
rect 171560 147988 173440 148016
rect 171560 147976 171566 147988
rect 173434 147976 173440 147988
rect 173492 147976 173498 148028
rect 181530 147636 181536 147688
rect 181588 147676 181594 147688
rect 197354 147676 197360 147688
rect 181588 147648 197360 147676
rect 181588 147636 181594 147648
rect 197354 147636 197360 147648
rect 197412 147636 197418 147688
rect 172330 147568 172336 147620
rect 172388 147608 172394 147620
rect 196802 147608 196808 147620
rect 172388 147580 196808 147608
rect 172388 147568 172394 147580
rect 196802 147568 196808 147580
rect 196860 147568 196866 147620
rect 371970 147568 371976 147620
rect 372028 147608 372034 147620
rect 380986 147608 380992 147620
rect 372028 147580 380992 147608
rect 372028 147568 372034 147580
rect 380986 147568 380992 147580
rect 381044 147568 381050 147620
rect 171686 147500 171692 147552
rect 171744 147540 171750 147552
rect 176102 147540 176108 147552
rect 171744 147512 176108 147540
rect 171744 147500 171750 147512
rect 176102 147500 176108 147512
rect 176160 147500 176166 147552
rect 371418 147500 371424 147552
rect 371476 147540 371482 147552
rect 378226 147540 378232 147552
rect 371476 147512 378232 147540
rect 371476 147500 371482 147512
rect 378226 147500 378232 147512
rect 378284 147500 378290 147552
rect 444374 146548 444380 146600
rect 444432 146588 444438 146600
rect 446122 146588 446128 146600
rect 444432 146560 446128 146588
rect 444432 146548 444438 146560
rect 446122 146548 446128 146560
rect 446180 146548 446186 146600
rect 172422 146208 172428 146260
rect 172480 146248 172486 146260
rect 183002 146248 183008 146260
rect 172480 146220 183008 146248
rect 172480 146208 172486 146220
rect 183002 146208 183008 146220
rect 183060 146208 183066 146260
rect 195330 146208 195336 146260
rect 195388 146248 195394 146260
rect 197998 146248 198004 146260
rect 195388 146220 198004 146248
rect 195388 146208 195394 146220
rect 197998 146208 198004 146220
rect 198056 146208 198062 146260
rect 302786 146208 302792 146260
rect 302844 146248 302850 146260
rect 358906 146248 358912 146260
rect 302844 146220 358912 146248
rect 302844 146208 302850 146220
rect 358906 146208 358912 146220
rect 358964 146208 358970 146260
rect 445662 146208 445668 146260
rect 445720 146248 445726 146260
rect 454126 146248 454132 146260
rect 445720 146220 454132 146248
rect 445720 146208 445726 146220
rect 454126 146208 454132 146220
rect 454184 146208 454190 146260
rect 171686 146140 171692 146192
rect 171744 146180 171750 146192
rect 181438 146180 181444 146192
rect 171744 146152 181444 146180
rect 171744 146140 171750 146152
rect 181438 146140 181444 146152
rect 181496 146140 181502 146192
rect 371418 146140 371424 146192
rect 371476 146180 371482 146192
rect 375926 146180 375932 146192
rect 371476 146152 375932 146180
rect 371476 146140 371482 146152
rect 375926 146140 375932 146152
rect 375984 146140 375990 146192
rect 371970 146072 371976 146124
rect 372028 146112 372034 146124
rect 376938 146112 376944 146124
rect 372028 146084 376944 146112
rect 372028 146072 372034 146084
rect 376938 146072 376944 146084
rect 376996 146072 377002 146124
rect 371418 145868 371424 145920
rect 371476 145908 371482 145920
rect 374362 145908 374368 145920
rect 371476 145880 374368 145908
rect 371476 145868 371482 145880
rect 374362 145868 374368 145880
rect 374420 145868 374426 145920
rect 172422 145732 172428 145784
rect 172480 145772 172486 145784
rect 178678 145772 178684 145784
rect 172480 145744 178684 145772
rect 172480 145732 172486 145744
rect 178678 145732 178684 145744
rect 178736 145732 178742 145784
rect 171686 144848 171692 144900
rect 171744 144888 171750 144900
rect 180150 144888 180156 144900
rect 171744 144860 180156 144888
rect 171744 144848 171750 144860
rect 180150 144848 180156 144860
rect 180208 144848 180214 144900
rect 445294 144780 445300 144832
rect 445352 144820 445358 144832
rect 450078 144820 450084 144832
rect 445352 144792 450084 144820
rect 445352 144780 445358 144792
rect 450078 144780 450084 144792
rect 450136 144780 450142 144832
rect 371418 144712 371424 144764
rect 371476 144752 371482 144764
rect 378134 144752 378140 144764
rect 371476 144724 378140 144752
rect 371476 144712 371482 144724
rect 378134 144712 378140 144724
rect 378192 144712 378198 144764
rect 371418 144236 371424 144288
rect 371476 144276 371482 144288
rect 375558 144276 375564 144288
rect 371476 144248 375564 144276
rect 371476 144236 371482 144248
rect 375558 144236 375564 144248
rect 375616 144236 375622 144288
rect 171870 144032 171876 144084
rect 171928 144072 171934 144084
rect 177298 144072 177304 144084
rect 171928 144044 177304 144072
rect 171928 144032 171934 144044
rect 177298 144032 177304 144044
rect 177356 144032 177362 144084
rect 371418 143896 371424 143948
rect 371476 143936 371482 143948
rect 375006 143936 375012 143948
rect 371476 143908 375012 143936
rect 371476 143896 371482 143908
rect 375006 143896 375012 143908
rect 375064 143896 375070 143948
rect 179414 143556 179420 143608
rect 179472 143596 179478 143608
rect 197354 143596 197360 143608
rect 179472 143568 197360 143596
rect 179472 143556 179478 143568
rect 197354 143556 197360 143568
rect 197412 143556 197418 143608
rect 172422 143488 172428 143540
rect 172480 143528 172486 143540
rect 184290 143528 184296 143540
rect 172480 143500 184296 143528
rect 172480 143488 172486 143500
rect 184290 143488 184296 143500
rect 184348 143488 184354 143540
rect 371970 143488 371976 143540
rect 372028 143528 372034 143540
rect 385218 143528 385224 143540
rect 372028 143500 385224 143528
rect 372028 143488 372034 143500
rect 385218 143488 385224 143500
rect 385276 143488 385282 143540
rect 371418 143420 371424 143472
rect 371476 143460 371482 143472
rect 378410 143460 378416 143472
rect 371476 143432 378416 143460
rect 371476 143420 371482 143432
rect 378410 143420 378416 143432
rect 378468 143420 378474 143472
rect 445202 142196 445208 142248
rect 445260 142236 445266 142248
rect 452838 142236 452844 142248
rect 445260 142208 452844 142236
rect 445260 142196 445266 142208
rect 452838 142196 452844 142208
rect 452896 142196 452902 142248
rect 172422 142060 172428 142112
rect 172480 142100 172486 142112
rect 196618 142100 196624 142112
rect 172480 142072 196624 142100
rect 172480 142060 172486 142072
rect 196618 142060 196624 142072
rect 196676 142060 196682 142112
rect 302786 142060 302792 142112
rect 302844 142100 302850 142112
rect 359550 142100 359556 142112
rect 302844 142072 359556 142100
rect 302844 142060 302850 142072
rect 359550 142060 359556 142072
rect 359608 142060 359614 142112
rect 371970 142060 371976 142112
rect 372028 142100 372034 142112
rect 383746 142100 383752 142112
rect 372028 142072 383752 142100
rect 372028 142060 372034 142072
rect 383746 142060 383752 142072
rect 383804 142060 383810 142112
rect 172330 141992 172336 142044
rect 172388 142032 172394 142044
rect 192478 142032 192484 142044
rect 172388 142004 192484 142032
rect 172388 141992 172394 142004
rect 192478 141992 192484 142004
rect 192536 141992 192542 142044
rect 372062 141992 372068 142044
rect 372120 142032 372126 142044
rect 382274 142032 382280 142044
rect 372120 142004 382280 142032
rect 372120 141992 372126 142004
rect 382274 141992 382280 142004
rect 382332 141992 382338 142044
rect 371418 141924 371424 141976
rect 371476 141964 371482 141976
rect 377030 141964 377036 141976
rect 371476 141936 377036 141964
rect 371476 141924 371482 141936
rect 377030 141924 377036 141936
rect 377088 141924 377094 141976
rect 445110 141924 445116 141976
rect 445168 141964 445174 141976
rect 448514 141964 448520 141976
rect 445168 141936 448520 141964
rect 445168 141924 445174 141936
rect 448514 141924 448520 141936
rect 448572 141924 448578 141976
rect 171870 141788 171876 141840
rect 171928 141828 171934 141840
rect 178770 141828 178776 141840
rect 171928 141800 178776 141828
rect 171928 141788 171934 141800
rect 178770 141788 178776 141800
rect 178828 141788 178834 141840
rect 178034 140768 178040 140820
rect 178092 140808 178098 140820
rect 197538 140808 197544 140820
rect 178092 140780 197544 140808
rect 178092 140768 178098 140780
rect 197538 140768 197544 140780
rect 197596 140768 197602 140820
rect 172422 140700 172428 140752
rect 172480 140740 172486 140752
rect 195330 140740 195336 140752
rect 172480 140712 195336 140740
rect 172480 140700 172486 140712
rect 195330 140700 195336 140712
rect 195388 140700 195394 140752
rect 371418 140632 371424 140684
rect 371476 140672 371482 140684
rect 376846 140672 376852 140684
rect 371476 140644 376852 140672
rect 371476 140632 371482 140644
rect 376846 140632 376852 140644
rect 376904 140632 376910 140684
rect 445110 140360 445116 140412
rect 445168 140400 445174 140412
rect 449986 140400 449992 140412
rect 445168 140372 449992 140400
rect 445168 140360 445174 140372
rect 449986 140360 449992 140372
rect 450044 140360 450050 140412
rect 172146 140292 172152 140344
rect 172204 140332 172210 140344
rect 173158 140332 173164 140344
rect 172204 140304 173164 140332
rect 172204 140292 172210 140304
rect 173158 140292 173164 140304
rect 173216 140292 173222 140344
rect 371970 140292 371976 140344
rect 372028 140332 372034 140344
rect 373166 140332 373172 140344
rect 372028 140304 373172 140332
rect 372028 140292 372034 140304
rect 373166 140292 373172 140304
rect 373224 140292 373230 140344
rect 171318 140020 171324 140072
rect 171376 140060 171382 140072
rect 198090 140060 198096 140072
rect 171376 140032 198096 140060
rect 171376 140020 171382 140032
rect 198090 140020 198096 140032
rect 198148 140020 198154 140072
rect 172422 139340 172428 139392
rect 172480 139380 172486 139392
rect 192570 139380 192576 139392
rect 172480 139352 192576 139380
rect 172480 139340 172486 139352
rect 192570 139340 192576 139352
rect 192628 139340 192634 139392
rect 302694 139340 302700 139392
rect 302752 139380 302758 139392
rect 359458 139380 359464 139392
rect 302752 139352 359464 139380
rect 302752 139340 302758 139352
rect 359458 139340 359464 139352
rect 359516 139340 359522 139392
rect 371418 139340 371424 139392
rect 371476 139380 371482 139392
rect 376754 139380 376760 139392
rect 371476 139352 376760 139380
rect 371476 139340 371482 139352
rect 376754 139340 376760 139352
rect 376812 139340 376818 139392
rect 548518 139340 548524 139392
rect 548576 139380 548582 139392
rect 580166 139380 580172 139392
rect 548576 139352 580172 139380
rect 548576 139340 548582 139352
rect 580166 139340 580172 139352
rect 580224 139340 580230 139392
rect 172330 139272 172336 139324
rect 172388 139312 172394 139324
rect 191098 139312 191104 139324
rect 172388 139284 191104 139312
rect 172388 139272 172394 139284
rect 191098 139272 191104 139284
rect 191156 139272 191162 139324
rect 172238 139204 172244 139256
rect 172296 139244 172302 139256
rect 177482 139244 177488 139256
rect 172296 139216 177488 139244
rect 172296 139204 172302 139216
rect 177482 139204 177488 139216
rect 177540 139204 177546 139256
rect 371970 139000 371976 139052
rect 372028 139040 372034 139052
rect 374178 139040 374184 139052
rect 372028 139012 374184 139040
rect 372028 139000 372034 139012
rect 374178 139000 374184 139012
rect 374236 139000 374242 139052
rect 371418 138660 371424 138712
rect 371476 138700 371482 138712
rect 375466 138700 375472 138712
rect 371476 138672 375472 138700
rect 371476 138660 371482 138672
rect 375466 138660 375472 138672
rect 375524 138660 375530 138712
rect 172054 137912 172060 137964
rect 172112 137952 172118 137964
rect 182818 137952 182824 137964
rect 172112 137924 182824 137952
rect 172112 137912 172118 137924
rect 182818 137912 182824 137924
rect 182876 137912 182882 137964
rect 444834 137912 444840 137964
rect 444892 137952 444898 137964
rect 448698 137952 448704 137964
rect 444892 137924 448704 137952
rect 444892 137912 444898 137924
rect 448698 137912 448704 137924
rect 448756 137912 448762 137964
rect 171686 137844 171692 137896
rect 171744 137884 171750 137896
rect 175918 137884 175924 137896
rect 171744 137856 175924 137884
rect 171744 137844 171750 137856
rect 175918 137844 175924 137856
rect 175976 137844 175982 137896
rect 176010 136620 176016 136672
rect 176068 136660 176074 136672
rect 197354 136660 197360 136672
rect 176068 136632 197360 136660
rect 176068 136620 176074 136632
rect 197354 136620 197360 136632
rect 197412 136620 197418 136672
rect 172238 136552 172244 136604
rect 172296 136592 172302 136604
rect 181530 136592 181536 136604
rect 172296 136564 181536 136592
rect 172296 136552 172302 136564
rect 181530 136552 181536 136564
rect 181588 136552 181594 136604
rect 172422 136484 172428 136536
rect 172480 136524 172486 136536
rect 174538 136524 174544 136536
rect 172480 136496 174544 136524
rect 172480 136484 172486 136496
rect 174538 136484 174544 136496
rect 174596 136484 174602 136536
rect 444374 136280 444380 136332
rect 444432 136320 444438 136332
rect 444558 136320 444564 136332
rect 444432 136292 444564 136320
rect 444432 136280 444438 136292
rect 444558 136280 444564 136292
rect 444616 136320 444622 136332
rect 447134 136320 447140 136332
rect 444616 136292 447140 136320
rect 444616 136280 444622 136292
rect 447134 136280 447140 136292
rect 447192 136280 447198 136332
rect 171870 136212 171876 136264
rect 171928 136252 171934 136264
rect 179414 136252 179420 136264
rect 171928 136224 179420 136252
rect 171928 136212 171934 136224
rect 179414 136212 179420 136224
rect 179472 136212 179478 136264
rect 172514 135872 172520 135924
rect 172572 135912 172578 135924
rect 197722 135912 197728 135924
rect 172572 135884 197728 135912
rect 172572 135872 172578 135884
rect 197722 135872 197728 135884
rect 197780 135872 197786 135924
rect 171686 135124 171692 135176
rect 171744 135164 171750 135176
rect 178034 135164 178040 135176
rect 171744 135136 178040 135164
rect 171744 135124 171750 135136
rect 178034 135124 178040 135136
rect 178092 135124 178098 135176
rect 172514 134512 172520 134564
rect 172572 134552 172578 134564
rect 197354 134552 197360 134564
rect 172572 134524 197360 134552
rect 172572 134512 172578 134524
rect 197354 134512 197360 134524
rect 197412 134512 197418 134564
rect 172054 134240 172060 134292
rect 172112 134280 172118 134292
rect 176010 134280 176016 134292
rect 172112 134252 176016 134280
rect 172112 134240 172118 134252
rect 176010 134240 176016 134252
rect 176068 134240 176074 134292
rect 444466 133152 444472 133204
rect 444524 133192 444530 133204
rect 458174 133192 458180 133204
rect 444524 133164 458180 133192
rect 444524 133152 444530 133164
rect 458174 133152 458180 133164
rect 458232 133152 458238 133204
rect 171134 132472 171140 132524
rect 171192 132512 171198 132524
rect 197354 132512 197360 132524
rect 171192 132484 197360 132512
rect 171192 132472 171198 132484
rect 197354 132472 197360 132484
rect 197412 132472 197418 132524
rect 445662 132404 445668 132456
rect 445720 132444 445726 132456
rect 454218 132444 454224 132456
rect 445720 132416 454224 132444
rect 445720 132404 445726 132416
rect 454218 132404 454224 132416
rect 454276 132404 454282 132456
rect 172422 131044 172428 131096
rect 172480 131084 172486 131096
rect 197354 131084 197360 131096
rect 172480 131056 197360 131084
rect 172480 131044 172486 131056
rect 197354 131044 197360 131056
rect 197412 131044 197418 131096
rect 444834 130432 444840 130484
rect 444892 130472 444898 130484
rect 451274 130472 451280 130484
rect 444892 130444 451280 130472
rect 444892 130432 444898 130444
rect 451274 130432 451280 130444
rect 451332 130432 451338 130484
rect 172422 130024 172428 130076
rect 172480 130064 172486 130076
rect 175274 130064 175280 130076
rect 172480 130036 175280 130064
rect 172480 130024 172486 130036
rect 175274 130024 175280 130036
rect 175332 130024 175338 130076
rect 171870 129752 171876 129804
rect 171928 129792 171934 129804
rect 176654 129792 176660 129804
rect 171928 129764 176660 129792
rect 171928 129752 171934 129764
rect 176654 129752 176660 129764
rect 176712 129752 176718 129804
rect 171502 129684 171508 129736
rect 171560 129724 171566 129736
rect 197354 129724 197360 129736
rect 171560 129696 197360 129724
rect 171560 129684 171566 129696
rect 197354 129684 197360 129696
rect 197412 129684 197418 129736
rect 444834 129684 444840 129736
rect 444892 129724 444898 129736
rect 456794 129724 456800 129736
rect 444892 129696 456800 129724
rect 444892 129684 444898 129696
rect 456794 129684 456800 129696
rect 456852 129684 456858 129736
rect 369854 129548 369860 129600
rect 369912 129588 369918 129600
rect 373994 129588 374000 129600
rect 369912 129560 374000 129588
rect 369912 129548 369918 129560
rect 373994 129548 374000 129560
rect 374052 129588 374058 129600
rect 375282 129588 375288 129600
rect 374052 129560 375288 129588
rect 374052 129548 374058 129560
rect 375282 129548 375288 129560
rect 375340 129548 375346 129600
rect 375282 129072 375288 129124
rect 375340 129112 375346 129124
rect 429194 129112 429200 129124
rect 375340 129084 429200 129112
rect 375340 129072 375346 129084
rect 429194 129072 429200 129084
rect 429252 129072 429258 129124
rect 370222 129004 370228 129056
rect 370280 129044 370286 129056
rect 371694 129044 371700 129056
rect 370280 129016 371700 129044
rect 370280 129004 370286 129016
rect 371694 129004 371700 129016
rect 371752 129044 371758 129056
rect 430574 129044 430580 129056
rect 371752 129016 430580 129044
rect 371752 129004 371758 129016
rect 430574 129004 430580 129016
rect 430632 129004 430638 129056
rect 171870 128528 171876 128580
rect 171928 128568 171934 128580
rect 174446 128568 174452 128580
rect 171928 128540 174452 128568
rect 171928 128528 171934 128540
rect 174446 128528 174452 128540
rect 174504 128528 174510 128580
rect 171502 128460 171508 128512
rect 171560 128500 171566 128512
rect 173158 128500 173164 128512
rect 171560 128472 173164 128500
rect 171560 128460 171566 128472
rect 173158 128460 173164 128472
rect 173216 128460 173222 128512
rect 174446 127576 174452 127628
rect 174504 127616 174510 127628
rect 197998 127616 198004 127628
rect 174504 127588 198004 127616
rect 174504 127576 174510 127588
rect 197998 127576 198004 127588
rect 198056 127576 198062 127628
rect 172422 127032 172428 127084
rect 172480 127072 172486 127084
rect 182818 127072 182824 127084
rect 172480 127044 182824 127072
rect 172480 127032 172486 127044
rect 182818 127032 182824 127044
rect 182876 127032 182882 127084
rect 171686 126964 171692 127016
rect 171744 127004 171750 127016
rect 191098 127004 191104 127016
rect 171744 126976 191104 127004
rect 171744 126964 171750 126976
rect 191098 126964 191104 126976
rect 191156 126964 191162 127016
rect 443638 126964 443644 127016
rect 443696 127004 443702 127016
rect 452654 127004 452660 127016
rect 443696 126976 452660 127004
rect 443696 126964 443702 126976
rect 452654 126964 452660 126976
rect 452712 126964 452718 127016
rect 176654 126896 176660 126948
rect 176712 126936 176718 126948
rect 198458 126936 198464 126948
rect 176712 126908 198464 126936
rect 176712 126896 176718 126908
rect 198458 126896 198464 126908
rect 198516 126896 198522 126948
rect 443270 126216 443276 126268
rect 443328 126256 443334 126268
rect 447226 126256 447232 126268
rect 443328 126228 447232 126256
rect 443328 126216 443334 126228
rect 447226 126216 447232 126228
rect 447284 126216 447290 126268
rect 371234 126012 371240 126064
rect 371292 126052 371298 126064
rect 441798 126052 441804 126064
rect 371292 126024 441804 126052
rect 371292 126012 371298 126024
rect 441798 126012 441804 126024
rect 441856 126012 441862 126064
rect 371786 125944 371792 125996
rect 371844 125984 371850 125996
rect 443638 125984 443644 125996
rect 371844 125956 443644 125984
rect 371844 125944 371850 125956
rect 443638 125944 443644 125956
rect 443696 125944 443702 125996
rect 371510 125876 371516 125928
rect 371568 125916 371574 125928
rect 442994 125916 443000 125928
rect 371568 125888 443000 125916
rect 371568 125876 371574 125888
rect 442994 125876 443000 125888
rect 443052 125876 443058 125928
rect 172330 125740 172336 125792
rect 172388 125780 172394 125792
rect 180058 125780 180064 125792
rect 172388 125752 180064 125780
rect 172388 125740 172394 125752
rect 180058 125740 180064 125752
rect 180116 125740 180122 125792
rect 172422 125672 172428 125724
rect 172480 125712 172486 125724
rect 178678 125712 178684 125724
rect 172480 125684 178684 125712
rect 172480 125672 172486 125684
rect 178678 125672 178684 125684
rect 178736 125672 178742 125724
rect 172054 125604 172060 125656
rect 172112 125644 172118 125656
rect 181438 125644 181444 125656
rect 172112 125616 181444 125644
rect 172112 125604 172118 125616
rect 181438 125604 181444 125616
rect 181496 125604 181502 125656
rect 175274 125536 175280 125588
rect 175332 125576 175338 125588
rect 197538 125576 197544 125588
rect 175332 125548 197544 125576
rect 175332 125536 175338 125548
rect 197538 125536 197544 125548
rect 197596 125536 197602 125588
rect 371234 125468 371240 125520
rect 371292 125508 371298 125520
rect 374086 125508 374092 125520
rect 371292 125480 374092 125508
rect 371292 125468 371298 125480
rect 374086 125468 374092 125480
rect 374144 125508 374150 125520
rect 441798 125508 441804 125520
rect 374144 125480 441804 125508
rect 374144 125468 374150 125480
rect 441798 125468 441804 125480
rect 441856 125468 441862 125520
rect 429194 125400 429200 125452
rect 429252 125440 429258 125452
rect 444558 125440 444564 125452
rect 429252 125412 444564 125440
rect 429252 125400 429258 125412
rect 444558 125400 444564 125412
rect 444616 125400 444622 125452
rect 430574 125332 430580 125384
rect 430632 125372 430638 125384
rect 444742 125372 444748 125384
rect 430632 125344 444748 125372
rect 430632 125332 430638 125344
rect 444742 125332 444748 125344
rect 444800 125332 444806 125384
rect 372522 125264 372528 125316
rect 372580 125304 372586 125316
rect 441890 125304 441896 125316
rect 372580 125276 441896 125304
rect 372580 125264 372586 125276
rect 441890 125264 441896 125276
rect 441948 125264 441954 125316
rect 302602 125196 302608 125248
rect 302660 125236 302666 125248
rect 370222 125236 370228 125248
rect 302660 125208 370228 125236
rect 302660 125196 302666 125208
rect 370222 125196 370228 125208
rect 370280 125196 370286 125248
rect 172422 125128 172428 125180
rect 172480 125168 172486 125180
rect 177298 125168 177304 125180
rect 172480 125140 177304 125168
rect 172480 125128 172486 125140
rect 177298 125128 177304 125140
rect 177356 125128 177362 125180
rect 302970 125128 302976 125180
rect 303028 125168 303034 125180
rect 369854 125168 369860 125180
rect 303028 125140 369860 125168
rect 303028 125128 303034 125140
rect 369854 125128 369860 125140
rect 369912 125128 369918 125180
rect 302786 125060 302792 125112
rect 302844 125100 302850 125112
rect 370038 125100 370044 125112
rect 302844 125072 370044 125100
rect 302844 125060 302850 125072
rect 370038 125060 370044 125072
rect 370096 125060 370102 125112
rect 302878 124992 302884 125044
rect 302936 125032 302942 125044
rect 369946 125032 369952 125044
rect 302936 125004 369952 125032
rect 302936 124992 302942 125004
rect 369946 124992 369952 125004
rect 370004 124992 370010 125044
rect 359458 124856 359464 124908
rect 359516 124896 359522 124908
rect 369302 124896 369308 124908
rect 359516 124868 369308 124896
rect 359516 124856 359522 124868
rect 369302 124856 369308 124868
rect 369360 124856 369366 124908
rect 372430 124856 372436 124908
rect 372488 124896 372494 124908
rect 441798 124896 441804 124908
rect 372488 124868 441804 124896
rect 372488 124856 372494 124868
rect 441798 124856 441804 124868
rect 441856 124896 441862 124908
rect 445846 124896 445852 124908
rect 441856 124868 445852 124896
rect 441856 124856 441862 124868
rect 445846 124856 445852 124868
rect 445904 124856 445910 124908
rect 171318 124584 171324 124636
rect 171376 124624 171382 124636
rect 175918 124624 175924 124636
rect 171376 124596 175924 124624
rect 171376 124584 171382 124596
rect 175918 124584 175924 124596
rect 175976 124584 175982 124636
rect 171962 124176 171968 124228
rect 172020 124216 172026 124228
rect 174538 124216 174544 124228
rect 172020 124188 174544 124216
rect 172020 124176 172026 124188
rect 174538 124176 174544 124188
rect 174596 124176 174602 124228
rect 302786 124108 302792 124160
rect 302844 124148 302850 124160
rect 371602 124148 371608 124160
rect 302844 124120 371608 124148
rect 302844 124108 302850 124120
rect 371602 124108 371608 124120
rect 371660 124148 371666 124160
rect 444466 124148 444472 124160
rect 371660 124120 444472 124148
rect 371660 124108 371666 124120
rect 444466 124108 444472 124120
rect 444524 124108 444530 124160
rect 367646 124040 367652 124092
rect 367704 124080 367710 124092
rect 369394 124080 369400 124092
rect 367704 124052 369400 124080
rect 367704 124040 367710 124052
rect 369394 124040 369400 124052
rect 369452 124040 369458 124092
rect 437198 124040 437204 124092
rect 437256 124080 437262 124092
rect 443178 124080 443184 124092
rect 437256 124052 443184 124080
rect 437256 124040 437262 124052
rect 443178 124040 443184 124052
rect 443236 124040 443242 124092
rect 302970 123564 302976 123616
rect 303028 123604 303034 123616
rect 370406 123604 370412 123616
rect 303028 123576 370412 123604
rect 303028 123564 303034 123576
rect 370406 123564 370412 123576
rect 370464 123564 370470 123616
rect 302878 123428 302884 123480
rect 302936 123468 302942 123480
rect 370222 123468 370228 123480
rect 302936 123440 370228 123468
rect 302936 123428 302942 123440
rect 370222 123428 370228 123440
rect 370280 123428 370286 123480
rect 162854 122884 162860 122936
rect 162912 122924 162918 122936
rect 188338 122924 188344 122936
rect 162912 122896 188344 122924
rect 162912 122884 162918 122896
rect 188338 122884 188344 122896
rect 188396 122884 188402 122936
rect 160922 122816 160928 122868
rect 160980 122856 160986 122868
rect 198826 122856 198832 122868
rect 160980 122828 198832 122856
rect 160980 122816 160986 122828
rect 198826 122816 198832 122828
rect 198884 122816 198890 122868
rect 166902 122748 166908 122800
rect 166960 122788 166966 122800
rect 170398 122788 170404 122800
rect 166960 122760 170404 122788
rect 166960 122748 166966 122760
rect 170398 122748 170404 122760
rect 170456 122748 170462 122800
rect 184198 122788 184204 122800
rect 171796 122760 184204 122788
rect 164878 122612 164884 122664
rect 164936 122652 164942 122664
rect 171796 122652 171824 122760
rect 184198 122748 184204 122760
rect 184256 122748 184262 122800
rect 322198 122748 322204 122800
rect 322256 122788 322262 122800
rect 438854 122788 438860 122800
rect 322256 122760 438860 122788
rect 322256 122748 322262 122760
rect 438854 122748 438860 122760
rect 438912 122748 438918 122800
rect 186958 122720 186964 122732
rect 164936 122624 171824 122652
rect 176626 122692 186964 122720
rect 164936 122612 164942 122624
rect 168926 122544 168932 122596
rect 168984 122584 168990 122596
rect 176626 122584 176654 122692
rect 186958 122680 186964 122692
rect 187016 122680 187022 122732
rect 320818 122680 320824 122732
rect 320876 122720 320882 122732
rect 366910 122720 366916 122732
rect 320876 122692 366916 122720
rect 320876 122680 320882 122692
rect 366910 122680 366916 122692
rect 366968 122680 366974 122732
rect 435174 122680 435180 122732
rect 435232 122720 435238 122732
rect 441706 122720 441712 122732
rect 435232 122692 441712 122720
rect 435232 122680 435238 122692
rect 441706 122680 441712 122692
rect 441764 122680 441770 122732
rect 168984 122556 176654 122584
rect 168984 122544 168990 122556
rect 173158 121388 173164 121440
rect 173216 121428 173222 121440
rect 197538 121428 197544 121440
rect 173216 121400 197544 121428
rect 173216 121388 173222 121400
rect 197538 121388 197544 121400
rect 197596 121388 197602 121440
rect 302510 121388 302516 121440
rect 302568 121428 302574 121440
rect 370314 121428 370320 121440
rect 302568 121400 370320 121428
rect 302568 121388 302574 121400
rect 370314 121388 370320 121400
rect 370372 121388 370378 121440
rect 171778 118600 171784 118652
rect 171836 118640 171842 118652
rect 197906 118640 197912 118652
rect 171836 118612 197912 118640
rect 171836 118600 171842 118612
rect 197906 118600 197912 118612
rect 197964 118600 197970 118652
rect 302786 117240 302792 117292
rect 302844 117280 302850 117292
rect 367646 117280 367652 117292
rect 302844 117252 367652 117280
rect 302844 117240 302850 117252
rect 367646 117240 367652 117252
rect 367704 117240 367710 117292
rect 191098 116628 191104 116680
rect 191156 116668 191162 116680
rect 198366 116668 198372 116680
rect 191156 116640 198372 116668
rect 191156 116628 191162 116640
rect 198366 116628 198372 116640
rect 198424 116628 198430 116680
rect 182818 114452 182824 114504
rect 182876 114492 182882 114504
rect 197354 114492 197360 114504
rect 182876 114464 197360 114492
rect 182876 114452 182882 114464
rect 197354 114452 197360 114464
rect 197412 114452 197418 114504
rect 307018 113092 307024 113144
rect 307076 113132 307082 113144
rect 579798 113132 579804 113144
rect 307076 113104 579804 113132
rect 307076 113092 307082 113104
rect 579798 113092 579804 113104
rect 579856 113092 579862 113144
rect 3418 111732 3424 111784
rect 3476 111772 3482 111784
rect 159358 111772 159364 111784
rect 3476 111744 159364 111772
rect 3476 111732 3482 111744
rect 159358 111732 159364 111744
rect 159416 111732 159422 111784
rect 181438 111732 181444 111784
rect 181496 111772 181502 111784
rect 197354 111772 197360 111784
rect 181496 111744 197360 111772
rect 181496 111732 181502 111744
rect 197354 111732 197360 111744
rect 197412 111732 197418 111784
rect 302786 111732 302792 111784
rect 302844 111772 302850 111784
rect 369946 111772 369952 111784
rect 302844 111744 369952 111772
rect 302844 111732 302850 111744
rect 369946 111732 369952 111744
rect 370004 111732 370010 111784
rect 180058 110372 180064 110424
rect 180116 110412 180122 110424
rect 197354 110412 197360 110424
rect 180116 110384 197360 110412
rect 180116 110372 180122 110384
rect 197354 110372 197360 110384
rect 197412 110372 197418 110424
rect 302786 108944 302792 108996
rect 302844 108984 302850 108996
rect 359458 108984 359464 108996
rect 302844 108956 359464 108984
rect 302844 108944 302850 108956
rect 359458 108944 359464 108956
rect 359516 108944 359522 108996
rect 178678 107584 178684 107636
rect 178736 107624 178742 107636
rect 198550 107624 198556 107636
rect 178736 107596 198556 107624
rect 178736 107584 178742 107596
rect 198550 107584 198556 107596
rect 198608 107584 198614 107636
rect 177298 106224 177304 106276
rect 177356 106264 177362 106276
rect 197538 106264 197544 106276
rect 177356 106236 197544 106264
rect 177356 106224 177362 106236
rect 197538 106224 197544 106236
rect 197596 106224 197602 106276
rect 175918 103436 175924 103488
rect 175976 103476 175982 103488
rect 197906 103476 197912 103488
rect 175976 103448 197912 103476
rect 175976 103436 175982 103448
rect 197906 103436 197912 103448
rect 197964 103436 197970 103488
rect 302786 102756 302792 102808
rect 302844 102796 302850 102808
rect 369854 102796 369860 102808
rect 302844 102768 369860 102796
rect 302844 102756 302850 102768
rect 369854 102756 369860 102768
rect 369912 102756 369918 102808
rect 174538 102076 174544 102128
rect 174596 102116 174602 102128
rect 197538 102116 197544 102128
rect 174596 102088 197544 102116
rect 174596 102076 174602 102088
rect 197538 102076 197544 102088
rect 197596 102076 197602 102128
rect 300210 101328 300216 101380
rect 300268 101368 300274 101380
rect 301498 101368 301504 101380
rect 300268 101340 301504 101368
rect 300268 101328 300274 101340
rect 301498 101328 301504 101340
rect 301556 101328 301562 101380
rect 316678 100648 316684 100700
rect 316736 100688 316742 100700
rect 580166 100688 580172 100700
rect 316736 100660 580172 100688
rect 316736 100648 316742 100660
rect 580166 100648 580172 100660
rect 580224 100648 580230 100700
rect 258166 100240 258172 100292
rect 258224 100280 258230 100292
rect 339494 100280 339500 100292
rect 258224 100252 339500 100280
rect 258224 100240 258230 100252
rect 339494 100240 339500 100252
rect 339552 100240 339558 100292
rect 255774 100172 255780 100224
rect 255832 100212 255838 100224
rect 323578 100212 323584 100224
rect 255832 100184 323584 100212
rect 255832 100172 255838 100184
rect 323578 100172 323584 100184
rect 323636 100172 323642 100224
rect 260742 100104 260748 100156
rect 260800 100144 260806 100156
rect 353938 100144 353944 100156
rect 260800 100116 353944 100144
rect 260800 100104 260806 100116
rect 353938 100104 353944 100116
rect 353996 100104 354002 100156
rect 195238 100036 195244 100088
rect 195296 100076 195302 100088
rect 299566 100076 299572 100088
rect 195296 100048 299572 100076
rect 195296 100036 195302 100048
rect 299566 100036 299572 100048
rect 299624 100036 299630 100088
rect 106182 99968 106188 100020
rect 106240 100008 106246 100020
rect 217962 100008 217968 100020
rect 106240 99980 217968 100008
rect 106240 99968 106246 99980
rect 217962 99968 217968 99980
rect 218020 99968 218026 100020
rect 264974 99968 264980 100020
rect 265032 100008 265038 100020
rect 376018 100008 376024 100020
rect 265032 99980 376024 100008
rect 265032 99968 265038 99980
rect 376018 99968 376024 99980
rect 376076 99968 376082 100020
rect 124858 99900 124864 99952
rect 124916 99940 124922 99952
rect 212810 99940 212816 99952
rect 124916 99912 212816 99940
rect 124916 99900 124922 99912
rect 212810 99900 212816 99912
rect 212868 99900 212874 99952
rect 270586 99900 270592 99952
rect 270644 99940 270650 99952
rect 412634 99940 412640 99952
rect 270644 99912 412640 99940
rect 270644 99900 270650 99912
rect 412634 99900 412640 99912
rect 412692 99900 412698 99952
rect 108298 99832 108304 99884
rect 108356 99872 108362 99884
rect 215202 99872 215208 99884
rect 108356 99844 215208 99872
rect 108356 99832 108362 99844
rect 215202 99832 215208 99844
rect 215260 99832 215266 99884
rect 271138 99832 271144 99884
rect 271196 99872 271202 99884
rect 414658 99872 414664 99884
rect 271196 99844 414664 99872
rect 271196 99832 271202 99844
rect 414658 99832 414664 99844
rect 414716 99832 414722 99884
rect 111058 99764 111064 99816
rect 111116 99804 111122 99816
rect 218422 99804 218428 99816
rect 111116 99776 218428 99804
rect 111116 99764 111122 99776
rect 218422 99764 218428 99776
rect 218480 99764 218486 99816
rect 272426 99764 272432 99816
rect 272484 99804 272490 99816
rect 423674 99804 423680 99816
rect 272484 99776 423680 99804
rect 272484 99764 272490 99776
rect 423674 99764 423680 99776
rect 423732 99764 423738 99816
rect 93118 99696 93124 99748
rect 93176 99736 93182 99748
rect 213362 99736 213368 99748
rect 93176 99708 213368 99736
rect 93176 99696 93182 99708
rect 213362 99696 213368 99708
rect 213420 99696 213426 99748
rect 273622 99696 273628 99748
rect 273680 99736 273686 99748
rect 430574 99736 430580 99748
rect 273680 99708 430580 99736
rect 273680 99696 273686 99708
rect 430574 99696 430580 99708
rect 430632 99696 430638 99748
rect 87598 99628 87604 99680
rect 87656 99668 87662 99680
rect 210786 99668 210792 99680
rect 87656 99640 210792 99668
rect 87656 99628 87662 99640
rect 210786 99628 210792 99640
rect 210844 99628 210850 99680
rect 274818 99628 274824 99680
rect 274876 99668 274882 99680
rect 435358 99668 435364 99680
rect 274876 99640 435364 99668
rect 274876 99628 274882 99640
rect 435358 99628 435364 99640
rect 435416 99628 435422 99680
rect 91002 99560 91008 99612
rect 91060 99600 91066 99612
rect 215386 99600 215392 99612
rect 91060 99572 215392 99600
rect 91060 99560 91066 99572
rect 215386 99560 215392 99572
rect 215444 99560 215450 99612
rect 275462 99560 275468 99612
rect 275520 99600 275526 99612
rect 440234 99600 440240 99612
rect 275520 99572 440240 99600
rect 275520 99560 275526 99572
rect 440234 99560 440240 99572
rect 440292 99560 440298 99612
rect 72418 99492 72424 99544
rect 72476 99532 72482 99544
rect 211154 99532 211160 99544
rect 72476 99504 211160 99532
rect 72476 99492 72482 99504
rect 211154 99492 211160 99504
rect 211212 99492 211218 99544
rect 276014 99492 276020 99544
rect 276072 99532 276078 99544
rect 442258 99532 442264 99544
rect 276072 99504 442264 99532
rect 276072 99492 276078 99504
rect 442258 99492 442264 99504
rect 442316 99492 442322 99544
rect 53098 99424 53104 99476
rect 53156 99464 53162 99476
rect 208394 99464 208400 99476
rect 53156 99436 208400 99464
rect 53156 99424 53162 99436
rect 208394 99424 208400 99436
rect 208452 99424 208458 99476
rect 278498 99424 278504 99476
rect 278556 99464 278562 99476
rect 457438 99464 457444 99476
rect 278556 99436 457444 99464
rect 278556 99424 278562 99436
rect 457438 99424 457444 99436
rect 457496 99424 457502 99476
rect 39298 99356 39304 99408
rect 39356 99396 39362 99408
rect 203702 99396 203708 99408
rect 39356 99368 203708 99396
rect 39356 99356 39362 99368
rect 203702 99356 203708 99368
rect 203760 99356 203766 99408
rect 279694 99356 279700 99408
rect 279752 99396 279758 99408
rect 464338 99396 464344 99408
rect 279752 99368 464344 99396
rect 279752 99356 279758 99368
rect 464338 99356 464344 99368
rect 464396 99356 464402 99408
rect 180702 99288 180708 99340
rect 180760 99328 180766 99340
rect 230750 99328 230756 99340
rect 180760 99300 230756 99328
rect 180760 99288 180766 99300
rect 230750 99288 230756 99300
rect 230808 99288 230814 99340
rect 282914 99288 282920 99340
rect 282972 99328 282978 99340
rect 316678 99328 316684 99340
rect 282972 99300 316684 99328
rect 282972 99288 282978 99300
rect 316678 99288 316684 99300
rect 316736 99288 316742 99340
rect 174538 99220 174544 99272
rect 174596 99260 174602 99272
rect 229554 99260 229560 99272
rect 174596 99232 229560 99260
rect 174596 99220 174602 99232
rect 229554 99220 229560 99232
rect 229612 99220 229618 99272
rect 265526 99220 265532 99272
rect 265584 99260 265590 99272
rect 311158 99260 311164 99272
rect 265584 99232 311164 99260
rect 265584 99220 265590 99232
rect 311158 99220 311164 99232
rect 311216 99220 311222 99272
rect 152550 99152 152556 99204
rect 152608 99192 152614 99204
rect 225322 99192 225328 99204
rect 152608 99164 225328 99192
rect 152608 99152 152614 99164
rect 225322 99152 225328 99164
rect 225380 99152 225386 99204
rect 253014 99152 253020 99204
rect 253072 99192 253078 99204
rect 309134 99192 309140 99204
rect 253072 99164 309140 99192
rect 253072 99152 253078 99164
rect 309134 99152 309140 99164
rect 309192 99152 309198 99204
rect 134518 99084 134524 99136
rect 134576 99124 134582 99136
rect 222286 99124 222292 99136
rect 134576 99096 222292 99124
rect 134576 99084 134582 99096
rect 222286 99084 222292 99096
rect 222344 99084 222350 99136
rect 253566 99084 253572 99136
rect 253624 99124 253630 99136
rect 312538 99124 312544 99136
rect 253624 99096 312544 99124
rect 253624 99084 253630 99096
rect 312538 99084 312544 99096
rect 312596 99084 312602 99136
rect 148318 99016 148324 99068
rect 148376 99056 148382 99068
rect 224494 99056 224500 99068
rect 148376 99028 224500 99056
rect 148376 99016 148382 99028
rect 224494 99016 224500 99028
rect 224552 99016 224558 99068
rect 255866 99016 255872 99068
rect 255924 99056 255930 99068
rect 324958 99056 324964 99068
rect 255924 99028 324964 99056
rect 255924 99016 255930 99028
rect 324958 99016 324964 99028
rect 325016 99016 325022 99068
rect 133782 98948 133788 99000
rect 133840 98988 133846 99000
rect 222654 98988 222660 99000
rect 133840 98960 222660 98988
rect 133840 98948 133846 98960
rect 222654 98948 222660 98960
rect 222712 98948 222718 99000
rect 263134 98948 263140 99000
rect 263192 98988 263198 99000
rect 360838 98988 360844 99000
rect 263192 98960 360844 98988
rect 263192 98948 263198 98960
rect 360838 98948 360844 98960
rect 360896 98948 360902 99000
rect 130378 98880 130384 98932
rect 130436 98920 130442 98932
rect 222102 98920 222108 98932
rect 130436 98892 222108 98920
rect 130436 98880 130442 98892
rect 222102 98880 222108 98892
rect 222160 98880 222166 98932
rect 279050 98880 279056 98932
rect 279108 98920 279114 98932
rect 460198 98920 460204 98932
rect 279108 98892 460204 98920
rect 279108 98880 279114 98892
rect 460198 98880 460204 98892
rect 460256 98880 460262 98932
rect 84102 98812 84108 98864
rect 84160 98852 84166 98864
rect 214190 98852 214196 98864
rect 84160 98824 214196 98852
rect 84160 98812 84166 98824
rect 214190 98812 214196 98824
rect 214248 98812 214254 98864
rect 292390 98812 292396 98864
rect 292448 98852 292454 98864
rect 485038 98852 485044 98864
rect 292448 98824 485044 98852
rect 292448 98812 292454 98824
rect 485038 98812 485044 98824
rect 485096 98812 485102 98864
rect 54478 98744 54484 98796
rect 54536 98784 54542 98796
rect 208762 98784 208768 98796
rect 54536 98756 208768 98784
rect 54536 98744 54542 98756
rect 208762 98744 208768 98756
rect 208820 98744 208826 98796
rect 286962 98744 286968 98796
rect 287020 98784 287026 98796
rect 507854 98784 507860 98796
rect 287020 98756 507860 98784
rect 287020 98744 287026 98756
rect 507854 98744 507860 98756
rect 507912 98744 507918 98796
rect 43438 98676 43444 98728
rect 43496 98716 43502 98728
rect 202506 98716 202512 98728
rect 43496 98688 202512 98716
rect 43496 98676 43502 98688
rect 202506 98676 202512 98688
rect 202564 98676 202570 98728
rect 287514 98676 287520 98728
rect 287572 98716 287578 98728
rect 511994 98716 512000 98728
rect 287572 98688 512000 98716
rect 287572 98676 287578 98688
rect 511994 98676 512000 98688
rect 512052 98676 512058 98728
rect 21358 98608 21364 98660
rect 21416 98648 21422 98660
rect 202874 98648 202880 98660
rect 21416 98620 202880 98648
rect 21416 98608 21422 98620
rect 202874 98608 202880 98620
rect 202932 98608 202938 98660
rect 290550 98608 290556 98660
rect 290608 98648 290614 98660
rect 529934 98648 529940 98660
rect 290608 98620 529940 98648
rect 290608 98608 290614 98620
rect 529934 98608 529940 98620
rect 529992 98608 529998 98660
rect 195882 98540 195888 98592
rect 195940 98580 195946 98592
rect 233418 98580 233424 98592
rect 195940 98552 233424 98580
rect 195940 98540 195946 98552
rect 233418 98540 233424 98552
rect 233476 98540 233482 98592
rect 198642 98472 198648 98524
rect 198700 98512 198706 98524
rect 234798 98512 234804 98524
rect 198700 98484 234804 98512
rect 198700 98472 198706 98484
rect 234798 98472 234804 98484
rect 234856 98472 234862 98524
rect 254946 98336 254952 98388
rect 255004 98376 255010 98388
rect 255004 98348 258074 98376
rect 255004 98336 255010 98348
rect 258046 98172 258074 98348
rect 320174 98172 320180 98184
rect 258046 98144 320180 98172
rect 320174 98132 320180 98144
rect 320232 98132 320238 98184
rect 333974 98104 333980 98116
rect 258046 98076 333980 98104
rect 188982 97996 188988 98048
rect 189040 98036 189046 98048
rect 212534 98036 212540 98048
rect 189040 98008 212540 98036
rect 189040 97996 189046 98008
rect 212534 97996 212540 98008
rect 212592 97996 212598 98048
rect 3418 97928 3424 97980
rect 3476 97968 3482 97980
rect 14458 97968 14464 97980
rect 3476 97940 14464 97968
rect 3476 97928 3482 97940
rect 14458 97928 14464 97940
rect 14516 97928 14522 97980
rect 191098 97928 191104 97980
rect 191156 97968 191162 97980
rect 214006 97968 214012 97980
rect 191156 97940 214012 97968
rect 191156 97928 191162 97940
rect 214006 97928 214012 97940
rect 214064 97928 214070 97980
rect 257246 97928 257252 97980
rect 257304 97968 257310 97980
rect 258046 97968 258074 98076
rect 333974 98064 333980 98076
rect 334032 98064 334038 98116
rect 358814 98036 358820 98048
rect 263520 98008 358820 98036
rect 257304 97940 258074 97968
rect 257304 97928 257310 97940
rect 261478 97928 261484 97980
rect 261536 97968 261542 97980
rect 263520 97968 263548 98008
rect 358814 97996 358820 98008
rect 358872 97996 358878 98048
rect 261536 97940 263548 97968
rect 261536 97928 261542 97940
rect 277578 97928 277584 97980
rect 277636 97968 277642 97980
rect 322198 97968 322204 97980
rect 277636 97940 322204 97968
rect 277636 97928 277642 97940
rect 322198 97928 322204 97940
rect 322256 97928 322262 97980
rect 184198 97860 184204 97912
rect 184256 97900 184262 97912
rect 217686 97900 217692 97912
rect 184256 97872 217692 97900
rect 184256 97860 184262 97872
rect 217686 97860 217692 97872
rect 217744 97860 217750 97912
rect 274634 97860 274640 97912
rect 274692 97900 274698 97912
rect 274692 97872 277394 97900
rect 274692 97860 274698 97872
rect 182818 97792 182824 97844
rect 182876 97832 182882 97844
rect 220078 97832 220084 97844
rect 182876 97804 220084 97832
rect 182876 97792 182882 97804
rect 220078 97792 220084 97804
rect 220136 97792 220142 97844
rect 268562 97792 268568 97844
rect 268620 97832 268626 97844
rect 277366 97832 277394 97872
rect 280706 97860 280712 97912
rect 280764 97900 280770 97912
rect 329098 97900 329104 97912
rect 280764 97872 329104 97900
rect 280764 97860 280770 97872
rect 329098 97860 329104 97872
rect 329156 97860 329162 97912
rect 335998 97832 336004 97844
rect 268620 97804 276888 97832
rect 277366 97804 336004 97832
rect 268620 97792 268626 97804
rect 173802 97724 173808 97776
rect 173860 97764 173866 97776
rect 206094 97764 206100 97776
rect 173860 97736 206100 97764
rect 173860 97724 173866 97736
rect 206094 97724 206100 97736
rect 206152 97724 206158 97776
rect 207750 97724 207756 97776
rect 207808 97764 207814 97776
rect 218882 97764 218888 97776
rect 207808 97736 218888 97764
rect 207808 97724 207814 97736
rect 218882 97724 218888 97736
rect 218940 97724 218946 97776
rect 238018 97724 238024 97776
rect 238076 97764 238082 97776
rect 239490 97764 239496 97776
rect 238076 97736 239496 97764
rect 238076 97724 238082 97736
rect 239490 97724 239496 97736
rect 239548 97724 239554 97776
rect 264330 97724 264336 97776
rect 264388 97764 264394 97776
rect 268378 97764 268384 97776
rect 264388 97736 268384 97764
rect 264388 97724 264394 97736
rect 268378 97724 268384 97736
rect 268436 97724 268442 97776
rect 269758 97724 269764 97776
rect 269816 97764 269822 97776
rect 269816 97736 274588 97764
rect 269816 97724 269822 97736
rect 121362 97656 121368 97708
rect 121420 97696 121426 97708
rect 220630 97696 220636 97708
rect 121420 97668 207888 97696
rect 121420 97656 121426 97668
rect 112438 97588 112444 97640
rect 112496 97628 112502 97640
rect 207750 97628 207756 97640
rect 112496 97600 207756 97628
rect 112496 97588 112502 97600
rect 207750 97588 207756 97600
rect 207808 97588 207814 97640
rect 207860 97628 207888 97668
rect 215266 97668 220636 97696
rect 215266 97628 215294 97668
rect 220630 97656 220636 97668
rect 220688 97656 220694 97708
rect 245562 97656 245568 97708
rect 245620 97696 245626 97708
rect 253290 97696 253296 97708
rect 245620 97668 253296 97696
rect 245620 97656 245626 97668
rect 253290 97656 253296 97668
rect 253348 97656 253354 97708
rect 262490 97656 262496 97708
rect 262548 97696 262554 97708
rect 271230 97696 271236 97708
rect 262548 97668 271236 97696
rect 262548 97656 262554 97668
rect 271230 97656 271236 97668
rect 271288 97656 271294 97708
rect 274560 97696 274588 97736
rect 276860 97696 276888 97804
rect 335998 97792 336004 97804
rect 336056 97792 336062 97844
rect 280798 97724 280804 97776
rect 280856 97764 280862 97776
rect 342898 97764 342904 97776
rect 280856 97736 342904 97764
rect 280856 97724 280862 97736
rect 342898 97724 342904 97736
rect 342956 97724 342962 97776
rect 393958 97696 393964 97708
rect 274560 97668 276704 97696
rect 276860 97668 393964 97696
rect 207860 97600 215294 97628
rect 218054 97588 218060 97640
rect 218112 97628 218118 97640
rect 228174 97628 228180 97640
rect 218112 97600 228180 97628
rect 218112 97588 218118 97600
rect 228174 97588 228180 97600
rect 228232 97588 228238 97640
rect 252370 97588 252376 97640
rect 252428 97628 252434 97640
rect 263778 97628 263784 97640
rect 252428 97600 263784 97628
rect 252428 97588 252434 97600
rect 263778 97588 263784 97600
rect 263836 97588 263842 97640
rect 270402 97588 270408 97640
rect 270460 97628 270466 97640
rect 276566 97628 276572 97640
rect 270460 97600 276572 97628
rect 270460 97588 270466 97600
rect 276566 97588 276572 97600
rect 276624 97588 276630 97640
rect 276676 97628 276704 97668
rect 393958 97656 393964 97668
rect 394016 97656 394022 97708
rect 400858 97628 400864 97640
rect 276676 97600 400864 97628
rect 400858 97588 400864 97600
rect 400916 97588 400922 97640
rect 97258 97520 97264 97572
rect 97316 97560 97322 97572
rect 216398 97560 216404 97572
rect 97316 97532 216404 97560
rect 97316 97520 97322 97532
rect 216398 97520 216404 97532
rect 216456 97520 216462 97572
rect 216766 97520 216772 97572
rect 216824 97560 216830 97572
rect 230014 97560 230020 97572
rect 216824 97532 230020 97560
rect 216824 97520 216830 97532
rect 230014 97520 230020 97532
rect 230072 97520 230078 97572
rect 247310 97520 247316 97572
rect 247368 97560 247374 97572
rect 255958 97560 255964 97572
rect 247368 97532 255964 97560
rect 247368 97520 247374 97532
rect 255958 97520 255964 97532
rect 256016 97520 256022 97572
rect 260834 97520 260840 97572
rect 260892 97560 260898 97572
rect 271506 97560 271512 97572
rect 260892 97532 271512 97560
rect 260892 97520 260898 97532
rect 271506 97520 271512 97532
rect 271564 97520 271570 97572
rect 275830 97520 275836 97572
rect 275888 97560 275894 97572
rect 436738 97560 436744 97572
rect 275888 97532 436744 97560
rect 275888 97520 275894 97532
rect 436738 97520 436744 97532
rect 436796 97520 436802 97572
rect 58618 97452 58624 97504
rect 58676 97492 58682 97504
rect 206738 97492 206744 97504
rect 58676 97464 206744 97492
rect 58676 97452 58682 97464
rect 206738 97452 206744 97464
rect 206796 97452 206802 97504
rect 218146 97452 218152 97504
rect 218204 97492 218210 97504
rect 230566 97492 230572 97504
rect 218204 97464 230572 97492
rect 218204 97452 218210 97464
rect 230566 97452 230572 97464
rect 230624 97452 230630 97504
rect 235810 97452 235816 97504
rect 235868 97492 235874 97504
rect 238846 97492 238852 97504
rect 235868 97464 238852 97492
rect 235868 97452 235874 97464
rect 238846 97452 238852 97464
rect 238904 97452 238910 97504
rect 266722 97452 266728 97504
rect 266780 97492 266786 97504
rect 271138 97492 271144 97504
rect 266780 97464 271144 97492
rect 266780 97452 266786 97464
rect 271138 97452 271144 97464
rect 271196 97452 271202 97504
rect 271598 97452 271604 97504
rect 271656 97492 271662 97504
rect 276106 97492 276112 97504
rect 271656 97464 276112 97492
rect 271656 97452 271662 97464
rect 276106 97452 276112 97464
rect 276164 97452 276170 97504
rect 277026 97452 277032 97504
rect 277084 97492 277090 97504
rect 443638 97492 443644 97504
rect 277084 97464 443644 97492
rect 277084 97452 277090 97464
rect 443638 97452 443644 97464
rect 443696 97452 443702 97504
rect 56502 97384 56508 97436
rect 56560 97424 56566 97436
rect 209590 97424 209596 97436
rect 56560 97396 209596 97424
rect 56560 97384 56566 97396
rect 209590 97384 209596 97396
rect 209648 97384 209654 97436
rect 210418 97384 210424 97436
rect 210476 97424 210482 97436
rect 221274 97424 221280 97436
rect 210476 97396 221280 97424
rect 210476 97384 210482 97396
rect 221274 97384 221280 97396
rect 221332 97384 221338 97436
rect 224862 97384 224868 97436
rect 224920 97424 224926 97436
rect 238294 97424 238300 97436
rect 224920 97396 238300 97424
rect 224920 97384 224926 97396
rect 238294 97384 238300 97396
rect 238352 97384 238358 97436
rect 249794 97384 249800 97436
rect 249852 97424 249858 97436
rect 266998 97424 267004 97436
rect 249852 97396 267004 97424
rect 249852 97384 249858 97396
rect 266998 97384 267004 97396
rect 267056 97384 267062 97436
rect 272150 97384 272156 97436
rect 272208 97424 272214 97436
rect 275370 97424 275376 97436
rect 272208 97396 275376 97424
rect 272208 97384 272214 97396
rect 275370 97384 275376 97396
rect 275428 97384 275434 97436
rect 278222 97384 278228 97436
rect 278280 97424 278286 97436
rect 447778 97424 447784 97436
rect 278280 97396 447784 97424
rect 278280 97384 278286 97396
rect 447778 97384 447784 97396
rect 447836 97384 447842 97436
rect 40678 97316 40684 97368
rect 40736 97356 40742 97368
rect 204070 97356 204076 97368
rect 40736 97328 204076 97356
rect 40736 97316 40742 97328
rect 204070 97316 204076 97328
rect 204128 97316 204134 97368
rect 209406 97316 209412 97368
rect 209464 97356 209470 97368
rect 227346 97356 227352 97368
rect 209464 97328 227352 97356
rect 209464 97316 209470 97328
rect 227346 97316 227352 97328
rect 227404 97316 227410 97368
rect 228542 97316 228548 97368
rect 228600 97356 228606 97368
rect 237006 97356 237012 97368
rect 228600 97328 237012 97356
rect 228600 97316 228606 97328
rect 237006 97316 237012 97328
rect 237064 97316 237070 97368
rect 242710 97316 242716 97368
rect 242768 97356 242774 97368
rect 263594 97356 263600 97368
rect 242768 97328 263600 97356
rect 242768 97316 242774 97328
rect 263594 97316 263600 97328
rect 263652 97316 263658 97368
rect 263686 97316 263692 97368
rect 263744 97356 263750 97368
rect 278038 97356 278044 97368
rect 263744 97328 278044 97356
rect 263744 97316 263750 97328
rect 278038 97316 278044 97328
rect 278096 97316 278102 97368
rect 279510 97316 279516 97368
rect 279568 97356 279574 97368
rect 450538 97356 450544 97368
rect 279568 97328 450544 97356
rect 279568 97316 279574 97328
rect 450538 97316 450544 97328
rect 450596 97316 450602 97368
rect 14550 97248 14556 97300
rect 14608 97288 14614 97300
rect 201034 97288 201040 97300
rect 14608 97260 201040 97288
rect 14608 97248 14614 97260
rect 201034 97248 201040 97260
rect 201092 97248 201098 97300
rect 205542 97288 205548 97300
rect 202800 97260 205548 97288
rect 192570 97180 192576 97232
rect 192628 97220 192634 97232
rect 202800 97220 202828 97260
rect 205542 97248 205548 97260
rect 205600 97248 205606 97300
rect 211154 97248 211160 97300
rect 211212 97288 211218 97300
rect 233602 97288 233608 97300
rect 211212 97260 233608 97288
rect 211212 97248 211218 97260
rect 233602 97248 233608 97260
rect 233660 97248 233666 97300
rect 247586 97248 247592 97300
rect 247644 97288 247650 97300
rect 269758 97288 269764 97300
rect 247644 97260 269764 97288
rect 247644 97248 247650 97260
rect 269758 97248 269764 97260
rect 269816 97248 269822 97300
rect 272794 97248 272800 97300
rect 272852 97288 272858 97300
rect 280798 97288 280804 97300
rect 272852 97260 280804 97288
rect 272852 97248 272858 97260
rect 280798 97248 280804 97260
rect 280856 97248 280862 97300
rect 280890 97248 280896 97300
rect 280948 97288 280954 97300
rect 281258 97288 281264 97300
rect 280948 97260 281264 97288
rect 280948 97248 280954 97260
rect 281258 97248 281264 97260
rect 281316 97248 281322 97300
rect 289354 97248 289360 97300
rect 289412 97288 289418 97300
rect 289722 97288 289728 97300
rect 289412 97260 289728 97288
rect 289412 97248 289418 97260
rect 289722 97248 289728 97260
rect 289780 97248 289786 97300
rect 291838 97248 291844 97300
rect 291896 97288 291902 97300
rect 454678 97288 454684 97300
rect 291896 97260 454684 97288
rect 291896 97248 291902 97260
rect 454678 97248 454684 97260
rect 454736 97248 454742 97300
rect 192628 97192 202828 97220
rect 192628 97180 192634 97192
rect 204898 97180 204904 97232
rect 204956 97220 204962 97232
rect 221458 97220 221464 97232
rect 204956 97192 221464 97220
rect 204956 97180 204962 97192
rect 221458 97180 221464 97192
rect 221516 97180 221522 97232
rect 235626 97180 235632 97232
rect 235684 97220 235690 97232
rect 239306 97220 239312 97232
rect 235684 97192 239312 97220
rect 235684 97180 235690 97192
rect 239306 97180 239312 97192
rect 239364 97180 239370 97232
rect 267366 97180 267372 97232
rect 267424 97220 267430 97232
rect 312630 97220 312636 97232
rect 267424 97192 312636 97220
rect 267424 97180 267430 97192
rect 312630 97180 312636 97192
rect 312688 97180 312694 97232
rect 199378 97112 199384 97164
rect 199436 97152 199442 97164
rect 212166 97152 212172 97164
rect 199436 97124 212172 97152
rect 199436 97112 199442 97124
rect 212166 97112 212172 97124
rect 212224 97112 212230 97164
rect 212534 97112 212540 97164
rect 212592 97152 212598 97164
rect 232222 97152 232228 97164
rect 212592 97124 232228 97152
rect 212592 97112 212598 97124
rect 232222 97112 232228 97124
rect 232280 97112 232286 97164
rect 243538 97112 243544 97164
rect 243596 97152 243602 97164
rect 249058 97152 249064 97164
rect 243596 97124 249064 97152
rect 243596 97112 243602 97124
rect 249058 97112 249064 97124
rect 249116 97112 249122 97164
rect 250346 97112 250352 97164
rect 250404 97152 250410 97164
rect 291746 97152 291752 97164
rect 250404 97124 291752 97152
rect 250404 97112 250410 97124
rect 291746 97112 291752 97124
rect 291804 97112 291810 97164
rect 293586 97112 293592 97164
rect 293644 97152 293650 97164
rect 293862 97152 293868 97164
rect 293644 97124 293868 97152
rect 293644 97112 293650 97124
rect 293862 97112 293868 97124
rect 293920 97112 293926 97164
rect 296254 97112 296260 97164
rect 296312 97152 296318 97164
rect 296438 97152 296444 97164
rect 296312 97124 296444 97152
rect 296312 97112 296318 97124
rect 296438 97112 296444 97124
rect 296496 97112 296502 97164
rect 197998 97044 198004 97096
rect 198056 97084 198062 97096
rect 210970 97084 210976 97096
rect 198056 97056 210976 97084
rect 198056 97044 198062 97056
rect 210970 97044 210976 97056
rect 211028 97044 211034 97096
rect 220630 97044 220636 97096
rect 220688 97084 220694 97096
rect 228726 97084 228732 97096
rect 220688 97056 228732 97084
rect 220688 97044 220694 97056
rect 228726 97044 228732 97056
rect 228784 97044 228790 97096
rect 232774 97044 232780 97096
rect 232832 97084 232838 97096
rect 238662 97084 238668 97096
rect 232832 97056 238668 97084
rect 232832 97044 232838 97056
rect 238662 97044 238668 97056
rect 238720 97044 238726 97096
rect 242894 97044 242900 97096
rect 242952 97084 242958 97096
rect 250438 97084 250444 97096
rect 242952 97056 250444 97084
rect 242952 97044 242958 97056
rect 250438 97044 250444 97056
rect 250496 97044 250502 97096
rect 259454 97044 259460 97096
rect 259512 97084 259518 97096
rect 260558 97084 260564 97096
rect 259512 97056 260564 97084
rect 259512 97044 259518 97056
rect 260558 97044 260564 97056
rect 260616 97044 260622 97096
rect 261846 97044 261852 97096
rect 261904 97084 261910 97096
rect 262122 97084 262128 97096
rect 261904 97056 262128 97084
rect 261904 97044 261910 97056
rect 262122 97044 262128 97056
rect 262180 97044 262186 97096
rect 273438 97044 273444 97096
rect 273496 97084 273502 97096
rect 275278 97084 275284 97096
rect 273496 97056 275284 97084
rect 273496 97044 273502 97056
rect 275278 97044 275284 97056
rect 275336 97044 275342 97096
rect 275370 97044 275376 97096
rect 275428 97084 275434 97096
rect 280706 97084 280712 97096
rect 275428 97056 280712 97084
rect 275428 97044 275434 97056
rect 280706 97044 280712 97056
rect 280764 97044 280770 97096
rect 281074 97044 281080 97096
rect 281132 97084 281138 97096
rect 281442 97084 281448 97096
rect 281132 97056 281448 97084
rect 281132 97044 281138 97056
rect 281442 97044 281448 97056
rect 281500 97044 281506 97096
rect 283926 97044 283932 97096
rect 283984 97084 283990 97096
rect 284202 97084 284208 97096
rect 283984 97056 284208 97084
rect 283984 97044 283990 97056
rect 284202 97044 284208 97056
rect 284260 97044 284266 97096
rect 304350 97084 304356 97096
rect 287026 97056 304356 97084
rect 203518 96976 203524 97028
rect 203576 97016 203582 97028
rect 207934 97016 207940 97028
rect 203576 96988 207940 97016
rect 203576 96976 203582 96988
rect 207934 96976 207940 96988
rect 207992 96976 207998 97028
rect 214558 96976 214564 97028
rect 214616 97016 214622 97028
rect 217042 97016 217048 97028
rect 214616 96988 217048 97016
rect 214616 96976 214622 96988
rect 217042 96976 217048 96988
rect 217100 96976 217106 97028
rect 223574 96976 223580 97028
rect 223632 97016 223638 97028
rect 225138 97016 225144 97028
rect 223632 96988 225144 97016
rect 223632 96976 223638 96988
rect 225138 96976 225144 96988
rect 225196 96976 225202 97028
rect 233510 96976 233516 97028
rect 233568 97016 233574 97028
rect 234338 97016 234344 97028
rect 233568 96988 234344 97016
rect 233568 96976 233574 96988
rect 234338 96976 234344 96988
rect 234396 96976 234402 97028
rect 242066 96976 242072 97028
rect 242124 97016 242130 97028
rect 242802 97016 242808 97028
rect 242124 96988 242808 97016
rect 242124 96976 242130 96988
rect 242802 96976 242808 96988
rect 242860 96976 242866 97028
rect 247954 96976 247960 97028
rect 248012 97016 248018 97028
rect 248138 97016 248144 97028
rect 248012 96988 248144 97016
rect 248012 96976 248018 96988
rect 248138 96976 248144 96988
rect 248196 96976 248202 97028
rect 248322 96976 248328 97028
rect 248380 97016 248386 97028
rect 280798 97016 280804 97028
rect 248380 96988 280804 97016
rect 248380 96976 248386 96988
rect 280798 96976 280804 96988
rect 280856 96976 280862 97028
rect 281718 96976 281724 97028
rect 281776 97016 281782 97028
rect 282730 97016 282736 97028
rect 281776 96988 282736 97016
rect 281776 96976 281782 96988
rect 282730 96976 282736 96988
rect 282788 96976 282794 97028
rect 283098 96976 283104 97028
rect 283156 97016 283162 97028
rect 284110 97016 284116 97028
rect 283156 96988 284116 97016
rect 283156 96976 283162 96988
rect 284110 96976 284116 96988
rect 284168 96976 284174 97028
rect 284294 96976 284300 97028
rect 284352 97016 284358 97028
rect 285398 97016 285404 97028
rect 284352 96988 285404 97016
rect 284352 96976 284358 96988
rect 285398 96976 285404 96988
rect 285456 96976 285462 97028
rect 285950 96976 285956 97028
rect 286008 97016 286014 97028
rect 286686 97016 286692 97028
rect 286008 96988 286692 97016
rect 286008 96976 286014 96988
rect 286686 96976 286692 96988
rect 286744 96976 286750 97028
rect 200390 96908 200396 96960
rect 200448 96948 200454 96960
rect 201126 96948 201132 96960
rect 200448 96920 201132 96948
rect 200448 96908 200454 96920
rect 201126 96908 201132 96920
rect 201184 96908 201190 96960
rect 201586 96908 201592 96960
rect 201644 96948 201650 96960
rect 202138 96948 202144 96960
rect 201644 96920 202144 96948
rect 201644 96908 201650 96920
rect 202138 96908 202144 96920
rect 202196 96908 202202 96960
rect 204622 96908 204628 96960
rect 204680 96948 204686 96960
rect 205174 96948 205180 96960
rect 204680 96920 205180 96948
rect 204680 96908 204686 96920
rect 205174 96908 205180 96920
rect 205232 96908 205238 96960
rect 218330 96908 218336 96960
rect 218388 96948 218394 96960
rect 219158 96948 219164 96960
rect 218388 96920 219164 96948
rect 218388 96908 218394 96920
rect 219158 96908 219164 96920
rect 219216 96908 219222 96960
rect 219802 96908 219808 96960
rect 219860 96948 219866 96960
rect 220354 96948 220360 96960
rect 219860 96920 220360 96948
rect 219860 96908 219866 96920
rect 220354 96908 220360 96920
rect 220412 96908 220418 96960
rect 222562 96908 222568 96960
rect 222620 96948 222626 96960
rect 223022 96948 223028 96960
rect 222620 96920 223028 96948
rect 222620 96908 222626 96920
rect 223022 96908 223028 96920
rect 223080 96908 223086 96960
rect 225230 96908 225236 96960
rect 225288 96948 225294 96960
rect 225598 96948 225604 96960
rect 225288 96920 225604 96948
rect 225288 96908 225294 96920
rect 225598 96908 225604 96920
rect 225656 96908 225662 96960
rect 226610 96908 226616 96960
rect 226668 96948 226674 96960
rect 226886 96948 226892 96960
rect 226668 96920 226892 96948
rect 226668 96908 226674 96920
rect 226886 96908 226892 96920
rect 226944 96908 226950 96960
rect 228082 96908 228088 96960
rect 228140 96948 228146 96960
rect 228450 96948 228456 96960
rect 228140 96920 228456 96948
rect 228140 96908 228146 96920
rect 228450 96908 228456 96920
rect 228508 96908 228514 96960
rect 229462 96908 229468 96960
rect 229520 96948 229526 96960
rect 230290 96948 230296 96960
rect 229520 96920 230296 96948
rect 229520 96908 229526 96920
rect 230290 96908 230296 96920
rect 230348 96908 230354 96960
rect 230842 96908 230848 96960
rect 230900 96948 230906 96960
rect 231486 96948 231492 96960
rect 230900 96920 231492 96948
rect 230900 96908 230906 96920
rect 231486 96908 231492 96920
rect 231544 96908 231550 96960
rect 233878 96908 233884 96960
rect 233936 96948 233942 96960
rect 234614 96948 234620 96960
rect 233936 96920 234620 96948
rect 233936 96908 233942 96920
rect 234614 96908 234620 96920
rect 234672 96908 234678 96960
rect 240134 96908 240140 96960
rect 240192 96948 240198 96960
rect 241054 96948 241060 96960
rect 240192 96920 241060 96948
rect 240192 96908 240198 96920
rect 241054 96908 241060 96920
rect 241112 96908 241118 96960
rect 241882 96908 241888 96960
rect 241940 96948 241946 96960
rect 242434 96948 242440 96960
rect 241940 96920 242440 96948
rect 241940 96908 241946 96920
rect 242434 96908 242440 96920
rect 242492 96908 242498 96960
rect 242618 96908 242624 96960
rect 242676 96948 242682 96960
rect 243262 96948 243268 96960
rect 242676 96920 243268 96948
rect 242676 96908 242682 96920
rect 243262 96908 243268 96920
rect 243320 96908 243326 96960
rect 244274 96908 244280 96960
rect 244332 96948 244338 96960
rect 245286 96948 245292 96960
rect 244332 96920 245292 96948
rect 244332 96908 244338 96920
rect 245286 96908 245292 96920
rect 245344 96908 245350 96960
rect 247770 96908 247776 96960
rect 247828 96948 247834 96960
rect 248230 96948 248236 96960
rect 247828 96920 248236 96948
rect 247828 96908 247834 96920
rect 248230 96908 248236 96920
rect 248288 96908 248294 96960
rect 248966 96908 248972 96960
rect 249024 96948 249030 96960
rect 249334 96948 249340 96960
rect 249024 96920 249340 96948
rect 249024 96908 249030 96920
rect 249334 96908 249340 96920
rect 249392 96908 249398 96960
rect 249426 96908 249432 96960
rect 249484 96948 249490 96960
rect 249610 96948 249616 96960
rect 249484 96920 249616 96948
rect 249484 96908 249490 96920
rect 249610 96908 249616 96920
rect 249668 96908 249674 96960
rect 249978 96908 249984 96960
rect 250036 96948 250042 96960
rect 250806 96948 250812 96960
rect 250036 96920 250812 96948
rect 250036 96908 250042 96920
rect 250806 96908 250812 96920
rect 250864 96908 250870 96960
rect 252002 96908 252008 96960
rect 252060 96948 252066 96960
rect 252186 96948 252192 96960
rect 252060 96920 252192 96948
rect 252060 96908 252066 96920
rect 252186 96908 252192 96920
rect 252244 96908 252250 96960
rect 253198 96908 253204 96960
rect 253256 96948 253262 96960
rect 253658 96948 253664 96960
rect 253256 96920 253664 96948
rect 253256 96908 253262 96920
rect 253658 96908 253664 96920
rect 253716 96908 253722 96960
rect 254210 96908 254216 96960
rect 254268 96948 254274 96960
rect 254854 96948 254860 96960
rect 254268 96920 254860 96948
rect 254268 96908 254274 96920
rect 254854 96908 254860 96920
rect 254912 96908 254918 96960
rect 256878 96908 256884 96960
rect 256936 96948 256942 96960
rect 257706 96948 257712 96960
rect 256936 96920 257712 96948
rect 256936 96908 256942 96920
rect 257706 96908 257712 96920
rect 257764 96908 257770 96960
rect 258258 96908 258264 96960
rect 258316 96948 258322 96960
rect 258902 96948 258908 96960
rect 258316 96920 258908 96948
rect 258316 96908 258322 96920
rect 258902 96908 258908 96920
rect 258960 96908 258966 96960
rect 259086 96908 259092 96960
rect 259144 96948 259150 96960
rect 259362 96948 259368 96960
rect 259144 96920 259368 96948
rect 259144 96908 259150 96920
rect 259362 96908 259368 96920
rect 259420 96908 259426 96960
rect 260098 96908 260104 96960
rect 260156 96948 260162 96960
rect 260466 96948 260472 96960
rect 260156 96920 260472 96948
rect 260156 96908 260162 96920
rect 260466 96908 260472 96920
rect 260524 96908 260530 96960
rect 261662 96908 261668 96960
rect 261720 96948 261726 96960
rect 262030 96948 262036 96960
rect 261720 96920 262036 96948
rect 261720 96908 261726 96920
rect 262030 96908 262036 96920
rect 262088 96908 262094 96960
rect 264146 96908 264152 96960
rect 264204 96948 264210 96960
rect 264698 96948 264704 96960
rect 264204 96920 264704 96948
rect 264204 96908 264210 96920
rect 264698 96908 264704 96920
rect 264756 96908 264762 96960
rect 265710 96908 265716 96960
rect 265768 96948 265774 96960
rect 265986 96948 265992 96960
rect 265768 96920 265992 96948
rect 265768 96908 265774 96920
rect 265986 96908 265992 96920
rect 266044 96908 266050 96960
rect 266354 96908 266360 96960
rect 266412 96948 266418 96960
rect 267366 96948 267372 96960
rect 266412 96920 267372 96948
rect 266412 96908 266418 96920
rect 267366 96908 267372 96920
rect 267424 96908 267430 96960
rect 268194 96908 268200 96960
rect 268252 96948 268258 96960
rect 268930 96948 268936 96960
rect 268252 96920 268936 96948
rect 268252 96908 268258 96920
rect 268930 96908 268936 96920
rect 268988 96908 268994 96960
rect 269390 96908 269396 96960
rect 269448 96948 269454 96960
rect 269942 96948 269948 96960
rect 269448 96920 269948 96948
rect 269448 96908 269454 96920
rect 269942 96908 269948 96920
rect 270000 96908 270006 96960
rect 271414 96908 271420 96960
rect 271472 96948 271478 96960
rect 271782 96948 271788 96960
rect 271472 96920 271788 96948
rect 271472 96908 271478 96920
rect 271782 96908 271788 96920
rect 271840 96908 271846 96960
rect 272610 96908 272616 96960
rect 272668 96948 272674 96960
rect 273070 96948 273076 96960
rect 272668 96920 273076 96948
rect 272668 96908 272674 96920
rect 273070 96908 273076 96920
rect 273128 96908 273134 96960
rect 273806 96908 273812 96960
rect 273864 96948 273870 96960
rect 274358 96948 274364 96960
rect 273864 96920 274364 96948
rect 273864 96908 273870 96920
rect 274358 96908 274364 96920
rect 274416 96908 274422 96960
rect 277578 96948 277584 96960
rect 275940 96920 277584 96948
rect 204438 96840 204444 96892
rect 204496 96880 204502 96892
rect 204990 96880 204996 96892
rect 204496 96852 204996 96880
rect 204496 96840 204502 96852
rect 204990 96840 204996 96852
rect 205048 96840 205054 96892
rect 219618 96840 219624 96892
rect 219676 96880 219682 96892
rect 220170 96880 220176 96892
rect 219676 96852 220176 96880
rect 219676 96840 219682 96852
rect 220170 96840 220176 96852
rect 220228 96840 220234 96892
rect 222378 96840 222384 96892
rect 222436 96880 222442 96892
rect 223390 96880 223396 96892
rect 222436 96852 223396 96880
rect 222436 96840 222442 96852
rect 223390 96840 223396 96852
rect 223448 96840 223454 96892
rect 225414 96840 225420 96892
rect 225472 96880 225478 96892
rect 226058 96880 226064 96892
rect 225472 96852 226064 96880
rect 225472 96840 225478 96852
rect 226058 96840 226064 96852
rect 226116 96840 226122 96892
rect 226794 96840 226800 96892
rect 226852 96880 226858 96892
rect 227438 96880 227444 96892
rect 226852 96852 227444 96880
rect 226852 96840 226858 96852
rect 227438 96840 227444 96852
rect 227496 96840 227502 96892
rect 227898 96840 227904 96892
rect 227956 96880 227962 96892
rect 228818 96880 228824 96892
rect 227956 96852 228824 96880
rect 227956 96840 227962 96852
rect 228818 96840 228824 96852
rect 228876 96840 228882 96892
rect 231026 96840 231032 96892
rect 231084 96880 231090 96892
rect 231302 96880 231308 96892
rect 231084 96852 231308 96880
rect 231084 96840 231090 96852
rect 231302 96840 231308 96852
rect 231360 96840 231366 96892
rect 233326 96840 233332 96892
rect 233384 96880 233390 96892
rect 234062 96880 234068 96892
rect 233384 96852 234068 96880
rect 233384 96840 233390 96852
rect 234062 96840 234068 96852
rect 234120 96840 234126 96892
rect 237374 96840 237380 96892
rect 237432 96880 237438 96892
rect 240502 96880 240508 96892
rect 237432 96852 240508 96880
rect 237432 96840 237438 96852
rect 240502 96840 240508 96852
rect 240560 96840 240566 96892
rect 242250 96840 242256 96892
rect 242308 96880 242314 96892
rect 242710 96880 242716 96892
rect 242308 96852 242716 96880
rect 242308 96840 242314 96852
rect 242710 96840 242716 96852
rect 242768 96840 242774 96892
rect 243078 96840 243084 96892
rect 243136 96880 243142 96892
rect 244090 96880 244096 96892
rect 243136 96852 244096 96880
rect 243136 96840 243142 96852
rect 244090 96840 244096 96852
rect 244148 96840 244154 96892
rect 244734 96840 244740 96892
rect 244792 96880 244798 96892
rect 245562 96880 245568 96892
rect 244792 96852 245568 96880
rect 244792 96840 244798 96852
rect 245562 96840 245568 96852
rect 245620 96840 245626 96892
rect 247126 96840 247132 96892
rect 247184 96880 247190 96892
rect 248138 96880 248144 96892
rect 247184 96852 248144 96880
rect 247184 96840 247190 96852
rect 248138 96840 248144 96852
rect 248196 96840 248202 96892
rect 251358 96840 251364 96892
rect 251416 96880 251422 96892
rect 252278 96880 252284 96892
rect 251416 96852 252284 96880
rect 251416 96840 251422 96852
rect 252278 96840 252284 96852
rect 252336 96840 252342 96892
rect 252830 96840 252836 96892
rect 252888 96880 252894 96892
rect 253566 96880 253572 96892
rect 252888 96852 253572 96880
rect 252888 96840 252894 96852
rect 253566 96840 253572 96852
rect 253624 96840 253630 96892
rect 254762 96840 254768 96892
rect 254820 96880 254826 96892
rect 255222 96880 255228 96892
rect 254820 96852 255228 96880
rect 254820 96840 254826 96852
rect 255222 96840 255228 96852
rect 255280 96840 255286 96892
rect 257062 96840 257068 96892
rect 257120 96880 257126 96892
rect 257890 96880 257896 96892
rect 257120 96852 257896 96880
rect 257120 96840 257126 96852
rect 257890 96840 257896 96852
rect 257948 96840 257954 96892
rect 260282 96840 260288 96892
rect 260340 96880 260346 96892
rect 260742 96880 260748 96892
rect 260340 96852 260748 96880
rect 260340 96840 260346 96852
rect 260742 96840 260748 96852
rect 260800 96840 260806 96892
rect 263870 96840 263876 96892
rect 263928 96880 263934 96892
rect 264882 96880 264888 96892
rect 263928 96852 264888 96880
rect 263928 96840 263934 96852
rect 264882 96840 264888 96852
rect 264940 96840 264946 96892
rect 265342 96840 265348 96892
rect 265400 96880 265406 96892
rect 266170 96880 266176 96892
rect 265400 96852 266176 96880
rect 265400 96840 265406 96852
rect 266170 96840 266176 96852
rect 266228 96840 266234 96892
rect 266906 96840 266912 96892
rect 266964 96880 266970 96892
rect 267642 96880 267648 96892
rect 266964 96852 267648 96880
rect 266964 96840 266970 96852
rect 267642 96840 267648 96852
rect 267700 96840 267706 96892
rect 270954 96840 270960 96892
rect 271012 96880 271018 96892
rect 271012 96852 271920 96880
rect 271012 96840 271018 96852
rect 200850 96772 200856 96824
rect 200908 96812 200914 96824
rect 207382 96812 207388 96824
rect 200908 96784 207388 96812
rect 200908 96772 200914 96784
rect 207382 96772 207388 96784
rect 207440 96772 207446 96824
rect 216858 96772 216864 96824
rect 216916 96812 216922 96824
rect 217134 96812 217140 96824
rect 216916 96784 217140 96812
rect 216916 96772 216922 96784
rect 217134 96772 217140 96784
rect 217192 96772 217198 96824
rect 229738 96772 229744 96824
rect 229796 96812 229802 96824
rect 233970 96812 233976 96824
rect 229796 96784 233976 96812
rect 229796 96772 229802 96784
rect 233970 96772 233976 96784
rect 234028 96772 234034 96824
rect 235074 96772 235080 96824
rect 235132 96812 235138 96824
rect 235534 96812 235540 96824
rect 235132 96784 235540 96812
rect 235132 96772 235138 96784
rect 235534 96772 235540 96784
rect 235592 96772 235598 96824
rect 236362 96772 236368 96824
rect 236420 96812 236426 96824
rect 237098 96812 237104 96824
rect 236420 96784 237104 96812
rect 236420 96772 236426 96784
rect 237098 96772 237104 96784
rect 237156 96772 237162 96824
rect 244550 96772 244556 96824
rect 244608 96812 244614 96824
rect 245102 96812 245108 96824
rect 244608 96784 245108 96812
rect 244608 96772 244614 96784
rect 245102 96772 245108 96784
rect 245160 96772 245166 96824
rect 248598 96772 248604 96824
rect 248656 96812 248662 96824
rect 249610 96812 249616 96824
rect 248656 96784 249616 96812
rect 248656 96772 248662 96784
rect 249610 96772 249616 96784
rect 249668 96772 249674 96824
rect 251542 96772 251548 96824
rect 251600 96812 251606 96824
rect 252370 96812 252376 96824
rect 251600 96784 252376 96812
rect 251600 96772 251606 96784
rect 252370 96772 252376 96784
rect 252428 96772 252434 96824
rect 252554 96772 252560 96824
rect 252612 96812 252618 96824
rect 253842 96812 253848 96824
rect 252612 96784 253848 96812
rect 252612 96772 252618 96784
rect 253842 96772 253848 96784
rect 253900 96772 253906 96824
rect 254026 96772 254032 96824
rect 254084 96812 254090 96824
rect 254946 96812 254952 96824
rect 254084 96784 254952 96812
rect 254084 96772 254090 96784
rect 254946 96772 254952 96784
rect 255004 96772 255010 96824
rect 257430 96772 257436 96824
rect 257488 96812 257494 96824
rect 257798 96812 257804 96824
rect 257488 96784 257804 96812
rect 257488 96772 257494 96784
rect 257798 96772 257804 96784
rect 257856 96772 257862 96824
rect 258626 96772 258632 96824
rect 258684 96812 258690 96824
rect 259086 96812 259092 96824
rect 258684 96784 259092 96812
rect 258684 96772 258690 96784
rect 259086 96772 259092 96784
rect 259144 96772 259150 96824
rect 259638 96772 259644 96824
rect 259696 96812 259702 96824
rect 260650 96812 260656 96824
rect 259696 96784 260656 96812
rect 259696 96772 259702 96784
rect 260650 96772 260656 96784
rect 260708 96772 260714 96824
rect 261110 96772 261116 96824
rect 261168 96812 261174 96824
rect 261938 96812 261944 96824
rect 261168 96784 261944 96812
rect 261168 96772 261174 96784
rect 261938 96772 261944 96784
rect 261996 96772 262002 96824
rect 262306 96772 262312 96824
rect 262364 96812 262370 96824
rect 263134 96812 263140 96824
rect 262364 96784 263140 96812
rect 262364 96772 262370 96784
rect 263134 96772 263140 96784
rect 263192 96772 263198 96824
rect 265158 96772 265164 96824
rect 265216 96812 265222 96824
rect 266262 96812 266268 96824
rect 265216 96784 266268 96812
rect 265216 96772 265222 96784
rect 266262 96772 266268 96784
rect 266320 96772 266326 96824
rect 266538 96772 266544 96824
rect 266596 96812 266602 96824
rect 267550 96812 267556 96824
rect 266596 96784 267556 96812
rect 266596 96772 266602 96784
rect 267550 96772 267556 96784
rect 267608 96772 267614 96824
rect 269574 96772 269580 96824
rect 269632 96812 269638 96824
rect 270310 96812 270316 96824
rect 269632 96784 270316 96812
rect 269632 96772 269638 96784
rect 270310 96772 270316 96784
rect 270368 96772 270374 96824
rect 270770 96772 270776 96824
rect 270828 96812 270834 96824
rect 271690 96812 271696 96824
rect 270828 96784 271696 96812
rect 270828 96772 270834 96784
rect 271690 96772 271696 96784
rect 271748 96772 271754 96824
rect 271892 96812 271920 96852
rect 271966 96840 271972 96892
rect 272024 96880 272030 96892
rect 272978 96880 272984 96892
rect 272024 96852 272984 96880
rect 272024 96840 272030 96852
rect 272978 96840 272984 96852
rect 273036 96840 273042 96892
rect 273990 96840 273996 96892
rect 274048 96880 274054 96892
rect 274542 96880 274548 96892
rect 274048 96852 274548 96880
rect 274048 96840 274054 96852
rect 274542 96840 274548 96852
rect 274600 96840 274606 96892
rect 275940 96880 275968 96920
rect 277578 96908 277584 96920
rect 277636 96908 277642 96960
rect 277670 96908 277676 96960
rect 277728 96948 277734 96960
rect 278314 96948 278320 96960
rect 277728 96920 278320 96948
rect 277728 96908 277734 96920
rect 278314 96908 278320 96920
rect 278372 96908 278378 96960
rect 278866 96908 278872 96960
rect 278924 96948 278930 96960
rect 279786 96948 279792 96960
rect 278924 96920 279792 96948
rect 278924 96908 278930 96920
rect 279786 96908 279792 96920
rect 279844 96908 279850 96960
rect 282270 96908 282276 96960
rect 282328 96948 282334 96960
rect 282638 96948 282644 96960
rect 282328 96920 282644 96948
rect 282328 96908 282334 96920
rect 282638 96908 282644 96920
rect 282696 96908 282702 96960
rect 283466 96908 283472 96960
rect 283524 96948 283530 96960
rect 283926 96948 283932 96960
rect 283524 96920 283932 96948
rect 283524 96908 283530 96920
rect 283926 96908 283932 96920
rect 283984 96908 283990 96960
rect 284754 96908 284760 96960
rect 284812 96948 284818 96960
rect 285306 96948 285312 96960
rect 284812 96920 285312 96948
rect 284812 96908 284818 96920
rect 285306 96908 285312 96920
rect 285364 96908 285370 96960
rect 286502 96908 286508 96960
rect 286560 96948 286566 96960
rect 286778 96948 286784 96960
rect 286560 96920 286784 96948
rect 286560 96908 286566 96920
rect 286778 96908 286784 96920
rect 286836 96908 286842 96960
rect 274928 96852 275968 96880
rect 274928 96812 274956 96852
rect 276106 96840 276112 96892
rect 276164 96880 276170 96892
rect 287026 96880 287054 97056
rect 304350 97044 304356 97056
rect 304408 97044 304414 97096
rect 287146 96976 287152 97028
rect 287204 97016 287210 97028
rect 288342 97016 288348 97028
rect 287204 96988 288348 97016
rect 287204 96976 287210 96988
rect 288342 96976 288348 96988
rect 288400 96976 288406 97028
rect 291562 96976 291568 97028
rect 291620 97016 291626 97028
rect 292390 97016 292396 97028
rect 291620 96988 292396 97016
rect 291620 96976 291626 96988
rect 292390 96976 292396 96988
rect 292448 96976 292454 97028
rect 292758 96976 292764 97028
rect 292816 97016 292822 97028
rect 293770 97016 293776 97028
rect 292816 96988 293776 97016
rect 292816 96976 292822 96988
rect 293770 96976 293776 96988
rect 293828 96976 293834 97028
rect 294046 96976 294052 97028
rect 294104 97016 294110 97028
rect 295058 97016 295064 97028
rect 294104 96988 295064 97016
rect 294104 96976 294110 96988
rect 295058 96976 295064 96988
rect 295116 96976 295122 97028
rect 287330 96908 287336 96960
rect 287388 96948 287394 96960
rect 287882 96948 287888 96960
rect 287388 96920 287888 96948
rect 287388 96908 287394 96920
rect 287882 96908 287888 96920
rect 287940 96908 287946 96960
rect 288986 96908 288992 96960
rect 289044 96948 289050 96960
rect 289538 96948 289544 96960
rect 289044 96920 289544 96948
rect 289044 96908 289050 96920
rect 289538 96908 289544 96920
rect 289596 96908 289602 96960
rect 290182 96908 290188 96960
rect 290240 96948 290246 96960
rect 291102 96948 291108 96960
rect 290240 96920 291108 96948
rect 290240 96908 290246 96920
rect 291102 96908 291108 96920
rect 291160 96908 291166 96960
rect 292022 96908 292028 96960
rect 292080 96948 292086 96960
rect 292298 96948 292304 96960
rect 292080 96920 292304 96948
rect 292080 96908 292086 96920
rect 292298 96908 292304 96920
rect 292356 96908 292362 96960
rect 293218 96908 293224 96960
rect 293276 96948 293282 96960
rect 293586 96948 293592 96960
rect 293276 96920 293592 96948
rect 293276 96908 293282 96920
rect 293586 96908 293592 96920
rect 293644 96908 293650 96960
rect 294414 96908 294420 96960
rect 294472 96948 294478 96960
rect 294874 96948 294880 96960
rect 294472 96920 294880 96948
rect 294472 96908 294478 96920
rect 294874 96908 294880 96920
rect 294932 96908 294938 96960
rect 295426 96908 295432 96960
rect 295484 96948 295490 96960
rect 298370 96948 298376 96960
rect 295484 96920 298376 96948
rect 295484 96908 295490 96920
rect 298370 96908 298376 96920
rect 298428 96908 298434 96960
rect 298462 96908 298468 96960
rect 298520 96948 298526 96960
rect 299014 96948 299020 96960
rect 298520 96920 299020 96948
rect 298520 96908 298526 96920
rect 299014 96908 299020 96920
rect 299072 96908 299078 96960
rect 276164 96852 287054 96880
rect 276164 96840 276170 96852
rect 287790 96840 287796 96892
rect 287848 96880 287854 96892
rect 288066 96880 288072 96892
rect 287848 96852 288072 96880
rect 287848 96840 287854 96852
rect 288066 96840 288072 96852
rect 288124 96840 288130 96892
rect 290826 96840 290832 96892
rect 290884 96880 290890 96892
rect 291010 96880 291016 96892
rect 290884 96852 291016 96880
rect 290884 96840 290890 96852
rect 291010 96840 291016 96852
rect 291068 96840 291074 96892
rect 291378 96840 291384 96892
rect 291436 96880 291442 96892
rect 292206 96880 292212 96892
rect 291436 96852 292212 96880
rect 291436 96840 291442 96852
rect 292206 96840 292212 96852
rect 292264 96840 292270 96892
rect 292574 96840 292580 96892
rect 292632 96880 292638 96892
rect 293402 96880 293408 96892
rect 292632 96852 293408 96880
rect 292632 96840 292638 96852
rect 293402 96840 293408 96852
rect 293460 96840 293466 96892
rect 294782 96840 294788 96892
rect 294840 96880 294846 96892
rect 295242 96880 295248 96892
rect 294840 96852 295248 96880
rect 294840 96840 294846 96852
rect 295242 96840 295248 96852
rect 295300 96840 295306 96892
rect 295794 96840 295800 96892
rect 295852 96880 295858 96892
rect 296530 96880 296536 96892
rect 295852 96852 296536 96880
rect 295852 96840 295858 96852
rect 296530 96840 296536 96852
rect 296588 96840 296594 96892
rect 298094 96840 298100 96892
rect 298152 96880 298158 96892
rect 301498 96880 301504 96892
rect 298152 96852 301504 96880
rect 298152 96840 298158 96852
rect 301498 96840 301504 96852
rect 301556 96840 301562 96892
rect 271892 96784 274956 96812
rect 275002 96772 275008 96824
rect 275060 96812 275066 96824
rect 275738 96812 275744 96824
rect 275060 96784 275744 96812
rect 275060 96772 275066 96784
rect 275738 96772 275744 96784
rect 275796 96772 275802 96824
rect 276198 96772 276204 96824
rect 276256 96812 276262 96824
rect 276934 96812 276940 96824
rect 276256 96784 276940 96812
rect 276256 96772 276262 96784
rect 276934 96772 276940 96784
rect 276992 96772 276998 96824
rect 277486 96772 277492 96824
rect 277544 96812 277550 96824
rect 278406 96812 278412 96824
rect 277544 96784 278412 96812
rect 277544 96772 277550 96784
rect 278406 96772 278412 96784
rect 278464 96772 278470 96824
rect 280430 96772 280436 96824
rect 280488 96812 280494 96824
rect 281258 96812 281264 96824
rect 280488 96784 281264 96812
rect 280488 96772 280494 96784
rect 281258 96772 281264 96784
rect 281316 96772 281322 96824
rect 286134 96772 286140 96824
rect 286192 96812 286198 96824
rect 286870 96812 286876 96824
rect 286192 96784 286876 96812
rect 286192 96772 286198 96784
rect 286870 96772 286876 96784
rect 286928 96772 286934 96824
rect 291838 96812 291844 96824
rect 287026 96784 291844 96812
rect 215938 96704 215944 96756
rect 215996 96744 216002 96756
rect 218238 96744 218244 96756
rect 215996 96716 218244 96744
rect 215996 96704 216002 96716
rect 218238 96704 218244 96716
rect 218296 96704 218302 96756
rect 231118 96704 231124 96756
rect 231176 96744 231182 96756
rect 236086 96744 236092 96756
rect 231176 96716 236092 96744
rect 231176 96704 231182 96716
rect 236086 96704 236092 96716
rect 236144 96704 236150 96756
rect 245746 96704 245752 96756
rect 245804 96744 245810 96756
rect 245804 96716 246896 96744
rect 245804 96704 245810 96716
rect 246868 96688 246896 96716
rect 250162 96704 250168 96756
rect 250220 96744 250226 96756
rect 250898 96744 250904 96756
rect 250220 96716 250904 96744
rect 250220 96704 250226 96716
rect 250898 96704 250904 96716
rect 250956 96704 250962 96756
rect 261294 96704 261300 96756
rect 261352 96744 261358 96756
rect 261846 96744 261852 96756
rect 261352 96716 261852 96744
rect 261352 96704 261358 96716
rect 261846 96704 261852 96716
rect 261904 96704 261910 96756
rect 267734 96704 267740 96756
rect 267792 96744 267798 96756
rect 268562 96744 268568 96756
rect 267792 96716 268568 96744
rect 267792 96704 267798 96716
rect 268562 96704 268568 96716
rect 268620 96704 268626 96756
rect 269206 96704 269212 96756
rect 269264 96744 269270 96756
rect 273898 96744 273904 96756
rect 269264 96716 273904 96744
rect 269264 96704 269270 96716
rect 273898 96704 273904 96716
rect 273956 96704 273962 96756
rect 275186 96704 275192 96756
rect 275244 96744 275250 96756
rect 275922 96744 275928 96756
rect 275244 96716 275928 96744
rect 275244 96704 275250 96716
rect 275922 96704 275928 96716
rect 275980 96704 275986 96756
rect 276658 96704 276664 96756
rect 276716 96744 276722 96756
rect 277302 96744 277308 96756
rect 276716 96716 277308 96744
rect 276716 96704 276722 96716
rect 277302 96704 277308 96716
rect 277360 96704 277366 96756
rect 280614 96704 280620 96756
rect 280672 96744 280678 96756
rect 287026 96744 287054 96784
rect 291838 96772 291844 96784
rect 291896 96772 291902 96824
rect 295610 96772 295616 96824
rect 295668 96812 295674 96824
rect 296346 96812 296352 96824
rect 295668 96784 296352 96812
rect 295668 96772 295674 96784
rect 296346 96772 296352 96784
rect 296404 96772 296410 96824
rect 280672 96716 287054 96744
rect 280672 96704 280678 96716
rect 290366 96704 290372 96756
rect 290424 96744 290430 96756
rect 291010 96744 291016 96756
rect 290424 96716 291016 96744
rect 290424 96704 290430 96716
rect 291010 96704 291016 96716
rect 291068 96704 291074 96756
rect 210510 96636 210516 96688
rect 210568 96676 210574 96688
rect 211614 96676 211620 96688
rect 210568 96648 211620 96676
rect 210568 96636 210574 96648
rect 211614 96636 211620 96648
rect 211672 96636 211678 96688
rect 233970 96636 233976 96688
rect 234028 96676 234034 96688
rect 238110 96676 238116 96688
rect 234028 96648 238116 96676
rect 234028 96636 234034 96648
rect 238110 96636 238116 96648
rect 238168 96636 238174 96688
rect 245930 96636 245936 96688
rect 245988 96676 245994 96688
rect 246758 96676 246764 96688
rect 245988 96648 246764 96676
rect 245988 96636 245994 96648
rect 246758 96636 246764 96648
rect 246816 96636 246822 96688
rect 246850 96636 246856 96688
rect 246908 96636 246914 96688
rect 267918 96636 267924 96688
rect 267976 96676 267982 96688
rect 269022 96676 269028 96688
rect 267976 96648 269028 96676
rect 267976 96636 267982 96648
rect 269022 96636 269028 96648
rect 269080 96636 269086 96688
rect 280246 96636 280252 96688
rect 280304 96676 280310 96688
rect 281442 96676 281448 96688
rect 280304 96648 281448 96676
rect 280304 96636 280310 96648
rect 281442 96636 281448 96648
rect 281500 96636 281506 96688
rect 288526 96636 288532 96688
rect 288584 96676 288590 96688
rect 289262 96676 289268 96688
rect 288584 96648 289268 96676
rect 288584 96636 288590 96648
rect 289262 96636 289268 96648
rect 289320 96636 289326 96688
rect 298278 96636 298284 96688
rect 298336 96676 298342 96688
rect 299198 96676 299204 96688
rect 298336 96648 299204 96676
rect 298336 96636 298342 96648
rect 299198 96636 299204 96648
rect 299256 96636 299262 96688
rect 191190 96568 191196 96620
rect 191248 96608 191254 96620
rect 232038 96608 232044 96620
rect 191248 96580 232044 96608
rect 191248 96568 191254 96580
rect 232038 96568 232044 96580
rect 232096 96568 232102 96620
rect 251174 96568 251180 96620
rect 251232 96608 251238 96620
rect 302326 96608 302332 96620
rect 251232 96580 302332 96608
rect 251232 96568 251238 96580
rect 302326 96568 302332 96580
rect 302384 96568 302390 96620
rect 176562 96500 176568 96552
rect 176620 96540 176626 96552
rect 216766 96540 216772 96552
rect 176620 96512 216772 96540
rect 176620 96500 176626 96512
rect 216766 96500 216772 96512
rect 216824 96500 216830 96552
rect 271506 96500 271512 96552
rect 271564 96540 271570 96552
rect 356054 96540 356060 96552
rect 271564 96512 356060 96540
rect 271564 96500 271570 96512
rect 356054 96500 356060 96512
rect 356112 96500 356118 96552
rect 186958 96432 186964 96484
rect 187016 96472 187022 96484
rect 231762 96472 231768 96484
rect 187016 96444 231768 96472
rect 187016 96432 187022 96444
rect 231762 96432 231768 96444
rect 231820 96432 231826 96484
rect 262122 96432 262128 96484
rect 262180 96472 262186 96484
rect 347038 96472 347044 96484
rect 262180 96444 347044 96472
rect 262180 96432 262186 96444
rect 347038 96432 347044 96444
rect 347096 96432 347102 96484
rect 161382 96364 161388 96416
rect 161440 96404 161446 96416
rect 209406 96404 209412 96416
rect 161440 96376 209412 96404
rect 161440 96364 161446 96376
rect 209406 96364 209412 96376
rect 209464 96364 209470 96416
rect 284202 96364 284208 96416
rect 284260 96404 284266 96416
rect 411898 96404 411904 96416
rect 284260 96376 411904 96404
rect 284260 96364 284266 96376
rect 411898 96364 411904 96376
rect 411956 96364 411962 96416
rect 169662 96296 169668 96348
rect 169720 96336 169726 96348
rect 220630 96336 220636 96348
rect 169720 96308 220636 96336
rect 169720 96296 169726 96308
rect 220630 96296 220636 96308
rect 220688 96296 220694 96348
rect 285122 96296 285128 96348
rect 285180 96336 285186 96348
rect 465718 96336 465724 96348
rect 285180 96308 465724 96336
rect 285180 96296 285186 96308
rect 465718 96296 465724 96308
rect 465776 96296 465782 96348
rect 165522 96228 165528 96280
rect 165580 96268 165586 96280
rect 218054 96268 218060 96280
rect 165580 96240 218060 96268
rect 165580 96228 165586 96240
rect 218054 96228 218060 96240
rect 218112 96228 218118 96280
rect 283282 96228 283288 96280
rect 283340 96268 283346 96280
rect 475378 96268 475384 96280
rect 283340 96240 475384 96268
rect 283340 96228 283346 96240
rect 475378 96228 475384 96240
rect 475436 96228 475442 96280
rect 173158 96160 173164 96212
rect 173216 96200 173222 96212
rect 229370 96200 229376 96212
rect 173216 96172 229376 96200
rect 173216 96160 173222 96172
rect 229370 96160 229376 96172
rect 229428 96160 229434 96212
rect 282086 96160 282092 96212
rect 282144 96200 282150 96212
rect 479518 96200 479524 96212
rect 282144 96172 479524 96200
rect 282144 96160 282150 96172
rect 479518 96160 479524 96172
rect 479576 96160 479582 96212
rect 166258 96092 166264 96144
rect 166316 96132 166322 96144
rect 225966 96132 225972 96144
rect 166316 96104 225972 96132
rect 166316 96092 166322 96104
rect 225966 96092 225972 96104
rect 226024 96092 226030 96144
rect 297450 96092 297456 96144
rect 297508 96132 297514 96144
rect 494054 96132 494060 96144
rect 297508 96104 494060 96132
rect 297508 96092 297514 96104
rect 494054 96092 494060 96104
rect 494112 96092 494118 96144
rect 126882 96024 126888 96076
rect 126940 96064 126946 96076
rect 204898 96064 204904 96076
rect 126940 96036 204904 96064
rect 126940 96024 126946 96036
rect 204898 96024 204904 96036
rect 204956 96024 204962 96076
rect 213178 96024 213184 96076
rect 213236 96064 213242 96076
rect 235994 96064 236000 96076
rect 213236 96036 236000 96064
rect 213236 96024 213242 96036
rect 235994 96024 236000 96036
rect 236052 96024 236058 96076
rect 243906 96024 243912 96076
rect 243964 96064 243970 96076
rect 269114 96064 269120 96076
rect 243964 96036 269120 96064
rect 243964 96024 243970 96036
rect 269114 96024 269120 96036
rect 269172 96024 269178 96076
rect 282822 96024 282828 96076
rect 282880 96064 282886 96076
rect 483014 96064 483020 96076
rect 282880 96036 483020 96064
rect 282880 96024 282886 96036
rect 483014 96024 483020 96036
rect 483072 96024 483078 96076
rect 37182 95956 37188 96008
rect 37240 95996 37246 96008
rect 173802 95996 173808 96008
rect 37240 95968 173808 95996
rect 37240 95956 37246 95968
rect 173802 95956 173808 95968
rect 173860 95956 173866 96008
rect 183462 95956 183468 96008
rect 183520 95996 183526 96008
rect 231210 95996 231216 96008
rect 183520 95968 231216 95996
rect 183520 95956 183526 95968
rect 231210 95956 231216 95968
rect 231268 95956 231274 96008
rect 237742 95956 237748 96008
rect 237800 95996 237806 96008
rect 238386 95996 238392 96008
rect 237800 95968 238392 95996
rect 237800 95956 237806 95968
rect 238386 95956 238392 95968
rect 238444 95956 238450 96008
rect 246298 95956 246304 96008
rect 246356 95996 246362 96008
rect 281534 95996 281540 96008
rect 246356 95968 281540 95996
rect 246356 95956 246362 95968
rect 281534 95956 281540 95968
rect 281592 95956 281598 96008
rect 285858 95956 285864 96008
rect 285916 95996 285922 96008
rect 500954 95996 500960 96008
rect 285916 95968 500960 95996
rect 285916 95956 285922 95968
rect 500954 95956 500960 95968
rect 501012 95956 501018 96008
rect 12250 95888 12256 95940
rect 12308 95928 12314 95940
rect 202046 95928 202052 95940
rect 12308 95900 202052 95928
rect 12308 95888 12314 95900
rect 202046 95888 202052 95900
rect 202104 95888 202110 95940
rect 202138 95888 202144 95940
rect 202196 95928 202202 95940
rect 234246 95928 234252 95940
rect 202196 95900 234252 95928
rect 202196 95888 202202 95900
rect 234246 95888 234252 95900
rect 234304 95888 234310 95940
rect 247954 95888 247960 95940
rect 248012 95928 248018 95940
rect 285766 95928 285772 95940
rect 248012 95900 285772 95928
rect 248012 95888 248018 95900
rect 285766 95888 285772 95900
rect 285824 95888 285830 95940
rect 291194 95888 291200 95940
rect 291252 95928 291258 95940
rect 532694 95928 532700 95940
rect 291252 95900 532700 95928
rect 291252 95888 291258 95900
rect 532694 95888 532700 95900
rect 532752 95888 532758 95940
rect 179322 95820 179328 95872
rect 179380 95860 179386 95872
rect 218146 95860 218152 95872
rect 179380 95832 218152 95860
rect 179380 95820 179386 95832
rect 218146 95820 218152 95832
rect 218204 95820 218210 95872
rect 231210 95820 231216 95872
rect 231268 95860 231274 95872
rect 236638 95860 236644 95872
rect 231268 95832 236644 95860
rect 231268 95820 231274 95832
rect 236638 95820 236644 95832
rect 236696 95820 236702 95872
rect 251818 95820 251824 95872
rect 251876 95860 251882 95872
rect 302234 95860 302240 95872
rect 251876 95832 302240 95860
rect 251876 95820 251882 95832
rect 302234 95820 302240 95832
rect 302292 95820 302298 95872
rect 195238 95752 195244 95804
rect 195296 95792 195302 95804
rect 232958 95792 232964 95804
rect 195296 95764 232964 95792
rect 195296 95752 195302 95764
rect 232958 95752 232964 95764
rect 233016 95752 233022 95804
rect 250530 95752 250536 95804
rect 250588 95792 250594 95804
rect 299566 95792 299572 95804
rect 250588 95764 299572 95792
rect 250588 95752 250594 95764
rect 299566 95752 299572 95764
rect 299624 95752 299630 95804
rect 197262 95684 197268 95736
rect 197320 95724 197326 95736
rect 211154 95724 211160 95736
rect 197320 95696 211160 95724
rect 197320 95684 197326 95696
rect 211154 95684 211160 95696
rect 211212 95684 211218 95736
rect 293862 95684 293868 95736
rect 293920 95724 293926 95736
rect 320818 95724 320824 95736
rect 293920 95696 320824 95724
rect 293920 95684 293926 95696
rect 320818 95684 320824 95696
rect 320876 95684 320882 95736
rect 235350 95412 235356 95464
rect 235408 95452 235414 95464
rect 235810 95452 235816 95464
rect 235408 95424 235816 95452
rect 235408 95412 235414 95424
rect 235810 95412 235816 95424
rect 235868 95412 235874 95464
rect 233142 95276 233148 95328
rect 233200 95316 233206 95328
rect 239674 95316 239680 95328
rect 233200 95288 239680 95316
rect 233200 95276 233206 95288
rect 239674 95276 239680 95288
rect 239732 95276 239738 95328
rect 162762 95140 162768 95192
rect 162820 95180 162826 95192
rect 227714 95180 227720 95192
rect 162820 95152 227720 95180
rect 162820 95140 162826 95152
rect 227714 95140 227720 95152
rect 227772 95140 227778 95192
rect 255406 95140 255412 95192
rect 255464 95180 255470 95192
rect 324406 95180 324412 95192
rect 255464 95152 324412 95180
rect 255464 95140 255470 95152
rect 324406 95140 324412 95152
rect 324464 95140 324470 95192
rect 158622 95072 158628 95124
rect 158680 95112 158686 95124
rect 226978 95112 226984 95124
rect 158680 95084 226984 95112
rect 158680 95072 158686 95084
rect 226978 95072 226984 95084
rect 227036 95072 227042 95124
rect 256050 95072 256056 95124
rect 256108 95112 256114 95124
rect 327074 95112 327080 95124
rect 256108 95084 327080 95112
rect 256108 95072 256114 95084
rect 327074 95072 327080 95084
rect 327132 95072 327138 95124
rect 155218 95004 155224 95056
rect 155276 95044 155282 95056
rect 226334 95044 226340 95056
rect 155276 95016 226340 95044
rect 155276 95004 155282 95016
rect 226334 95004 226340 95016
rect 226392 95004 226398 95056
rect 258442 95004 258448 95056
rect 258500 95044 258506 95056
rect 340874 95044 340880 95056
rect 258500 95016 340880 95044
rect 258500 95004 258506 95016
rect 340874 95004 340880 95016
rect 340932 95004 340938 95056
rect 147582 94936 147588 94988
rect 147640 94976 147646 94988
rect 223574 94976 223580 94988
rect 147640 94948 223580 94976
rect 147640 94936 147646 94948
rect 223574 94936 223580 94948
rect 223632 94936 223638 94988
rect 262674 94936 262680 94988
rect 262732 94976 262738 94988
rect 364978 94976 364984 94988
rect 262732 94948 364984 94976
rect 262732 94936 262738 94948
rect 364978 94936 364984 94948
rect 365036 94936 365042 94988
rect 146202 94868 146208 94920
rect 146260 94908 146266 94920
rect 224954 94908 224960 94920
rect 146260 94880 224960 94908
rect 146260 94868 146266 94880
rect 224954 94868 224960 94880
rect 225012 94868 225018 94920
rect 276474 94868 276480 94920
rect 276532 94908 276538 94920
rect 385678 94908 385684 94920
rect 276532 94880 385684 94908
rect 276532 94868 276538 94880
rect 385678 94868 385684 94880
rect 385736 94868 385742 94920
rect 137278 94800 137284 94852
rect 137336 94840 137342 94852
rect 223298 94840 223304 94852
rect 137336 94812 223304 94840
rect 137336 94800 137342 94812
rect 223298 94800 223304 94812
rect 223356 94800 223362 94852
rect 279234 94800 279240 94852
rect 279292 94840 279298 94852
rect 429838 94840 429844 94852
rect 279292 94812 429844 94840
rect 279292 94800 279298 94812
rect 429838 94800 429844 94812
rect 429896 94800 429902 94852
rect 114462 94732 114468 94784
rect 114520 94772 114526 94784
rect 219434 94772 219440 94784
rect 114520 94744 219440 94772
rect 114520 94732 114526 94744
rect 219434 94732 219440 94744
rect 219492 94732 219498 94784
rect 277854 94732 277860 94784
rect 277912 94772 277918 94784
rect 453298 94772 453304 94784
rect 277912 94744 453304 94772
rect 277912 94732 277918 94744
rect 453298 94732 453304 94744
rect 453356 94732 453362 94784
rect 79318 94664 79324 94716
rect 79376 94704 79382 94716
rect 205634 94704 205640 94716
rect 79376 94676 205640 94704
rect 79376 94664 79382 94676
rect 205634 94664 205640 94676
rect 205692 94664 205698 94716
rect 209130 94704 209136 94716
rect 205744 94676 209136 94704
rect 53742 94596 53748 94648
rect 53800 94636 53806 94648
rect 205744 94636 205772 94676
rect 209130 94664 209136 94676
rect 209188 94664 209194 94716
rect 288158 94664 288164 94716
rect 288216 94704 288222 94716
rect 489178 94704 489184 94716
rect 288216 94676 489184 94704
rect 288216 94664 288222 94676
rect 489178 94664 489184 94676
rect 489236 94664 489242 94716
rect 208578 94636 208584 94648
rect 53800 94608 205772 94636
rect 205836 94608 208584 94636
rect 53800 94596 53806 94608
rect 50982 94528 50988 94580
rect 51040 94568 51046 94580
rect 205836 94568 205864 94608
rect 208578 94596 208584 94608
rect 208636 94596 208642 94648
rect 240686 94596 240692 94648
rect 240744 94636 240750 94648
rect 251266 94636 251272 94648
rect 240744 94608 251272 94636
rect 240744 94596 240750 94608
rect 251266 94596 251272 94608
rect 251324 94596 251330 94648
rect 286318 94596 286324 94648
rect 286376 94636 286382 94648
rect 502978 94636 502984 94648
rect 286376 94608 502984 94636
rect 286376 94596 286382 94608
rect 502978 94596 502984 94608
rect 503036 94596 503042 94648
rect 51040 94540 205864 94568
rect 51040 94528 51046 94540
rect 209958 94528 209964 94580
rect 210016 94568 210022 94580
rect 210326 94568 210332 94580
rect 210016 94540 210332 94568
rect 210016 94528 210022 94540
rect 210326 94528 210332 94540
rect 210384 94528 210390 94580
rect 211430 94528 211436 94580
rect 211488 94568 211494 94580
rect 211890 94568 211896 94580
rect 211488 94540 211896 94568
rect 211488 94528 211494 94540
rect 211890 94528 211896 94540
rect 211948 94528 211954 94580
rect 212902 94528 212908 94580
rect 212960 94568 212966 94580
rect 213730 94568 213736 94580
rect 212960 94540 213736 94568
rect 212960 94528 212966 94540
rect 213730 94528 213736 94540
rect 213788 94528 213794 94580
rect 228358 94528 228364 94580
rect 228416 94568 228422 94580
rect 234798 94568 234804 94580
rect 228416 94540 234804 94568
rect 228416 94528 228422 94540
rect 234798 94528 234804 94540
rect 234856 94528 234862 94580
rect 237558 94528 237564 94580
rect 237616 94568 237622 94580
rect 237926 94568 237932 94580
rect 237616 94540 237932 94568
rect 237616 94528 237622 94540
rect 237926 94528 237932 94540
rect 237984 94528 237990 94580
rect 288802 94528 288808 94580
rect 288860 94568 288866 94580
rect 518894 94568 518900 94580
rect 288860 94540 518900 94568
rect 288860 94528 288866 94540
rect 518894 94528 518900 94540
rect 518952 94528 518958 94580
rect 48222 94460 48228 94512
rect 48280 94500 48286 94512
rect 208118 94500 208124 94512
rect 48280 94472 208124 94500
rect 48280 94460 48286 94472
rect 208118 94460 208124 94472
rect 208176 94460 208182 94512
rect 226978 94460 226984 94512
rect 227036 94500 227042 94512
rect 237650 94500 237656 94512
rect 227036 94472 237656 94500
rect 227036 94460 227042 94472
rect 237650 94460 237656 94472
rect 237708 94460 237714 94512
rect 248782 94460 248788 94512
rect 248840 94500 248846 94512
rect 288434 94500 288440 94512
rect 248840 94472 288440 94500
rect 248840 94460 248846 94472
rect 288434 94460 288440 94472
rect 288492 94460 288498 94512
rect 289722 94460 289728 94512
rect 289780 94500 289786 94512
rect 520918 94500 520924 94512
rect 289780 94472 520924 94500
rect 289780 94460 289786 94472
rect 520918 94460 520924 94472
rect 520976 94460 520982 94512
rect 177942 94392 177948 94444
rect 178000 94432 178006 94444
rect 230198 94432 230204 94444
rect 178000 94404 230204 94432
rect 178000 94392 178006 94404
rect 230198 94392 230204 94404
rect 230256 94392 230262 94444
rect 254394 94392 254400 94444
rect 254452 94432 254458 94444
rect 317414 94432 317420 94444
rect 254452 94404 317420 94432
rect 254452 94392 254458 94404
rect 317414 94392 317420 94404
rect 317472 94392 317478 94444
rect 192478 94324 192484 94376
rect 192536 94364 192542 94376
rect 232590 94364 232596 94376
rect 192536 94336 232596 94364
rect 192536 94324 192542 94336
rect 232590 94324 232596 94336
rect 232648 94324 232654 94376
rect 263778 94324 263784 94376
rect 263836 94364 263842 94376
rect 306374 94364 306380 94376
rect 263836 94336 306380 94364
rect 263836 94324 263842 94336
rect 306374 94324 306380 94336
rect 306432 94324 306438 94376
rect 200022 94256 200028 94308
rect 200080 94296 200086 94308
rect 235166 94296 235172 94308
rect 200080 94268 235172 94296
rect 200080 94256 200086 94268
rect 235166 94256 235172 94268
rect 235224 94256 235230 94308
rect 263502 94256 263508 94308
rect 263560 94296 263566 94308
rect 304258 94296 304264 94308
rect 263560 94268 304264 94296
rect 263560 94256 263566 94268
rect 304258 94256 304264 94268
rect 304316 94256 304322 94308
rect 205634 94188 205640 94240
rect 205692 94228 205698 94240
rect 212994 94228 213000 94240
rect 205692 94200 213000 94228
rect 205692 94188 205698 94200
rect 212994 94188 213000 94200
rect 213052 94188 213058 94240
rect 205818 94120 205824 94172
rect 205876 94160 205882 94172
rect 206830 94160 206836 94172
rect 205876 94132 206836 94160
rect 205876 94120 205882 94132
rect 206830 94120 206836 94132
rect 206888 94120 206894 94172
rect 235902 93848 235908 93900
rect 235960 93888 235966 93900
rect 240226 93888 240232 93900
rect 235960 93860 240232 93888
rect 235960 93848 235966 93860
rect 240226 93848 240232 93860
rect 240284 93848 240290 93900
rect 181438 93780 181444 93832
rect 181496 93820 181502 93832
rect 229646 93820 229652 93832
rect 181496 93792 229652 93820
rect 181496 93780 181502 93792
rect 229646 93780 229652 93792
rect 229704 93780 229710 93832
rect 259362 93780 259368 93832
rect 259420 93820 259426 93832
rect 345014 93820 345020 93832
rect 259420 93792 345020 93820
rect 259420 93780 259426 93792
rect 345014 93780 345020 93792
rect 345072 93780 345078 93832
rect 170398 93712 170404 93764
rect 170456 93752 170462 93764
rect 227898 93752 227904 93764
rect 170456 93724 227904 93752
rect 170456 93712 170462 93724
rect 227898 93712 227904 93724
rect 227956 93712 227962 93764
rect 260742 93712 260748 93764
rect 260800 93752 260806 93764
rect 351914 93752 351920 93764
rect 260800 93724 351920 93752
rect 260800 93712 260806 93724
rect 351914 93712 351920 93724
rect 351972 93712 351978 93764
rect 166902 93644 166908 93696
rect 166960 93684 166966 93696
rect 228266 93684 228272 93696
rect 166960 93656 228272 93684
rect 166960 93644 166966 93656
rect 228266 93644 228272 93656
rect 228324 93644 228330 93696
rect 261754 93644 261760 93696
rect 261812 93684 261818 93696
rect 362954 93684 362960 93696
rect 261812 93656 362960 93684
rect 261812 93644 261818 93656
rect 362954 93644 362960 93656
rect 363012 93644 363018 93696
rect 142062 93576 142068 93628
rect 142120 93616 142126 93628
rect 224126 93616 224132 93628
rect 142120 93588 224132 93616
rect 142120 93576 142126 93588
rect 224126 93576 224132 93588
rect 224184 93576 224190 93628
rect 266262 93576 266268 93628
rect 266320 93616 266326 93628
rect 378778 93616 378784 93628
rect 266320 93588 378784 93616
rect 266320 93576 266326 93588
rect 378778 93576 378784 93588
rect 378836 93576 378842 93628
rect 135162 93508 135168 93560
rect 135220 93548 135226 93560
rect 222746 93548 222752 93560
rect 135220 93520 222752 93548
rect 135220 93508 135226 93520
rect 222746 93508 222752 93520
rect 222804 93508 222810 93560
rect 268930 93508 268936 93560
rect 268988 93548 268994 93560
rect 398834 93548 398840 93560
rect 268988 93520 398840 93548
rect 268988 93508 268994 93520
rect 398834 93508 398840 93520
rect 398892 93508 398898 93560
rect 128262 93440 128268 93492
rect 128320 93480 128326 93492
rect 221734 93480 221740 93492
rect 128320 93452 221740 93480
rect 128320 93440 128326 93452
rect 221734 93440 221740 93452
rect 221792 93440 221798 93492
rect 277302 93440 277308 93492
rect 277360 93480 277366 93492
rect 448514 93480 448520 93492
rect 277360 93452 448520 93480
rect 277360 93440 277366 93452
rect 448514 93440 448520 93452
rect 448572 93440 448578 93492
rect 65518 93372 65524 93424
rect 65576 93412 65582 93424
rect 210050 93412 210056 93424
rect 65576 93384 210056 93412
rect 65576 93372 65582 93384
rect 210050 93372 210056 93384
rect 210108 93372 210114 93424
rect 279878 93372 279884 93424
rect 279936 93412 279942 93424
rect 466454 93412 466460 93424
rect 279936 93384 466460 93412
rect 279936 93372 279942 93384
rect 466454 93372 466460 93384
rect 466512 93372 466518 93424
rect 61378 93304 61384 93356
rect 61436 93344 61442 93356
rect 209222 93344 209228 93356
rect 61436 93316 209228 93344
rect 61436 93304 61442 93316
rect 209222 93304 209228 93316
rect 209280 93304 209286 93356
rect 291930 93304 291936 93356
rect 291988 93344 291994 93356
rect 524414 93344 524420 93356
rect 291988 93316 524420 93344
rect 291988 93304 291994 93316
rect 524414 93304 524420 93316
rect 524472 93304 524478 93356
rect 33042 93236 33048 93288
rect 33100 93276 33106 93288
rect 192570 93276 192576 93288
rect 33100 93248 192576 93276
rect 33100 93236 33106 93248
rect 192570 93236 192576 93248
rect 192628 93236 192634 93288
rect 194502 93236 194508 93288
rect 194560 93276 194566 93288
rect 234062 93276 234068 93288
rect 194560 93248 234068 93276
rect 194560 93236 194566 93248
rect 234062 93236 234068 93248
rect 234120 93236 234126 93288
rect 291102 93236 291108 93288
rect 291160 93276 291166 93288
rect 525058 93276 525064 93288
rect 291160 93248 525064 93276
rect 291160 93236 291166 93248
rect 525058 93236 525064 93248
rect 525116 93236 525122 93288
rect 25498 93168 25504 93220
rect 25556 93208 25562 93220
rect 200482 93208 200488 93220
rect 25556 93180 200488 93208
rect 25556 93168 25562 93180
rect 200482 93168 200488 93180
rect 200540 93168 200546 93220
rect 296622 93168 296628 93220
rect 296680 93208 296686 93220
rect 538858 93208 538864 93220
rect 296680 93180 538864 93208
rect 296680 93168 296686 93180
rect 538858 93168 538864 93180
rect 538916 93168 538922 93220
rect 15838 93100 15844 93152
rect 15896 93140 15902 93152
rect 201494 93140 201500 93152
rect 15896 93112 201500 93140
rect 15896 93100 15902 93112
rect 201494 93100 201500 93112
rect 201552 93100 201558 93152
rect 228450 93100 228456 93152
rect 228508 93140 228514 93152
rect 237926 93140 237932 93152
rect 228508 93112 237932 93140
rect 228508 93100 228514 93112
rect 237926 93100 237932 93112
rect 237984 93100 237990 93152
rect 238662 93100 238668 93152
rect 238720 93140 238726 93152
rect 241698 93140 241704 93152
rect 238720 93112 241704 93140
rect 238720 93100 238726 93112
rect 241698 93100 241704 93112
rect 241756 93100 241762 93152
rect 245470 93100 245476 93152
rect 245528 93140 245534 93152
rect 255958 93140 255964 93152
rect 245528 93112 255964 93140
rect 245528 93100 245534 93112
rect 255958 93100 255964 93112
rect 256016 93100 256022 93152
rect 295242 93100 295248 93152
rect 295300 93140 295306 93152
rect 554774 93140 554780 93152
rect 295300 93112 554780 93140
rect 295300 93100 295306 93112
rect 554774 93100 554780 93112
rect 554832 93100 554838 93152
rect 184842 93032 184848 93084
rect 184900 93072 184906 93084
rect 231026 93072 231032 93084
rect 184900 93044 231032 93072
rect 184900 93032 184906 93044
rect 231026 93032 231032 93044
rect 231084 93032 231090 93084
rect 257982 93032 257988 93084
rect 258040 93072 258046 93084
rect 338114 93072 338120 93084
rect 258040 93044 338120 93072
rect 258040 93032 258046 93044
rect 338114 93032 338120 93044
rect 338172 93032 338178 93084
rect 188338 92964 188344 93016
rect 188396 93004 188402 93016
rect 231946 93004 231952 93016
rect 188396 92976 231952 93004
rect 188396 92964 188402 92976
rect 231946 92964 231952 92976
rect 232004 92964 232010 93016
rect 256510 92964 256516 93016
rect 256568 93004 256574 93016
rect 331214 93004 331220 93016
rect 256568 92976 331220 93004
rect 256568 92964 256574 92976
rect 331214 92964 331220 92976
rect 331272 92964 331278 93016
rect 197170 92896 197176 92948
rect 197228 92936 197234 92948
rect 233694 92936 233700 92948
rect 197228 92908 233700 92936
rect 197228 92896 197234 92908
rect 233694 92896 233700 92908
rect 233752 92896 233758 92948
rect 253842 92896 253848 92948
rect 253900 92936 253906 92948
rect 307018 92936 307024 92948
rect 253900 92908 307024 92936
rect 253900 92896 253906 92908
rect 307018 92896 307024 92908
rect 307076 92896 307082 92948
rect 234522 92488 234528 92540
rect 234580 92528 234586 92540
rect 239950 92528 239956 92540
rect 234580 92500 239956 92528
rect 234580 92488 234586 92500
rect 239950 92488 239956 92500
rect 240008 92488 240014 92540
rect 164142 92420 164148 92472
rect 164200 92460 164206 92472
rect 227990 92460 227996 92472
rect 164200 92432 227996 92460
rect 164200 92420 164206 92432
rect 227990 92420 227996 92432
rect 228048 92420 228054 92472
rect 263318 92420 263324 92472
rect 263376 92460 263382 92472
rect 369854 92460 369860 92472
rect 263376 92432 369860 92460
rect 263376 92420 263382 92432
rect 369854 92420 369860 92432
rect 369912 92420 369918 92472
rect 160002 92352 160008 92404
rect 160060 92392 160066 92404
rect 227070 92392 227076 92404
rect 160060 92364 227076 92392
rect 160060 92352 160066 92364
rect 227070 92352 227076 92364
rect 227128 92352 227134 92404
rect 264606 92352 264612 92404
rect 264664 92392 264670 92404
rect 374638 92392 374644 92404
rect 264664 92364 374644 92392
rect 264664 92352 264670 92364
rect 374638 92352 374644 92364
rect 374696 92352 374702 92404
rect 156690 92284 156696 92336
rect 156748 92324 156754 92336
rect 226886 92324 226892 92336
rect 156748 92296 226892 92324
rect 156748 92284 156754 92296
rect 226886 92284 226892 92296
rect 226944 92284 226950 92336
rect 269022 92284 269028 92336
rect 269080 92324 269086 92336
rect 381538 92324 381544 92336
rect 269080 92296 381544 92324
rect 269080 92284 269086 92296
rect 381538 92284 381544 92296
rect 381596 92284 381602 92336
rect 148962 92216 148968 92268
rect 149020 92256 149026 92268
rect 225506 92256 225512 92268
rect 149020 92228 225512 92256
rect 149020 92216 149026 92228
rect 225506 92216 225512 92228
rect 225564 92216 225570 92268
rect 252186 92216 252192 92268
rect 252244 92256 252250 92268
rect 303614 92256 303620 92268
rect 252244 92228 303620 92256
rect 252244 92216 252250 92228
rect 303614 92216 303620 92228
rect 303672 92216 303678 92268
rect 304350 92216 304356 92268
rect 304408 92256 304414 92268
rect 418154 92256 418160 92268
rect 304408 92228 418160 92256
rect 304408 92216 304414 92228
rect 418154 92216 418160 92228
rect 418212 92216 418218 92268
rect 144822 92148 144828 92200
rect 144880 92188 144886 92200
rect 224586 92188 224592 92200
rect 144880 92160 224592 92188
rect 144880 92148 144886 92160
rect 224586 92148 224592 92160
rect 224644 92148 224650 92200
rect 265986 92148 265992 92200
rect 266044 92188 266050 92200
rect 382918 92188 382924 92200
rect 266044 92160 382924 92188
rect 266044 92148 266050 92160
rect 382918 92148 382924 92160
rect 382976 92148 382982 92200
rect 142798 92080 142804 92132
rect 142856 92120 142862 92132
rect 222378 92120 222384 92132
rect 142856 92092 222384 92120
rect 142856 92080 142862 92092
rect 222378 92080 222384 92092
rect 222436 92080 222442 92132
rect 267366 92080 267372 92132
rect 267424 92120 267430 92132
rect 387794 92120 387800 92132
rect 267424 92092 387800 92120
rect 267424 92080 267430 92092
rect 387794 92080 387800 92092
rect 387852 92080 387858 92132
rect 98638 92012 98644 92064
rect 98696 92052 98702 92064
rect 216674 92052 216680 92064
rect 98696 92024 216680 92052
rect 98696 92012 98702 92024
rect 216674 92012 216680 92024
rect 216732 92012 216738 92064
rect 267642 92012 267648 92064
rect 267700 92052 267706 92064
rect 389818 92052 389824 92064
rect 267700 92024 389824 92052
rect 267700 92012 267706 92024
rect 389818 92012 389824 92024
rect 389876 92012 389882 92064
rect 71038 91944 71044 91996
rect 71096 91984 71102 91996
rect 210602 91984 210608 91996
rect 71096 91956 210608 91984
rect 71096 91944 71102 91956
rect 210602 91944 210608 91956
rect 210660 91944 210666 91996
rect 269942 91944 269948 91996
rect 270000 91984 270006 91996
rect 405734 91984 405740 91996
rect 270000 91956 405740 91984
rect 270000 91944 270006 91956
rect 405734 91944 405740 91956
rect 405792 91944 405798 91996
rect 70302 91876 70308 91928
rect 70360 91916 70366 91928
rect 211798 91916 211804 91928
rect 70360 91888 211804 91916
rect 70360 91876 70366 91888
rect 211798 91876 211804 91888
rect 211856 91876 211862 91928
rect 272886 91876 272892 91928
rect 272944 91916 272950 91928
rect 421558 91916 421564 91928
rect 272944 91888 421564 91916
rect 272944 91876 272950 91888
rect 421558 91876 421564 91888
rect 421616 91876 421622 91928
rect 46842 91808 46848 91860
rect 46900 91848 46906 91860
rect 203518 91848 203524 91860
rect 46900 91820 203524 91848
rect 46900 91808 46906 91820
rect 203518 91808 203524 91820
rect 203576 91808 203582 91860
rect 243998 91808 244004 91860
rect 244056 91848 244062 91860
rect 263686 91848 263692 91860
rect 244056 91820 263692 91848
rect 244056 91808 244062 91820
rect 263686 91808 263692 91820
rect 263744 91808 263750 91860
rect 281074 91808 281080 91860
rect 281132 91848 281138 91860
rect 471238 91848 471244 91860
rect 281132 91820 471244 91848
rect 281132 91808 281138 91820
rect 471238 91808 471244 91820
rect 471296 91808 471302 91860
rect 34422 91740 34428 91792
rect 34480 91780 34486 91792
rect 205726 91780 205732 91792
rect 34480 91752 205732 91780
rect 34480 91740 34486 91752
rect 205726 91740 205732 91752
rect 205784 91740 205790 91792
rect 222838 91740 222844 91792
rect 222896 91780 222902 91792
rect 235718 91780 235724 91792
rect 222896 91752 235724 91780
rect 222896 91740 222902 91752
rect 235718 91740 235724 91752
rect 235776 91740 235782 91792
rect 245562 91740 245568 91792
rect 245620 91780 245626 91792
rect 266446 91780 266452 91792
rect 245620 91752 266452 91780
rect 245620 91740 245626 91752
rect 266446 91740 266452 91752
rect 266504 91740 266510 91792
rect 290918 91740 290924 91792
rect 290976 91780 290982 91792
rect 529198 91780 529204 91792
rect 290976 91752 529204 91780
rect 290976 91740 290982 91752
rect 529198 91740 529204 91752
rect 529256 91740 529262 91792
rect 171042 91672 171048 91724
rect 171100 91712 171106 91724
rect 229186 91712 229192 91724
rect 171100 91684 229192 91712
rect 171100 91672 171106 91684
rect 229186 91672 229192 91684
rect 229244 91672 229250 91724
rect 257706 91672 257712 91724
rect 257764 91712 257770 91724
rect 330478 91712 330484 91724
rect 257764 91684 330484 91712
rect 257764 91672 257770 91684
rect 330478 91672 330484 91684
rect 330536 91672 330542 91724
rect 182082 91604 182088 91656
rect 182140 91644 182146 91656
rect 230934 91644 230940 91656
rect 182140 91616 230940 91644
rect 182140 91604 182146 91616
rect 230934 91604 230940 91616
rect 230992 91604 230998 91656
rect 231302 91060 231308 91112
rect 231360 91100 231366 91112
rect 236178 91100 236184 91112
rect 231360 91072 236184 91100
rect 231360 91060 231366 91072
rect 236178 91060 236184 91072
rect 236236 91060 236242 91112
rect 187050 90992 187056 91044
rect 187108 91032 187114 91044
rect 230842 91032 230848 91044
rect 187108 91004 230848 91032
rect 187108 90992 187114 91004
rect 230842 90992 230848 91004
rect 230900 90992 230906 91044
rect 267458 90992 267464 91044
rect 267516 91032 267522 91044
rect 394694 91032 394700 91044
rect 267516 91004 394700 91032
rect 267516 90992 267522 91004
rect 394694 90992 394700 91004
rect 394752 90992 394758 91044
rect 169018 90924 169024 90976
rect 169076 90964 169082 90976
rect 228082 90964 228088 90976
rect 169076 90936 228088 90964
rect 169076 90924 169082 90936
rect 228082 90924 228088 90936
rect 228140 90924 228146 90976
rect 268746 90924 268752 90976
rect 268804 90964 268810 90976
rect 396718 90964 396724 90976
rect 268804 90936 396724 90964
rect 268804 90924 268810 90936
rect 396718 90924 396724 90936
rect 396776 90924 396782 90976
rect 139302 90856 139308 90908
rect 139360 90896 139366 90908
rect 223758 90896 223764 90908
rect 139360 90868 223764 90896
rect 139360 90856 139366 90868
rect 223758 90856 223764 90868
rect 223816 90856 223822 90908
rect 270218 90856 270224 90908
rect 270276 90896 270282 90908
rect 407758 90896 407764 90908
rect 270276 90868 407764 90896
rect 270276 90856 270282 90868
rect 407758 90856 407764 90868
rect 407816 90856 407822 90908
rect 137370 90788 137376 90840
rect 137428 90828 137434 90840
rect 222562 90828 222568 90840
rect 137428 90800 222568 90828
rect 137428 90788 137434 90800
rect 222562 90788 222568 90800
rect 222620 90788 222626 90840
rect 271598 90788 271604 90840
rect 271656 90828 271662 90840
rect 417418 90828 417424 90840
rect 271656 90800 417424 90828
rect 271656 90788 271662 90800
rect 417418 90788 417424 90800
rect 417476 90788 417482 90840
rect 116578 90720 116584 90772
rect 116636 90760 116642 90772
rect 219710 90760 219716 90772
rect 116636 90732 219716 90760
rect 116636 90720 116642 90732
rect 219710 90720 219716 90732
rect 219768 90720 219774 90772
rect 274266 90720 274272 90772
rect 274324 90760 274330 90772
rect 432598 90760 432604 90772
rect 274324 90732 432604 90760
rect 274324 90720 274330 90732
rect 432598 90720 432604 90732
rect 432656 90720 432662 90772
rect 95142 90652 95148 90704
rect 95200 90692 95206 90704
rect 215754 90692 215760 90704
rect 95200 90664 215760 90692
rect 95200 90652 95206 90664
rect 215754 90652 215760 90664
rect 215812 90652 215818 90704
rect 277118 90652 277124 90704
rect 277176 90692 277182 90704
rect 446398 90692 446404 90704
rect 277176 90664 446404 90692
rect 277176 90652 277182 90664
rect 446398 90652 446404 90664
rect 446456 90652 446462 90704
rect 86862 90584 86868 90636
rect 86920 90624 86926 90636
rect 214742 90624 214748 90636
rect 86920 90596 214748 90624
rect 86920 90584 86926 90596
rect 214742 90584 214748 90596
rect 214800 90584 214806 90636
rect 281442 90584 281448 90636
rect 281500 90624 281506 90636
rect 467098 90624 467104 90636
rect 281500 90596 467104 90624
rect 281500 90584 281506 90596
rect 467098 90584 467104 90596
rect 467156 90584 467162 90636
rect 80698 90516 80704 90568
rect 80756 90556 80762 90568
rect 213454 90556 213460 90568
rect 80756 90528 213460 90556
rect 80756 90516 80762 90528
rect 213454 90516 213460 90528
rect 213512 90516 213518 90568
rect 283926 90516 283932 90568
rect 283984 90556 283990 90568
rect 486418 90556 486424 90568
rect 283984 90528 486424 90556
rect 283984 90516 283990 90528
rect 486418 90516 486424 90528
rect 486476 90516 486482 90568
rect 76558 90448 76564 90500
rect 76616 90488 76622 90500
rect 212258 90488 212264 90500
rect 76616 90460 212264 90488
rect 76616 90448 76622 90460
rect 212258 90448 212264 90460
rect 212316 90448 212322 90500
rect 253290 90448 253296 90500
rect 253348 90488 253354 90500
rect 266354 90488 266360 90500
rect 253348 90460 266360 90488
rect 253348 90448 253354 90460
rect 266354 90448 266360 90460
rect 266412 90448 266418 90500
rect 288342 90448 288348 90500
rect 288400 90488 288406 90500
rect 504358 90488 504364 90500
rect 288400 90460 504364 90488
rect 288400 90448 288406 90460
rect 504358 90448 504364 90460
rect 504416 90448 504422 90500
rect 57882 90380 57888 90432
rect 57940 90420 57946 90432
rect 209682 90420 209688 90432
rect 57940 90392 209688 90420
rect 57940 90380 57946 90392
rect 209682 90380 209688 90392
rect 209740 90380 209746 90432
rect 246206 90380 246212 90432
rect 246264 90420 246270 90432
rect 268378 90420 268384 90432
rect 246264 90392 268384 90420
rect 246264 90380 246270 90392
rect 268378 90380 268384 90392
rect 268436 90380 268442 90432
rect 293402 90380 293408 90432
rect 293460 90420 293466 90432
rect 540238 90420 540244 90432
rect 293460 90392 540244 90420
rect 293460 90380 293466 90392
rect 540238 90380 540244 90392
rect 540296 90380 540302 90432
rect 45462 90312 45468 90364
rect 45520 90352 45526 90364
rect 207474 90352 207480 90364
rect 45520 90324 207480 90352
rect 45520 90312 45526 90324
rect 207474 90312 207480 90324
rect 207532 90312 207538 90364
rect 248138 90312 248144 90364
rect 248196 90352 248202 90364
rect 280246 90352 280252 90364
rect 248196 90324 280252 90352
rect 248196 90312 248202 90324
rect 280246 90312 280252 90324
rect 280304 90312 280310 90364
rect 297174 90312 297180 90364
rect 297232 90352 297238 90364
rect 566458 90352 566464 90364
rect 297232 90324 566464 90352
rect 297232 90312 297238 90324
rect 566458 90312 566464 90324
rect 566516 90312 566522 90364
rect 193122 90244 193128 90296
rect 193180 90284 193186 90296
rect 232130 90284 232136 90296
rect 193180 90256 232136 90284
rect 193180 90244 193186 90256
rect 232130 90244 232136 90256
rect 232188 90244 232194 90296
rect 255130 90244 255136 90296
rect 255188 90284 255194 90296
rect 321554 90284 321560 90296
rect 255188 90256 321560 90284
rect 255188 90244 255194 90256
rect 321554 90244 321560 90256
rect 321612 90244 321618 90296
rect 253566 90176 253572 90228
rect 253624 90216 253630 90228
rect 309226 90216 309232 90228
rect 253624 90188 309232 90216
rect 253624 90176 253630 90188
rect 309226 90176 309232 90188
rect 309284 90176 309290 90228
rect 250806 89972 250812 90024
rect 250864 90012 250870 90024
rect 253198 90012 253204 90024
rect 250864 89984 253204 90012
rect 250864 89972 250870 89984
rect 253198 89972 253204 89984
rect 253256 89972 253262 90024
rect 256234 89632 256240 89684
rect 256292 89672 256298 89684
rect 328454 89672 328460 89684
rect 256292 89644 328460 89672
rect 256292 89632 256298 89644
rect 328454 89632 328460 89644
rect 328512 89632 328518 89684
rect 266078 89564 266084 89616
rect 266136 89604 266142 89616
rect 377398 89604 377404 89616
rect 266136 89576 377404 89604
rect 266136 89564 266142 89576
rect 377398 89564 377404 89576
rect 377456 89564 377462 89616
rect 275738 89496 275744 89548
rect 275796 89536 275802 89548
rect 438854 89536 438860 89548
rect 275796 89508 438860 89536
rect 275796 89496 275802 89508
rect 438854 89496 438860 89508
rect 438912 89496 438918 89548
rect 122742 89428 122748 89480
rect 122800 89468 122806 89480
rect 220998 89468 221004 89480
rect 122800 89440 221004 89468
rect 122800 89428 122806 89440
rect 220998 89428 221004 89440
rect 221056 89428 221062 89480
rect 281166 89428 281172 89480
rect 281224 89468 281230 89480
rect 476114 89468 476120 89480
rect 281224 89440 476120 89468
rect 281224 89428 281230 89440
rect 476114 89428 476120 89440
rect 476172 89428 476178 89480
rect 119982 89360 119988 89412
rect 120040 89400 120046 89412
rect 219618 89400 219624 89412
rect 120040 89372 219624 89400
rect 120040 89360 120046 89372
rect 219618 89360 219624 89372
rect 219676 89360 219682 89412
rect 282638 89360 282644 89412
rect 282696 89400 282702 89412
rect 481634 89400 481640 89412
rect 282696 89372 481640 89400
rect 282696 89360 282702 89372
rect 481634 89360 481640 89372
rect 481692 89360 481698 89412
rect 115198 89292 115204 89344
rect 115256 89332 115262 89344
rect 218974 89332 218980 89344
rect 115256 89304 218980 89332
rect 115256 89292 115262 89304
rect 218974 89292 218980 89304
rect 219032 89292 219038 89344
rect 284018 89292 284024 89344
rect 284076 89332 284082 89344
rect 490558 89332 490564 89344
rect 284076 89304 490564 89332
rect 284076 89292 284082 89304
rect 490558 89292 490564 89304
rect 490616 89292 490622 89344
rect 104802 89224 104808 89276
rect 104860 89264 104866 89276
rect 217778 89264 217784 89276
rect 104860 89236 217784 89264
rect 104860 89224 104866 89236
rect 217778 89224 217784 89236
rect 217836 89224 217842 89276
rect 285306 89224 285312 89276
rect 285364 89264 285370 89276
rect 493318 89264 493324 89276
rect 285364 89236 493324 89264
rect 285364 89224 285370 89236
rect 493318 89224 493324 89236
rect 493376 89224 493382 89276
rect 102042 89156 102048 89208
rect 102100 89196 102106 89208
rect 216950 89196 216956 89208
rect 102100 89168 216956 89196
rect 102100 89156 102106 89168
rect 216950 89156 216956 89168
rect 217008 89156 217014 89208
rect 285214 89156 285220 89208
rect 285272 89196 285278 89208
rect 497458 89196 497464 89208
rect 285272 89168 497464 89196
rect 285272 89156 285278 89168
rect 497458 89156 497464 89168
rect 497516 89156 497522 89208
rect 37090 89088 37096 89140
rect 37148 89128 37154 89140
rect 206186 89128 206192 89140
rect 37148 89100 206192 89128
rect 37148 89088 37154 89100
rect 206186 89088 206192 89100
rect 206244 89088 206250 89140
rect 286686 89088 286692 89140
rect 286744 89128 286750 89140
rect 500218 89128 500224 89140
rect 286744 89100 500224 89128
rect 286744 89088 286750 89100
rect 500218 89088 500224 89100
rect 500276 89088 500282 89140
rect 27522 89020 27528 89072
rect 27580 89060 27586 89072
rect 204530 89060 204536 89072
rect 27580 89032 204536 89060
rect 27580 89020 27586 89032
rect 204530 89020 204536 89032
rect 204588 89020 204594 89072
rect 242434 89020 242440 89072
rect 242492 89060 242498 89072
rect 252646 89060 252652 89072
rect 242492 89032 252652 89060
rect 242492 89020 242498 89032
rect 252646 89020 252652 89032
rect 252704 89020 252710 89072
rect 289446 89020 289452 89072
rect 289504 89060 289510 89072
rect 522298 89060 522304 89072
rect 289504 89032 522304 89060
rect 289504 89020 289510 89032
rect 522298 89020 522304 89032
rect 522356 89020 522362 89072
rect 18598 88952 18604 89004
rect 18656 88992 18662 89004
rect 201586 88992 201592 89004
rect 18656 88964 201592 88992
rect 18656 88952 18662 88964
rect 201586 88952 201592 88964
rect 201644 88952 201650 89004
rect 249334 88952 249340 89004
rect 249392 88992 249398 89004
rect 285674 88992 285680 89004
rect 249392 88964 285680 88992
rect 249392 88952 249398 88964
rect 285674 88952 285680 88964
rect 285732 88952 285738 89004
rect 294874 88952 294880 89004
rect 294932 88992 294938 89004
rect 553394 88992 553400 89004
rect 294932 88964 553400 88992
rect 294932 88952 294938 88964
rect 553394 88952 553400 88964
rect 553452 88952 553458 89004
rect 253658 88884 253664 88936
rect 253716 88924 253722 88936
rect 310514 88924 310520 88936
rect 253716 88896 310520 88924
rect 253716 88884 253722 88896
rect 310514 88884 310520 88896
rect 310572 88884 310578 88936
rect 257798 88272 257804 88324
rect 257856 88312 257862 88324
rect 335354 88312 335360 88324
rect 257856 88284 335360 88312
rect 257856 88272 257862 88284
rect 335354 88272 335360 88284
rect 335412 88272 335418 88324
rect 260374 88204 260380 88256
rect 260432 88244 260438 88256
rect 353294 88244 353300 88256
rect 260432 88216 353300 88244
rect 260432 88204 260438 88216
rect 353294 88204 353300 88216
rect 353352 88204 353358 88256
rect 292206 88136 292212 88188
rect 292264 88176 292270 88188
rect 428458 88176 428464 88188
rect 292264 88148 428464 88176
rect 292264 88136 292270 88148
rect 428458 88136 428464 88148
rect 428516 88136 428522 88188
rect 105538 88068 105544 88120
rect 105596 88108 105602 88120
rect 215478 88108 215484 88120
rect 105596 88080 215484 88108
rect 105596 88068 105602 88080
rect 215478 88068 215484 88080
rect 215536 88068 215542 88120
rect 272978 88068 272984 88120
rect 273036 88108 273042 88120
rect 420914 88108 420920 88120
rect 273036 88080 420920 88108
rect 273036 88068 273042 88080
rect 420914 88068 420920 88080
rect 420972 88068 420978 88120
rect 88978 88000 88984 88052
rect 89036 88040 89042 88052
rect 208854 88040 208860 88052
rect 89036 88012 208860 88040
rect 89036 88000 89042 88012
rect 208854 88000 208860 88012
rect 208912 88000 208918 88052
rect 286778 88000 286784 88052
rect 286836 88040 286842 88052
rect 506474 88040 506480 88052
rect 286836 88012 506480 88040
rect 286836 88000 286842 88012
rect 506474 88000 506480 88012
rect 506532 88000 506538 88052
rect 71682 87932 71688 87984
rect 71740 87972 71746 87984
rect 199378 87972 199384 87984
rect 71740 87944 199384 87972
rect 71740 87932 71746 87944
rect 199378 87932 199384 87944
rect 199436 87932 199442 87984
rect 288066 87932 288072 87984
rect 288124 87972 288130 87984
rect 511258 87972 511264 87984
rect 288124 87944 511264 87972
rect 288124 87932 288130 87944
rect 511258 87932 511264 87944
rect 511316 87932 511322 87984
rect 75178 87864 75184 87916
rect 75236 87904 75242 87916
rect 212718 87904 212724 87916
rect 75236 87876 212724 87904
rect 75236 87864 75242 87876
rect 212718 87864 212724 87876
rect 212776 87864 212782 87916
rect 300302 87864 300308 87916
rect 300360 87904 300366 87916
rect 525794 87904 525800 87916
rect 300360 87876 525800 87904
rect 300360 87864 300366 87876
rect 525794 87864 525800 87876
rect 525852 87864 525858 87916
rect 61470 87796 61476 87848
rect 61528 87836 61534 87848
rect 210142 87836 210148 87848
rect 61528 87808 210148 87836
rect 61528 87796 61534 87808
rect 210142 87796 210148 87808
rect 210200 87796 210206 87848
rect 288250 87796 288256 87848
rect 288308 87836 288314 87848
rect 515398 87836 515404 87848
rect 288308 87808 515404 87836
rect 288308 87796 288314 87808
rect 515398 87796 515404 87808
rect 515456 87796 515462 87848
rect 41322 87728 41328 87780
rect 41380 87768 41386 87780
rect 205818 87768 205824 87780
rect 41380 87740 205824 87768
rect 41380 87728 41386 87740
rect 205818 87728 205824 87740
rect 205876 87728 205882 87780
rect 289538 87728 289544 87780
rect 289596 87768 289602 87780
rect 518158 87768 518164 87780
rect 289596 87740 518164 87768
rect 289596 87728 289602 87740
rect 518158 87728 518164 87740
rect 518216 87728 518222 87780
rect 28902 87660 28908 87712
rect 28960 87700 28966 87712
rect 196618 87700 196624 87712
rect 28960 87672 196624 87700
rect 28960 87660 28966 87672
rect 196618 87660 196624 87672
rect 196676 87660 196682 87712
rect 293586 87660 293592 87712
rect 293644 87700 293650 87712
rect 542998 87700 543004 87712
rect 293644 87672 543004 87700
rect 293644 87660 293650 87672
rect 542998 87660 543004 87672
rect 543056 87660 543062 87712
rect 30282 87592 30288 87644
rect 30340 87632 30346 87644
rect 204438 87632 204444 87644
rect 30340 87604 204444 87632
rect 30340 87592 30346 87604
rect 204438 87592 204444 87604
rect 204496 87592 204502 87644
rect 209038 87592 209044 87644
rect 209096 87632 209102 87644
rect 233510 87632 233516 87644
rect 209096 87604 233516 87632
rect 209096 87592 209102 87604
rect 233510 87592 233516 87604
rect 233568 87592 233574 87644
rect 248230 87592 248236 87644
rect 248288 87632 248294 87644
rect 287054 87632 287060 87644
rect 248288 87604 287060 87632
rect 248288 87592 248294 87604
rect 287054 87592 287060 87604
rect 287112 87592 287118 87644
rect 297910 87592 297916 87644
rect 297968 87632 297974 87644
rect 569954 87632 569960 87644
rect 297968 87604 569960 87632
rect 297968 87592 297974 87604
rect 569954 87592 569960 87604
rect 570012 87592 570018 87644
rect 254946 87524 254952 87576
rect 255004 87564 255010 87576
rect 316126 87564 316132 87576
rect 255004 87536 316132 87564
rect 255004 87524 255010 87536
rect 316126 87524 316132 87536
rect 316184 87524 316190 87576
rect 253750 87456 253756 87508
rect 253808 87496 253814 87508
rect 314010 87496 314016 87508
rect 253808 87468 314016 87496
rect 253808 87456 253814 87468
rect 314010 87456 314016 87468
rect 314068 87456 314074 87508
rect 259086 86912 259092 86964
rect 259144 86952 259150 86964
rect 342254 86952 342260 86964
rect 259144 86924 342260 86952
rect 259144 86912 259150 86924
rect 342254 86912 342260 86924
rect 342312 86912 342318 86964
rect 342898 86912 342904 86964
rect 342956 86952 342962 86964
rect 425054 86952 425060 86964
rect 342956 86924 425060 86952
rect 342956 86912 342962 86924
rect 425054 86912 425060 86924
rect 425112 86912 425118 86964
rect 259178 86844 259184 86896
rect 259236 86884 259242 86896
rect 346394 86884 346400 86896
rect 259236 86856 346400 86884
rect 259236 86844 259242 86856
rect 346394 86844 346400 86856
rect 346452 86844 346458 86896
rect 271230 86776 271236 86828
rect 271288 86816 271294 86828
rect 365806 86816 365812 86828
rect 271288 86788 365812 86816
rect 271288 86776 271294 86788
rect 365806 86776 365812 86788
rect 365864 86776 365870 86828
rect 261938 86708 261944 86760
rect 261996 86748 262002 86760
rect 357434 86748 357440 86760
rect 261996 86720 357440 86748
rect 261996 86708 262002 86720
rect 357434 86708 357440 86720
rect 357492 86708 357498 86760
rect 267550 86640 267556 86692
rect 267608 86680 267614 86692
rect 392026 86680 392032 86692
rect 267608 86652 392032 86680
rect 267608 86640 267614 86652
rect 392026 86640 392032 86652
rect 392084 86640 392090 86692
rect 123478 86572 123484 86624
rect 123536 86612 123542 86624
rect 219894 86612 219900 86624
rect 123536 86584 219900 86612
rect 123536 86572 123542 86584
rect 219894 86572 219900 86584
rect 219952 86572 219958 86624
rect 275830 86572 275836 86624
rect 275888 86612 275894 86624
rect 441614 86612 441620 86624
rect 275888 86584 441620 86612
rect 275888 86572 275894 86584
rect 441614 86572 441620 86584
rect 441672 86572 441678 86624
rect 106918 86504 106924 86556
rect 106976 86544 106982 86556
rect 210050 86544 210056 86556
rect 106976 86516 210056 86544
rect 106976 86504 106982 86516
rect 210050 86504 210056 86516
rect 210108 86504 210114 86556
rect 292298 86504 292304 86556
rect 292356 86544 292362 86556
rect 536098 86544 536104 86556
rect 292356 86516 536104 86544
rect 292356 86504 292362 86516
rect 536098 86504 536104 86516
rect 536156 86504 536162 86556
rect 111150 86436 111156 86488
rect 111208 86476 111214 86488
rect 218514 86476 218520 86488
rect 111208 86448 218520 86476
rect 111208 86436 111214 86448
rect 218514 86436 218520 86448
rect 218572 86436 218578 86488
rect 293678 86436 293684 86488
rect 293736 86476 293742 86488
rect 547138 86476 547144 86488
rect 293736 86448 547144 86476
rect 293736 86436 293742 86448
rect 547138 86436 547144 86448
rect 547196 86436 547202 86488
rect 86218 86368 86224 86420
rect 86276 86408 86282 86420
rect 214098 86408 214104 86420
rect 86276 86380 214104 86408
rect 86276 86368 86282 86380
rect 214098 86368 214104 86380
rect 214156 86368 214162 86420
rect 244090 86368 244096 86420
rect 244148 86408 244154 86420
rect 258074 86408 258080 86420
rect 244148 86380 258080 86408
rect 244148 86368 244154 86380
rect 258074 86368 258080 86380
rect 258132 86368 258138 86420
rect 294966 86368 294972 86420
rect 295024 86408 295030 86420
rect 556154 86408 556160 86420
rect 295024 86380 556160 86408
rect 295024 86368 295030 86380
rect 556154 86368 556160 86380
rect 556212 86368 556218 86420
rect 79410 86300 79416 86352
rect 79468 86340 79474 86352
rect 213086 86340 213092 86352
rect 79468 86312 213092 86340
rect 79468 86300 79474 86312
rect 213086 86300 213092 86312
rect 213144 86300 213150 86352
rect 249426 86300 249432 86352
rect 249484 86340 249490 86352
rect 291286 86340 291292 86352
rect 249484 86312 291292 86340
rect 249484 86300 249490 86312
rect 291286 86300 291292 86312
rect 291344 86300 291350 86352
rect 296346 86300 296352 86352
rect 296404 86340 296410 86352
rect 560386 86340 560392 86352
rect 296404 86312 560392 86340
rect 296404 86300 296410 86312
rect 560386 86300 560392 86312
rect 560444 86300 560450 86352
rect 68278 86232 68284 86284
rect 68336 86272 68342 86284
rect 211706 86272 211712 86284
rect 68336 86244 211712 86272
rect 68336 86232 68342 86244
rect 211706 86232 211712 86244
rect 211764 86232 211770 86284
rect 250898 86232 250904 86284
rect 250956 86272 250962 86284
rect 295334 86272 295340 86284
rect 250956 86244 295340 86272
rect 250956 86232 250962 86244
rect 295334 86232 295340 86244
rect 295392 86232 295398 86284
rect 299106 86232 299112 86284
rect 299164 86272 299170 86284
rect 582742 86272 582748 86284
rect 299164 86244 582748 86272
rect 299164 86232 299170 86244
rect 582742 86232 582748 86244
rect 582800 86232 582806 86284
rect 3142 85484 3148 85536
rect 3200 85524 3206 85536
rect 152458 85524 152464 85536
rect 3200 85496 152464 85524
rect 3200 85484 3206 85496
rect 152458 85484 152464 85496
rect 152516 85484 152522 85536
rect 262030 85416 262036 85468
rect 262088 85456 262094 85468
rect 360194 85456 360200 85468
rect 262088 85428 360200 85456
rect 262088 85416 262094 85428
rect 360194 85416 360200 85428
rect 360252 85416 360258 85468
rect 263134 85348 263140 85400
rect 263192 85388 263198 85400
rect 364334 85388 364340 85400
rect 263192 85360 364340 85388
rect 263192 85348 263198 85360
rect 364334 85348 364340 85360
rect 364392 85348 364398 85400
rect 263226 85280 263232 85332
rect 263284 85320 263290 85332
rect 367094 85320 367100 85332
rect 263284 85292 367100 85320
rect 263284 85280 263290 85292
rect 367094 85280 367100 85292
rect 367152 85280 367158 85332
rect 266170 85212 266176 85264
rect 266228 85252 266234 85264
rect 382366 85252 382372 85264
rect 266228 85224 382372 85252
rect 266228 85212 266234 85224
rect 382366 85212 382372 85224
rect 382424 85212 382430 85264
rect 268838 85144 268844 85196
rect 268896 85184 268902 85196
rect 402974 85184 402980 85196
rect 268896 85156 402980 85184
rect 268896 85144 268902 85156
rect 402974 85144 402980 85156
rect 403032 85144 403038 85196
rect 153102 85076 153108 85128
rect 153160 85116 153166 85128
rect 225414 85116 225420 85128
rect 153160 85088 225420 85116
rect 153160 85076 153166 85088
rect 225414 85076 225420 85088
rect 225472 85076 225478 85128
rect 278406 85076 278412 85128
rect 278464 85116 278470 85128
rect 452654 85116 452660 85128
rect 278464 85088 452660 85116
rect 278464 85076 278470 85088
rect 452654 85076 452660 85088
rect 452712 85076 452718 85128
rect 124122 85008 124128 85060
rect 124180 85048 124186 85060
rect 221090 85048 221096 85060
rect 124180 85020 221096 85048
rect 124180 85008 124186 85020
rect 221090 85008 221096 85020
rect 221148 85008 221154 85060
rect 291010 85008 291016 85060
rect 291068 85048 291074 85060
rect 528554 85048 528560 85060
rect 291068 85020 528560 85048
rect 291068 85008 291074 85020
rect 528554 85008 528560 85020
rect 528612 85008 528618 85060
rect 95050 84940 95056 84992
rect 95108 84980 95114 84992
rect 216122 84980 216128 84992
rect 95108 84952 216128 84980
rect 95108 84940 95114 84952
rect 216122 84940 216128 84952
rect 216180 84940 216186 84992
rect 300118 84940 300124 84992
rect 300176 84980 300182 84992
rect 565814 84980 565820 84992
rect 300176 84952 565820 84980
rect 300176 84940 300182 84952
rect 565814 84940 565820 84952
rect 565872 84940 565878 84992
rect 88242 84872 88248 84924
rect 88300 84912 88306 84924
rect 214926 84912 214932 84924
rect 88300 84884 214932 84912
rect 88300 84872 88306 84884
rect 214926 84872 214932 84884
rect 214984 84872 214990 84924
rect 245286 84872 245292 84924
rect 245344 84912 245350 84924
rect 262214 84912 262220 84924
rect 245344 84884 262220 84912
rect 245344 84872 245350 84884
rect 262214 84872 262220 84884
rect 262272 84872 262278 84924
rect 296438 84872 296444 84924
rect 296496 84912 296502 84924
rect 564526 84912 564532 84924
rect 296496 84884 564532 84912
rect 296496 84872 296502 84884
rect 564526 84872 564532 84884
rect 564584 84872 564590 84924
rect 10962 84804 10968 84856
rect 11020 84844 11026 84856
rect 201770 84844 201776 84856
rect 11020 84816 201776 84844
rect 11020 84804 11026 84816
rect 201770 84804 201776 84816
rect 201828 84804 201834 84856
rect 252278 84804 252284 84856
rect 252336 84844 252342 84856
rect 299474 84844 299480 84856
rect 252336 84816 299480 84844
rect 252336 84804 252342 84816
rect 299474 84804 299480 84816
rect 299532 84804 299538 84856
rect 301498 84804 301504 84856
rect 301556 84844 301562 84856
rect 572806 84844 572812 84856
rect 301556 84816 572812 84844
rect 301556 84804 301562 84816
rect 572806 84804 572812 84816
rect 572864 84804 572870 84856
rect 260466 83988 260472 84040
rect 260524 84028 260530 84040
rect 327718 84028 327724 84040
rect 260524 84000 327724 84028
rect 260524 83988 260530 84000
rect 327718 83988 327724 84000
rect 327776 83988 327782 84040
rect 264698 83920 264704 83972
rect 264756 83960 264762 83972
rect 374086 83960 374092 83972
rect 264756 83932 374092 83960
rect 264756 83920 264762 83932
rect 374086 83920 374092 83932
rect 374144 83920 374150 83972
rect 264790 83852 264796 83904
rect 264848 83892 264854 83904
rect 378134 83892 378140 83904
rect 264848 83864 378140 83892
rect 264848 83852 264854 83864
rect 378134 83852 378140 83864
rect 378192 83852 378198 83904
rect 265894 83784 265900 83836
rect 265952 83824 265958 83836
rect 385034 83824 385040 83836
rect 265952 83796 385040 83824
rect 265952 83784 265958 83796
rect 385034 83784 385040 83796
rect 385092 83784 385098 83836
rect 267274 83716 267280 83768
rect 267332 83756 267338 83768
rect 391934 83756 391940 83768
rect 267332 83728 391940 83756
rect 267332 83716 267338 83728
rect 391934 83716 391940 83728
rect 391992 83716 391998 83768
rect 268562 83648 268568 83700
rect 268620 83688 268626 83700
rect 396074 83688 396080 83700
rect 268620 83660 396080 83688
rect 268620 83648 268626 83660
rect 396074 83648 396080 83660
rect 396132 83648 396138 83700
rect 270310 83580 270316 83632
rect 270368 83620 270374 83632
rect 409966 83620 409972 83632
rect 270368 83592 409972 83620
rect 270368 83580 270374 83592
rect 409966 83580 409972 83592
rect 410024 83580 410030 83632
rect 45370 83512 45376 83564
rect 45428 83552 45434 83564
rect 207474 83552 207480 83564
rect 45428 83524 207480 83552
rect 45428 83512 45434 83524
rect 207474 83512 207480 83524
rect 207532 83512 207538 83564
rect 274358 83512 274364 83564
rect 274416 83552 274422 83564
rect 432046 83552 432052 83564
rect 274416 83524 432052 83552
rect 274416 83512 274422 83524
rect 432046 83512 432052 83524
rect 432104 83512 432110 83564
rect 35158 83444 35164 83496
rect 35216 83484 35222 83496
rect 204714 83484 204720 83496
rect 35216 83456 204720 83484
rect 35216 83444 35222 83456
rect 204714 83444 204720 83456
rect 204772 83444 204778 83496
rect 246574 83444 246580 83496
rect 246632 83484 246638 83496
rect 260098 83484 260104 83496
rect 246632 83456 260104 83484
rect 246632 83444 246638 83456
rect 260098 83444 260104 83456
rect 260156 83444 260162 83496
rect 281258 83444 281264 83496
rect 281316 83484 281322 83496
rect 470594 83484 470600 83496
rect 281316 83456 470600 83484
rect 281316 83444 281322 83456
rect 470594 83444 470600 83456
rect 470652 83444 470658 83496
rect 268654 82560 268660 82612
rect 268712 82600 268718 82612
rect 398926 82600 398932 82612
rect 268712 82572 398932 82600
rect 268712 82560 268718 82572
rect 398926 82560 398932 82572
rect 398984 82560 398990 82612
rect 270402 82492 270408 82544
rect 270460 82532 270466 82544
rect 409874 82532 409880 82544
rect 270460 82504 409880 82532
rect 270460 82492 270466 82504
rect 409874 82492 409880 82504
rect 409932 82492 409938 82544
rect 271690 82424 271696 82476
rect 271748 82464 271754 82476
rect 414014 82464 414020 82476
rect 271748 82436 414020 82464
rect 271748 82424 271754 82436
rect 414014 82424 414020 82436
rect 414072 82424 414078 82476
rect 273070 82356 273076 82408
rect 273128 82396 273134 82408
rect 423766 82396 423772 82408
rect 273128 82368 423772 82396
rect 273128 82356 273134 82368
rect 423766 82356 423772 82368
rect 423824 82356 423830 82408
rect 276934 82288 276940 82340
rect 276992 82328 276998 82340
rect 445754 82328 445760 82340
rect 276992 82300 445760 82328
rect 276992 82288 276998 82300
rect 445754 82288 445760 82300
rect 445812 82288 445818 82340
rect 5442 82220 5448 82272
rect 5500 82260 5506 82272
rect 200942 82260 200948 82272
rect 5500 82232 200948 82260
rect 5500 82220 5506 82232
rect 200942 82220 200948 82232
rect 201000 82220 201006 82272
rect 278498 82220 278504 82272
rect 278556 82260 278562 82272
rect 456886 82260 456892 82272
rect 278556 82232 456892 82260
rect 278556 82220 278562 82232
rect 456886 82220 456892 82232
rect 456944 82220 456950 82272
rect 21450 82152 21456 82204
rect 21508 82192 21514 82204
rect 203150 82192 203156 82204
rect 21508 82164 203156 82192
rect 21508 82152 21514 82164
rect 203150 82152 203156 82164
rect 203208 82152 203214 82204
rect 246666 82152 246672 82204
rect 246724 82192 246730 82204
rect 271230 82192 271236 82204
rect 246724 82164 271236 82192
rect 246724 82152 246730 82164
rect 271230 82152 271236 82164
rect 271288 82152 271294 82204
rect 284110 82152 284116 82204
rect 284168 82192 284174 82204
rect 485774 82192 485780 82204
rect 284168 82164 485780 82192
rect 284168 82152 284174 82164
rect 485774 82152 485780 82164
rect 485832 82152 485838 82204
rect 200758 82084 200764 82136
rect 200816 82124 200822 82136
rect 226794 82124 226800 82136
rect 200816 82096 226800 82124
rect 200816 82084 200822 82096
rect 226794 82084 226800 82096
rect 226852 82084 226858 82136
rect 249518 82084 249524 82136
rect 249576 82124 249582 82136
rect 278130 82124 278136 82136
rect 249576 82096 278136 82124
rect 249576 82084 249582 82096
rect 278130 82084 278136 82096
rect 278188 82084 278194 82136
rect 298002 82084 298008 82136
rect 298060 82124 298066 82136
rect 571334 82124 571340 82136
rect 298060 82096 571340 82124
rect 298060 82084 298066 82096
rect 571334 82084 571340 82096
rect 571392 82084 571398 82136
rect 255038 81132 255044 81184
rect 255096 81172 255102 81184
rect 318058 81172 318064 81184
rect 255096 81144 318064 81172
rect 255096 81132 255102 81144
rect 318058 81132 318064 81144
rect 318116 81132 318122 81184
rect 271782 81064 271788 81116
rect 271840 81104 271846 81116
rect 416774 81104 416780 81116
rect 271840 81076 416780 81104
rect 271840 81064 271846 81076
rect 416774 81064 416780 81076
rect 416832 81064 416838 81116
rect 273162 80996 273168 81048
rect 273220 81036 273226 81048
rect 427814 81036 427820 81048
rect 273220 81008 427820 81036
rect 273220 80996 273226 81008
rect 427814 80996 427820 81008
rect 427872 80996 427878 81048
rect 274450 80928 274456 80980
rect 274508 80968 274514 80980
rect 434714 80968 434720 80980
rect 274508 80940 434720 80968
rect 274508 80928 274514 80940
rect 434714 80928 434720 80940
rect 434772 80928 434778 80980
rect 278590 80860 278596 80912
rect 278648 80900 278654 80912
rect 459554 80900 459560 80912
rect 278648 80872 459560 80900
rect 278648 80860 278654 80872
rect 459554 80860 459560 80872
rect 459612 80860 459618 80912
rect 282730 80792 282736 80844
rect 282788 80832 282794 80844
rect 477494 80832 477500 80844
rect 282788 80804 477500 80832
rect 282788 80792 282794 80804
rect 477494 80792 477500 80804
rect 477552 80792 477558 80844
rect 286870 80724 286876 80776
rect 286928 80764 286934 80776
rect 503714 80764 503720 80776
rect 286928 80736 503720 80764
rect 286928 80724 286934 80736
rect 503714 80724 503720 80736
rect 503772 80724 503778 80776
rect 299198 80656 299204 80708
rect 299256 80696 299262 80708
rect 574094 80696 574100 80708
rect 299256 80668 574100 80696
rect 299256 80656 299262 80668
rect 574094 80656 574100 80668
rect 574152 80656 574158 80708
rect 257890 79704 257896 79756
rect 257948 79744 257954 79756
rect 331858 79744 331864 79756
rect 257948 79716 331864 79744
rect 257948 79704 257954 79716
rect 331858 79704 331864 79716
rect 331916 79704 331922 79756
rect 260558 79636 260564 79688
rect 260616 79676 260622 79688
rect 347774 79676 347780 79688
rect 260616 79648 347780 79676
rect 260616 79636 260622 79648
rect 347774 79636 347780 79648
rect 347832 79636 347838 79688
rect 277026 79568 277032 79620
rect 277084 79608 277090 79620
rect 448606 79608 448612 79620
rect 277084 79580 448612 79608
rect 277084 79568 277090 79580
rect 448606 79568 448612 79580
rect 448664 79568 448670 79620
rect 281350 79500 281356 79552
rect 281408 79540 281414 79552
rect 472618 79540 472624 79552
rect 281408 79512 472624 79540
rect 281408 79500 281414 79512
rect 472618 79500 472624 79512
rect 472676 79500 472682 79552
rect 282546 79432 282552 79484
rect 282604 79472 282610 79484
rect 481726 79472 481732 79484
rect 282604 79444 481732 79472
rect 282604 79432 282610 79444
rect 481726 79432 481732 79444
rect 481784 79432 481790 79484
rect 286594 79364 286600 79416
rect 286652 79404 286658 79416
rect 506566 79404 506572 79416
rect 286652 79376 506572 79404
rect 286652 79364 286658 79376
rect 506566 79364 506572 79376
rect 506624 79364 506630 79416
rect 256050 79296 256056 79348
rect 256108 79336 256114 79348
rect 276014 79336 276020 79348
rect 256108 79308 276020 79336
rect 256108 79296 256114 79308
rect 276014 79296 276020 79308
rect 276072 79296 276078 79348
rect 290826 79296 290832 79348
rect 290884 79336 290890 79348
rect 530578 79336 530584 79348
rect 290884 79308 530584 79336
rect 290884 79296 290890 79308
rect 530578 79296 530584 79308
rect 530636 79296 530642 79348
rect 258902 78276 258908 78328
rect 258960 78316 258966 78328
rect 340966 78316 340972 78328
rect 258960 78288 340972 78316
rect 258960 78276 258966 78288
rect 340966 78276 340972 78288
rect 341024 78276 341030 78328
rect 261846 78208 261852 78260
rect 261904 78248 261910 78260
rect 357526 78248 357532 78260
rect 261904 78220 357532 78248
rect 261904 78208 261910 78220
rect 357526 78208 357532 78220
rect 357584 78208 357590 78260
rect 283834 78140 283840 78192
rect 283892 78180 283898 78192
rect 490006 78180 490012 78192
rect 283892 78152 490012 78180
rect 283892 78140 283898 78152
rect 490006 78140 490012 78152
rect 490064 78140 490070 78192
rect 285398 78072 285404 78124
rect 285456 78112 285462 78124
rect 492674 78112 492680 78124
rect 285456 78084 492680 78112
rect 285456 78072 285462 78084
rect 492674 78072 492680 78084
rect 492732 78072 492738 78124
rect 287882 78004 287888 78056
rect 287940 78044 287946 78056
rect 510614 78044 510620 78056
rect 287940 78016 510620 78044
rect 287940 78004 287946 78016
rect 510614 78004 510620 78016
rect 510672 78004 510678 78056
rect 293770 77936 293776 77988
rect 293828 77976 293834 77988
rect 542354 77976 542360 77988
rect 293828 77948 542360 77976
rect 293828 77936 293834 77948
rect 542354 77936 542360 77948
rect 542412 77936 542418 77988
rect 276658 76712 276664 76764
rect 276716 76752 276722 76764
rect 411254 76752 411260 76764
rect 276716 76724 411260 76752
rect 276716 76712 276722 76724
rect 411254 76712 411260 76724
rect 411312 76712 411318 76764
rect 289262 76644 289268 76696
rect 289320 76684 289326 76696
rect 517514 76684 517520 76696
rect 289320 76656 517520 76684
rect 289320 76644 289326 76656
rect 517514 76644 517520 76656
rect 517572 76644 517578 76696
rect 292390 76576 292396 76628
rect 292448 76616 292454 76628
rect 535454 76616 535460 76628
rect 292448 76588 535460 76616
rect 292448 76576 292454 76588
rect 535454 76576 535460 76588
rect 535512 76576 535518 76628
rect 295058 76508 295064 76560
rect 295116 76548 295122 76560
rect 548518 76548 548524 76560
rect 295116 76520 548524 76548
rect 295116 76508 295122 76520
rect 548518 76508 548524 76520
rect 548576 76508 548582 76560
rect 275278 75284 275284 75336
rect 275336 75324 275342 75336
rect 429194 75324 429200 75336
rect 275336 75296 429200 75324
rect 275336 75284 275342 75296
rect 429194 75284 429200 75296
rect 429252 75284 429258 75336
rect 296530 75216 296536 75268
rect 296588 75256 296594 75268
rect 560294 75256 560300 75268
rect 296588 75228 560300 75256
rect 296588 75216 296594 75228
rect 560294 75216 560300 75228
rect 560352 75216 560358 75268
rect 250990 75148 250996 75200
rect 251048 75188 251054 75200
rect 298094 75188 298100 75200
rect 251048 75160 298100 75188
rect 251048 75148 251054 75160
rect 298094 75148 298100 75160
rect 298152 75148 298158 75200
rect 299290 75148 299296 75200
rect 299348 75188 299354 75200
rect 578234 75188 578240 75200
rect 299348 75160 578240 75188
rect 299348 75148 299354 75160
rect 578234 75148 578240 75160
rect 578292 75148 578298 75200
rect 279970 73856 279976 73908
rect 280028 73896 280034 73908
rect 467834 73896 467840 73908
rect 280028 73868 467840 73896
rect 280028 73856 280034 73868
rect 467834 73856 467840 73868
rect 467892 73856 467898 73908
rect 299382 73788 299388 73840
rect 299440 73828 299446 73840
rect 582926 73828 582932 73840
rect 299440 73800 582932 73828
rect 299440 73788 299446 73800
rect 582926 73788 582932 73800
rect 582984 73788 582990 73840
rect 305638 73108 305644 73160
rect 305696 73148 305702 73160
rect 579982 73148 579988 73160
rect 305696 73120 579988 73148
rect 305696 73108 305702 73120
rect 579982 73108 579988 73120
rect 580040 73108 580046 73160
rect 3418 71680 3424 71732
rect 3476 71720 3482 71732
rect 157978 71720 157984 71732
rect 3476 71692 157984 71720
rect 3476 71680 3482 71692
rect 157978 71680 157984 71692
rect 158036 71680 158042 71732
rect 158070 71000 158076 71052
rect 158128 71040 158134 71052
rect 226702 71040 226708 71052
rect 158128 71012 226708 71040
rect 158128 71000 158134 71012
rect 226702 71000 226708 71012
rect 226760 71000 226766 71052
rect 68922 69640 68928 69692
rect 68980 69680 68986 69692
rect 210510 69680 210516 69692
rect 68980 69652 210516 69680
rect 68980 69640 68986 69652
rect 210510 69640 210516 69652
rect 210568 69640 210574 69692
rect 278314 69640 278320 69692
rect 278372 69680 278378 69692
rect 454034 69680 454040 69692
rect 278372 69652 454040 69680
rect 278372 69640 278378 69652
rect 454034 69640 454040 69652
rect 454092 69640 454098 69692
rect 313918 60664 313924 60716
rect 313976 60704 313982 60716
rect 580166 60704 580172 60716
rect 313976 60676 580172 60704
rect 313976 60664 313982 60676
rect 580166 60664 580172 60676
rect 580224 60664 580230 60716
rect 3050 59304 3056 59356
rect 3108 59344 3114 59356
rect 146938 59344 146944 59356
rect 3108 59316 146944 59344
rect 3108 59304 3114 59316
rect 146938 59304 146944 59316
rect 146996 59304 147002 59356
rect 3418 45500 3424 45552
rect 3476 45540 3482 45552
rect 151078 45540 151084 45552
rect 3476 45512 151084 45540
rect 3476 45500 3482 45512
rect 151078 45500 151084 45512
rect 151136 45500 151142 45552
rect 249610 39312 249616 39364
rect 249668 39352 249674 39364
rect 284294 39352 284300 39364
rect 249668 39324 284300 39352
rect 249668 39312 249674 39324
rect 284294 39312 284300 39324
rect 284352 39312 284358 39364
rect 242526 37884 242532 37936
rect 242584 37924 242590 37936
rect 248414 37924 248420 37936
rect 242584 37896 248420 37924
rect 242584 37884 242590 37896
rect 248414 37884 248420 37896
rect 248472 37884 248478 37936
rect 89070 35164 89076 35216
rect 89128 35204 89134 35216
rect 214282 35204 214288 35216
rect 89128 35176 214288 35204
rect 89128 35164 89134 35176
rect 214282 35164 214288 35176
rect 214340 35164 214346 35216
rect 580258 33940 580264 33992
rect 580316 33980 580322 33992
rect 582558 33980 582564 33992
rect 580316 33952 582564 33980
rect 580316 33940 580322 33952
rect 582558 33940 582564 33952
rect 582616 33940 582622 33992
rect 275922 33736 275928 33788
rect 275980 33776 275986 33788
rect 440326 33776 440332 33788
rect 275980 33748 440332 33776
rect 275980 33736 275986 33748
rect 440326 33736 440332 33748
rect 440384 33736 440390 33788
rect 2866 33056 2872 33108
rect 2924 33096 2930 33108
rect 156598 33096 156604 33108
rect 2924 33068 156604 33096
rect 2924 33056 2930 33068
rect 156598 33056 156604 33068
rect 156656 33056 156662 33108
rect 273898 32376 273904 32428
rect 273956 32416 273962 32428
rect 404354 32416 404360 32428
rect 273956 32388 404360 32416
rect 273956 32376 273962 32388
rect 404354 32376 404360 32388
rect 404412 32376 404418 32428
rect 248046 31016 248052 31068
rect 248104 31056 248110 31068
rect 280154 31056 280160 31068
rect 248104 31028 280160 31056
rect 248104 31016 248110 31028
rect 280154 31016 280160 31028
rect 280212 31016 280218 31068
rect 280982 31016 280988 31068
rect 281040 31056 281046 31068
rect 474734 31056 474740 31068
rect 281040 31028 474740 31056
rect 281040 31016 281046 31028
rect 474734 31016 474740 31028
rect 474792 31016 474798 31068
rect 257614 29656 257620 29708
rect 257672 29696 257678 29708
rect 336090 29696 336096 29708
rect 257672 29668 336096 29696
rect 257672 29656 257678 29668
rect 336090 29656 336096 29668
rect 336148 29656 336154 29708
rect 335998 29588 336004 29640
rect 336056 29628 336062 29640
rect 436094 29628 436100 29640
rect 336056 29600 436100 29628
rect 336056 29588 336062 29600
rect 436094 29588 436100 29600
rect 436152 29588 436158 29640
rect 258994 28228 259000 28280
rect 259052 28268 259058 28280
rect 342898 28268 342904 28280
rect 259052 28240 342904 28268
rect 259052 28228 259058 28240
rect 342898 28228 342904 28240
rect 342956 28228 342962 28280
rect 256326 26868 256332 26920
rect 256384 26908 256390 26920
rect 329834 26908 329840 26920
rect 256384 26880 329840 26908
rect 256384 26868 256390 26880
rect 329834 26868 329840 26880
rect 329892 26868 329898 26920
rect 113082 25508 113088 25560
rect 113140 25548 113146 25560
rect 218330 25548 218336 25560
rect 113140 25520 218336 25548
rect 113140 25508 113146 25520
rect 218330 25508 218336 25520
rect 218388 25508 218394 25560
rect 295150 25508 295156 25560
rect 295208 25548 295214 25560
rect 556246 25548 556252 25560
rect 295208 25520 556252 25548
rect 295208 25508 295214 25520
rect 556246 25508 556252 25520
rect 556304 25508 556310 25560
rect 253474 24080 253480 24132
rect 253532 24120 253538 24132
rect 311894 24120 311900 24132
rect 253532 24092 311900 24120
rect 253532 24080 253538 24092
rect 311894 24080 311900 24092
rect 311952 24080 311958 24132
rect 312630 24080 312636 24132
rect 312688 24120 312694 24132
rect 393314 24120 393320 24132
rect 312688 24092 393320 24120
rect 312688 24080 312694 24092
rect 393314 24080 393320 24092
rect 393372 24080 393378 24132
rect 26142 22720 26148 22772
rect 26200 22760 26206 22772
rect 35250 22760 35256 22772
rect 26200 22732 35256 22760
rect 26200 22720 26206 22732
rect 35250 22720 35256 22732
rect 35308 22720 35314 22772
rect 252370 22720 252376 22772
rect 252428 22760 252434 22772
rect 300854 22760 300860 22772
rect 252428 22732 300860 22760
rect 252428 22720 252434 22732
rect 300854 22720 300860 22732
rect 300912 22720 300918 22772
rect 44082 21360 44088 21412
rect 44140 21400 44146 21412
rect 200850 21400 200856 21412
rect 44140 21372 200856 21400
rect 44140 21360 44146 21372
rect 200850 21360 200856 21372
rect 200908 21360 200914 21412
rect 3418 20612 3424 20664
rect 3476 20652 3482 20664
rect 144178 20652 144184 20664
rect 3476 20624 144184 20652
rect 3476 20612 3482 20624
rect 144178 20612 144184 20624
rect 144236 20612 144242 20664
rect 177850 19932 177856 19984
rect 177908 19972 177914 19984
rect 229462 19972 229468 19984
rect 177908 19944 229468 19972
rect 177908 19932 177914 19944
rect 229462 19932 229468 19944
rect 229520 19932 229526 19984
rect 296254 19932 296260 19984
rect 296312 19972 296318 19984
rect 564618 19972 564624 19984
rect 296312 19944 564624 19972
rect 296312 19932 296318 19944
rect 564618 19932 564624 19944
rect 564676 19932 564682 19984
rect 246758 18708 246764 18760
rect 246816 18748 246822 18760
rect 257338 18748 257344 18760
rect 246816 18720 257344 18748
rect 246816 18708 246822 18720
rect 257338 18708 257344 18720
rect 257396 18708 257402 18760
rect 243906 18640 243912 18692
rect 243964 18680 243970 18692
rect 255314 18680 255320 18692
rect 243964 18652 255320 18680
rect 243964 18640 243970 18652
rect 255314 18640 255320 18652
rect 255372 18640 255378 18692
rect 143442 18572 143448 18624
rect 143500 18612 143506 18624
rect 224034 18612 224040 18624
rect 143500 18584 224040 18612
rect 143500 18572 143506 18584
rect 224034 18572 224040 18584
rect 224092 18572 224098 18624
rect 245378 18572 245384 18624
rect 245436 18612 245442 18624
rect 260190 18612 260196 18624
rect 245436 18584 260196 18612
rect 245436 18572 245442 18584
rect 260190 18572 260196 18584
rect 260248 18572 260254 18624
rect 268470 18572 268476 18624
rect 268528 18612 268534 18624
rect 375374 18612 375380 18624
rect 268528 18584 375380 18612
rect 268528 18572 268534 18584
rect 375374 18572 375380 18584
rect 375432 18572 375438 18624
rect 232590 17892 232596 17944
rect 232648 17932 232654 17944
rect 236730 17932 236736 17944
rect 232648 17904 236736 17932
rect 232648 17892 232654 17904
rect 236730 17892 236736 17904
rect 236788 17892 236794 17944
rect 250438 17892 250444 17944
rect 250496 17932 250502 17944
rect 251174 17932 251180 17944
rect 250496 17904 251180 17932
rect 250496 17892 250502 17904
rect 251174 17892 251180 17904
rect 251232 17892 251238 17944
rect 249058 17824 249064 17876
rect 249116 17864 249122 17876
rect 253934 17864 253940 17876
rect 249116 17836 253940 17864
rect 249116 17824 249122 17836
rect 253934 17824 253940 17836
rect 253992 17824 253998 17876
rect 97350 17212 97356 17264
rect 97408 17252 97414 17264
rect 215570 17252 215576 17264
rect 97408 17224 215576 17252
rect 97408 17212 97414 17224
rect 215570 17212 215576 17224
rect 215628 17212 215634 17264
rect 254762 17212 254768 17264
rect 254820 17252 254826 17264
rect 322934 17252 322940 17264
rect 254820 17224 322940 17252
rect 254820 17212 254826 17224
rect 322934 17212 322940 17224
rect 322992 17212 322998 17264
rect 436738 17212 436744 17264
rect 436796 17252 436802 17264
rect 442994 17252 443000 17264
rect 436796 17224 443000 17252
rect 436796 17212 436802 17224
rect 442994 17212 443000 17224
rect 443052 17212 443058 17264
rect 454678 17212 454684 17264
rect 454736 17252 454742 17264
rect 471974 17252 471980 17264
rect 454736 17224 471980 17252
rect 454736 17212 454742 17224
rect 471974 17212 471980 17224
rect 472032 17212 472038 17264
rect 39390 15852 39396 15904
rect 39448 15892 39454 15904
rect 206278 15892 206284 15904
rect 39448 15864 206284 15892
rect 39448 15852 39454 15864
rect 206278 15852 206284 15864
rect 206336 15852 206342 15904
rect 227622 15852 227628 15904
rect 227680 15892 227686 15904
rect 232498 15892 232504 15904
rect 227680 15864 232504 15892
rect 227680 15852 227686 15864
rect 232498 15852 232504 15864
rect 232556 15852 232562 15904
rect 293494 15852 293500 15904
rect 293552 15892 293558 15904
rect 546678 15892 546684 15904
rect 293552 15864 546684 15892
rect 293552 15852 293558 15864
rect 546678 15852 546684 15864
rect 546736 15852 546742 15904
rect 236638 15172 236644 15224
rect 236696 15212 236702 15224
rect 239030 15212 239036 15224
rect 236696 15184 239036 15212
rect 236696 15172 236702 15184
rect 239030 15172 239036 15184
rect 239088 15172 239094 15224
rect 245102 14492 245108 14544
rect 245160 14532 245166 14544
rect 258718 14532 258724 14544
rect 245160 14504 258724 14532
rect 245160 14492 245166 14504
rect 258718 14492 258724 14504
rect 258776 14492 258782 14544
rect 119890 14424 119896 14476
rect 119948 14464 119954 14476
rect 219802 14464 219808 14476
rect 119948 14436 219808 14464
rect 119948 14424 119954 14436
rect 219802 14424 219808 14436
rect 219860 14424 219866 14476
rect 246850 14424 246856 14476
rect 246908 14464 246914 14476
rect 267734 14464 267740 14476
rect 246908 14436 267740 14464
rect 246908 14424 246914 14436
rect 267734 14424 267740 14436
rect 267792 14424 267798 14476
rect 287974 14424 287980 14476
rect 288032 14464 288038 14476
rect 514754 14464 514760 14476
rect 288032 14436 514760 14464
rect 288032 14424 288038 14436
rect 514754 14424 514760 14436
rect 514812 14424 514818 14476
rect 234062 13812 234068 13864
rect 234120 13852 234126 13864
rect 235074 13852 235080 13864
rect 234120 13824 235080 13852
rect 234120 13812 234126 13824
rect 235074 13812 235080 13824
rect 235132 13812 235138 13864
rect 64782 13064 64788 13116
rect 64840 13104 64846 13116
rect 197998 13104 198004 13116
rect 64840 13076 198004 13104
rect 64840 13064 64846 13076
rect 197998 13064 198004 13076
rect 198056 13064 198062 13116
rect 285490 13064 285496 13116
rect 285548 13104 285554 13116
rect 500218 13104 500224 13116
rect 285548 13076 500224 13104
rect 285548 13064 285554 13076
rect 500218 13064 500224 13076
rect 500276 13064 500282 13116
rect 357526 11772 357532 11824
rect 357584 11812 357590 11824
rect 358722 11812 358728 11824
rect 357584 11784 358728 11812
rect 357584 11772 357590 11784
rect 358722 11772 358728 11784
rect 358780 11772 358786 11824
rect 398926 11772 398932 11824
rect 398984 11812 398990 11824
rect 400122 11812 400128 11824
rect 398984 11784 400128 11812
rect 398984 11772 398990 11784
rect 400122 11772 400128 11784
rect 400180 11772 400186 11824
rect 35802 11704 35808 11756
rect 35860 11744 35866 11756
rect 206002 11744 206008 11756
rect 35860 11716 206008 11744
rect 35860 11704 35866 11716
rect 206002 11704 206008 11716
rect 206060 11704 206066 11756
rect 219342 11704 219348 11756
rect 219400 11744 219406 11756
rect 236362 11744 236368 11756
rect 219400 11716 236368 11744
rect 219400 11704 219406 11716
rect 236362 11704 236368 11716
rect 236420 11704 236426 11756
rect 242618 11704 242624 11756
rect 242676 11744 242682 11756
rect 252554 11744 252560 11756
rect 242676 11716 252560 11744
rect 242676 11704 242682 11716
rect 252554 11704 252560 11716
rect 252612 11704 252618 11756
rect 329098 11704 329104 11756
rect 329156 11744 329162 11756
rect 422570 11744 422576 11756
rect 329156 11716 422576 11744
rect 329156 11704 329162 11716
rect 422570 11704 422576 11716
rect 422628 11704 422634 11756
rect 423766 11704 423772 11756
rect 423824 11744 423830 11756
rect 424962 11744 424968 11756
rect 423824 11716 424968 11744
rect 423824 11704 423830 11716
rect 424962 11704 424968 11716
rect 425020 11704 425026 11756
rect 448606 11704 448612 11756
rect 448664 11744 448670 11756
rect 449802 11744 449808 11756
rect 448664 11716 449808 11744
rect 448664 11704 448670 11716
rect 449802 11704 449808 11716
rect 449860 11704 449866 11756
rect 223482 10344 223488 10396
rect 223540 10384 223546 10396
rect 233970 10384 233976 10396
rect 223540 10356 233976 10384
rect 223540 10344 223546 10356
rect 233970 10344 233976 10356
rect 234028 10344 234034 10396
rect 81342 10276 81348 10328
rect 81400 10316 81406 10328
rect 212902 10316 212908 10328
rect 81400 10288 212908 10316
rect 81400 10276 81406 10288
rect 212902 10276 212908 10288
rect 212960 10276 212966 10328
rect 217962 10276 217968 10328
rect 218020 10316 218026 10328
rect 228542 10316 228548 10328
rect 218020 10288 228548 10316
rect 218020 10276 218026 10288
rect 228542 10276 228548 10288
rect 228600 10276 228606 10328
rect 266998 10276 267004 10328
rect 267056 10316 267062 10328
rect 291194 10316 291200 10328
rect 267056 10288 291200 10316
rect 267056 10276 267062 10288
rect 291194 10276 291200 10288
rect 291252 10276 291258 10328
rect 292022 10276 292028 10328
rect 292080 10316 292086 10328
rect 539594 10316 539600 10328
rect 292080 10288 539600 10316
rect 292080 10276 292086 10288
rect 539594 10276 539600 10288
rect 539652 10276 539658 10328
rect 234154 9868 234160 9920
rect 234212 9908 234218 9920
rect 237834 9908 237840 9920
rect 234212 9880 237840 9908
rect 234212 9868 234218 9880
rect 237834 9868 237840 9880
rect 237892 9868 237898 9920
rect 234798 9596 234804 9648
rect 234856 9636 234862 9648
rect 237742 9636 237748 9648
rect 234856 9608 237748 9636
rect 234856 9596 234862 9608
rect 237742 9596 237748 9608
rect 237800 9596 237806 9648
rect 70210 8916 70216 8968
rect 70268 8956 70274 8968
rect 211430 8956 211436 8968
rect 70268 8928 211436 8956
rect 70268 8916 70274 8928
rect 211430 8916 211436 8928
rect 211488 8916 211494 8968
rect 227530 8916 227536 8968
rect 227588 8956 227594 8968
rect 235350 8956 235356 8968
rect 227588 8928 235356 8956
rect 227588 8916 227594 8928
rect 235350 8916 235356 8928
rect 235408 8916 235414 8968
rect 285122 8916 285128 8968
rect 285180 8956 285186 8968
rect 497090 8956 497096 8968
rect 285180 8928 497096 8956
rect 285180 8916 285186 8928
rect 497090 8916 497096 8928
rect 497148 8916 497154 8968
rect 233418 8372 233424 8424
rect 233476 8412 233482 8424
rect 239122 8412 239128 8424
rect 233476 8384 239128 8412
rect 233476 8372 233482 8384
rect 239122 8372 239128 8384
rect 239180 8372 239186 8424
rect 242710 8236 242716 8288
rect 242768 8276 242774 8288
rect 245654 8276 245660 8288
rect 242768 8248 245660 8276
rect 242768 8236 242774 8248
rect 245654 8236 245660 8248
rect 245712 8236 245718 8288
rect 393958 8236 393964 8288
rect 394016 8276 394022 8288
rect 401318 8276 401324 8288
rect 394016 8248 401324 8276
rect 394016 8236 394022 8248
rect 401318 8236 401324 8248
rect 401376 8236 401382 8288
rect 443638 8236 443644 8288
rect 443696 8276 443702 8288
rect 450906 8276 450912 8288
rect 443696 8248 450912 8276
rect 443696 8236 443702 8248
rect 450906 8236 450912 8248
rect 450964 8236 450970 8288
rect 202690 7692 202696 7744
rect 202748 7732 202754 7744
rect 233878 7732 233884 7744
rect 202748 7704 233884 7732
rect 202748 7692 202754 7704
rect 233878 7692 233884 7704
rect 233936 7692 233942 7744
rect 124674 7624 124680 7676
rect 124732 7664 124738 7676
rect 210418 7664 210424 7676
rect 124732 7636 210424 7664
rect 124732 7624 124738 7636
rect 210418 7624 210424 7636
rect 210476 7624 210482 7676
rect 102226 7556 102232 7608
rect 102284 7596 102290 7608
rect 217502 7596 217508 7608
rect 102284 7568 217508 7596
rect 102284 7556 102290 7568
rect 217502 7556 217508 7568
rect 217560 7556 217566 7608
rect 400858 7556 400864 7608
rect 400916 7596 400922 7608
rect 408402 7596 408408 7608
rect 400916 7568 408408 7596
rect 400916 7556 400922 7568
rect 408402 7556 408408 7568
rect 408460 7556 408466 7608
rect 450538 7556 450544 7608
rect 450596 7596 450602 7608
rect 465166 7596 465172 7608
rect 450596 7568 465172 7596
rect 450596 7556 450602 7568
rect 465166 7556 465172 7568
rect 465224 7556 465230 7608
rect 229830 7420 229836 7472
rect 229888 7460 229894 7472
rect 235258 7460 235264 7472
rect 229888 7432 235264 7460
rect 229888 7420 229894 7432
rect 235258 7420 235264 7432
rect 235316 7420 235322 7472
rect 3418 6808 3424 6860
rect 3476 6848 3482 6860
rect 128998 6848 129004 6860
rect 3476 6820 129004 6848
rect 3476 6808 3482 6820
rect 128998 6808 129004 6820
rect 129056 6808 129062 6860
rect 199102 6264 199108 6316
rect 199160 6304 199166 6316
rect 229738 6304 229744 6316
rect 199160 6276 229744 6304
rect 199160 6264 199166 6276
rect 229738 6264 229744 6276
rect 229796 6264 229802 6316
rect 131758 6196 131764 6248
rect 131816 6236 131822 6248
rect 222470 6236 222476 6248
rect 131816 6208 222476 6236
rect 131816 6196 131822 6208
rect 222470 6196 222476 6208
rect 222528 6196 222534 6248
rect 107010 6128 107016 6180
rect 107068 6168 107074 6180
rect 215938 6168 215944 6180
rect 107068 6140 215944 6168
rect 107068 6128 107074 6140
rect 215938 6128 215944 6140
rect 215996 6128 216002 6180
rect 249242 6128 249248 6180
rect 249300 6168 249306 6180
rect 287790 6168 287796 6180
rect 249300 6140 287796 6168
rect 249300 6128 249306 6140
rect 287790 6128 287796 6140
rect 287848 6128 287854 6180
rect 289354 6128 289360 6180
rect 289412 6168 289418 6180
rect 521838 6168 521844 6180
rect 289412 6140 521844 6168
rect 289412 6128 289418 6140
rect 521838 6128 521844 6140
rect 521896 6128 521902 6180
rect 241330 5516 241336 5568
rect 241388 5556 241394 5568
rect 241698 5556 241704 5568
rect 241388 5528 241704 5556
rect 241388 5516 241394 5528
rect 241698 5516 241704 5528
rect 241756 5516 241762 5568
rect 242802 5516 242808 5568
rect 242860 5556 242866 5568
rect 246390 5556 246396 5568
rect 242860 5528 246396 5556
rect 242860 5516 242866 5528
rect 246390 5516 246396 5528
rect 246448 5516 246454 5568
rect 245194 5448 245200 5500
rect 245252 5488 245258 5500
rect 251082 5488 251088 5500
rect 245252 5460 251088 5488
rect 245252 5448 245258 5460
rect 251082 5448 251088 5460
rect 251140 5448 251146 5500
rect 250714 4972 250720 5024
rect 250772 5012 250778 5024
rect 297266 5012 297272 5024
rect 250772 4984 297272 5012
rect 250772 4972 250778 4984
rect 297266 4972 297272 4984
rect 297324 4972 297330 5024
rect 212166 4904 212172 4956
rect 212224 4944 212230 4956
rect 231118 4944 231124 4956
rect 212224 4916 231124 4944
rect 212224 4904 212230 4916
rect 231118 4904 231124 4916
rect 231176 4904 231182 4956
rect 278038 4904 278044 4956
rect 278096 4944 278102 4956
rect 372890 4944 372896 4956
rect 278096 4916 372896 4944
rect 278096 4904 278102 4916
rect 372890 4904 372896 4916
rect 372948 4904 372954 4956
rect 99834 4836 99840 4888
rect 99892 4876 99898 4888
rect 214558 4876 214564 4888
rect 99892 4848 214564 4876
rect 99892 4836 99898 4848
rect 214558 4836 214564 4848
rect 214616 4836 214622 4888
rect 271138 4836 271144 4888
rect 271196 4876 271202 4888
rect 390646 4876 390652 4888
rect 271196 4848 390652 4876
rect 271196 4836 271202 4848
rect 390646 4836 390652 4848
rect 390704 4836 390710 4888
rect 98730 4768 98736 4820
rect 98788 4808 98794 4820
rect 217134 4808 217140 4820
rect 98788 4780 217140 4808
rect 98788 4768 98794 4780
rect 217134 4768 217140 4780
rect 217192 4768 217198 4820
rect 269758 4768 269764 4820
rect 269816 4808 269822 4820
rect 278314 4808 278320 4820
rect 269816 4780 278320 4808
rect 269816 4768 269822 4780
rect 278314 4768 278320 4780
rect 278372 4768 278378 4820
rect 294782 4768 294788 4820
rect 294840 4808 294846 4820
rect 553762 4808 553768 4820
rect 294840 4780 553768 4808
rect 294840 4768 294846 4780
rect 553762 4768 553768 4780
rect 553820 4768 553826 4820
rect 152476 4168 152688 4196
rect 15930 4088 15936 4140
rect 15988 4128 15994 4140
rect 17218 4128 17224 4140
rect 15988 4100 17224 4128
rect 15988 4088 15994 4100
rect 17218 4088 17224 4100
rect 17276 4088 17282 4140
rect 20622 4088 20628 4140
rect 20680 4128 20686 4140
rect 21450 4128 21456 4140
rect 20680 4100 21456 4128
rect 20680 4088 20686 4100
rect 21450 4088 21456 4100
rect 21508 4088 21514 4140
rect 72602 4088 72608 4140
rect 72660 4128 72666 4140
rect 76558 4128 76564 4140
rect 72660 4100 76564 4128
rect 72660 4088 72666 4100
rect 76558 4088 76564 4100
rect 76616 4088 76622 4140
rect 148962 4088 148968 4140
rect 149020 4128 149026 4140
rect 149514 4128 149520 4140
rect 149020 4100 149520 4128
rect 149020 4088 149026 4100
rect 149514 4088 149520 4100
rect 149572 4088 149578 4140
rect 17034 4020 17040 4072
rect 17092 4060 17098 4072
rect 21358 4060 21364 4072
rect 17092 4032 21364 4060
rect 17092 4020 17098 4032
rect 21358 4020 21364 4032
rect 21416 4020 21422 4072
rect 58434 4020 58440 4072
rect 58492 4060 58498 4072
rect 65518 4060 65524 4072
rect 58492 4032 65524 4060
rect 58492 4020 58498 4032
rect 65518 4020 65524 4032
rect 65576 4020 65582 4072
rect 78582 4020 78588 4072
rect 78640 4060 78646 4072
rect 93118 4060 93124 4072
rect 78640 4032 93124 4060
rect 78640 4020 78646 4032
rect 93118 4020 93124 4032
rect 93176 4020 93182 4072
rect 105538 4060 105544 4072
rect 93826 4032 105544 4060
rect 13538 3952 13544 4004
rect 13596 3992 13602 4004
rect 18598 3992 18604 4004
rect 13596 3964 18604 3992
rect 13596 3952 13602 3964
rect 18598 3952 18604 3964
rect 18656 3952 18662 4004
rect 24210 3952 24216 4004
rect 24268 3992 24274 4004
rect 24268 3964 26234 3992
rect 24268 3952 24274 3964
rect 14660 3896 17448 3924
rect 14550 3720 14556 3732
rect 6886 3692 14556 3720
rect 6454 3612 6460 3664
rect 6512 3652 6518 3664
rect 6886 3652 6914 3692
rect 14550 3680 14556 3692
rect 14608 3680 14614 3732
rect 6512 3624 6914 3652
rect 6512 3612 6518 3624
rect 11146 3612 11152 3664
rect 11204 3652 11210 3664
rect 12250 3652 12256 3664
rect 11204 3624 12256 3652
rect 11204 3612 11210 3624
rect 12250 3612 12256 3624
rect 12308 3612 12314 3664
rect 2866 3544 2872 3596
rect 2924 3584 2930 3596
rect 14660 3584 14688 3896
rect 17420 3856 17448 3896
rect 19426 3884 19432 3936
rect 19484 3924 19490 3936
rect 19484 3896 25728 3924
rect 19484 3884 19490 3896
rect 17420 3828 22094 3856
rect 22066 3788 22094 3828
rect 25498 3788 25504 3800
rect 22066 3760 25504 3788
rect 25498 3748 25504 3760
rect 25556 3748 25562 3800
rect 25700 3788 25728 3896
rect 26206 3856 26234 3964
rect 54938 3952 54944 4004
rect 54996 3992 55002 4004
rect 61378 3992 61384 4004
rect 54996 3964 61384 3992
rect 54996 3952 55002 3964
rect 61378 3952 61384 3964
rect 61436 3952 61442 4004
rect 63218 3952 63224 4004
rect 63276 3992 63282 4004
rect 87598 3992 87604 4004
rect 63276 3964 87604 3992
rect 63276 3952 63282 3964
rect 87598 3952 87604 3964
rect 87656 3952 87662 4004
rect 91646 3952 91652 4004
rect 91704 3992 91710 4004
rect 93826 3992 93854 4032
rect 105538 4020 105544 4032
rect 105596 4020 105602 4072
rect 111610 4020 111616 4072
rect 111668 4060 111674 4072
rect 115198 4060 115204 4072
rect 111668 4032 115204 4060
rect 111668 4020 111674 4032
rect 115198 4020 115204 4032
rect 115256 4020 115262 4072
rect 117590 4020 117596 4072
rect 117648 4060 117654 4072
rect 152476 4060 152504 4168
rect 152660 4128 152688 4168
rect 241422 4156 241428 4208
rect 241480 4196 241486 4208
rect 242894 4196 242900 4208
rect 241480 4168 242900 4196
rect 241480 4156 241486 4168
rect 242894 4156 242900 4168
rect 242952 4156 242958 4208
rect 152660 4100 152780 4128
rect 117648 4032 152504 4060
rect 152752 4060 152780 4100
rect 154206 4088 154212 4140
rect 154264 4128 154270 4140
rect 155218 4128 155224 4140
rect 154264 4100 155224 4128
rect 154264 4088 154270 4100
rect 155218 4088 155224 4100
rect 155276 4088 155282 4140
rect 155402 4088 155408 4140
rect 155460 4128 155466 4140
rect 156690 4128 156696 4140
rect 155460 4100 156696 4128
rect 155460 4088 155466 4100
rect 156690 4088 156696 4100
rect 156748 4088 156754 4140
rect 160094 4088 160100 4140
rect 160152 4128 160158 4140
rect 161382 4128 161388 4140
rect 160152 4100 161388 4128
rect 160152 4088 160158 4100
rect 161382 4088 161388 4100
rect 161440 4088 161446 4140
rect 161474 4088 161480 4140
rect 161532 4128 161538 4140
rect 200758 4128 200764 4140
rect 161532 4100 200764 4128
rect 161532 4088 161538 4100
rect 200758 4088 200764 4100
rect 200816 4088 200822 4140
rect 219250 4088 219256 4140
rect 219308 4128 219314 4140
rect 228450 4128 228456 4140
rect 219308 4100 228456 4128
rect 219308 4088 219314 4100
rect 228450 4088 228456 4100
rect 228508 4088 228514 4140
rect 265342 4128 265348 4140
rect 258046 4100 265348 4128
rect 172146 4060 172152 4072
rect 152752 4032 172152 4060
rect 117648 4020 117654 4032
rect 172146 4020 172152 4032
rect 172204 4020 172210 4072
rect 189718 4020 189724 4072
rect 189776 4060 189782 4072
rect 191190 4060 191196 4072
rect 189776 4032 191196 4060
rect 189776 4020 189782 4032
rect 191190 4020 191196 4032
rect 191248 4020 191254 4072
rect 198642 4020 198648 4072
rect 198700 4060 198706 4072
rect 203886 4060 203892 4072
rect 198700 4032 203892 4060
rect 198700 4020 198706 4032
rect 203886 4020 203892 4032
rect 203944 4020 203950 4072
rect 209774 4020 209780 4072
rect 209832 4060 209838 4072
rect 222838 4060 222844 4072
rect 209832 4032 222844 4060
rect 209832 4020 209838 4032
rect 222838 4020 222844 4032
rect 222896 4020 222902 4072
rect 255958 4020 255964 4072
rect 256016 4060 256022 4072
rect 258046 4060 258074 4100
rect 265342 4088 265348 4100
rect 265400 4088 265406 4140
rect 353938 4088 353944 4140
rect 353996 4128 354002 4140
rect 355226 4128 355232 4140
rect 353996 4100 355232 4128
rect 353996 4088 354002 4100
rect 355226 4088 355232 4100
rect 355284 4088 355290 4140
rect 382918 4088 382924 4140
rect 382976 4128 382982 4140
rect 384758 4128 384764 4140
rect 382976 4100 384764 4128
rect 382976 4088 382982 4100
rect 384758 4088 384764 4100
rect 384816 4088 384822 4140
rect 460198 4088 460204 4140
rect 460256 4128 460262 4140
rect 462774 4128 462780 4140
rect 460256 4100 462780 4128
rect 460256 4088 460262 4100
rect 462774 4088 462780 4100
rect 462832 4088 462838 4140
rect 479518 4088 479524 4140
rect 479576 4128 479582 4140
rect 480530 4128 480536 4140
rect 479576 4100 480536 4128
rect 479576 4088 479582 4100
rect 480530 4088 480536 4100
rect 480588 4088 480594 4140
rect 547138 4088 547144 4140
rect 547196 4128 547202 4140
rect 549070 4128 549076 4140
rect 547196 4100 549076 4128
rect 547196 4088 547202 4100
rect 549070 4088 549076 4100
rect 549128 4088 549134 4140
rect 566550 4088 566556 4140
rect 566608 4128 566614 4140
rect 568022 4128 568028 4140
rect 566608 4100 568028 4128
rect 566608 4088 566614 4100
rect 568022 4088 568028 4100
rect 568080 4088 568086 4140
rect 256016 4032 258074 4060
rect 256016 4020 256022 4032
rect 260834 4020 260840 4072
rect 260892 4060 260898 4072
rect 263594 4060 263600 4072
rect 260892 4032 263600 4060
rect 260892 4020 260898 4032
rect 263594 4020 263600 4032
rect 263652 4020 263658 4072
rect 276014 4020 276020 4072
rect 276072 4060 276078 4072
rect 280246 4060 280252 4072
rect 276072 4032 280252 4060
rect 276072 4020 276078 4032
rect 280246 4020 280252 4032
rect 280304 4020 280310 4072
rect 347038 4020 347044 4072
rect 347096 4060 347102 4072
rect 362310 4060 362316 4072
rect 347096 4032 362316 4060
rect 347096 4020 347102 4032
rect 362310 4020 362316 4032
rect 362368 4020 362374 4072
rect 91704 3964 93854 3992
rect 91704 3952 91710 3964
rect 93946 3952 93952 4004
rect 94004 3992 94010 4004
rect 108298 3992 108304 4004
rect 94004 3964 108304 3992
rect 94004 3952 94010 3964
rect 108298 3952 108304 3964
rect 108356 3952 108362 4004
rect 130562 3952 130568 4004
rect 130620 3992 130626 4004
rect 134518 3992 134524 4004
rect 130620 3964 134524 3992
rect 130620 3952 130626 3964
rect 134518 3952 134524 3964
rect 134576 3952 134582 4004
rect 137646 3952 137652 4004
rect 137704 3992 137710 4004
rect 142798 3992 142804 4004
rect 137704 3964 142804 3992
rect 137704 3952 137710 3964
rect 142798 3952 142804 3964
rect 142856 3952 142862 4004
rect 148318 3952 148324 4004
rect 148376 3992 148382 4004
rect 152550 3992 152556 4004
rect 148376 3964 152556 3992
rect 148376 3952 148382 3964
rect 152550 3952 152556 3964
rect 152608 3952 152614 4004
rect 152642 3952 152648 4004
rect 152700 3992 152706 4004
rect 225230 3992 225236 4004
rect 152700 3964 225236 3992
rect 152700 3952 152706 3964
rect 225230 3952 225236 3964
rect 225288 3952 225294 4004
rect 225322 3952 225328 4004
rect 225380 3992 225386 4004
rect 228358 3992 228364 4004
rect 225380 3964 228364 3992
rect 225380 3952 225386 3964
rect 228358 3952 228364 3964
rect 228416 3952 228422 4004
rect 228726 3952 228732 4004
rect 228784 3992 228790 4004
rect 236638 3992 236644 4004
rect 228784 3964 236644 3992
rect 228784 3952 228790 3964
rect 236638 3952 236644 3964
rect 236696 3952 236702 4004
rect 257338 3952 257344 4004
rect 257396 3992 257402 4004
rect 268838 3992 268844 4004
rect 257396 3964 268844 3992
rect 257396 3952 257402 3964
rect 268838 3952 268844 3964
rect 268896 3952 268902 4004
rect 279510 3952 279516 4004
rect 279568 3992 279574 4004
rect 287054 3992 287060 4004
rect 279568 3964 287060 3992
rect 279568 3952 279574 3964
rect 287054 3952 287060 3964
rect 287112 3952 287118 4004
rect 327718 3952 327724 4004
rect 327776 3992 327782 4004
rect 351638 3992 351644 4004
rect 327776 3964 351644 3992
rect 327776 3952 327782 3964
rect 351638 3952 351644 3964
rect 351696 3952 351702 4004
rect 360838 3952 360844 4004
rect 360896 3992 360902 4004
rect 369394 3992 369400 4004
rect 360896 3964 369400 3992
rect 360896 3952 360902 3964
rect 369394 3952 369400 3964
rect 369452 3952 369458 4004
rect 377398 3952 377404 4004
rect 377456 3992 377462 4004
rect 387150 3992 387156 4004
rect 377456 3964 387156 3992
rect 377456 3952 377462 3964
rect 387150 3952 387156 3964
rect 387208 3952 387214 4004
rect 52546 3884 52552 3936
rect 52604 3924 52610 3936
rect 88978 3924 88984 3936
rect 52604 3896 88984 3924
rect 52604 3884 52610 3896
rect 88978 3884 88984 3896
rect 89036 3884 89042 3936
rect 92750 3884 92756 3936
rect 92808 3924 92814 3936
rect 97350 3924 97356 3936
rect 92808 3896 97356 3924
rect 92808 3884 92814 3896
rect 97350 3884 97356 3896
rect 97408 3884 97414 3936
rect 103330 3884 103336 3936
rect 103388 3924 103394 3936
rect 184198 3924 184204 3936
rect 103388 3896 184204 3924
rect 103388 3884 103394 3896
rect 184198 3884 184204 3896
rect 184256 3884 184262 3936
rect 200022 3884 200028 3936
rect 200080 3924 200086 3936
rect 207382 3924 207388 3936
rect 200080 3896 207388 3924
rect 200080 3884 200086 3896
rect 207382 3884 207388 3896
rect 207440 3884 207446 3936
rect 214466 3884 214472 3936
rect 214524 3924 214530 3936
rect 231210 3924 231216 3936
rect 214524 3896 231216 3924
rect 214524 3884 214530 3896
rect 231210 3884 231216 3896
rect 231268 3884 231274 3936
rect 257062 3884 257068 3936
rect 257120 3924 257126 3936
rect 269114 3924 269120 3936
rect 257120 3896 269120 3924
rect 257120 3884 257126 3896
rect 269114 3884 269120 3896
rect 269172 3884 269178 3936
rect 271322 3884 271328 3936
rect 271380 3924 271386 3936
rect 281534 3924 281540 3936
rect 271380 3896 281540 3924
rect 271380 3884 271386 3896
rect 281534 3884 281540 3896
rect 281592 3884 281598 3936
rect 304258 3884 304264 3936
rect 304316 3924 304322 3936
rect 371694 3924 371700 3936
rect 304316 3896 371700 3924
rect 304316 3884 304322 3896
rect 371694 3884 371700 3896
rect 371752 3884 371758 3936
rect 385678 3884 385684 3936
rect 385736 3924 385742 3936
rect 447410 3924 447416 3936
rect 385736 3896 447416 3924
rect 385736 3884 385742 3896
rect 447410 3884 447416 3896
rect 447468 3884 447474 3936
rect 475470 3884 475476 3936
rect 475528 3924 475534 3936
rect 487614 3924 487620 3936
rect 475528 3896 487620 3924
rect 475528 3884 475534 3896
rect 487614 3884 487620 3896
rect 487672 3884 487678 3936
rect 40678 3856 40684 3868
rect 26206 3828 40684 3856
rect 40678 3816 40684 3828
rect 40736 3816 40742 3868
rect 60826 3816 60832 3868
rect 60884 3856 60890 3868
rect 106918 3856 106924 3868
rect 60884 3828 106924 3856
rect 60884 3816 60890 3828
rect 106918 3816 106924 3828
rect 106976 3816 106982 3868
rect 140038 3816 140044 3868
rect 140096 3856 140102 3868
rect 223850 3856 223856 3868
rect 140096 3828 223856 3856
rect 140096 3816 140102 3828
rect 223850 3816 223856 3828
rect 223908 3816 223914 3868
rect 225138 3816 225144 3868
rect 225196 3856 225202 3868
rect 234798 3856 234804 3868
rect 225196 3828 234804 3856
rect 225196 3816 225202 3828
rect 234798 3816 234804 3828
rect 234856 3816 234862 3868
rect 260098 3816 260104 3868
rect 260156 3856 260162 3868
rect 273622 3856 273628 3868
rect 260156 3828 273628 3856
rect 260156 3816 260162 3828
rect 273622 3816 273628 3828
rect 273680 3816 273686 3868
rect 278130 3816 278136 3868
rect 278188 3856 278194 3868
rect 288986 3856 288992 3868
rect 278188 3828 288992 3856
rect 278188 3816 278194 3828
rect 288986 3816 288992 3828
rect 289044 3816 289050 3868
rect 292574 3856 292580 3868
rect 289832 3828 292580 3856
rect 29638 3788 29644 3800
rect 25700 3760 29644 3788
rect 29638 3748 29644 3760
rect 29696 3748 29702 3800
rect 39574 3748 39580 3800
rect 39632 3788 39638 3800
rect 58618 3788 58624 3800
rect 39632 3760 58624 3788
rect 39632 3748 39638 3760
rect 58618 3748 58624 3760
rect 58676 3748 58682 3800
rect 74994 3748 75000 3800
rect 75052 3788 75058 3800
rect 124858 3788 124864 3800
rect 75052 3760 124864 3788
rect 75052 3748 75058 3760
rect 124858 3748 124864 3760
rect 124916 3748 124922 3800
rect 150618 3748 150624 3800
rect 150676 3788 150682 3800
rect 152642 3788 152648 3800
rect 150676 3760 152648 3788
rect 150676 3748 150682 3760
rect 152642 3748 152648 3760
rect 152700 3748 152706 3800
rect 172146 3748 172152 3800
rect 172204 3788 172210 3800
rect 182818 3788 182824 3800
rect 172204 3760 182824 3788
rect 172204 3748 172210 3760
rect 182818 3748 182824 3760
rect 182876 3748 182882 3800
rect 221550 3748 221556 3800
rect 221608 3788 221614 3800
rect 234154 3788 234160 3800
rect 221608 3760 234160 3788
rect 221608 3748 221614 3760
rect 234154 3748 234160 3760
rect 234212 3748 234218 3800
rect 245194 3748 245200 3800
rect 245252 3788 245258 3800
rect 252646 3788 252652 3800
rect 245252 3760 252652 3788
rect 245252 3748 245258 3760
rect 252646 3748 252652 3760
rect 252704 3748 252710 3800
rect 253198 3748 253204 3800
rect 253256 3788 253262 3800
rect 289832 3788 289860 3828
rect 292574 3816 292580 3828
rect 292632 3816 292638 3868
rect 311158 3816 311164 3868
rect 311216 3856 311222 3868
rect 383562 3856 383568 3868
rect 311216 3828 383568 3856
rect 311216 3816 311222 3828
rect 383562 3816 383568 3828
rect 383620 3816 383626 3868
rect 411898 3816 411904 3868
rect 411956 3856 411962 3868
rect 491110 3856 491116 3868
rect 411956 3828 491116 3856
rect 411956 3816 411962 3828
rect 491110 3816 491116 3828
rect 491168 3816 491174 3868
rect 518158 3816 518164 3868
rect 518216 3856 518222 3868
rect 520734 3856 520740 3868
rect 518216 3828 520740 3856
rect 518216 3816 518222 3828
rect 520734 3816 520740 3828
rect 520792 3816 520798 3868
rect 536098 3816 536104 3868
rect 536156 3856 536162 3868
rect 538398 3856 538404 3868
rect 536156 3828 538404 3856
rect 536156 3816 536162 3828
rect 538398 3816 538404 3828
rect 538456 3816 538462 3868
rect 253256 3760 289860 3788
rect 253256 3748 253262 3760
rect 290182 3748 290188 3800
rect 290240 3788 290246 3800
rect 291286 3788 291292 3800
rect 290240 3760 291292 3788
rect 290240 3748 290246 3760
rect 291286 3748 291292 3760
rect 291344 3748 291350 3800
rect 296070 3748 296076 3800
rect 296128 3788 296134 3800
rect 299566 3788 299572 3800
rect 296128 3760 299572 3788
rect 296128 3748 296134 3760
rect 299566 3748 299572 3760
rect 299624 3748 299630 3800
rect 322198 3748 322204 3800
rect 322256 3788 322262 3800
rect 415486 3788 415492 3800
rect 322256 3760 415492 3788
rect 322256 3748 322262 3760
rect 415486 3748 415492 3760
rect 415544 3748 415550 3800
rect 429838 3748 429844 3800
rect 429896 3788 429902 3800
rect 463970 3788 463976 3800
rect 429896 3760 463976 3788
rect 429896 3748 429902 3760
rect 463970 3748 463976 3760
rect 464028 3748 464034 3800
rect 465718 3748 465724 3800
rect 465776 3788 465782 3800
rect 498194 3788 498200 3800
rect 465776 3760 498200 3788
rect 465776 3748 465782 3760
rect 498194 3748 498200 3760
rect 498252 3748 498258 3800
rect 538186 3760 547874 3788
rect 14734 3680 14740 3732
rect 14792 3720 14798 3732
rect 43438 3720 43444 3732
rect 14792 3692 43444 3720
rect 14792 3680 14798 3692
rect 43438 3680 43444 3692
rect 43496 3680 43502 3732
rect 62022 3680 62028 3732
rect 62080 3720 62086 3732
rect 71038 3720 71044 3732
rect 62080 3692 71044 3720
rect 62080 3680 62086 3692
rect 71038 3680 71044 3692
rect 71096 3680 71102 3732
rect 82078 3680 82084 3732
rect 82136 3720 82142 3732
rect 191098 3720 191104 3732
rect 82136 3692 191104 3720
rect 82136 3680 82142 3692
rect 191098 3680 191104 3692
rect 191156 3680 191162 3732
rect 215662 3680 215668 3732
rect 215720 3720 215726 3732
rect 232590 3720 232596 3732
rect 215720 3692 232596 3720
rect 215720 3680 215726 3692
rect 232590 3680 232596 3692
rect 232648 3680 232654 3732
rect 251082 3680 251088 3732
rect 251140 3720 251146 3732
rect 262950 3720 262956 3732
rect 251140 3692 262956 3720
rect 251140 3680 251146 3692
rect 262950 3680 262956 3692
rect 263008 3680 263014 3732
rect 264882 3680 264888 3732
rect 264940 3720 264946 3732
rect 374086 3720 374092 3732
rect 264940 3692 374092 3720
rect 264940 3680 264946 3692
rect 374086 3680 374092 3692
rect 374144 3680 374150 3732
rect 381538 3680 381544 3732
rect 381596 3720 381602 3732
rect 397730 3720 397736 3732
rect 381596 3692 397736 3720
rect 381596 3680 381602 3692
rect 397730 3680 397736 3692
rect 397788 3680 397794 3732
rect 421558 3680 421564 3732
rect 421616 3720 421622 3732
rect 427262 3720 427268 3732
rect 421616 3692 427268 3720
rect 421616 3680 421622 3692
rect 427262 3680 427268 3692
rect 427320 3680 427326 3732
rect 428458 3680 428464 3732
rect 428516 3720 428522 3732
rect 534902 3720 534908 3732
rect 428516 3692 534908 3720
rect 428516 3680 428522 3692
rect 534902 3680 534908 3692
rect 534960 3680 534966 3732
rect 21818 3612 21824 3664
rect 21876 3652 21882 3664
rect 39298 3652 39304 3664
rect 21876 3624 39304 3652
rect 21876 3612 21882 3624
rect 39298 3612 39304 3624
rect 39356 3612 39362 3664
rect 41874 3612 41880 3664
rect 41932 3652 41938 3664
rect 207290 3652 207296 3664
rect 41932 3624 207296 3652
rect 41932 3612 41938 3624
rect 207290 3612 207296 3624
rect 207348 3612 207354 3664
rect 213362 3612 213368 3664
rect 213420 3652 213426 3664
rect 231302 3652 231308 3664
rect 213420 3624 231308 3652
rect 213420 3612 213426 3624
rect 231302 3612 231308 3624
rect 231360 3612 231366 3664
rect 249978 3612 249984 3664
rect 250036 3652 250042 3664
rect 260834 3652 260840 3664
rect 250036 3624 260840 3652
rect 250036 3612 250042 3624
rect 260834 3612 260840 3624
rect 260892 3612 260898 3664
rect 261754 3612 261760 3664
rect 261812 3652 261818 3664
rect 266446 3652 266452 3664
rect 261812 3624 266452 3652
rect 261812 3612 261818 3624
rect 266446 3612 266452 3624
rect 266504 3612 266510 3664
rect 274542 3612 274548 3664
rect 274600 3652 274606 3664
rect 433242 3652 433248 3664
rect 274600 3624 433248 3652
rect 274600 3612 274606 3624
rect 433242 3612 433248 3624
rect 433300 3612 433306 3664
rect 447778 3612 447784 3664
rect 447836 3652 447842 3664
rect 458082 3652 458088 3664
rect 447836 3624 458088 3652
rect 447836 3612 447842 3624
rect 458082 3612 458088 3624
rect 458140 3612 458146 3664
rect 458818 3612 458824 3664
rect 458876 3652 458882 3664
rect 538186 3652 538214 3760
rect 458876 3624 538214 3652
rect 458876 3612 458882 3624
rect 538858 3612 538864 3664
rect 538916 3652 538922 3664
rect 547846 3652 547874 3760
rect 572714 3652 572720 3664
rect 538916 3624 540928 3652
rect 547846 3624 572720 3652
rect 538916 3612 538922 3624
rect 2924 3556 14688 3584
rect 2924 3544 2930 3556
rect 25314 3544 25320 3596
rect 25372 3584 25378 3596
rect 26142 3584 26148 3596
rect 25372 3556 26148 3584
rect 25372 3544 25378 3556
rect 26142 3544 26148 3556
rect 26200 3544 26206 3596
rect 26510 3544 26516 3596
rect 26568 3584 26574 3596
rect 27522 3584 27528 3596
rect 26568 3556 27528 3584
rect 26568 3544 26574 3556
rect 27522 3544 27528 3556
rect 27580 3544 27586 3596
rect 32398 3544 32404 3596
rect 32456 3584 32462 3596
rect 33042 3584 33048 3596
rect 32456 3556 33048 3584
rect 32456 3544 32462 3556
rect 33042 3544 33048 3556
rect 33100 3544 33106 3596
rect 33594 3544 33600 3596
rect 33652 3584 33658 3596
rect 34422 3584 34428 3596
rect 33652 3556 34428 3584
rect 33652 3544 33658 3556
rect 34422 3544 34428 3556
rect 34480 3544 34486 3596
rect 34790 3544 34796 3596
rect 34848 3584 34854 3596
rect 35802 3584 35808 3596
rect 34848 3556 35808 3584
rect 34848 3544 34854 3556
rect 35802 3544 35808 3556
rect 35860 3544 35866 3596
rect 35986 3544 35992 3596
rect 36044 3584 36050 3596
rect 37090 3584 37096 3596
rect 36044 3556 37096 3584
rect 36044 3544 36050 3556
rect 37090 3544 37096 3556
rect 37148 3544 37154 3596
rect 38378 3544 38384 3596
rect 38436 3584 38442 3596
rect 39390 3584 39396 3596
rect 38436 3556 39396 3584
rect 38436 3544 38442 3556
rect 39390 3544 39396 3556
rect 39448 3544 39454 3596
rect 40678 3544 40684 3596
rect 40736 3584 40742 3596
rect 41322 3584 41328 3596
rect 40736 3556 41328 3584
rect 40736 3544 40742 3556
rect 41322 3544 41328 3556
rect 41380 3544 41386 3596
rect 43070 3544 43076 3596
rect 43128 3584 43134 3596
rect 44082 3584 44088 3596
rect 43128 3556 44088 3584
rect 43128 3544 43134 3556
rect 44082 3544 44088 3556
rect 44140 3544 44146 3596
rect 44266 3544 44272 3596
rect 44324 3584 44330 3596
rect 45370 3584 45376 3596
rect 44324 3556 45376 3584
rect 44324 3544 44330 3556
rect 45370 3544 45376 3556
rect 45428 3544 45434 3596
rect 50154 3544 50160 3596
rect 50212 3584 50218 3596
rect 50982 3584 50988 3596
rect 50212 3556 50988 3584
rect 50212 3544 50218 3556
rect 50982 3544 50988 3556
rect 51040 3544 51046 3596
rect 51350 3544 51356 3596
rect 51408 3584 51414 3596
rect 54478 3584 54484 3596
rect 51408 3556 54484 3584
rect 51408 3544 51414 3556
rect 54478 3544 54484 3556
rect 54536 3544 54542 3596
rect 56042 3544 56048 3596
rect 56100 3584 56106 3596
rect 56502 3584 56508 3596
rect 56100 3556 56508 3584
rect 56100 3544 56106 3556
rect 56502 3544 56508 3556
rect 56560 3544 56566 3596
rect 57238 3544 57244 3596
rect 57296 3584 57302 3596
rect 57882 3584 57888 3596
rect 57296 3556 57888 3584
rect 57296 3544 57302 3556
rect 57882 3544 57888 3556
rect 57940 3544 57946 3596
rect 59630 3544 59636 3596
rect 59688 3584 59694 3596
rect 61470 3584 61476 3596
rect 59688 3556 61476 3584
rect 59688 3544 59694 3556
rect 61470 3544 61476 3556
rect 61528 3544 61534 3596
rect 64322 3544 64328 3596
rect 64380 3584 64386 3596
rect 64782 3584 64788 3596
rect 64380 3556 64788 3584
rect 64380 3544 64386 3556
rect 64782 3544 64788 3556
rect 64840 3544 64846 3596
rect 67910 3544 67916 3596
rect 67968 3584 67974 3596
rect 68922 3584 68928 3596
rect 67968 3556 68928 3584
rect 67968 3544 67974 3556
rect 68922 3544 68928 3556
rect 68980 3544 68986 3596
rect 69106 3544 69112 3596
rect 69164 3584 69170 3596
rect 70302 3584 70308 3596
rect 69164 3556 70308 3584
rect 69164 3544 69170 3556
rect 70302 3544 70308 3556
rect 70360 3544 70366 3596
rect 79686 3544 79692 3596
rect 79744 3584 79750 3596
rect 80698 3584 80704 3596
rect 79744 3556 80704 3584
rect 79744 3544 79750 3556
rect 80698 3544 80704 3556
rect 80756 3544 80762 3596
rect 80882 3544 80888 3596
rect 80940 3584 80946 3596
rect 81342 3584 81348 3596
rect 80940 3556 81348 3584
rect 80940 3544 80946 3556
rect 81342 3544 81348 3556
rect 81400 3544 81406 3596
rect 83274 3544 83280 3596
rect 83332 3584 83338 3596
rect 84102 3584 84108 3596
rect 83332 3556 84108 3584
rect 83332 3544 83338 3556
rect 84102 3544 84108 3556
rect 84160 3544 84166 3596
rect 84470 3544 84476 3596
rect 84528 3584 84534 3596
rect 86218 3584 86224 3596
rect 84528 3556 86224 3584
rect 84528 3544 84534 3556
rect 86218 3544 86224 3556
rect 86276 3544 86282 3596
rect 90358 3544 90364 3596
rect 90416 3584 90422 3596
rect 91002 3584 91008 3596
rect 90416 3556 91008 3584
rect 90416 3544 90422 3556
rect 91002 3544 91008 3556
rect 91060 3544 91066 3596
rect 91554 3544 91560 3596
rect 91612 3584 91618 3596
rect 93854 3584 93860 3596
rect 91612 3556 93860 3584
rect 91612 3544 91618 3556
rect 93854 3544 93860 3556
rect 93912 3544 93918 3596
rect 93946 3544 93952 3596
rect 94004 3584 94010 3596
rect 95050 3584 95056 3596
rect 94004 3556 95056 3584
rect 94004 3544 94010 3556
rect 95050 3544 95056 3556
rect 95108 3544 95114 3596
rect 97442 3544 97448 3596
rect 97500 3584 97506 3596
rect 98638 3584 98644 3596
rect 97500 3556 98644 3584
rect 97500 3544 97506 3556
rect 98638 3544 98644 3556
rect 98696 3544 98702 3596
rect 101030 3544 101036 3596
rect 101088 3584 101094 3596
rect 102042 3584 102048 3596
rect 101088 3556 102048 3584
rect 101088 3544 101094 3556
rect 102042 3544 102048 3556
rect 102100 3544 102106 3596
rect 105722 3544 105728 3596
rect 105780 3584 105786 3596
rect 106182 3584 106188 3596
rect 105780 3556 106188 3584
rect 105780 3544 105786 3556
rect 106182 3544 106188 3556
rect 106240 3544 106246 3596
rect 109310 3544 109316 3596
rect 109368 3584 109374 3596
rect 111150 3584 111156 3596
rect 109368 3556 111156 3584
rect 109368 3544 109374 3556
rect 111150 3544 111156 3556
rect 111208 3544 111214 3596
rect 114002 3544 114008 3596
rect 114060 3584 114066 3596
rect 114462 3584 114468 3596
rect 114060 3556 114468 3584
rect 114060 3544 114066 3556
rect 114462 3544 114468 3556
rect 114520 3544 114526 3596
rect 115198 3544 115204 3596
rect 115256 3584 115262 3596
rect 116578 3584 116584 3596
rect 115256 3556 116584 3584
rect 115256 3544 115262 3556
rect 116578 3544 116584 3556
rect 116636 3544 116642 3596
rect 122282 3544 122288 3596
rect 122340 3584 122346 3596
rect 122742 3584 122748 3596
rect 122340 3556 122748 3584
rect 122340 3544 122346 3556
rect 122742 3544 122748 3556
rect 122800 3544 122806 3596
rect 123478 3544 123484 3596
rect 123536 3584 123542 3596
rect 124122 3584 124128 3596
rect 123536 3556 124128 3584
rect 123536 3544 123542 3556
rect 124122 3544 124128 3556
rect 124180 3544 124186 3596
rect 125870 3544 125876 3596
rect 125928 3584 125934 3596
rect 126882 3584 126888 3596
rect 125928 3556 126888 3584
rect 125928 3544 125934 3556
rect 126882 3544 126888 3556
rect 126940 3544 126946 3596
rect 129366 3544 129372 3596
rect 129424 3584 129430 3596
rect 130378 3584 130384 3596
rect 129424 3556 130384 3584
rect 129424 3544 129430 3556
rect 130378 3544 130384 3556
rect 130436 3544 130442 3596
rect 132954 3544 132960 3596
rect 133012 3584 133018 3596
rect 133782 3584 133788 3596
rect 133012 3556 133788 3584
rect 133012 3544 133018 3556
rect 133782 3544 133788 3556
rect 133840 3544 133846 3596
rect 134150 3544 134156 3596
rect 134208 3584 134214 3596
rect 135162 3584 135168 3596
rect 134208 3556 135168 3584
rect 134208 3544 134214 3556
rect 135162 3544 135168 3556
rect 135220 3544 135226 3596
rect 136450 3544 136456 3596
rect 136508 3584 136514 3596
rect 137278 3584 137284 3596
rect 136508 3556 137284 3584
rect 136508 3544 136514 3556
rect 137278 3544 137284 3556
rect 137336 3544 137342 3596
rect 138842 3544 138848 3596
rect 138900 3584 138906 3596
rect 139302 3584 139308 3596
rect 138900 3556 139308 3584
rect 138900 3544 138906 3556
rect 139302 3544 139308 3556
rect 139360 3544 139366 3596
rect 141234 3544 141240 3596
rect 141292 3584 141298 3596
rect 142062 3584 142068 3596
rect 141292 3556 142068 3584
rect 141292 3544 141298 3556
rect 142062 3544 142068 3556
rect 142120 3544 142126 3596
rect 142430 3544 142436 3596
rect 142488 3584 142494 3596
rect 143442 3584 143448 3596
rect 142488 3556 143448 3584
rect 142488 3544 142494 3556
rect 143442 3544 143448 3556
rect 143500 3544 143506 3596
rect 147122 3544 147128 3596
rect 147180 3584 147186 3596
rect 147582 3584 147588 3596
rect 147180 3556 147588 3584
rect 147180 3544 147186 3556
rect 147582 3544 147588 3556
rect 147640 3544 147646 3596
rect 157794 3544 157800 3596
rect 157852 3584 157858 3596
rect 158622 3584 158628 3596
rect 157852 3556 158628 3584
rect 157852 3544 157858 3556
rect 158622 3544 158628 3556
rect 158680 3544 158686 3596
rect 158898 3544 158904 3596
rect 158956 3584 158962 3596
rect 160002 3584 160008 3596
rect 158956 3556 160008 3584
rect 158956 3544 158962 3556
rect 160002 3544 160008 3556
rect 160060 3544 160066 3596
rect 163682 3544 163688 3596
rect 163740 3584 163746 3596
rect 164142 3584 164148 3596
rect 163740 3556 164148 3584
rect 163740 3544 163746 3556
rect 164142 3544 164148 3556
rect 164200 3544 164206 3596
rect 164878 3544 164884 3596
rect 164936 3584 164942 3596
rect 165522 3584 165528 3596
rect 164936 3556 165528 3584
rect 164936 3544 164942 3556
rect 165522 3544 165528 3556
rect 165580 3544 165586 3596
rect 166074 3544 166080 3596
rect 166132 3584 166138 3596
rect 166902 3584 166908 3596
rect 166132 3556 166908 3584
rect 166132 3544 166138 3556
rect 166902 3544 166908 3556
rect 166960 3544 166966 3596
rect 167178 3544 167184 3596
rect 167236 3584 167242 3596
rect 169018 3584 169024 3596
rect 167236 3556 169024 3584
rect 167236 3544 167242 3556
rect 169018 3544 169024 3556
rect 169076 3544 169082 3596
rect 169570 3544 169576 3596
rect 169628 3584 169634 3596
rect 170398 3584 170404 3596
rect 169628 3556 170404 3584
rect 169628 3544 169634 3556
rect 170398 3544 170404 3556
rect 170456 3544 170462 3596
rect 171962 3544 171968 3596
rect 172020 3584 172026 3596
rect 173158 3584 173164 3596
rect 172020 3556 173164 3584
rect 172020 3544 172026 3556
rect 173158 3544 173164 3556
rect 173216 3544 173222 3596
rect 175458 3544 175464 3596
rect 175516 3584 175522 3596
rect 176562 3584 176568 3596
rect 175516 3556 176568 3584
rect 175516 3544 175522 3556
rect 176562 3544 176568 3556
rect 176620 3544 176626 3596
rect 176654 3544 176660 3596
rect 176712 3584 176718 3596
rect 177942 3584 177948 3596
rect 176712 3556 177948 3584
rect 176712 3544 176718 3556
rect 177942 3544 177948 3556
rect 178000 3544 178006 3596
rect 180242 3544 180248 3596
rect 180300 3584 180306 3596
rect 180702 3584 180708 3596
rect 180300 3556 180708 3584
rect 180300 3544 180306 3556
rect 180702 3544 180708 3556
rect 180760 3544 180766 3596
rect 181438 3544 181444 3596
rect 181496 3584 181502 3596
rect 182082 3584 182088 3596
rect 181496 3556 182088 3584
rect 181496 3544 181502 3556
rect 182082 3544 182088 3556
rect 182140 3544 182146 3596
rect 182542 3544 182548 3596
rect 182600 3584 182606 3596
rect 183462 3584 183468 3596
rect 182600 3556 183468 3584
rect 182600 3544 182606 3556
rect 183462 3544 183468 3556
rect 183520 3544 183526 3596
rect 183738 3544 183744 3596
rect 183796 3584 183802 3596
rect 184842 3584 184848 3596
rect 183796 3556 184848 3584
rect 183796 3544 183802 3556
rect 184842 3544 184848 3556
rect 184900 3544 184906 3596
rect 186130 3544 186136 3596
rect 186188 3584 186194 3596
rect 186958 3584 186964 3596
rect 186188 3556 186964 3584
rect 186188 3544 186194 3556
rect 186958 3544 186964 3556
rect 187016 3544 187022 3596
rect 187326 3544 187332 3596
rect 187384 3584 187390 3596
rect 188338 3584 188344 3596
rect 187384 3556 188344 3584
rect 187384 3544 187390 3556
rect 188338 3544 188344 3556
rect 188396 3544 188402 3596
rect 188522 3544 188528 3596
rect 188580 3584 188586 3596
rect 188982 3584 188988 3596
rect 188580 3556 188988 3584
rect 188580 3544 188586 3556
rect 188982 3544 188988 3556
rect 189040 3544 189046 3596
rect 192018 3544 192024 3596
rect 192076 3584 192082 3596
rect 193122 3584 193128 3596
rect 192076 3556 193128 3584
rect 192076 3544 192082 3556
rect 193122 3544 193128 3556
rect 193180 3544 193186 3596
rect 193214 3544 193220 3596
rect 193272 3584 193278 3596
rect 195238 3584 195244 3596
rect 193272 3556 195244 3584
rect 193272 3544 193278 3556
rect 195238 3544 195244 3556
rect 195296 3544 195302 3596
rect 197170 3544 197176 3596
rect 197228 3584 197234 3596
rect 197906 3584 197912 3596
rect 197228 3556 197912 3584
rect 197228 3544 197234 3556
rect 197906 3544 197912 3556
rect 197964 3544 197970 3596
rect 200390 3584 200396 3596
rect 200086 3556 200396 3584
rect 566 3476 572 3528
rect 624 3516 630 3528
rect 1302 3516 1308 3528
rect 624 3488 1308 3516
rect 624 3476 630 3488
rect 1302 3476 1308 3488
rect 1360 3476 1366 3528
rect 9950 3476 9956 3528
rect 10008 3516 10014 3528
rect 10962 3516 10968 3528
rect 10008 3488 10968 3516
rect 10008 3476 10014 3488
rect 10962 3476 10968 3488
rect 11020 3476 11026 3528
rect 200086 3516 200114 3556
rect 200390 3544 200396 3556
rect 200448 3544 200454 3596
rect 205082 3544 205088 3596
rect 205140 3584 205146 3596
rect 225322 3584 225328 3596
rect 205140 3556 225328 3584
rect 205140 3544 205146 3556
rect 225322 3544 225328 3556
rect 225380 3544 225386 3596
rect 226334 3544 226340 3596
rect 226392 3584 226398 3596
rect 227622 3584 227628 3596
rect 226392 3556 227628 3584
rect 226392 3544 226398 3556
rect 227622 3544 227628 3556
rect 227680 3544 227686 3596
rect 234062 3584 234068 3596
rect 229066 3556 234068 3584
rect 11164 3488 200114 3516
rect 1670 3408 1676 3460
rect 1728 3448 1734 3460
rect 1728 3420 6914 3448
rect 1728 3408 1734 3420
rect 6886 3312 6914 3420
rect 7650 3340 7656 3392
rect 7708 3380 7714 3392
rect 11164 3380 11192 3488
rect 200298 3476 200304 3528
rect 200356 3516 200362 3528
rect 202138 3516 202144 3528
rect 200356 3488 202144 3516
rect 200356 3476 200362 3488
rect 202138 3476 202144 3488
rect 202196 3476 202202 3528
rect 208578 3476 208584 3528
rect 208636 3516 208642 3528
rect 229066 3516 229094 3556
rect 234062 3544 234068 3556
rect 234120 3544 234126 3596
rect 252094 3544 252100 3596
rect 252152 3584 252158 3596
rect 299382 3584 299388 3596
rect 252152 3556 299388 3584
rect 252152 3544 252158 3556
rect 299382 3544 299388 3556
rect 299440 3544 299446 3596
rect 299474 3544 299480 3596
rect 299532 3584 299538 3596
rect 300762 3584 300768 3596
rect 299532 3556 300768 3584
rect 299532 3544 299538 3556
rect 300762 3544 300768 3556
rect 300820 3544 300826 3596
rect 307018 3544 307024 3596
rect 307076 3584 307082 3596
rect 307938 3584 307944 3596
rect 307076 3556 307944 3584
rect 307076 3544 307082 3556
rect 307938 3544 307944 3556
rect 307996 3544 308002 3596
rect 309134 3544 309140 3596
rect 309192 3584 309198 3596
rect 310238 3584 310244 3596
rect 309192 3556 310244 3584
rect 309192 3544 309198 3556
rect 310238 3544 310244 3556
rect 310296 3544 310302 3596
rect 312538 3544 312544 3596
rect 312596 3584 312602 3596
rect 313826 3584 313832 3596
rect 312596 3556 313832 3584
rect 312596 3544 312602 3556
rect 313826 3544 313832 3556
rect 313884 3544 313890 3596
rect 314010 3544 314016 3596
rect 314068 3584 314074 3596
rect 315022 3584 315028 3596
rect 314068 3556 315028 3584
rect 314068 3544 314074 3556
rect 315022 3544 315028 3556
rect 315080 3544 315086 3596
rect 316678 3544 316684 3596
rect 316736 3584 316742 3596
rect 485222 3584 485228 3596
rect 316736 3556 485228 3584
rect 316736 3544 316742 3556
rect 485222 3544 485228 3556
rect 485280 3544 485286 3596
rect 485332 3556 488948 3584
rect 208636 3488 229094 3516
rect 208636 3476 208642 3488
rect 232222 3476 232228 3528
rect 232280 3516 232286 3528
rect 233142 3516 233148 3528
rect 232280 3488 233148 3516
rect 232280 3476 232286 3488
rect 233142 3476 233148 3488
rect 233200 3476 233206 3528
rect 238662 3476 238668 3528
rect 238720 3516 238726 3528
rect 244090 3516 244096 3528
rect 238720 3488 244096 3516
rect 238720 3476 238726 3488
rect 244090 3476 244096 3488
rect 244148 3476 244154 3528
rect 246482 3476 246488 3528
rect 246540 3516 246546 3528
rect 246540 3488 268240 3516
rect 246540 3476 246546 3488
rect 200206 3448 200212 3460
rect 7708 3352 11192 3380
rect 12406 3420 200212 3448
rect 7708 3340 7714 3352
rect 12406 3312 12434 3420
rect 200206 3408 200212 3420
rect 200264 3408 200270 3460
rect 206186 3408 206192 3460
rect 206244 3448 206250 3460
rect 234890 3448 234896 3460
rect 206244 3420 234896 3448
rect 206244 3408 206250 3420
rect 234890 3408 234896 3420
rect 234948 3408 234954 3460
rect 238110 3408 238116 3460
rect 238168 3448 238174 3460
rect 251266 3448 251272 3460
rect 238168 3420 251272 3448
rect 238168 3408 238174 3420
rect 251266 3408 251272 3420
rect 251324 3408 251330 3460
rect 254854 3408 254860 3460
rect 254912 3448 254918 3460
rect 254912 3420 258074 3448
rect 254912 3408 254918 3420
rect 66714 3340 66720 3392
rect 66772 3380 66778 3392
rect 68278 3380 68284 3392
rect 66772 3352 68284 3380
rect 66772 3340 66778 3352
rect 68278 3340 68284 3352
rect 68336 3340 68342 3392
rect 85666 3340 85672 3392
rect 85724 3380 85730 3392
rect 89070 3380 89076 3392
rect 85724 3352 89076 3380
rect 85724 3340 85730 3352
rect 89070 3340 89076 3352
rect 89128 3340 89134 3392
rect 89162 3340 89168 3392
rect 89220 3380 89226 3392
rect 91554 3380 91560 3392
rect 89220 3352 91560 3380
rect 89220 3340 89226 3352
rect 91554 3340 91560 3352
rect 91612 3340 91618 3392
rect 96246 3340 96252 3392
rect 96304 3380 96310 3392
rect 97258 3380 97264 3392
rect 96304 3352 97264 3380
rect 96304 3340 96310 3352
rect 97258 3340 97264 3352
rect 97316 3340 97322 3392
rect 110506 3340 110512 3392
rect 110564 3380 110570 3392
rect 112438 3380 112444 3392
rect 110564 3352 112444 3380
rect 110564 3340 110570 3352
rect 112438 3340 112444 3352
rect 112496 3340 112502 3392
rect 135254 3340 135260 3392
rect 135312 3380 135318 3392
rect 137370 3380 137376 3392
rect 135312 3352 137376 3380
rect 135312 3340 135318 3352
rect 137370 3340 137376 3352
rect 137428 3340 137434 3392
rect 156598 3340 156604 3392
rect 156656 3380 156662 3392
rect 158070 3380 158076 3392
rect 156656 3352 158076 3380
rect 156656 3340 156662 3352
rect 158070 3340 158076 3352
rect 158128 3340 158134 3392
rect 168374 3340 168380 3392
rect 168432 3380 168438 3392
rect 169662 3380 169668 3392
rect 168432 3352 169668 3380
rect 168432 3340 168438 3352
rect 169662 3340 169668 3352
rect 169720 3340 169726 3392
rect 173158 3340 173164 3392
rect 173216 3380 173222 3392
rect 174538 3380 174544 3392
rect 173216 3352 174544 3380
rect 173216 3340 173222 3352
rect 174538 3340 174544 3352
rect 174596 3340 174602 3392
rect 184934 3340 184940 3392
rect 184992 3380 184998 3392
rect 187050 3380 187056 3392
rect 184992 3352 187056 3380
rect 184992 3340 184998 3352
rect 187050 3340 187056 3352
rect 187108 3340 187114 3392
rect 190822 3340 190828 3392
rect 190880 3380 190886 3392
rect 192478 3380 192484 3392
rect 190880 3352 192484 3380
rect 190880 3340 190886 3352
rect 192478 3340 192484 3352
rect 192536 3340 192542 3392
rect 196802 3340 196808 3392
rect 196860 3380 196866 3392
rect 197262 3380 197268 3392
rect 196860 3352 197268 3380
rect 196860 3340 196866 3352
rect 197262 3340 197268 3352
rect 197320 3340 197326 3392
rect 210970 3340 210976 3392
rect 211028 3380 211034 3392
rect 213178 3380 213184 3392
rect 211028 3352 213184 3380
rect 211028 3340 211034 3352
rect 213178 3340 213184 3352
rect 213236 3340 213242 3392
rect 216858 3340 216864 3392
rect 216916 3380 216922 3392
rect 217962 3380 217968 3392
rect 216916 3352 217968 3380
rect 216916 3340 216922 3352
rect 217962 3340 217968 3352
rect 218020 3340 218026 3392
rect 218054 3340 218060 3392
rect 218112 3380 218118 3392
rect 219342 3380 219348 3392
rect 218112 3352 219348 3380
rect 218112 3340 218118 3352
rect 219342 3340 219348 3352
rect 219400 3340 219406 3392
rect 6886 3284 12434 3312
rect 65518 3272 65524 3324
rect 65576 3312 65582 3324
rect 72418 3312 72424 3324
rect 65576 3284 72424 3312
rect 65576 3272 65582 3284
rect 72418 3272 72424 3284
rect 72476 3272 72482 3324
rect 108114 3272 108120 3324
rect 108172 3312 108178 3324
rect 111058 3312 111064 3324
rect 108172 3284 111064 3312
rect 108172 3272 108178 3284
rect 111058 3272 111064 3284
rect 111116 3272 111122 3324
rect 116394 3272 116400 3324
rect 116452 3312 116458 3324
rect 123386 3312 123392 3324
rect 116452 3284 123392 3312
rect 116452 3272 116458 3284
rect 123386 3272 123392 3284
rect 123444 3272 123450 3324
rect 151814 3272 151820 3324
rect 151872 3312 151878 3324
rect 166258 3312 166264 3324
rect 151872 3284 166264 3312
rect 151872 3272 151878 3284
rect 166258 3272 166264 3284
rect 166316 3272 166322 3324
rect 258046 3312 258074 3420
rect 258718 3408 258724 3460
rect 258776 3448 258782 3460
rect 260650 3448 260656 3460
rect 258776 3420 260656 3448
rect 258776 3408 258782 3420
rect 260650 3408 260656 3420
rect 260708 3408 260714 3460
rect 258258 3340 258264 3392
rect 258316 3380 258322 3392
rect 263686 3380 263692 3392
rect 258316 3352 263692 3380
rect 258316 3340 258322 3352
rect 263686 3340 263692 3352
rect 263744 3340 263750 3392
rect 268212 3380 268240 3488
rect 268378 3476 268384 3528
rect 268436 3516 268442 3528
rect 270034 3516 270040 3528
rect 268436 3488 270040 3516
rect 268436 3476 268442 3488
rect 270034 3476 270040 3488
rect 270092 3476 270098 3528
rect 279786 3476 279792 3528
rect 279844 3516 279850 3528
rect 461578 3516 461584 3528
rect 279844 3488 461584 3516
rect 279844 3476 279850 3488
rect 461578 3476 461584 3488
rect 461636 3476 461642 3528
rect 464338 3476 464344 3528
rect 464396 3516 464402 3528
rect 466270 3516 466276 3528
rect 464396 3488 466276 3516
rect 464396 3476 464402 3488
rect 466270 3476 466276 3488
rect 466328 3476 466334 3528
rect 466380 3488 472572 3516
rect 317322 3448 317328 3460
rect 277366 3420 317328 3448
rect 272426 3380 272432 3392
rect 268212 3352 272432 3380
rect 272426 3340 272432 3352
rect 272484 3340 272490 3392
rect 277366 3312 277394 3420
rect 317322 3408 317328 3420
rect 317380 3408 317386 3460
rect 320818 3408 320824 3460
rect 320876 3448 320882 3460
rect 320876 3420 451274 3448
rect 320876 3408 320882 3420
rect 285398 3340 285404 3392
rect 285456 3380 285462 3392
rect 288434 3380 288440 3392
rect 285456 3352 288440 3380
rect 285456 3340 285462 3352
rect 288434 3340 288440 3352
rect 288492 3340 288498 3392
rect 293678 3340 293684 3392
rect 293736 3380 293742 3392
rect 295334 3380 295340 3392
rect 293736 3352 295340 3380
rect 293736 3340 293742 3352
rect 295334 3340 295340 3352
rect 295392 3340 295398 3392
rect 299382 3340 299388 3392
rect 299440 3380 299446 3392
rect 305546 3380 305552 3392
rect 299440 3352 305552 3380
rect 299440 3340 299446 3352
rect 305546 3340 305552 3352
rect 305604 3340 305610 3392
rect 323578 3340 323584 3392
rect 323636 3380 323642 3392
rect 325602 3380 325608 3392
rect 323636 3352 325608 3380
rect 323636 3340 323642 3352
rect 325602 3340 325608 3352
rect 325660 3340 325666 3392
rect 331858 3340 331864 3392
rect 331916 3380 331922 3392
rect 333882 3380 333888 3392
rect 331916 3352 333888 3380
rect 331916 3340 331922 3352
rect 333882 3340 333888 3352
rect 333940 3340 333946 3392
rect 340874 3340 340880 3392
rect 340932 3380 340938 3392
rect 342162 3380 342168 3392
rect 340932 3352 342168 3380
rect 340932 3340 340938 3352
rect 342162 3340 342168 3352
rect 342220 3340 342226 3392
rect 364978 3340 364984 3392
rect 365036 3380 365042 3392
rect 367002 3380 367008 3392
rect 365036 3352 367008 3380
rect 365036 3340 365042 3352
rect 367002 3340 367008 3352
rect 367060 3340 367066 3392
rect 378778 3340 378784 3392
rect 378836 3380 378842 3392
rect 381170 3380 381176 3392
rect 378836 3352 381176 3380
rect 378836 3340 378842 3352
rect 381170 3340 381176 3352
rect 381228 3340 381234 3392
rect 389818 3340 389824 3392
rect 389876 3380 389882 3392
rect 391842 3380 391848 3392
rect 389876 3352 391848 3380
rect 389876 3340 389882 3352
rect 391842 3340 391848 3352
rect 391900 3340 391906 3392
rect 396718 3340 396724 3392
rect 396776 3380 396782 3392
rect 402514 3380 402520 3392
rect 396776 3352 402520 3380
rect 396776 3340 396782 3352
rect 402514 3340 402520 3352
rect 402572 3340 402578 3392
rect 407758 3340 407764 3392
rect 407816 3380 407822 3392
rect 409598 3380 409604 3392
rect 407816 3352 409604 3380
rect 407816 3340 407822 3352
rect 409598 3340 409604 3352
rect 409656 3340 409662 3392
rect 414658 3340 414664 3392
rect 414716 3380 414722 3392
rect 416682 3380 416688 3392
rect 414716 3352 416688 3380
rect 414716 3340 414722 3352
rect 416682 3340 416688 3352
rect 416740 3340 416746 3392
rect 440234 3340 440240 3392
rect 440292 3380 440298 3392
rect 441522 3380 441528 3392
rect 440292 3352 441528 3380
rect 440292 3340 440298 3352
rect 441522 3340 441528 3352
rect 441580 3340 441586 3392
rect 258046 3284 277394 3312
rect 281902 3272 281908 3324
rect 281960 3312 281966 3324
rect 285766 3312 285772 3324
rect 281960 3284 285772 3312
rect 281960 3272 281966 3284
rect 285766 3272 285772 3284
rect 285824 3272 285830 3324
rect 291838 3272 291844 3324
rect 291896 3312 291902 3324
rect 294874 3312 294880 3324
rect 291896 3284 294880 3312
rect 291896 3272 291902 3284
rect 294874 3272 294880 3284
rect 294932 3272 294938 3324
rect 318150 3272 318156 3324
rect 318208 3312 318214 3324
rect 319714 3312 319720 3324
rect 318208 3284 319720 3312
rect 318208 3272 318214 3284
rect 319714 3272 319720 3284
rect 319772 3272 319778 3324
rect 330478 3272 330484 3324
rect 330536 3312 330542 3324
rect 332686 3312 332692 3324
rect 330536 3284 332692 3312
rect 330536 3272 330542 3284
rect 332686 3272 332692 3284
rect 332744 3272 332750 3324
rect 336090 3272 336096 3324
rect 336148 3312 336154 3324
rect 337470 3312 337476 3324
rect 336148 3284 337476 3312
rect 336148 3272 336154 3284
rect 337470 3272 337476 3284
rect 337528 3272 337534 3324
rect 376110 3272 376116 3324
rect 376168 3312 376174 3324
rect 379974 3312 379980 3324
rect 376168 3284 379980 3312
rect 376168 3272 376174 3284
rect 379974 3272 379980 3284
rect 380032 3272 380038 3324
rect 407206 3272 407212 3324
rect 407264 3312 407270 3324
rect 409966 3312 409972 3324
rect 407264 3284 409972 3312
rect 407264 3272 407270 3284
rect 409966 3272 409972 3284
rect 410024 3272 410030 3324
rect 451246 3312 451274 3420
rect 453298 3408 453304 3460
rect 453356 3448 453362 3460
rect 455690 3448 455696 3460
rect 453356 3420 455696 3448
rect 453356 3408 453362 3420
rect 455690 3408 455696 3420
rect 455748 3408 455754 3460
rect 457438 3408 457444 3460
rect 457496 3448 457502 3460
rect 459186 3448 459192 3460
rect 457496 3420 459192 3448
rect 457496 3408 457502 3420
rect 459186 3408 459192 3420
rect 459244 3408 459250 3460
rect 461670 3340 461676 3392
rect 461728 3380 461734 3392
rect 466380 3380 466408 3488
rect 472544 3380 472572 3488
rect 472618 3476 472624 3528
rect 472676 3516 472682 3528
rect 474550 3516 474556 3528
rect 472676 3488 474556 3516
rect 472676 3476 472682 3488
rect 474550 3476 474556 3488
rect 474608 3476 474614 3528
rect 485038 3476 485044 3528
rect 485096 3516 485102 3528
rect 485332 3516 485360 3556
rect 485096 3488 485360 3516
rect 485096 3476 485102 3488
rect 486418 3476 486424 3528
rect 486476 3516 486482 3528
rect 488810 3516 488816 3528
rect 486476 3488 488816 3516
rect 486476 3476 486482 3488
rect 488810 3476 488816 3488
rect 488868 3476 488874 3528
rect 488920 3516 488948 3556
rect 489178 3544 489184 3596
rect 489236 3584 489242 3596
rect 515030 3584 515036 3596
rect 489236 3556 515036 3584
rect 489236 3544 489242 3556
rect 515030 3544 515036 3556
rect 515088 3544 515094 3596
rect 515398 3544 515404 3596
rect 515456 3584 515462 3596
rect 517146 3584 517152 3596
rect 515456 3556 517152 3584
rect 515456 3544 515462 3556
rect 517146 3544 517152 3556
rect 517204 3544 517210 3596
rect 522298 3544 522304 3596
rect 522356 3584 522362 3596
rect 524230 3584 524236 3596
rect 522356 3556 524236 3584
rect 522356 3544 522362 3556
rect 524230 3544 524236 3556
rect 524288 3544 524294 3596
rect 540790 3584 540796 3596
rect 528526 3556 540796 3584
rect 528526 3516 528554 3556
rect 540790 3544 540796 3556
rect 540848 3544 540854 3596
rect 540900 3584 540928 3624
rect 572714 3612 572720 3624
rect 572772 3612 572778 3664
rect 540900 3556 563192 3584
rect 488920 3488 528554 3516
rect 530578 3476 530584 3528
rect 530636 3516 530642 3528
rect 532510 3516 532516 3528
rect 530636 3488 532516 3516
rect 530636 3476 530642 3488
rect 532510 3476 532516 3488
rect 532568 3476 532574 3528
rect 540238 3476 540244 3528
rect 540296 3516 540302 3528
rect 541986 3516 541992 3528
rect 540296 3488 541992 3516
rect 540296 3476 540302 3488
rect 541986 3476 541992 3488
rect 542044 3476 542050 3528
rect 548518 3476 548524 3528
rect 548576 3516 548582 3528
rect 550266 3516 550272 3528
rect 548576 3488 550272 3516
rect 548576 3476 548582 3488
rect 550266 3476 550272 3488
rect 550324 3476 550330 3528
rect 552658 3476 552664 3528
rect 552716 3516 552722 3528
rect 553394 3516 553400 3528
rect 552716 3488 553400 3516
rect 552716 3476 552722 3488
rect 553394 3476 553400 3488
rect 553452 3476 553458 3528
rect 559742 3476 559748 3528
rect 559800 3516 559806 3528
rect 560478 3516 560484 3528
rect 559800 3488 560484 3516
rect 559800 3476 559806 3488
rect 560478 3476 560484 3488
rect 560536 3476 560542 3528
rect 563164 3516 563192 3556
rect 563238 3544 563244 3596
rect 563296 3584 563302 3596
rect 564526 3584 564532 3596
rect 563296 3556 564532 3584
rect 563296 3544 563302 3556
rect 564526 3544 564532 3556
rect 564584 3544 564590 3596
rect 577406 3544 577412 3596
rect 577464 3584 577470 3596
rect 582742 3584 582748 3596
rect 577464 3556 582748 3584
rect 577464 3544 577470 3556
rect 582742 3544 582748 3556
rect 582800 3544 582806 3596
rect 565630 3516 565636 3528
rect 563164 3488 565636 3516
rect 565630 3476 565636 3488
rect 565688 3476 565694 3528
rect 582190 3476 582196 3528
rect 582248 3516 582254 3528
rect 582926 3516 582932 3528
rect 582248 3488 582932 3516
rect 582248 3476 582254 3488
rect 582926 3476 582932 3488
rect 582984 3476 582990 3528
rect 547874 3448 547880 3460
rect 480226 3420 547880 3448
rect 479334 3380 479340 3392
rect 461728 3352 466408 3380
rect 466472 3352 470594 3380
rect 472544 3352 479340 3380
rect 461728 3340 461734 3352
rect 466472 3312 466500 3352
rect 451246 3284 466500 3312
rect 467190 3272 467196 3324
rect 467248 3312 467254 3324
rect 469858 3312 469864 3324
rect 467248 3284 469864 3312
rect 467248 3272 467254 3284
rect 469858 3272 469864 3284
rect 469916 3272 469922 3324
rect 470566 3312 470594 3352
rect 479334 3340 479340 3352
rect 479392 3340 479398 3392
rect 480226 3312 480254 3420
rect 547874 3408 547880 3420
rect 547932 3408 547938 3460
rect 580994 3408 581000 3460
rect 581052 3448 581058 3460
rect 582834 3448 582840 3460
rect 581052 3420 582840 3448
rect 581052 3408 581058 3420
rect 582834 3408 582840 3420
rect 582892 3408 582898 3460
rect 490558 3340 490564 3392
rect 490616 3380 490622 3392
rect 492306 3380 492312 3392
rect 490616 3352 492312 3380
rect 490616 3340 490622 3352
rect 492306 3340 492312 3352
rect 492364 3340 492370 3392
rect 497458 3340 497464 3392
rect 497516 3380 497522 3392
rect 499390 3380 499396 3392
rect 497516 3352 499396 3380
rect 497516 3340 497522 3352
rect 499390 3340 499396 3352
rect 499448 3340 499454 3392
rect 502978 3340 502984 3392
rect 503036 3380 503042 3392
rect 505370 3380 505376 3392
rect 503036 3352 505376 3380
rect 503036 3340 503042 3352
rect 505370 3340 505376 3352
rect 505428 3340 505434 3392
rect 520918 3340 520924 3392
rect 520976 3380 520982 3392
rect 523034 3380 523040 3392
rect 520976 3352 523040 3380
rect 520976 3340 520982 3352
rect 523034 3340 523040 3352
rect 523092 3340 523098 3392
rect 470566 3284 480254 3312
rect 204622 3244 204628 3256
rect 45526 3216 204628 3244
rect 18230 3136 18236 3188
rect 18288 3176 18294 3188
rect 22738 3176 22744 3188
rect 18288 3148 22744 3176
rect 18288 3136 18294 3148
rect 22738 3136 22744 3148
rect 22796 3136 22802 3188
rect 31294 3068 31300 3120
rect 31352 3108 31358 3120
rect 45526 3108 45554 3216
rect 204622 3204 204628 3216
rect 204680 3204 204686 3256
rect 221182 3244 221188 3256
rect 219406 3216 221188 3244
rect 48958 3136 48964 3188
rect 49016 3176 49022 3188
rect 53098 3176 53104 3188
rect 49016 3148 53104 3176
rect 49016 3136 49022 3148
rect 53098 3136 53104 3148
rect 53156 3136 53162 3188
rect 126974 3136 126980 3188
rect 127032 3176 127038 3188
rect 219406 3176 219434 3216
rect 221182 3204 221188 3216
rect 221240 3204 221246 3256
rect 324958 3204 324964 3256
rect 325016 3244 325022 3256
rect 326798 3244 326804 3256
rect 325016 3216 326804 3244
rect 325016 3204 325022 3216
rect 326798 3204 326804 3216
rect 326856 3204 326862 3256
rect 500310 3204 500316 3256
rect 500368 3244 500374 3256
rect 502978 3244 502984 3256
rect 500368 3216 502984 3244
rect 500368 3204 500374 3216
rect 502978 3204 502984 3216
rect 503036 3204 503042 3256
rect 127032 3148 219434 3176
rect 127032 3136 127038 3148
rect 220446 3136 220452 3188
rect 220504 3176 220510 3188
rect 226978 3176 226984 3188
rect 220504 3148 226984 3176
rect 220504 3136 220510 3148
rect 226978 3136 226984 3148
rect 227036 3136 227042 3188
rect 260190 3136 260196 3188
rect 260248 3176 260254 3188
rect 264146 3176 264152 3188
rect 260248 3148 264152 3176
rect 260248 3136 260254 3148
rect 264146 3136 264152 3148
rect 264204 3136 264210 3188
rect 271230 3136 271236 3188
rect 271288 3176 271294 3188
rect 274818 3176 274824 3188
rect 271288 3148 274824 3176
rect 271288 3136 271294 3148
rect 274818 3136 274824 3148
rect 274876 3136 274882 3188
rect 299658 3136 299664 3188
rect 299716 3176 299722 3188
rect 302326 3176 302332 3188
rect 299716 3148 302332 3176
rect 299716 3136 299722 3148
rect 302326 3136 302332 3148
rect 302384 3136 302390 3188
rect 389450 3136 389456 3188
rect 389508 3176 389514 3188
rect 392026 3176 392032 3188
rect 389508 3148 392032 3176
rect 389508 3136 389514 3148
rect 392026 3136 392032 3148
rect 392084 3136 392090 3188
rect 31352 3080 45554 3108
rect 31352 3068 31358 3080
rect 143534 3068 143540 3120
rect 143592 3108 143598 3120
rect 148226 3108 148232 3120
rect 143592 3080 148232 3108
rect 143592 3068 143598 3080
rect 148226 3068 148232 3080
rect 148284 3068 148290 3120
rect 231026 3068 231032 3120
rect 231084 3108 231090 3120
rect 238018 3108 238024 3120
rect 231084 3080 238024 3108
rect 231084 3068 231090 3080
rect 238018 3068 238024 3080
rect 238076 3068 238082 3120
rect 239306 3068 239312 3120
rect 239364 3108 239370 3120
rect 240594 3108 240600 3120
rect 239364 3080 240600 3108
rect 239364 3068 239370 3080
rect 240594 3068 240600 3080
rect 240652 3068 240658 3120
rect 542998 3068 543004 3120
rect 543056 3108 543062 3120
rect 545482 3108 545488 3120
rect 543056 3080 545488 3108
rect 543056 3068 543062 3080
rect 545482 3068 545488 3080
rect 545540 3068 545546 3120
rect 8754 3000 8760 3052
rect 8812 3040 8818 3052
rect 15838 3040 15844 3052
rect 8812 3012 15844 3040
rect 8812 3000 8818 3012
rect 15838 3000 15844 3012
rect 15896 3000 15902 3052
rect 27706 3000 27712 3052
rect 27764 3040 27770 3052
rect 35158 3040 35164 3052
rect 27764 3012 35164 3040
rect 27764 3000 27770 3012
rect 35158 3000 35164 3012
rect 35216 3000 35222 3052
rect 73798 3000 73804 3052
rect 73856 3040 73862 3052
rect 75178 3040 75184 3052
rect 73856 3012 75184 3040
rect 73856 3000 73862 3012
rect 75178 3000 75184 3012
rect 75236 3000 75242 3052
rect 118786 3000 118792 3052
rect 118844 3040 118850 3052
rect 119982 3040 119988 3052
rect 118844 3012 119988 3040
rect 118844 3000 118850 3012
rect 119982 3000 119988 3012
rect 120040 3000 120046 3052
rect 174262 3000 174268 3052
rect 174320 3040 174326 3052
rect 181346 3040 181352 3052
rect 174320 3012 181352 3040
rect 174320 3000 174326 3012
rect 181346 3000 181352 3012
rect 181404 3000 181410 3052
rect 252370 3000 252376 3052
rect 252428 3040 252434 3052
rect 258074 3040 258080 3052
rect 252428 3012 258080 3040
rect 252428 3000 252434 3012
rect 258074 3000 258080 3012
rect 258132 3000 258138 3052
rect 259454 3000 259460 3052
rect 259512 3040 259518 3052
rect 262214 3040 262220 3052
rect 259512 3012 262220 3040
rect 259512 3000 259518 3012
rect 262214 3000 262220 3012
rect 262272 3000 262278 3052
rect 280798 3000 280804 3052
rect 280856 3040 280862 3052
rect 283098 3040 283104 3052
rect 280856 3012 283104 3040
rect 280856 3000 280862 3012
rect 283098 3000 283104 3012
rect 283156 3000 283162 3052
rect 342990 3000 342996 3052
rect 343048 3040 343054 3052
rect 344554 3040 344560 3052
rect 343048 3012 344560 3040
rect 343048 3000 343054 3012
rect 344554 3000 344560 3012
rect 344612 3000 344618 3052
rect 374638 3000 374644 3052
rect 374696 3040 374702 3052
rect 377674 3040 377680 3052
rect 374696 3012 377680 3040
rect 374696 3000 374702 3012
rect 377674 3000 377680 3012
rect 377732 3000 377738 3052
rect 446398 3000 446404 3052
rect 446456 3040 446462 3052
rect 452102 3040 452108 3052
rect 446456 3012 452108 3040
rect 446456 3000 446462 3012
rect 452102 3000 452108 3012
rect 452160 3000 452166 3052
rect 493318 3000 493324 3052
rect 493376 3040 493382 3052
rect 495894 3040 495900 3052
rect 493376 3012 495900 3040
rect 493376 3000 493382 3012
rect 495894 3000 495900 3012
rect 495952 3000 495958 3052
rect 504358 3000 504364 3052
rect 504416 3040 504422 3052
rect 510062 3040 510068 3052
rect 504416 3012 510068 3040
rect 504416 3000 504422 3012
rect 510062 3000 510068 3012
rect 510120 3000 510126 3052
rect 511258 3000 511264 3052
rect 511316 3040 511322 3052
rect 513558 3040 513564 3052
rect 511316 3012 513564 3040
rect 511316 3000 511322 3012
rect 513558 3000 513564 3012
rect 513616 3000 513622 3052
rect 529198 3000 529204 3052
rect 529256 3040 529262 3052
rect 531314 3040 531320 3052
rect 529256 3012 531320 3040
rect 529256 3000 529262 3012
rect 531314 3000 531320 3012
rect 531372 3000 531378 3052
rect 23014 2932 23020 2984
rect 23072 2972 23078 2984
rect 28258 2972 28264 2984
rect 23072 2944 28264 2972
rect 23072 2932 23078 2944
rect 28258 2932 28264 2944
rect 28316 2932 28322 2984
rect 76190 2932 76196 2984
rect 76248 2972 76254 2984
rect 79318 2972 79324 2984
rect 76248 2944 79324 2972
rect 76248 2932 76254 2944
rect 79318 2932 79324 2944
rect 79376 2932 79382 2984
rect 222746 2932 222752 2984
rect 222804 2972 222810 2984
rect 223482 2972 223488 2984
rect 222804 2944 223488 2972
rect 222804 2932 222810 2944
rect 223482 2932 223488 2944
rect 223540 2932 223546 2984
rect 245654 2932 245660 2984
rect 245712 2972 245718 2984
rect 247586 2972 247592 2984
rect 245712 2944 247592 2972
rect 245712 2932 245718 2944
rect 247586 2932 247592 2944
rect 247644 2932 247650 2984
rect 435358 2932 435364 2984
rect 435416 2972 435422 2984
rect 437934 2972 437940 2984
rect 435416 2944 437940 2972
rect 435416 2932 435422 2944
rect 437934 2932 437940 2944
rect 437992 2932 437998 2984
rect 525150 2932 525156 2984
rect 525208 2972 525214 2984
rect 527818 2972 527824 2984
rect 525208 2944 527824 2972
rect 525208 2932 525214 2944
rect 527818 2932 527824 2944
rect 527876 2932 527882 2984
rect 77386 2864 77392 2916
rect 77444 2904 77450 2916
rect 79410 2904 79416 2916
rect 77444 2876 79416 2904
rect 77444 2864 77450 2876
rect 79410 2864 79416 2876
rect 79468 2864 79474 2916
rect 201494 2864 201500 2916
rect 201552 2904 201558 2916
rect 209038 2904 209044 2916
rect 201552 2876 209044 2904
rect 201552 2864 201558 2876
rect 209038 2864 209044 2876
rect 209096 2864 209102 2916
rect 223942 2864 223948 2916
rect 224000 2904 224006 2916
rect 224862 2904 224868 2916
rect 224000 2876 224868 2904
rect 224000 2864 224006 2876
rect 224862 2864 224868 2876
rect 224920 2864 224926 2916
rect 417510 2864 417516 2916
rect 417568 2904 417574 2916
rect 420178 2904 420184 2916
rect 417568 2876 420184 2904
rect 417568 2864 417574 2876
rect 420178 2864 420184 2876
rect 420236 2864 420242 2916
rect 432598 2864 432604 2916
rect 432656 2904 432662 2916
rect 434438 2904 434444 2916
rect 432656 2876 434444 2904
rect 432656 2864 432662 2876
rect 434438 2864 434444 2876
rect 434496 2864 434502 2916
rect 442350 2864 442356 2916
rect 442408 2904 442414 2916
rect 445018 2904 445024 2916
rect 442408 2876 445024 2904
rect 442408 2864 442414 2876
rect 445018 2864 445024 2876
rect 445076 2864 445082 2916
rect 471238 2864 471244 2916
rect 471296 2904 471302 2916
rect 473446 2904 473452 2916
rect 471296 2876 473452 2904
rect 471296 2864 471302 2876
rect 473446 2864 473452 2876
rect 473504 2864 473510 2916
rect 515030 2796 515036 2848
rect 515088 2836 515094 2848
rect 515950 2836 515956 2848
rect 515088 2808 515956 2836
rect 515088 2796 515094 2808
rect 515950 2796 515956 2808
rect 516008 2796 516014 2848
<< via1 >>
rect 331220 702992 331272 703044
rect 332508 702992 332560 703044
rect 170312 700884 170364 700936
rect 171048 700884 171100 700936
rect 252468 700612 252520 700664
rect 283840 700612 283892 700664
rect 246948 700544 247000 700596
rect 413652 700544 413704 700596
rect 72976 700476 73028 700528
rect 258080 700476 258132 700528
rect 40500 700408 40552 700460
rect 41328 700408 41380 700460
rect 235172 700408 235224 700460
rect 242164 700408 242216 700460
rect 244188 700408 244240 700460
rect 478512 700408 478564 700460
rect 24308 700340 24360 700392
rect 260104 700340 260156 700392
rect 479524 700340 479576 700392
rect 527180 700340 527232 700392
rect 218980 700272 219032 700324
rect 222844 700272 222896 700324
rect 241428 700272 241480 700324
rect 543464 700272 543516 700324
rect 105452 699660 105504 699712
rect 106188 699660 106240 699712
rect 154120 699660 154172 699712
rect 155224 699660 155276 699712
rect 347044 699660 347096 699712
rect 348792 699660 348844 699712
rect 359464 699660 359516 699712
rect 364984 699660 365036 699712
rect 396724 699660 396776 699712
rect 397460 699660 397512 699712
rect 249064 698912 249116 698964
rect 462320 698912 462372 698964
rect 266360 697552 266412 697604
rect 267648 697552 267700 697604
rect 238668 696940 238720 696992
rect 580172 696940 580224 696992
rect 3424 683204 3476 683256
rect 262220 683204 262272 683256
rect 238576 683136 238628 683188
rect 580172 683136 580224 683188
rect 237288 670692 237340 670744
rect 580172 670692 580224 670744
rect 3516 656888 3568 656940
rect 263692 656888 263744 656940
rect 235908 643084 235960 643136
rect 580172 643084 580224 643136
rect 3516 632068 3568 632120
rect 264980 632068 265032 632120
rect 237196 630640 237248 630692
rect 580172 630640 580224 630692
rect 3516 618264 3568 618316
rect 217324 618264 217376 618316
rect 234528 616836 234580 616888
rect 580172 616836 580224 616888
rect 250996 607860 251048 607912
rect 266360 607860 266412 607912
rect 3516 605820 3568 605872
rect 266360 605820 266412 605872
rect 233148 590656 233200 590708
rect 579804 590656 579856 590708
rect 3332 579640 3384 579692
rect 267740 579640 267792 579692
rect 234436 576852 234488 576904
rect 580172 576852 580224 576904
rect 3240 565836 3292 565888
rect 215944 565836 215996 565888
rect 231768 563048 231820 563100
rect 579804 563048 579856 563100
rect 3332 553392 3384 553444
rect 267832 553392 267884 553444
rect 230388 536800 230440 536852
rect 580172 536800 580224 536852
rect 2964 527144 3016 527196
rect 270500 527144 270552 527196
rect 231676 524424 231728 524476
rect 580172 524424 580224 524476
rect 3516 514768 3568 514820
rect 269764 514768 269816 514820
rect 229008 510620 229060 510672
rect 580172 510620 580224 510672
rect 3056 500964 3108 501016
rect 270592 500964 270644 501016
rect 227628 484372 227680 484424
rect 580172 484372 580224 484424
rect 3056 474716 3108 474768
rect 273260 474716 273312 474768
rect 228916 470568 228968 470620
rect 579988 470568 580040 470620
rect 3516 462340 3568 462392
rect 214564 462340 214616 462392
rect 227536 456764 227588 456816
rect 580172 456764 580224 456816
rect 3148 448536 3200 448588
rect 273352 448536 273404 448588
rect 224868 430584 224920 430636
rect 580172 430584 580224 430636
rect 3516 422288 3568 422340
rect 276020 422288 276072 422340
rect 226248 418140 226300 418192
rect 580172 418140 580224 418192
rect 2872 409844 2924 409896
rect 213184 409844 213236 409896
rect 224776 404336 224828 404388
rect 580172 404336 580224 404388
rect 3516 397468 3568 397520
rect 276112 397468 276164 397520
rect 3516 371220 3568 371272
rect 277400 371220 277452 371272
rect 371608 368908 371660 368960
rect 374184 368908 374236 368960
rect 445208 368500 445260 368552
rect 454040 368500 454092 368552
rect 371608 367140 371660 367192
rect 378140 367140 378192 367192
rect 371700 367072 371752 367124
rect 383660 367072 383712 367124
rect 445668 367072 445720 367124
rect 449900 367072 449952 367124
rect 371608 365848 371660 365900
rect 376944 365848 376996 365900
rect 371240 365780 371292 365832
rect 382280 365780 382332 365832
rect 371516 365712 371568 365764
rect 385040 365712 385092 365764
rect 445300 365712 445352 365764
rect 456800 365712 456852 365764
rect 371240 364624 371292 364676
rect 375564 364624 375616 364676
rect 371608 364352 371660 364404
rect 382372 364352 382424 364404
rect 445668 364352 445720 364404
rect 452752 364352 452804 364404
rect 371608 363060 371660 363112
rect 378324 363060 378376 363112
rect 371700 362924 371752 362976
rect 374276 362924 374328 362976
rect 444932 362924 444984 362976
rect 448612 362924 448664 362976
rect 371608 361632 371660 361684
rect 377036 361632 377088 361684
rect 371700 361564 371752 361616
rect 380992 361564 381044 361616
rect 445208 361564 445260 361616
rect 454132 361564 454184 361616
rect 371608 361496 371660 361548
rect 375380 361496 375432 361548
rect 445116 360748 445168 360800
rect 449992 360748 450044 360800
rect 371608 360408 371660 360460
rect 374460 360408 374512 360460
rect 371424 360340 371476 360392
rect 378232 360340 378284 360392
rect 444564 360272 444616 360324
rect 452660 360272 452712 360324
rect 371884 359524 371936 359576
rect 379520 359524 379572 359576
rect 372068 359456 372120 359508
rect 372896 359456 372948 359508
rect 371700 357484 371752 357536
rect 376760 357484 376812 357536
rect 3148 357416 3200 357468
rect 253204 357416 253256 357468
rect 371608 357416 371660 357468
rect 382556 357416 382608 357468
rect 444564 357416 444616 357468
rect 448520 357416 448572 357468
rect 371608 356192 371660 356244
rect 375656 356192 375708 356244
rect 444380 356192 444432 356244
rect 447140 356192 447192 356244
rect 371240 356124 371292 356176
rect 381084 356124 381136 356176
rect 371516 356056 371568 356108
rect 385224 356056 385276 356108
rect 444748 355036 444800 355088
rect 450084 355036 450136 355088
rect 371516 354764 371568 354816
rect 376852 354764 376904 354816
rect 371608 354696 371660 354748
rect 380900 354696 380952 354748
rect 371976 353948 372028 354000
rect 383752 353948 383804 354000
rect 371332 353336 371384 353388
rect 375472 353336 375524 353388
rect 371700 353268 371752 353320
rect 374092 353268 374144 353320
rect 372160 352588 372212 352640
rect 378416 352588 378468 352640
rect 372344 352520 372396 352572
rect 379612 352520 379664 352572
rect 444748 352452 444800 352504
rect 448704 352452 448756 352504
rect 444472 351976 444524 352028
rect 447232 351976 447284 352028
rect 371608 349256 371660 349308
rect 374000 349256 374052 349308
rect 371608 348168 371660 348220
rect 374368 348168 374420 348220
rect 445668 347760 445720 347812
rect 454224 347760 454276 347812
rect 444656 346400 444708 346452
rect 447508 346400 447560 346452
rect 445300 345108 445352 345160
rect 452844 345108 452896 345160
rect 3332 345040 3384 345092
rect 278780 345040 278832 345092
rect 445668 345040 445720 345092
rect 456892 345040 456944 345092
rect 445668 343680 445720 343732
rect 451280 343680 451332 343732
rect 445024 342252 445076 342304
rect 458180 342252 458232 342304
rect 444564 341232 444616 341284
rect 447416 341232 447468 341284
rect 369952 340552 370004 340604
rect 370136 340552 370188 340604
rect 444564 340144 444616 340196
rect 446036 340144 446088 340196
rect 300768 337424 300820 337476
rect 438952 337424 439004 337476
rect 198556 337356 198608 337408
rect 366916 337356 366968 337408
rect 441252 336744 441304 336796
rect 441620 336744 441672 336796
rect 369032 335316 369084 335368
rect 369308 335316 369360 335368
rect 137928 326340 137980 326392
rect 255320 326340 255372 326392
rect 220728 324300 220780 324352
rect 580172 324300 580224 324352
rect 3332 318792 3384 318844
rect 280896 318792 280948 318844
rect 220636 311856 220688 311908
rect 580172 311856 580224 311908
rect 245476 309748 245528 309800
rect 396724 309748 396776 309800
rect 3424 308388 3476 308440
rect 263232 308388 263284 308440
rect 253204 307504 253256 307556
rect 280344 307504 280396 307556
rect 217324 307436 217376 307488
rect 267280 307436 267332 307488
rect 215944 307368 215996 307420
rect 269948 307368 270000 307420
rect 213184 307300 213236 307352
rect 277768 307300 277820 307352
rect 249432 307232 249484 307284
rect 347044 307232 347096 307284
rect 89628 307164 89680 307216
rect 256240 307164 256292 307216
rect 8208 307096 8260 307148
rect 258080 307096 258132 307148
rect 222936 307028 222988 307080
rect 582472 307028 582524 307080
rect 222844 306076 222896 306128
rect 254308 306076 254360 306128
rect 214564 306008 214616 306060
rect 275100 306008 275152 306060
rect 248420 305940 248472 305992
rect 331220 305940 331272 305992
rect 155224 305872 155276 305924
rect 256884 305872 256936 305924
rect 41328 305804 41380 305856
rect 260380 305804 260432 305856
rect 240324 305736 240376 305788
rect 479524 305736 479576 305788
rect 222108 305668 222160 305720
rect 582380 305668 582432 305720
rect 221188 305600 221240 305652
rect 582564 305600 582616 305652
rect 3240 304988 3292 305040
rect 282828 304988 282880 305040
rect 242164 304784 242216 304836
rect 252560 304784 252612 304836
rect 249892 304716 249944 304768
rect 299480 304716 299532 304768
rect 202788 304648 202840 304700
rect 251824 304648 251876 304700
rect 171048 304580 171100 304632
rect 255136 304580 255188 304632
rect 247316 304512 247368 304564
rect 359464 304512 359516 304564
rect 106188 304444 106240 304496
rect 257712 304444 257764 304496
rect 244740 304376 244792 304428
rect 429200 304376 429252 304428
rect 242072 304308 242124 304360
rect 494060 304308 494112 304360
rect 239496 304240 239548 304292
rect 558920 304240 558972 304292
rect 129004 303696 129056 303748
rect 297732 303696 297784 303748
rect 202052 303628 202104 303680
rect 582472 303628 582524 303680
rect 242992 303492 243044 303544
rect 249064 303492 249116 303544
rect 256240 303288 256292 303340
rect 259460 303288 259512 303340
rect 209872 303084 209924 303136
rect 548524 303084 548576 303136
rect 258080 303016 258132 303068
rect 261208 303016 261260 303068
rect 237748 302948 237800 303000
rect 238668 302948 238720 303000
rect 251640 302948 251692 303000
rect 252468 302948 252520 303000
rect 260104 302948 260156 303000
rect 262128 302948 262180 303000
rect 263232 302948 263284 303000
rect 264704 302948 264756 303000
rect 269764 302948 269816 303000
rect 272524 302948 272576 303000
rect 211620 302880 211672 302932
rect 311164 302880 311216 302932
rect 209044 302812 209096 302864
rect 309784 302812 309836 302864
rect 180064 302744 180116 302796
rect 285588 302744 285640 302796
rect 299480 302744 299532 302796
rect 300768 302744 300820 302796
rect 212540 302676 212592 302728
rect 318064 302676 318116 302728
rect 204720 302608 204772 302660
rect 313924 302608 313976 302660
rect 207296 302540 207348 302592
rect 316684 302540 316736 302592
rect 166264 302472 166316 302524
rect 288164 302472 288216 302524
rect 148324 302404 148376 302456
rect 290832 302404 290884 302456
rect 215116 302336 215168 302388
rect 443644 302336 443696 302388
rect 14464 302268 14516 302320
rect 293408 302268 293460 302320
rect 251824 302200 251876 302252
rect 253388 302200 253440 302252
rect 285680 302200 285732 302252
rect 289912 302200 289964 302252
rect 223856 302064 223908 302116
rect 224776 302064 224828 302116
rect 228180 302064 228232 302116
rect 228916 302064 228968 302116
rect 230756 302064 230808 302116
rect 231676 302064 231728 302116
rect 233424 302064 233476 302116
rect 234436 302064 234488 302116
rect 235172 302064 235224 302116
rect 235908 302064 235960 302116
rect 236000 302064 236052 302116
rect 237196 302064 237248 302116
rect 216036 301588 216088 301640
rect 301504 301588 301556 301640
rect 199384 301520 199436 301572
rect 286416 301520 286468 301572
rect 206468 301452 206520 301504
rect 307024 301452 307076 301504
rect 174544 301384 174596 301436
rect 284668 301384 284720 301436
rect 152464 301316 152516 301368
rect 292488 301316 292540 301368
rect 156604 301248 156656 301300
rect 296904 301248 296956 301300
rect 144184 301180 144236 301232
rect 298652 301180 298704 301232
rect 90364 301112 90416 301164
rect 283840 301112 283892 301164
rect 210792 301044 210844 301096
rect 582932 301044 582984 301096
rect 202972 300976 203024 301028
rect 582656 300976 582708 301028
rect 200396 300908 200448 300960
rect 582380 300908 582432 300960
rect 201224 300840 201276 300892
rect 583116 300840 583168 300892
rect 213368 300296 213420 300348
rect 219348 300296 219400 300348
rect 219440 300296 219492 300348
rect 220728 300296 220780 300348
rect 226432 300296 226484 300348
rect 227536 300296 227588 300348
rect 196624 300228 196676 300280
rect 282092 300228 282144 300280
rect 203800 300160 203852 300212
rect 305644 300160 305696 300212
rect 159364 300092 159416 300144
rect 291660 300092 291712 300144
rect 155224 300024 155276 300076
rect 287152 300024 287204 300076
rect 157984 299956 158036 300008
rect 293960 299956 294012 300008
rect 151084 299888 151136 299940
rect 294788 299888 294840 299940
rect 146944 299820 146996 299872
rect 295708 299820 295760 299872
rect 88984 299752 89036 299804
rect 288716 299752 288768 299804
rect 218888 299684 218940 299736
rect 579896 299684 579948 299736
rect 219348 299616 219400 299668
rect 583024 299616 583076 299668
rect 208308 299548 208360 299600
rect 582840 299548 582892 299600
rect 205640 299480 205692 299532
rect 582564 299480 582616 299532
rect 216772 299412 216824 299464
rect 214656 299344 214708 299396
rect 216772 299276 216824 299328
rect 217416 299276 217468 299328
rect 217692 299276 217744 299328
rect 3424 298800 3476 298852
rect 199844 298256 199896 298308
rect 217968 299344 218020 299396
rect 218060 299276 218112 299328
rect 285680 299276 285732 299328
rect 580264 298732 580316 298784
rect 302792 298324 302844 298376
rect 323584 298324 323636 298376
rect 359464 298256 359516 298308
rect 312544 298188 312596 298240
rect 442264 298120 442316 298172
rect 436100 297644 436152 297696
rect 443000 297644 443052 297696
rect 434720 297576 434772 297628
rect 441712 297576 441764 297628
rect 373264 297440 373316 297492
rect 379520 297440 379572 297492
rect 374184 297372 374236 297424
rect 385132 297372 385184 297424
rect 450176 297372 450228 297424
rect 454040 297372 454092 297424
rect 445668 297032 445720 297084
rect 450176 297032 450228 297084
rect 302976 296760 303028 296812
rect 369492 296760 369544 296812
rect 373264 296760 373316 296812
rect 302884 296692 302936 296744
rect 369400 296692 369452 296744
rect 374184 296692 374236 296744
rect 370136 296080 370188 296132
rect 378140 296080 378192 296132
rect 372896 296012 372948 296064
rect 379520 296012 379572 296064
rect 369400 295944 369452 295996
rect 327724 295876 327776 295928
rect 352564 295808 352616 295860
rect 369400 295808 369452 295860
rect 383660 295944 383712 295996
rect 445760 295944 445812 295996
rect 458272 295944 458324 295996
rect 302792 295332 302844 295384
rect 322204 295332 322256 295384
rect 371240 295264 371292 295316
rect 376944 295264 376996 295316
rect 385408 295264 385460 295316
rect 445668 295264 445720 295316
rect 449900 295264 449952 295316
rect 449900 294652 449952 294704
rect 454040 294652 454092 294704
rect 371700 294584 371752 294636
rect 382280 294584 382332 294636
rect 445668 294584 445720 294636
rect 448796 294584 448848 294636
rect 456800 294584 456852 294636
rect 170404 293972 170456 294024
rect 197912 293972 197964 294024
rect 371700 293972 371752 294024
rect 376944 293972 376996 294024
rect 385040 293972 385092 294024
rect 3056 293904 3108 293956
rect 196624 293904 196676 293956
rect 373356 293904 373408 293956
rect 375564 293904 375616 293956
rect 372160 293428 372212 293480
rect 373356 293428 373408 293480
rect 371700 293224 371752 293276
rect 376024 293224 376076 293276
rect 382372 293224 382424 293276
rect 445668 293224 445720 293276
rect 452752 293224 452804 293276
rect 456800 293224 456852 293276
rect 371240 292408 371292 292460
rect 378324 292408 378376 292460
rect 371700 292340 371752 292392
rect 374184 292340 374236 292392
rect 378324 292000 378376 292052
rect 382372 292000 382424 292052
rect 372160 291932 372212 291984
rect 372712 291932 372764 291984
rect 378508 291932 378560 291984
rect 302240 291456 302292 291508
rect 304264 291456 304316 291508
rect 175924 291184 175976 291236
rect 197544 291184 197596 291236
rect 445668 291184 445720 291236
rect 448612 291184 448664 291236
rect 452752 291184 452804 291236
rect 371240 290504 371292 290556
rect 377036 290504 377088 290556
rect 371700 290436 371752 290488
rect 380992 290436 381044 290488
rect 445760 290436 445812 290488
rect 454132 290436 454184 290488
rect 371700 289552 371752 289604
rect 375380 289552 375432 289604
rect 375564 289552 375616 289604
rect 445668 289144 445720 289196
rect 449992 289144 450044 289196
rect 454132 289144 454184 289196
rect 371700 289076 371752 289128
rect 378232 289076 378284 289128
rect 371700 288464 371752 288516
rect 374460 288464 374512 288516
rect 302700 288396 302752 288448
rect 320824 288396 320876 288448
rect 371700 288328 371752 288380
rect 379612 288328 379664 288380
rect 371700 287648 371752 287700
rect 378416 287648 378468 287700
rect 449992 287376 450044 287428
rect 452660 287376 452712 287428
rect 445484 287240 445536 287292
rect 445852 287240 445904 287292
rect 452660 287240 452712 287292
rect 445668 287104 445720 287156
rect 449992 287104 450044 287156
rect 176016 287036 176068 287088
rect 197544 287036 197596 287088
rect 379612 287036 379664 287088
rect 385316 287036 385368 287088
rect 371700 286968 371752 287020
rect 376760 286968 376812 287020
rect 371976 286628 372028 286680
rect 372160 286628 372212 286680
rect 371608 286492 371660 286544
rect 371976 286492 372028 286544
rect 371608 286356 371660 286408
rect 374644 286356 374696 286408
rect 382556 286356 382608 286408
rect 371240 286288 371292 286340
rect 383752 286288 383804 286340
rect 445668 285948 445720 286000
rect 448520 285948 448572 286000
rect 302792 285676 302844 285728
rect 324964 285676 325016 285728
rect 376760 285676 376812 285728
rect 381268 285676 381320 285728
rect 371700 285608 371752 285660
rect 381084 285608 381136 285660
rect 371608 285472 371660 285524
rect 375380 285472 375432 285524
rect 375656 285472 375708 285524
rect 445392 284792 445444 284844
rect 447140 284792 447192 284844
rect 381084 284384 381136 284436
rect 382280 284384 382332 284436
rect 371608 284316 371660 284368
rect 377404 284316 377456 284368
rect 385224 284316 385276 284368
rect 447140 284316 447192 284368
rect 447324 284316 447376 284368
rect 371700 283636 371752 283688
rect 376760 283636 376812 283688
rect 371608 283568 371660 283620
rect 380900 283568 380952 283620
rect 445668 283568 445720 283620
rect 450084 283568 450136 283620
rect 178684 282888 178736 282940
rect 197360 282888 197412 282940
rect 380900 282888 380952 282940
rect 381176 282888 381228 282940
rect 371608 282684 371660 282736
rect 375472 282684 375524 282736
rect 371608 282140 371660 282192
rect 374092 282140 374144 282192
rect 374276 282140 374328 282192
rect 181444 281528 181496 281580
rect 197360 281528 197412 281580
rect 302516 281528 302568 281580
rect 353944 281528 353996 281580
rect 445668 281324 445720 281376
rect 448704 281324 448756 281376
rect 445024 280236 445076 280288
rect 447232 280236 447284 280288
rect 444380 279624 444432 279676
rect 444656 279624 444708 279676
rect 371976 278944 372028 278996
rect 374092 278944 374144 278996
rect 173164 278740 173216 278792
rect 197728 278740 197780 278792
rect 302792 278740 302844 278792
rect 356704 278740 356756 278792
rect 369124 278604 369176 278656
rect 369400 278604 369452 278656
rect 371700 277312 371752 277364
rect 374000 277312 374052 277364
rect 445668 276632 445720 276684
rect 454224 276632 454276 276684
rect 371700 276088 371752 276140
rect 374368 276088 374420 276140
rect 375104 276088 375156 276140
rect 169668 276020 169720 276072
rect 197360 276020 197412 276072
rect 302792 276020 302844 276072
rect 360200 276020 360252 276072
rect 360660 276020 360712 276072
rect 374000 276020 374052 276072
rect 374552 276020 374604 276072
rect 445668 275952 445720 276004
rect 447508 275952 447560 276004
rect 369216 275340 369268 275392
rect 369400 275340 369452 275392
rect 447508 275272 447560 275324
rect 458364 275272 458416 275324
rect 372620 274728 372672 274780
rect 373080 274728 373132 274780
rect 196624 274660 196676 274712
rect 198648 274660 198700 274712
rect 370320 274660 370372 274712
rect 372896 274660 372948 274712
rect 445668 274592 445720 274644
rect 446404 274592 446456 274644
rect 452844 274592 452896 274644
rect 445024 273912 445076 273964
rect 453304 273912 453356 273964
rect 456892 273912 456944 273964
rect 442264 273164 442316 273216
rect 579896 273164 579948 273216
rect 445668 272484 445720 272536
rect 451280 272484 451332 272536
rect 456892 272484 456944 272536
rect 177304 271872 177356 271924
rect 197544 271872 197596 271924
rect 195244 270512 195296 270564
rect 197728 270512 197780 270564
rect 445668 270512 445720 270564
rect 451372 270512 451424 270564
rect 458180 270512 458232 270564
rect 447232 270444 447284 270496
rect 447416 270444 447468 270496
rect 445392 269764 445444 269816
rect 447232 269764 447284 269816
rect 369032 268744 369084 268796
rect 444564 268676 444616 268728
rect 446036 268676 446088 268728
rect 369124 268404 369176 268456
rect 303252 268336 303304 268388
rect 327724 268336 327776 268388
rect 192484 268132 192536 268184
rect 197820 268132 197872 268184
rect 3516 267656 3568 267708
rect 90364 267656 90416 267708
rect 323584 267656 323636 267708
rect 438860 267656 438912 267708
rect 191104 266432 191156 266484
rect 197360 266432 197412 266484
rect 359464 266296 359516 266348
rect 366916 266296 366968 266348
rect 362868 266228 362920 266280
rect 435180 266296 435232 266348
rect 441620 266296 441672 266348
rect 324964 266160 325016 266212
rect 364892 266160 364944 266212
rect 437388 266228 437440 266280
rect 443000 266228 443052 266280
rect 368480 266092 368532 266144
rect 360200 265684 360252 265736
rect 360936 265684 360988 265736
rect 431960 265684 432012 265736
rect 432604 265684 432656 265736
rect 368480 265616 368532 265668
rect 369308 265616 369360 265668
rect 440884 265616 440936 265668
rect 302792 264868 302844 264920
rect 352564 264868 352616 264920
rect 188436 263576 188488 263628
rect 197360 263576 197412 263628
rect 187056 262216 187108 262268
rect 197360 262216 197412 262268
rect 302792 262148 302844 262200
rect 370136 262148 370188 262200
rect 184296 259428 184348 259480
rect 197728 259428 197780 259480
rect 182824 256708 182876 256760
rect 197544 256708 197596 256760
rect 302792 256708 302844 256760
rect 370504 256708 370556 256760
rect 181536 255280 181588 255332
rect 197912 255280 197964 255332
rect 3148 255212 3200 255264
rect 180064 255212 180116 255264
rect 302332 253920 302384 253972
rect 359464 253920 359516 253972
rect 180064 252560 180116 252612
rect 197544 252560 197596 252612
rect 178776 251200 178828 251252
rect 197360 251200 197412 251252
rect 370228 249704 370280 249756
rect 373356 249704 373408 249756
rect 171784 248412 171836 248464
rect 197636 248412 197688 248464
rect 302792 248412 302844 248464
rect 370228 248412 370280 248464
rect 301504 245556 301556 245608
rect 580172 245556 580224 245608
rect 173256 244264 173308 244316
rect 197360 244264 197412 244316
rect 191196 241476 191248 241528
rect 197912 241476 197964 241528
rect 3516 241408 3568 241460
rect 174544 241408 174596 241460
rect 180156 240116 180208 240168
rect 197728 240116 197780 240168
rect 302976 239368 303028 239420
rect 370320 239368 370372 239420
rect 192576 237396 192628 237448
rect 197544 237396 197596 237448
rect 195336 236104 195388 236156
rect 197728 236104 197780 236156
rect 193864 233792 193916 233844
rect 197728 233792 197780 233844
rect 312544 233180 312596 233232
rect 579988 233180 580040 233232
rect 196716 231888 196768 231940
rect 198372 231888 198424 231940
rect 303068 231072 303120 231124
rect 369584 231072 369636 231124
rect 374184 231072 374236 231124
rect 303160 229712 303212 229764
rect 372804 229712 372856 229764
rect 177396 229100 177448 229152
rect 197636 229100 197688 229152
rect 311164 228352 311216 228404
rect 580264 228352 580316 228404
rect 186964 227740 187016 227792
rect 197360 227740 197412 227792
rect 303252 226992 303304 227044
rect 372620 226992 372672 227044
rect 440884 226244 440936 226296
rect 443000 226244 443052 226296
rect 437388 226176 437440 226228
rect 441712 226176 441764 226228
rect 371608 225700 371660 225752
rect 372344 225700 372396 225752
rect 372988 225700 373040 225752
rect 373540 225700 373592 225752
rect 378416 225700 378468 225752
rect 372252 225632 372304 225684
rect 373264 225632 373316 225684
rect 381084 225632 381136 225684
rect 302884 225564 302936 225616
rect 369860 225564 369912 225616
rect 371608 225564 371660 225616
rect 385132 225564 385184 225616
rect 359648 225292 359700 225344
rect 372988 225292 373040 225344
rect 372804 225224 372856 225276
rect 373172 225224 373224 225276
rect 359372 225156 359424 225208
rect 374368 225156 374420 225208
rect 378324 225156 378376 225208
rect 359556 225088 359608 225140
rect 383752 225088 383804 225140
rect 371240 225020 371292 225072
rect 372804 225020 372856 225072
rect 441804 225020 441856 225072
rect 184204 224952 184256 225004
rect 197360 224952 197412 225004
rect 372528 224952 372580 225004
rect 372988 224952 373040 225004
rect 444564 224952 444616 225004
rect 449900 224952 449952 225004
rect 450176 224952 450228 225004
rect 359464 224408 359516 224460
rect 369400 224408 369452 224460
rect 302792 224340 302844 224392
rect 369952 224340 370004 224392
rect 302700 224272 302752 224324
rect 370228 224272 370280 224324
rect 371332 224272 371384 224324
rect 379520 224272 379572 224324
rect 302976 224204 303028 224256
rect 370412 224204 370464 224256
rect 371608 224204 371660 224256
rect 383660 224204 383712 224256
rect 359740 223932 359792 223984
rect 385316 223932 385368 223984
rect 359464 223864 359516 223916
rect 374460 223864 374512 223916
rect 441804 224204 441856 224256
rect 458272 224204 458324 224256
rect 374000 223796 374052 223848
rect 302792 223524 302844 223576
rect 359372 223524 359424 223576
rect 378324 223524 378376 223576
rect 382464 223524 382516 223576
rect 444564 223524 444616 223576
rect 454040 223524 454092 223576
rect 371608 222844 371660 222896
rect 374920 222844 374972 222896
rect 378140 222844 378192 222896
rect 371240 222368 371292 222420
rect 375656 222368 375708 222420
rect 376944 222368 376996 222420
rect 371608 222300 371660 222352
rect 372344 222300 372396 222352
rect 374000 222300 374052 222352
rect 371332 222232 371384 222284
rect 378324 222232 378376 222284
rect 188344 222164 188396 222216
rect 197360 222164 197412 222216
rect 445668 222096 445720 222148
rect 448612 222096 448664 222148
rect 448796 222096 448848 222148
rect 370136 221416 370188 221468
rect 385040 221416 385092 221468
rect 371240 220872 371292 220924
rect 382464 220872 382516 220924
rect 385408 220872 385460 220924
rect 302792 220736 302844 220788
rect 359464 220736 359516 220788
rect 369860 220736 369912 220788
rect 376024 220736 376076 220788
rect 380900 220736 380952 220788
rect 456800 220736 456852 220788
rect 456984 220736 457036 220788
rect 371240 220668 371292 220720
rect 372804 220668 372856 220720
rect 373172 220668 373224 220720
rect 382372 220668 382424 220720
rect 372068 220600 372120 220652
rect 445116 220056 445168 220108
rect 456984 220056 457036 220108
rect 445668 219580 445720 219632
rect 452752 219580 452804 219632
rect 372620 219376 372672 219428
rect 380992 219376 381044 219428
rect 443644 219376 443696 219428
rect 579896 219376 579948 219428
rect 370412 218696 370464 218748
rect 378508 218696 378560 218748
rect 378232 218220 378284 218272
rect 378508 218220 378560 218272
rect 371056 218084 371108 218136
rect 375932 218084 375984 218136
rect 377036 218084 377088 218136
rect 174544 218016 174596 218068
rect 197544 218016 197596 218068
rect 445760 218016 445812 218068
rect 446128 218016 446180 218068
rect 302516 217948 302568 218000
rect 359740 217948 359792 218000
rect 370228 217948 370280 218000
rect 375564 217948 375616 218000
rect 445668 217268 445720 217320
rect 454132 217268 454184 217320
rect 371608 217132 371660 217184
rect 372252 217132 372304 217184
rect 371608 216996 371660 217048
rect 374368 216996 374420 217048
rect 174636 216656 174688 216708
rect 197360 216656 197412 216708
rect 375564 216656 375616 216708
rect 376944 216656 376996 216708
rect 445668 216112 445720 216164
rect 449992 216112 450044 216164
rect 371332 215976 371384 216028
rect 374460 215976 374512 216028
rect 378140 215976 378192 216028
rect 371608 215908 371660 215960
rect 375564 215908 375616 215960
rect 385224 215908 385276 215960
rect 372344 215432 372396 215484
rect 373540 215432 373592 215484
rect 375012 215432 375064 215484
rect 449992 215296 450044 215348
rect 450176 215296 450228 215348
rect 3332 215228 3384 215280
rect 199384 215228 199436 215280
rect 302792 215228 302844 215280
rect 359648 215228 359700 215280
rect 371608 215228 371660 215280
rect 383752 215160 383804 215212
rect 385224 215160 385276 215212
rect 378416 214344 378468 214396
rect 381268 214344 381320 214396
rect 445668 214004 445720 214056
rect 452660 214004 452712 214056
rect 452844 214004 452896 214056
rect 174728 213936 174780 213988
rect 197544 213936 197596 213988
rect 371608 213936 371660 213988
rect 378416 213936 378468 213988
rect 445668 213868 445720 213920
rect 448520 213868 448572 213920
rect 372068 213732 372120 213784
rect 377404 213732 377456 213784
rect 382556 213732 382608 213784
rect 371332 213256 371384 213308
rect 374644 213256 374696 213308
rect 377036 213256 377088 213308
rect 371608 213188 371660 213240
rect 375380 213188 375432 213240
rect 383752 213188 383804 213240
rect 371332 213120 371384 213172
rect 372252 213120 372304 213172
rect 445300 212780 445352 212832
rect 447324 212780 447376 212832
rect 170496 212508 170548 212560
rect 197360 212508 197412 212560
rect 376852 212440 376904 212492
rect 381176 212440 381228 212492
rect 372252 211760 372304 211812
rect 373172 211760 373224 211812
rect 382280 211760 382332 211812
rect 445668 211556 445720 211608
rect 450084 211556 450136 211608
rect 371608 211216 371660 211268
rect 376760 211216 376812 211268
rect 370412 211148 370464 211200
rect 376852 211148 376904 211200
rect 302792 211080 302844 211132
rect 359556 211080 359608 211132
rect 374736 211080 374788 211132
rect 375472 211080 375524 211132
rect 445852 211080 445904 211132
rect 446036 211080 446088 211132
rect 371608 210604 371660 210656
rect 374736 210604 374788 210656
rect 444564 210468 444616 210520
rect 446036 210468 446088 210520
rect 372712 210060 372764 210112
rect 374276 210060 374328 210112
rect 182916 209788 182968 209840
rect 197360 209788 197412 209840
rect 375840 209788 375892 209840
rect 376760 209788 376812 209840
rect 445668 209176 445720 209228
rect 448704 209176 448756 209228
rect 160008 209040 160060 209092
rect 198096 209040 198148 209092
rect 369676 208700 369728 208752
rect 372988 208700 373040 208752
rect 445116 208156 445168 208208
rect 447140 208156 447192 208208
rect 302332 207000 302384 207052
rect 359464 207000 359516 207052
rect 369768 206932 369820 206984
rect 374092 206932 374144 206984
rect 369308 206456 369360 206508
rect 369216 206252 369268 206304
rect 369124 206116 369176 206168
rect 369400 206116 369452 206168
rect 371608 205776 371660 205828
rect 372620 205776 372672 205828
rect 373264 205776 373316 205828
rect 181628 205640 181680 205692
rect 197360 205640 197412 205692
rect 445300 205572 445352 205624
rect 454224 205572 454276 205624
rect 458180 205572 458232 205624
rect 371608 205300 371660 205352
rect 374552 205300 374604 205352
rect 371608 204756 371660 204808
rect 372896 204756 372948 204808
rect 302700 204280 302752 204332
rect 359556 204280 359608 204332
rect 371608 204212 371660 204264
rect 374000 204212 374052 204264
rect 375104 204212 375156 204264
rect 454224 204212 454276 204264
rect 458364 204212 458416 204264
rect 369584 204008 369636 204060
rect 369584 203804 369636 203856
rect 445024 202852 445076 202904
rect 454224 202852 454276 202904
rect 3056 202784 3108 202836
rect 166264 202784 166316 202836
rect 372068 202784 372120 202836
rect 373080 202784 373132 202836
rect 373356 202784 373408 202836
rect 371240 202444 371292 202496
rect 374644 202444 374696 202496
rect 370044 201560 370096 201612
rect 374000 201560 374052 201612
rect 180248 201492 180300 201544
rect 197360 201492 197412 201544
rect 302792 201492 302844 201544
rect 360108 201492 360160 201544
rect 445668 201492 445720 201544
rect 446404 201492 446456 201544
rect 451280 201492 451332 201544
rect 445668 200744 445720 200796
rect 453304 200744 453356 200796
rect 456800 200744 456852 200796
rect 445668 199384 445720 199436
rect 452660 199384 452712 199436
rect 456892 199384 456944 199436
rect 445668 198772 445720 198824
rect 451372 198772 451424 198824
rect 193956 198704 194008 198756
rect 198280 198704 198332 198756
rect 445392 197616 445444 197668
rect 447232 197616 447284 197668
rect 173348 197344 173400 197396
rect 197360 197344 197412 197396
rect 302792 197344 302844 197396
rect 441344 197276 441396 197328
rect 443000 197276 443052 197328
rect 360108 197208 360160 197260
rect 383752 197208 383804 197260
rect 382556 197140 382608 197192
rect 359464 197072 359516 197124
rect 378416 197072 378468 197124
rect 359556 197004 359608 197056
rect 377036 197004 377088 197056
rect 382280 196732 382332 196784
rect 382556 196732 382608 196784
rect 302884 195984 302936 196036
rect 369492 195984 369544 196036
rect 302332 195916 302384 195968
rect 371240 195916 371292 195968
rect 374092 195916 374144 195968
rect 373172 195848 373224 195900
rect 302976 195236 303028 195288
rect 372620 195236 372672 195288
rect 374184 195236 374236 195288
rect 173440 194556 173492 194608
rect 197636 194556 197688 194608
rect 304264 194488 304316 194540
rect 366916 194488 366968 194540
rect 436008 194488 436060 194540
rect 441620 194488 441672 194540
rect 437204 194420 437256 194472
rect 441712 194420 441764 194472
rect 443184 194420 443236 194472
rect 301504 193808 301556 193860
rect 438952 193808 439004 193860
rect 435180 193672 435232 193724
rect 436008 193672 436060 193724
rect 176108 193196 176160 193248
rect 197360 193196 197412 193248
rect 171876 193128 171928 193180
rect 173256 193128 173308 193180
rect 302792 193128 302844 193180
rect 370412 193128 370464 193180
rect 191288 191632 191340 191684
rect 198188 191632 198240 191684
rect 172428 190136 172480 190188
rect 178684 190136 178736 190188
rect 183008 189048 183060 189100
rect 197360 189048 197412 189100
rect 3516 188980 3568 189032
rect 155224 188980 155276 189032
rect 172060 188980 172112 189032
rect 181444 188980 181496 189032
rect 302792 188980 302844 189032
rect 375840 188980 375892 189032
rect 172152 187620 172204 187672
rect 173164 187620 173216 187672
rect 178684 186328 178736 186380
rect 197360 186328 197412 186380
rect 302700 186260 302752 186312
rect 374736 186260 374788 186312
rect 375288 186260 375340 186312
rect 171968 185512 172020 185564
rect 180156 185512 180208 185564
rect 195428 185172 195480 185224
rect 198096 185172 198148 185224
rect 172428 184832 172480 184884
rect 196624 184832 196676 184884
rect 171692 184764 171744 184816
rect 177304 184764 177356 184816
rect 196808 184152 196860 184204
rect 198372 184152 198424 184204
rect 172428 183472 172480 183524
rect 195244 183472 195296 183524
rect 181444 182792 181496 182844
rect 197360 182792 197412 182844
rect 172060 182112 172112 182164
rect 192484 182112 192536 182164
rect 436008 181636 436060 181688
rect 441712 181636 441764 181688
rect 172428 180752 172480 180804
rect 191104 180752 191156 180804
rect 302792 180072 302844 180124
rect 370320 180072 370372 180124
rect 192484 179392 192536 179444
rect 198372 179392 198424 179444
rect 172428 179324 172480 179376
rect 188436 179324 188488 179376
rect 318064 179324 318116 179376
rect 580172 179324 580224 179376
rect 188528 178032 188580 178084
rect 197360 178032 197412 178084
rect 172428 177964 172480 178016
rect 187056 177964 187108 178016
rect 172336 177896 172388 177948
rect 184296 177896 184348 177948
rect 172244 176604 172296 176656
rect 182824 176604 182876 176656
rect 302792 175924 302844 175976
rect 370136 175924 370188 175976
rect 370780 175924 370832 175976
rect 177304 175244 177356 175296
rect 197636 175244 197688 175296
rect 172428 175176 172480 175228
rect 181536 175176 181588 175228
rect 370596 175176 370648 175228
rect 375748 175176 375800 175228
rect 448612 175176 448664 175228
rect 184296 173884 184348 173936
rect 197360 173884 197412 173936
rect 172428 173612 172480 173664
rect 180064 173612 180116 173664
rect 180156 173136 180208 173188
rect 198096 173136 198148 173188
rect 374552 172456 374604 172508
rect 450176 172456 450228 172508
rect 172428 172388 172480 172440
rect 178776 172388 178828 172440
rect 369676 171096 369728 171148
rect 374552 171096 374604 171148
rect 172244 171028 172296 171080
rect 198004 171028 198056 171080
rect 302792 170348 302844 170400
rect 370596 170348 370648 170400
rect 172244 168988 172296 169040
rect 193864 168988 193916 169040
rect 172428 168308 172480 168360
rect 191196 168308 191248 168360
rect 370044 168308 370096 168360
rect 446128 168376 446180 168428
rect 369124 167900 369176 167952
rect 370044 167900 370096 167952
rect 369308 166948 369360 167000
rect 370504 166948 370556 167000
rect 449992 167016 450044 167068
rect 178776 166336 178828 166388
rect 197728 166336 197780 166388
rect 171784 166268 171836 166320
rect 192484 166268 192536 166320
rect 172060 165520 172112 165572
rect 192576 165520 192628 165572
rect 192484 164500 192536 164552
rect 197544 164500 197596 164552
rect 448704 164228 448756 164280
rect 3240 164160 3292 164212
rect 88984 164160 89036 164212
rect 172428 164160 172480 164212
rect 195336 164160 195388 164212
rect 370228 164160 370280 164212
rect 370504 164160 370556 164212
rect 370596 164160 370648 164212
rect 372896 164160 372948 164212
rect 452844 164160 452896 164212
rect 172152 162800 172204 162852
rect 196624 162800 196676 162852
rect 198188 162800 198240 162852
rect 196716 162732 196768 162784
rect 373264 162120 373316 162172
rect 454132 162120 454184 162172
rect 303068 161372 303120 161424
rect 369768 161372 369820 161424
rect 370228 161372 370280 161424
rect 172428 161168 172480 161220
rect 177396 161168 177448 161220
rect 169208 160760 169260 160812
rect 175924 160760 175976 160812
rect 165160 160488 165212 160540
rect 198740 160692 198792 160744
rect 372620 160692 372672 160744
rect 373356 160692 373408 160744
rect 445944 160692 445996 160744
rect 177488 160080 177540 160132
rect 197544 160080 197596 160132
rect 192576 158788 192628 158840
rect 197360 158788 197412 158840
rect 162860 158652 162912 158704
rect 176016 158652 176068 158704
rect 369400 158652 369452 158704
rect 373908 158652 373960 158704
rect 448520 158652 448572 158704
rect 166908 157972 166960 158024
rect 195244 157972 195296 158024
rect 372068 156680 372120 156732
rect 444472 156680 444524 156732
rect 171968 156612 172020 156664
rect 188528 156612 188580 156664
rect 309784 156612 309836 156664
rect 579620 156612 579672 156664
rect 191104 155932 191156 155984
rect 197820 155932 197872 155984
rect 302884 155864 302936 155916
rect 369584 155864 369636 155916
rect 370872 155864 370924 155916
rect 444564 155864 444616 155916
rect 447324 155864 447376 155916
rect 182824 154572 182876 154624
rect 197360 154572 197412 154624
rect 374644 154572 374696 154624
rect 444564 154572 444616 154624
rect 171600 154504 171652 154556
rect 174544 154504 174596 154556
rect 371976 154504 372028 154556
rect 385132 154504 385184 154556
rect 371424 154436 371476 154488
rect 381084 154436 381136 154488
rect 444932 154028 444984 154080
rect 449900 154028 449952 154080
rect 171692 153756 171744 153808
rect 174636 153756 174688 153808
rect 370872 153280 370924 153332
rect 444380 153348 444432 153400
rect 452752 153348 452804 153400
rect 370228 153212 370280 153264
rect 441804 153212 441856 153264
rect 445300 153212 445352 153264
rect 171600 153144 171652 153196
rect 174728 153144 174780 153196
rect 302516 153144 302568 153196
rect 302608 153076 302660 153128
rect 302792 153008 302844 153060
rect 369308 153144 369360 153196
rect 369584 153144 369636 153196
rect 370136 153144 370188 153196
rect 370596 153144 370648 153196
rect 371884 153144 371936 153196
rect 383660 153144 383712 153196
rect 445668 153144 445720 153196
rect 458272 153144 458324 153196
rect 371424 153076 371476 153128
rect 379520 153076 379572 153128
rect 370044 153008 370096 153060
rect 369676 152872 369728 152924
rect 369308 152804 369360 152856
rect 359464 152124 359516 152176
rect 369124 152124 369176 152176
rect 372620 152124 372672 152176
rect 358912 152056 358964 152108
rect 369216 152056 369268 152108
rect 374644 152056 374696 152108
rect 360108 151988 360160 152040
rect 369400 151988 369452 152040
rect 359556 151920 359608 151972
rect 369584 151920 369636 151972
rect 175924 151784 175976 151836
rect 197360 151784 197412 151836
rect 172244 151716 172296 151768
rect 191288 151716 191340 151768
rect 302700 151716 302752 151768
rect 370136 151852 370188 151904
rect 371424 151716 371476 151768
rect 374920 151716 374972 151768
rect 444932 151716 444984 151768
rect 454040 151716 454092 151768
rect 172428 151648 172480 151700
rect 182916 151648 182968 151700
rect 171692 151580 171744 151632
rect 181628 151580 181680 151632
rect 371976 151580 372028 151632
rect 378324 151580 378376 151632
rect 371424 150900 371476 150952
rect 375656 150900 375708 150952
rect 3516 150356 3568 150408
rect 148324 150356 148376 150408
rect 172428 150356 172480 150408
rect 193956 150356 194008 150408
rect 371976 150356 372028 150408
rect 385040 150356 385092 150408
rect 371424 150288 371476 150340
rect 382464 150288 382516 150340
rect 444932 150152 444984 150204
rect 448612 150152 448664 150204
rect 171508 149744 171560 149796
rect 180248 149744 180300 149796
rect 174544 149064 174596 149116
rect 197360 149064 197412 149116
rect 302332 148996 302384 149048
rect 360108 148996 360160 149048
rect 371976 148996 372028 149048
rect 382372 148996 382424 149048
rect 445300 148996 445352 149048
rect 456984 148996 457036 149048
rect 371424 148928 371476 148980
rect 380900 148928 380952 148980
rect 172428 148860 172480 148912
rect 195428 148860 195480 148912
rect 171692 148316 171744 148368
rect 173348 148316 173400 148368
rect 173164 148248 173216 148300
rect 198096 148316 198148 148368
rect 171508 147976 171560 148028
rect 173440 147976 173492 148028
rect 181536 147636 181588 147688
rect 197360 147636 197412 147688
rect 172336 147568 172388 147620
rect 196808 147568 196860 147620
rect 371976 147568 372028 147620
rect 380992 147568 381044 147620
rect 171692 147500 171744 147552
rect 176108 147500 176160 147552
rect 371424 147500 371476 147552
rect 378232 147500 378284 147552
rect 444380 146548 444432 146600
rect 446128 146548 446180 146600
rect 172428 146208 172480 146260
rect 183008 146208 183060 146260
rect 195336 146208 195388 146260
rect 198004 146208 198056 146260
rect 302792 146208 302844 146260
rect 358912 146208 358964 146260
rect 445668 146208 445720 146260
rect 454132 146208 454184 146260
rect 171692 146140 171744 146192
rect 181444 146140 181496 146192
rect 371424 146140 371476 146192
rect 375932 146140 375984 146192
rect 371976 146072 372028 146124
rect 376944 146072 376996 146124
rect 371424 145868 371476 145920
rect 374368 145868 374420 145920
rect 172428 145732 172480 145784
rect 178684 145732 178736 145784
rect 171692 144848 171744 144900
rect 180156 144848 180208 144900
rect 445300 144780 445352 144832
rect 450084 144780 450136 144832
rect 371424 144712 371476 144764
rect 378140 144712 378192 144764
rect 371424 144236 371476 144288
rect 375564 144236 375616 144288
rect 171876 144032 171928 144084
rect 177304 144032 177356 144084
rect 371424 143896 371476 143948
rect 375012 143896 375064 143948
rect 179420 143556 179472 143608
rect 197360 143556 197412 143608
rect 172428 143488 172480 143540
rect 184296 143488 184348 143540
rect 371976 143488 372028 143540
rect 385224 143488 385276 143540
rect 371424 143420 371476 143472
rect 378416 143420 378468 143472
rect 445208 142196 445260 142248
rect 452844 142196 452896 142248
rect 172428 142060 172480 142112
rect 196624 142060 196676 142112
rect 302792 142060 302844 142112
rect 359556 142060 359608 142112
rect 371976 142060 372028 142112
rect 383752 142060 383804 142112
rect 172336 141992 172388 142044
rect 192484 141992 192536 142044
rect 372068 141992 372120 142044
rect 382280 141992 382332 142044
rect 371424 141924 371476 141976
rect 377036 141924 377088 141976
rect 445116 141924 445168 141976
rect 448520 141924 448572 141976
rect 171876 141788 171928 141840
rect 178776 141788 178828 141840
rect 178040 140768 178092 140820
rect 197544 140768 197596 140820
rect 172428 140700 172480 140752
rect 195336 140700 195388 140752
rect 371424 140632 371476 140684
rect 376852 140632 376904 140684
rect 445116 140360 445168 140412
rect 449992 140360 450044 140412
rect 172152 140292 172204 140344
rect 173164 140292 173216 140344
rect 371976 140292 372028 140344
rect 373172 140292 373224 140344
rect 171324 140020 171376 140072
rect 198096 140020 198148 140072
rect 172428 139340 172480 139392
rect 192576 139340 192628 139392
rect 302700 139340 302752 139392
rect 359464 139340 359516 139392
rect 371424 139340 371476 139392
rect 376760 139340 376812 139392
rect 548524 139340 548576 139392
rect 580172 139340 580224 139392
rect 172336 139272 172388 139324
rect 191104 139272 191156 139324
rect 172244 139204 172296 139256
rect 177488 139204 177540 139256
rect 371976 139000 372028 139052
rect 374184 139000 374236 139052
rect 371424 138660 371476 138712
rect 375472 138660 375524 138712
rect 172060 137912 172112 137964
rect 182824 137912 182876 137964
rect 444840 137912 444892 137964
rect 448704 137912 448756 137964
rect 171692 137844 171744 137896
rect 175924 137844 175976 137896
rect 176016 136620 176068 136672
rect 197360 136620 197412 136672
rect 172244 136552 172296 136604
rect 181536 136552 181588 136604
rect 172428 136484 172480 136536
rect 174544 136484 174596 136536
rect 444380 136280 444432 136332
rect 444564 136280 444616 136332
rect 447140 136280 447192 136332
rect 171876 136212 171928 136264
rect 179420 136212 179472 136264
rect 172520 135872 172572 135924
rect 197728 135872 197780 135924
rect 171692 135124 171744 135176
rect 178040 135124 178092 135176
rect 172520 134512 172572 134564
rect 197360 134512 197412 134564
rect 172060 134240 172112 134292
rect 176016 134240 176068 134292
rect 444472 133152 444524 133204
rect 458180 133152 458232 133204
rect 171140 132472 171192 132524
rect 197360 132472 197412 132524
rect 445668 132404 445720 132456
rect 454224 132404 454276 132456
rect 172428 131044 172480 131096
rect 197360 131044 197412 131096
rect 444840 130432 444892 130484
rect 451280 130432 451332 130484
rect 172428 130024 172480 130076
rect 175280 130024 175332 130076
rect 171876 129752 171928 129804
rect 176660 129752 176712 129804
rect 171508 129684 171560 129736
rect 197360 129684 197412 129736
rect 444840 129684 444892 129736
rect 456800 129684 456852 129736
rect 369860 129548 369912 129600
rect 374000 129548 374052 129600
rect 375288 129548 375340 129600
rect 375288 129072 375340 129124
rect 429200 129072 429252 129124
rect 370228 129004 370280 129056
rect 371700 129004 371752 129056
rect 430580 129004 430632 129056
rect 171876 128528 171928 128580
rect 174452 128528 174504 128580
rect 171508 128460 171560 128512
rect 173164 128460 173216 128512
rect 174452 127576 174504 127628
rect 198004 127576 198056 127628
rect 172428 127032 172480 127084
rect 182824 127032 182876 127084
rect 171692 126964 171744 127016
rect 191104 126964 191156 127016
rect 443644 126964 443696 127016
rect 452660 126964 452712 127016
rect 176660 126896 176712 126948
rect 198464 126896 198516 126948
rect 443276 126216 443328 126268
rect 447232 126216 447284 126268
rect 371240 126012 371292 126064
rect 441804 126012 441856 126064
rect 371792 125944 371844 125996
rect 443644 125944 443696 125996
rect 371516 125876 371568 125928
rect 443000 125876 443052 125928
rect 172336 125740 172388 125792
rect 180064 125740 180116 125792
rect 172428 125672 172480 125724
rect 178684 125672 178736 125724
rect 172060 125604 172112 125656
rect 181444 125604 181496 125656
rect 175280 125536 175332 125588
rect 197544 125536 197596 125588
rect 371240 125468 371292 125520
rect 374092 125468 374144 125520
rect 441804 125468 441856 125520
rect 429200 125400 429252 125452
rect 444564 125400 444616 125452
rect 430580 125332 430632 125384
rect 444748 125332 444800 125384
rect 372528 125264 372580 125316
rect 441896 125264 441948 125316
rect 302608 125196 302660 125248
rect 370228 125196 370280 125248
rect 172428 125128 172480 125180
rect 177304 125128 177356 125180
rect 302976 125128 303028 125180
rect 369860 125128 369912 125180
rect 302792 125060 302844 125112
rect 370044 125060 370096 125112
rect 302884 124992 302936 125044
rect 369952 124992 370004 125044
rect 359464 124856 359516 124908
rect 369308 124856 369360 124908
rect 372436 124856 372488 124908
rect 441804 124856 441856 124908
rect 445852 124856 445904 124908
rect 171324 124584 171376 124636
rect 175924 124584 175976 124636
rect 171968 124176 172020 124228
rect 174544 124176 174596 124228
rect 302792 124108 302844 124160
rect 371608 124108 371660 124160
rect 444472 124108 444524 124160
rect 367652 124040 367704 124092
rect 369400 124040 369452 124092
rect 437204 124040 437256 124092
rect 443184 124040 443236 124092
rect 302976 123564 303028 123616
rect 370412 123564 370464 123616
rect 302884 123428 302936 123480
rect 370228 123428 370280 123480
rect 162860 122884 162912 122936
rect 188344 122884 188396 122936
rect 160928 122816 160980 122868
rect 198832 122816 198884 122868
rect 166908 122748 166960 122800
rect 170404 122748 170456 122800
rect 164884 122612 164936 122664
rect 184204 122748 184256 122800
rect 322204 122748 322256 122800
rect 438860 122748 438912 122800
rect 168932 122544 168984 122596
rect 186964 122680 187016 122732
rect 320824 122680 320876 122732
rect 366916 122680 366968 122732
rect 435180 122680 435232 122732
rect 441712 122680 441764 122732
rect 173164 121388 173216 121440
rect 197544 121388 197596 121440
rect 302516 121388 302568 121440
rect 370320 121388 370372 121440
rect 171784 118600 171836 118652
rect 197912 118600 197964 118652
rect 302792 117240 302844 117292
rect 367652 117240 367704 117292
rect 191104 116628 191156 116680
rect 198372 116628 198424 116680
rect 182824 114452 182876 114504
rect 197360 114452 197412 114504
rect 307024 113092 307076 113144
rect 579804 113092 579856 113144
rect 3424 111732 3476 111784
rect 159364 111732 159416 111784
rect 181444 111732 181496 111784
rect 197360 111732 197412 111784
rect 302792 111732 302844 111784
rect 369952 111732 370004 111784
rect 180064 110372 180116 110424
rect 197360 110372 197412 110424
rect 302792 108944 302844 108996
rect 359464 108944 359516 108996
rect 178684 107584 178736 107636
rect 198556 107584 198608 107636
rect 177304 106224 177356 106276
rect 197544 106224 197596 106276
rect 175924 103436 175976 103488
rect 197912 103436 197964 103488
rect 302792 102756 302844 102808
rect 369860 102756 369912 102808
rect 174544 102076 174596 102128
rect 197544 102076 197596 102128
rect 300216 101328 300268 101380
rect 301504 101328 301556 101380
rect 316684 100648 316736 100700
rect 580172 100648 580224 100700
rect 258172 100240 258224 100292
rect 339500 100240 339552 100292
rect 255780 100172 255832 100224
rect 323584 100172 323636 100224
rect 260748 100104 260800 100156
rect 353944 100104 353996 100156
rect 195244 100036 195296 100088
rect 299572 100036 299624 100088
rect 106188 99968 106240 100020
rect 217968 99968 218020 100020
rect 264980 99968 265032 100020
rect 376024 99968 376076 100020
rect 124864 99900 124916 99952
rect 212816 99900 212868 99952
rect 270592 99900 270644 99952
rect 412640 99900 412692 99952
rect 108304 99832 108356 99884
rect 215208 99832 215260 99884
rect 271144 99832 271196 99884
rect 414664 99832 414716 99884
rect 111064 99764 111116 99816
rect 218428 99764 218480 99816
rect 272432 99764 272484 99816
rect 423680 99764 423732 99816
rect 93124 99696 93176 99748
rect 213368 99696 213420 99748
rect 273628 99696 273680 99748
rect 430580 99696 430632 99748
rect 87604 99628 87656 99680
rect 210792 99628 210844 99680
rect 274824 99628 274876 99680
rect 435364 99628 435416 99680
rect 91008 99560 91060 99612
rect 215392 99560 215444 99612
rect 275468 99560 275520 99612
rect 440240 99560 440292 99612
rect 72424 99492 72476 99544
rect 211160 99492 211212 99544
rect 276020 99492 276072 99544
rect 442264 99492 442316 99544
rect 53104 99424 53156 99476
rect 208400 99424 208452 99476
rect 278504 99424 278556 99476
rect 457444 99424 457496 99476
rect 39304 99356 39356 99408
rect 203708 99356 203760 99408
rect 279700 99356 279752 99408
rect 464344 99356 464396 99408
rect 180708 99288 180760 99340
rect 230756 99288 230808 99340
rect 282920 99288 282972 99340
rect 316684 99288 316736 99340
rect 174544 99220 174596 99272
rect 229560 99220 229612 99272
rect 265532 99220 265584 99272
rect 311164 99220 311216 99272
rect 152556 99152 152608 99204
rect 225328 99152 225380 99204
rect 253020 99152 253072 99204
rect 309140 99152 309192 99204
rect 134524 99084 134576 99136
rect 222292 99084 222344 99136
rect 253572 99084 253624 99136
rect 312544 99084 312596 99136
rect 148324 99016 148376 99068
rect 224500 99016 224552 99068
rect 255872 99016 255924 99068
rect 324964 99016 325016 99068
rect 133788 98948 133840 99000
rect 222660 98948 222712 99000
rect 263140 98948 263192 99000
rect 360844 98948 360896 99000
rect 130384 98880 130436 98932
rect 222108 98880 222160 98932
rect 279056 98880 279108 98932
rect 460204 98880 460256 98932
rect 84108 98812 84160 98864
rect 214196 98812 214248 98864
rect 292396 98812 292448 98864
rect 485044 98812 485096 98864
rect 54484 98744 54536 98796
rect 208768 98744 208820 98796
rect 286968 98744 287020 98796
rect 507860 98744 507912 98796
rect 43444 98676 43496 98728
rect 202512 98676 202564 98728
rect 287520 98676 287572 98728
rect 512000 98676 512052 98728
rect 21364 98608 21416 98660
rect 202880 98608 202932 98660
rect 290556 98608 290608 98660
rect 529940 98608 529992 98660
rect 195888 98540 195940 98592
rect 233424 98540 233476 98592
rect 198648 98472 198700 98524
rect 234804 98472 234856 98524
rect 254952 98336 255004 98388
rect 320180 98132 320232 98184
rect 188988 97996 189040 98048
rect 212540 97996 212592 98048
rect 3424 97928 3476 97980
rect 14464 97928 14516 97980
rect 191104 97928 191156 97980
rect 214012 97928 214064 97980
rect 257252 97928 257304 97980
rect 333980 98064 334032 98116
rect 261484 97928 261536 97980
rect 358820 97996 358872 98048
rect 277584 97928 277636 97980
rect 322204 97928 322256 97980
rect 184204 97860 184256 97912
rect 217692 97860 217744 97912
rect 274640 97860 274692 97912
rect 182824 97792 182876 97844
rect 220084 97792 220136 97844
rect 268568 97792 268620 97844
rect 280712 97860 280764 97912
rect 329104 97860 329156 97912
rect 173808 97724 173860 97776
rect 206100 97724 206152 97776
rect 207756 97724 207808 97776
rect 218888 97724 218940 97776
rect 238024 97724 238076 97776
rect 239496 97724 239548 97776
rect 264336 97724 264388 97776
rect 268384 97724 268436 97776
rect 269764 97724 269816 97776
rect 121368 97656 121420 97708
rect 112444 97588 112496 97640
rect 207756 97588 207808 97640
rect 220636 97656 220688 97708
rect 245568 97656 245620 97708
rect 253296 97656 253348 97708
rect 262496 97656 262548 97708
rect 271236 97656 271288 97708
rect 336004 97792 336056 97844
rect 280804 97724 280856 97776
rect 342904 97724 342956 97776
rect 218060 97588 218112 97640
rect 228180 97588 228232 97640
rect 252376 97588 252428 97640
rect 263784 97588 263836 97640
rect 270408 97588 270460 97640
rect 276572 97588 276624 97640
rect 393964 97656 394016 97708
rect 400864 97588 400916 97640
rect 97264 97520 97316 97572
rect 216404 97520 216456 97572
rect 216772 97520 216824 97572
rect 230020 97520 230072 97572
rect 247316 97520 247368 97572
rect 255964 97520 256016 97572
rect 260840 97520 260892 97572
rect 271512 97520 271564 97572
rect 275836 97520 275888 97572
rect 436744 97520 436796 97572
rect 58624 97452 58676 97504
rect 206744 97452 206796 97504
rect 218152 97452 218204 97504
rect 230572 97452 230624 97504
rect 235816 97452 235868 97504
rect 238852 97452 238904 97504
rect 266728 97452 266780 97504
rect 271144 97452 271196 97504
rect 271604 97452 271656 97504
rect 276112 97452 276164 97504
rect 277032 97452 277084 97504
rect 443644 97452 443696 97504
rect 56508 97384 56560 97436
rect 209596 97384 209648 97436
rect 210424 97384 210476 97436
rect 221280 97384 221332 97436
rect 224868 97384 224920 97436
rect 238300 97384 238352 97436
rect 249800 97384 249852 97436
rect 267004 97384 267056 97436
rect 272156 97384 272208 97436
rect 275376 97384 275428 97436
rect 278228 97384 278280 97436
rect 447784 97384 447836 97436
rect 40684 97316 40736 97368
rect 204076 97316 204128 97368
rect 209412 97316 209464 97368
rect 227352 97316 227404 97368
rect 228548 97316 228600 97368
rect 237012 97316 237064 97368
rect 242716 97316 242768 97368
rect 263600 97316 263652 97368
rect 263692 97316 263744 97368
rect 278044 97316 278096 97368
rect 279516 97316 279568 97368
rect 450544 97316 450596 97368
rect 14556 97248 14608 97300
rect 201040 97248 201092 97300
rect 192576 97180 192628 97232
rect 205548 97248 205600 97300
rect 211160 97248 211212 97300
rect 233608 97248 233660 97300
rect 247592 97248 247644 97300
rect 269764 97248 269816 97300
rect 272800 97248 272852 97300
rect 280804 97248 280856 97300
rect 280896 97248 280948 97300
rect 281264 97248 281316 97300
rect 289360 97248 289412 97300
rect 289728 97248 289780 97300
rect 291844 97248 291896 97300
rect 454684 97248 454736 97300
rect 204904 97180 204956 97232
rect 221464 97180 221516 97232
rect 235632 97180 235684 97232
rect 239312 97180 239364 97232
rect 267372 97180 267424 97232
rect 312636 97180 312688 97232
rect 199384 97112 199436 97164
rect 212172 97112 212224 97164
rect 212540 97112 212592 97164
rect 232228 97112 232280 97164
rect 243544 97112 243596 97164
rect 249064 97112 249116 97164
rect 250352 97112 250404 97164
rect 291752 97112 291804 97164
rect 293592 97112 293644 97164
rect 293868 97112 293920 97164
rect 296260 97112 296312 97164
rect 296444 97112 296496 97164
rect 198004 97044 198056 97096
rect 210976 97044 211028 97096
rect 220636 97044 220688 97096
rect 228732 97044 228784 97096
rect 232780 97044 232832 97096
rect 238668 97044 238720 97096
rect 242900 97044 242952 97096
rect 250444 97044 250496 97096
rect 259460 97044 259512 97096
rect 260564 97044 260616 97096
rect 261852 97044 261904 97096
rect 262128 97044 262180 97096
rect 273444 97044 273496 97096
rect 275284 97044 275336 97096
rect 275376 97044 275428 97096
rect 280712 97044 280764 97096
rect 281080 97044 281132 97096
rect 281448 97044 281500 97096
rect 283932 97044 283984 97096
rect 284208 97044 284260 97096
rect 203524 96976 203576 97028
rect 207940 96976 207992 97028
rect 214564 96976 214616 97028
rect 217048 96976 217100 97028
rect 223580 96976 223632 97028
rect 225144 96976 225196 97028
rect 233516 96976 233568 97028
rect 234344 96976 234396 97028
rect 242072 96976 242124 97028
rect 242808 96976 242860 97028
rect 247960 96976 248012 97028
rect 248144 96976 248196 97028
rect 248328 96976 248380 97028
rect 280804 96976 280856 97028
rect 281724 96976 281776 97028
rect 282736 96976 282788 97028
rect 283104 96976 283156 97028
rect 284116 96976 284168 97028
rect 284300 96976 284352 97028
rect 285404 96976 285456 97028
rect 285956 96976 286008 97028
rect 286692 96976 286744 97028
rect 200396 96908 200448 96960
rect 201132 96908 201184 96960
rect 201592 96908 201644 96960
rect 202144 96908 202196 96960
rect 204628 96908 204680 96960
rect 205180 96908 205232 96960
rect 218336 96908 218388 96960
rect 219164 96908 219216 96960
rect 219808 96908 219860 96960
rect 220360 96908 220412 96960
rect 222568 96908 222620 96960
rect 223028 96908 223080 96960
rect 225236 96908 225288 96960
rect 225604 96908 225656 96960
rect 226616 96908 226668 96960
rect 226892 96908 226944 96960
rect 228088 96908 228140 96960
rect 228456 96908 228508 96960
rect 229468 96908 229520 96960
rect 230296 96908 230348 96960
rect 230848 96908 230900 96960
rect 231492 96908 231544 96960
rect 233884 96908 233936 96960
rect 234620 96908 234672 96960
rect 240140 96908 240192 96960
rect 241060 96908 241112 96960
rect 241888 96908 241940 96960
rect 242440 96908 242492 96960
rect 242624 96908 242676 96960
rect 243268 96908 243320 96960
rect 244280 96908 244332 96960
rect 245292 96908 245344 96960
rect 247776 96908 247828 96960
rect 248236 96908 248288 96960
rect 248972 96908 249024 96960
rect 249340 96908 249392 96960
rect 249432 96908 249484 96960
rect 249616 96908 249668 96960
rect 249984 96908 250036 96960
rect 250812 96908 250864 96960
rect 252008 96908 252060 96960
rect 252192 96908 252244 96960
rect 253204 96908 253256 96960
rect 253664 96908 253716 96960
rect 254216 96908 254268 96960
rect 254860 96908 254912 96960
rect 256884 96908 256936 96960
rect 257712 96908 257764 96960
rect 258264 96908 258316 96960
rect 258908 96908 258960 96960
rect 259092 96908 259144 96960
rect 259368 96908 259420 96960
rect 260104 96908 260156 96960
rect 260472 96908 260524 96960
rect 261668 96908 261720 96960
rect 262036 96908 262088 96960
rect 264152 96908 264204 96960
rect 264704 96908 264756 96960
rect 265716 96908 265768 96960
rect 265992 96908 266044 96960
rect 266360 96908 266412 96960
rect 267372 96908 267424 96960
rect 268200 96908 268252 96960
rect 268936 96908 268988 96960
rect 269396 96908 269448 96960
rect 269948 96908 270000 96960
rect 271420 96908 271472 96960
rect 271788 96908 271840 96960
rect 272616 96908 272668 96960
rect 273076 96908 273128 96960
rect 273812 96908 273864 96960
rect 274364 96908 274416 96960
rect 204444 96840 204496 96892
rect 204996 96840 205048 96892
rect 219624 96840 219676 96892
rect 220176 96840 220228 96892
rect 222384 96840 222436 96892
rect 223396 96840 223448 96892
rect 225420 96840 225472 96892
rect 226064 96840 226116 96892
rect 226800 96840 226852 96892
rect 227444 96840 227496 96892
rect 227904 96840 227956 96892
rect 228824 96840 228876 96892
rect 231032 96840 231084 96892
rect 231308 96840 231360 96892
rect 233332 96840 233384 96892
rect 234068 96840 234120 96892
rect 237380 96840 237432 96892
rect 240508 96840 240560 96892
rect 242256 96840 242308 96892
rect 242716 96840 242768 96892
rect 243084 96840 243136 96892
rect 244096 96840 244148 96892
rect 244740 96840 244792 96892
rect 245568 96840 245620 96892
rect 247132 96840 247184 96892
rect 248144 96840 248196 96892
rect 251364 96840 251416 96892
rect 252284 96840 252336 96892
rect 252836 96840 252888 96892
rect 253572 96840 253624 96892
rect 254768 96840 254820 96892
rect 255228 96840 255280 96892
rect 257068 96840 257120 96892
rect 257896 96840 257948 96892
rect 260288 96840 260340 96892
rect 260748 96840 260800 96892
rect 263876 96840 263928 96892
rect 264888 96840 264940 96892
rect 265348 96840 265400 96892
rect 266176 96840 266228 96892
rect 266912 96840 266964 96892
rect 267648 96840 267700 96892
rect 270960 96840 271012 96892
rect 200856 96772 200908 96824
rect 207388 96772 207440 96824
rect 216864 96772 216916 96824
rect 217140 96772 217192 96824
rect 229744 96772 229796 96824
rect 233976 96772 234028 96824
rect 235080 96772 235132 96824
rect 235540 96772 235592 96824
rect 236368 96772 236420 96824
rect 237104 96772 237156 96824
rect 244556 96772 244608 96824
rect 245108 96772 245160 96824
rect 248604 96772 248656 96824
rect 249616 96772 249668 96824
rect 251548 96772 251600 96824
rect 252376 96772 252428 96824
rect 252560 96772 252612 96824
rect 253848 96772 253900 96824
rect 254032 96772 254084 96824
rect 254952 96772 255004 96824
rect 257436 96772 257488 96824
rect 257804 96772 257856 96824
rect 258632 96772 258684 96824
rect 259092 96772 259144 96824
rect 259644 96772 259696 96824
rect 260656 96772 260708 96824
rect 261116 96772 261168 96824
rect 261944 96772 261996 96824
rect 262312 96772 262364 96824
rect 263140 96772 263192 96824
rect 265164 96772 265216 96824
rect 266268 96772 266320 96824
rect 266544 96772 266596 96824
rect 267556 96772 267608 96824
rect 269580 96772 269632 96824
rect 270316 96772 270368 96824
rect 270776 96772 270828 96824
rect 271696 96772 271748 96824
rect 271972 96840 272024 96892
rect 272984 96840 273036 96892
rect 273996 96840 274048 96892
rect 274548 96840 274600 96892
rect 277584 96908 277636 96960
rect 277676 96908 277728 96960
rect 278320 96908 278372 96960
rect 278872 96908 278924 96960
rect 279792 96908 279844 96960
rect 282276 96908 282328 96960
rect 282644 96908 282696 96960
rect 283472 96908 283524 96960
rect 283932 96908 283984 96960
rect 284760 96908 284812 96960
rect 285312 96908 285364 96960
rect 286508 96908 286560 96960
rect 286784 96908 286836 96960
rect 276112 96840 276164 96892
rect 304356 97044 304408 97096
rect 287152 96976 287204 97028
rect 288348 96976 288400 97028
rect 291568 96976 291620 97028
rect 292396 96976 292448 97028
rect 292764 96976 292816 97028
rect 293776 96976 293828 97028
rect 294052 96976 294104 97028
rect 295064 96976 295116 97028
rect 287336 96908 287388 96960
rect 287888 96908 287940 96960
rect 288992 96908 289044 96960
rect 289544 96908 289596 96960
rect 290188 96908 290240 96960
rect 291108 96908 291160 96960
rect 292028 96908 292080 96960
rect 292304 96908 292356 96960
rect 293224 96908 293276 96960
rect 293592 96908 293644 96960
rect 294420 96908 294472 96960
rect 294880 96908 294932 96960
rect 295432 96908 295484 96960
rect 298376 96908 298428 96960
rect 298468 96908 298520 96960
rect 299020 96908 299072 96960
rect 287796 96840 287848 96892
rect 288072 96840 288124 96892
rect 290832 96840 290884 96892
rect 291016 96840 291068 96892
rect 291384 96840 291436 96892
rect 292212 96840 292264 96892
rect 292580 96840 292632 96892
rect 293408 96840 293460 96892
rect 294788 96840 294840 96892
rect 295248 96840 295300 96892
rect 295800 96840 295852 96892
rect 296536 96840 296588 96892
rect 298100 96840 298152 96892
rect 301504 96840 301556 96892
rect 275008 96772 275060 96824
rect 275744 96772 275796 96824
rect 276204 96772 276256 96824
rect 276940 96772 276992 96824
rect 277492 96772 277544 96824
rect 278412 96772 278464 96824
rect 280436 96772 280488 96824
rect 281264 96772 281316 96824
rect 286140 96772 286192 96824
rect 286876 96772 286928 96824
rect 215944 96704 215996 96756
rect 218244 96704 218296 96756
rect 231124 96704 231176 96756
rect 236092 96704 236144 96756
rect 245752 96704 245804 96756
rect 250168 96704 250220 96756
rect 250904 96704 250956 96756
rect 261300 96704 261352 96756
rect 261852 96704 261904 96756
rect 267740 96704 267792 96756
rect 268568 96704 268620 96756
rect 269212 96704 269264 96756
rect 273904 96704 273956 96756
rect 275192 96704 275244 96756
rect 275928 96704 275980 96756
rect 276664 96704 276716 96756
rect 277308 96704 277360 96756
rect 280620 96704 280672 96756
rect 291844 96772 291896 96824
rect 295616 96772 295668 96824
rect 296352 96772 296404 96824
rect 290372 96704 290424 96756
rect 291016 96704 291068 96756
rect 210516 96636 210568 96688
rect 211620 96636 211672 96688
rect 233976 96636 234028 96688
rect 238116 96636 238168 96688
rect 245936 96636 245988 96688
rect 246764 96636 246816 96688
rect 246856 96636 246908 96688
rect 267924 96636 267976 96688
rect 269028 96636 269080 96688
rect 280252 96636 280304 96688
rect 281448 96636 281500 96688
rect 288532 96636 288584 96688
rect 289268 96636 289320 96688
rect 298284 96636 298336 96688
rect 299204 96636 299256 96688
rect 191196 96568 191248 96620
rect 232044 96568 232096 96620
rect 251180 96568 251232 96620
rect 302332 96568 302384 96620
rect 176568 96500 176620 96552
rect 216772 96500 216824 96552
rect 271512 96500 271564 96552
rect 356060 96500 356112 96552
rect 186964 96432 187016 96484
rect 231768 96432 231820 96484
rect 262128 96432 262180 96484
rect 347044 96432 347096 96484
rect 161388 96364 161440 96416
rect 209412 96364 209464 96416
rect 284208 96364 284260 96416
rect 411904 96364 411956 96416
rect 169668 96296 169720 96348
rect 220636 96296 220688 96348
rect 285128 96296 285180 96348
rect 465724 96296 465776 96348
rect 165528 96228 165580 96280
rect 218060 96228 218112 96280
rect 283288 96228 283340 96280
rect 475384 96228 475436 96280
rect 173164 96160 173216 96212
rect 229376 96160 229428 96212
rect 282092 96160 282144 96212
rect 479524 96160 479576 96212
rect 166264 96092 166316 96144
rect 225972 96092 226024 96144
rect 297456 96092 297508 96144
rect 494060 96092 494112 96144
rect 126888 96024 126940 96076
rect 204904 96024 204956 96076
rect 213184 96024 213236 96076
rect 236000 96024 236052 96076
rect 243912 96024 243964 96076
rect 269120 96024 269172 96076
rect 282828 96024 282880 96076
rect 483020 96024 483072 96076
rect 37188 95956 37240 96008
rect 173808 95956 173860 96008
rect 183468 95956 183520 96008
rect 231216 95956 231268 96008
rect 237748 95956 237800 96008
rect 238392 95956 238444 96008
rect 246304 95956 246356 96008
rect 281540 95956 281592 96008
rect 285864 95956 285916 96008
rect 500960 95956 501012 96008
rect 12256 95888 12308 95940
rect 202052 95888 202104 95940
rect 202144 95888 202196 95940
rect 234252 95888 234304 95940
rect 247960 95888 248012 95940
rect 285772 95888 285824 95940
rect 291200 95888 291252 95940
rect 532700 95888 532752 95940
rect 179328 95820 179380 95872
rect 218152 95820 218204 95872
rect 231216 95820 231268 95872
rect 236644 95820 236696 95872
rect 251824 95820 251876 95872
rect 302240 95820 302292 95872
rect 195244 95752 195296 95804
rect 232964 95752 233016 95804
rect 250536 95752 250588 95804
rect 299572 95752 299624 95804
rect 197268 95684 197320 95736
rect 211160 95684 211212 95736
rect 293868 95684 293920 95736
rect 320824 95684 320876 95736
rect 235356 95412 235408 95464
rect 235816 95412 235868 95464
rect 233148 95276 233200 95328
rect 239680 95276 239732 95328
rect 162768 95140 162820 95192
rect 227720 95140 227772 95192
rect 255412 95140 255464 95192
rect 324412 95140 324464 95192
rect 158628 95072 158680 95124
rect 226984 95072 227036 95124
rect 256056 95072 256108 95124
rect 327080 95072 327132 95124
rect 155224 95004 155276 95056
rect 226340 95004 226392 95056
rect 258448 95004 258500 95056
rect 340880 95004 340932 95056
rect 147588 94936 147640 94988
rect 223580 94936 223632 94988
rect 262680 94936 262732 94988
rect 364984 94936 365036 94988
rect 146208 94868 146260 94920
rect 224960 94868 225012 94920
rect 276480 94868 276532 94920
rect 385684 94868 385736 94920
rect 137284 94800 137336 94852
rect 223304 94800 223356 94852
rect 279240 94800 279292 94852
rect 429844 94800 429896 94852
rect 114468 94732 114520 94784
rect 219440 94732 219492 94784
rect 277860 94732 277912 94784
rect 453304 94732 453356 94784
rect 79324 94664 79376 94716
rect 205640 94664 205692 94716
rect 53748 94596 53800 94648
rect 209136 94664 209188 94716
rect 288164 94664 288216 94716
rect 489184 94664 489236 94716
rect 50988 94528 51040 94580
rect 208584 94596 208636 94648
rect 240692 94596 240744 94648
rect 251272 94596 251324 94648
rect 286324 94596 286376 94648
rect 502984 94596 503036 94648
rect 209964 94528 210016 94580
rect 210332 94528 210384 94580
rect 211436 94528 211488 94580
rect 211896 94528 211948 94580
rect 212908 94528 212960 94580
rect 213736 94528 213788 94580
rect 228364 94528 228416 94580
rect 234804 94528 234856 94580
rect 237564 94528 237616 94580
rect 237932 94528 237984 94580
rect 288808 94528 288860 94580
rect 518900 94528 518952 94580
rect 48228 94460 48280 94512
rect 208124 94460 208176 94512
rect 226984 94460 227036 94512
rect 237656 94460 237708 94512
rect 248788 94460 248840 94512
rect 288440 94460 288492 94512
rect 289728 94460 289780 94512
rect 520924 94460 520976 94512
rect 177948 94392 178000 94444
rect 230204 94392 230256 94444
rect 254400 94392 254452 94444
rect 317420 94392 317472 94444
rect 192484 94324 192536 94376
rect 232596 94324 232648 94376
rect 263784 94324 263836 94376
rect 306380 94324 306432 94376
rect 200028 94256 200080 94308
rect 235172 94256 235224 94308
rect 263508 94256 263560 94308
rect 304264 94256 304316 94308
rect 205640 94188 205692 94240
rect 213000 94188 213052 94240
rect 205824 94120 205876 94172
rect 206836 94120 206888 94172
rect 235908 93848 235960 93900
rect 240232 93848 240284 93900
rect 181444 93780 181496 93832
rect 229652 93780 229704 93832
rect 259368 93780 259420 93832
rect 345020 93780 345072 93832
rect 170404 93712 170456 93764
rect 227904 93712 227956 93764
rect 260748 93712 260800 93764
rect 351920 93712 351972 93764
rect 166908 93644 166960 93696
rect 228272 93644 228324 93696
rect 261760 93644 261812 93696
rect 362960 93644 363012 93696
rect 142068 93576 142120 93628
rect 224132 93576 224184 93628
rect 266268 93576 266320 93628
rect 378784 93576 378836 93628
rect 135168 93508 135220 93560
rect 222752 93508 222804 93560
rect 268936 93508 268988 93560
rect 398840 93508 398892 93560
rect 128268 93440 128320 93492
rect 221740 93440 221792 93492
rect 277308 93440 277360 93492
rect 448520 93440 448572 93492
rect 65524 93372 65576 93424
rect 210056 93372 210108 93424
rect 279884 93372 279936 93424
rect 466460 93372 466512 93424
rect 61384 93304 61436 93356
rect 209228 93304 209280 93356
rect 291936 93304 291988 93356
rect 524420 93304 524472 93356
rect 33048 93236 33100 93288
rect 192576 93236 192628 93288
rect 194508 93236 194560 93288
rect 234068 93236 234120 93288
rect 291108 93236 291160 93288
rect 525064 93236 525116 93288
rect 25504 93168 25556 93220
rect 200488 93168 200540 93220
rect 296628 93168 296680 93220
rect 538864 93168 538916 93220
rect 15844 93100 15896 93152
rect 201500 93100 201552 93152
rect 228456 93100 228508 93152
rect 237932 93100 237984 93152
rect 238668 93100 238720 93152
rect 241704 93100 241756 93152
rect 245476 93100 245528 93152
rect 255964 93100 256016 93152
rect 295248 93100 295300 93152
rect 554780 93100 554832 93152
rect 184848 93032 184900 93084
rect 231032 93032 231084 93084
rect 257988 93032 258040 93084
rect 338120 93032 338172 93084
rect 188344 92964 188396 93016
rect 231952 92964 232004 93016
rect 256516 92964 256568 93016
rect 331220 92964 331272 93016
rect 197176 92896 197228 92948
rect 233700 92896 233752 92948
rect 253848 92896 253900 92948
rect 307024 92896 307076 92948
rect 234528 92488 234580 92540
rect 239956 92488 240008 92540
rect 164148 92420 164200 92472
rect 227996 92420 228048 92472
rect 263324 92420 263376 92472
rect 369860 92420 369912 92472
rect 160008 92352 160060 92404
rect 227076 92352 227128 92404
rect 264612 92352 264664 92404
rect 374644 92352 374696 92404
rect 156696 92284 156748 92336
rect 226892 92284 226944 92336
rect 269028 92284 269080 92336
rect 381544 92284 381596 92336
rect 148968 92216 149020 92268
rect 225512 92216 225564 92268
rect 252192 92216 252244 92268
rect 303620 92216 303672 92268
rect 304356 92216 304408 92268
rect 418160 92216 418212 92268
rect 144828 92148 144880 92200
rect 224592 92148 224644 92200
rect 265992 92148 266044 92200
rect 382924 92148 382976 92200
rect 142804 92080 142856 92132
rect 222384 92080 222436 92132
rect 267372 92080 267424 92132
rect 387800 92080 387852 92132
rect 98644 92012 98696 92064
rect 216680 92012 216732 92064
rect 267648 92012 267700 92064
rect 389824 92012 389876 92064
rect 71044 91944 71096 91996
rect 210608 91944 210660 91996
rect 269948 91944 270000 91996
rect 405740 91944 405792 91996
rect 70308 91876 70360 91928
rect 211804 91876 211856 91928
rect 272892 91876 272944 91928
rect 421564 91876 421616 91928
rect 46848 91808 46900 91860
rect 203524 91808 203576 91860
rect 244004 91808 244056 91860
rect 263692 91808 263744 91860
rect 281080 91808 281132 91860
rect 471244 91808 471296 91860
rect 34428 91740 34480 91792
rect 205732 91740 205784 91792
rect 222844 91740 222896 91792
rect 235724 91740 235776 91792
rect 245568 91740 245620 91792
rect 266452 91740 266504 91792
rect 290924 91740 290976 91792
rect 529204 91740 529256 91792
rect 171048 91672 171100 91724
rect 229192 91672 229244 91724
rect 257712 91672 257764 91724
rect 330484 91672 330536 91724
rect 182088 91604 182140 91656
rect 230940 91604 230992 91656
rect 231308 91060 231360 91112
rect 236184 91060 236236 91112
rect 187056 90992 187108 91044
rect 230848 90992 230900 91044
rect 267464 90992 267516 91044
rect 394700 90992 394752 91044
rect 169024 90924 169076 90976
rect 228088 90924 228140 90976
rect 268752 90924 268804 90976
rect 396724 90924 396776 90976
rect 139308 90856 139360 90908
rect 223764 90856 223816 90908
rect 270224 90856 270276 90908
rect 407764 90856 407816 90908
rect 137376 90788 137428 90840
rect 222568 90788 222620 90840
rect 271604 90788 271656 90840
rect 417424 90788 417476 90840
rect 116584 90720 116636 90772
rect 219716 90720 219768 90772
rect 274272 90720 274324 90772
rect 432604 90720 432656 90772
rect 95148 90652 95200 90704
rect 215760 90652 215812 90704
rect 277124 90652 277176 90704
rect 446404 90652 446456 90704
rect 86868 90584 86920 90636
rect 214748 90584 214800 90636
rect 281448 90584 281500 90636
rect 467104 90584 467156 90636
rect 80704 90516 80756 90568
rect 213460 90516 213512 90568
rect 283932 90516 283984 90568
rect 486424 90516 486476 90568
rect 76564 90448 76616 90500
rect 212264 90448 212316 90500
rect 253296 90448 253348 90500
rect 266360 90448 266412 90500
rect 288348 90448 288400 90500
rect 504364 90448 504416 90500
rect 57888 90380 57940 90432
rect 209688 90380 209740 90432
rect 246212 90380 246264 90432
rect 268384 90380 268436 90432
rect 293408 90380 293460 90432
rect 540244 90380 540296 90432
rect 45468 90312 45520 90364
rect 207480 90312 207532 90364
rect 248144 90312 248196 90364
rect 280252 90312 280304 90364
rect 297180 90312 297232 90364
rect 566464 90312 566516 90364
rect 193128 90244 193180 90296
rect 232136 90244 232188 90296
rect 255136 90244 255188 90296
rect 321560 90244 321612 90296
rect 253572 90176 253624 90228
rect 309232 90176 309284 90228
rect 250812 89972 250864 90024
rect 253204 89972 253256 90024
rect 256240 89632 256292 89684
rect 328460 89632 328512 89684
rect 266084 89564 266136 89616
rect 377404 89564 377456 89616
rect 275744 89496 275796 89548
rect 438860 89496 438912 89548
rect 122748 89428 122800 89480
rect 221004 89428 221056 89480
rect 281172 89428 281224 89480
rect 476120 89428 476172 89480
rect 119988 89360 120040 89412
rect 219624 89360 219676 89412
rect 282644 89360 282696 89412
rect 481640 89360 481692 89412
rect 115204 89292 115256 89344
rect 218980 89292 219032 89344
rect 284024 89292 284076 89344
rect 490564 89292 490616 89344
rect 104808 89224 104860 89276
rect 217784 89224 217836 89276
rect 285312 89224 285364 89276
rect 493324 89224 493376 89276
rect 102048 89156 102100 89208
rect 216956 89156 217008 89208
rect 285220 89156 285272 89208
rect 497464 89156 497516 89208
rect 37096 89088 37148 89140
rect 206192 89088 206244 89140
rect 286692 89088 286744 89140
rect 500224 89088 500276 89140
rect 27528 89020 27580 89072
rect 204536 89020 204588 89072
rect 242440 89020 242492 89072
rect 252652 89020 252704 89072
rect 289452 89020 289504 89072
rect 522304 89020 522356 89072
rect 18604 88952 18656 89004
rect 201592 88952 201644 89004
rect 249340 88952 249392 89004
rect 285680 88952 285732 89004
rect 294880 88952 294932 89004
rect 553400 88952 553452 89004
rect 253664 88884 253716 88936
rect 310520 88884 310572 88936
rect 257804 88272 257856 88324
rect 335360 88272 335412 88324
rect 260380 88204 260432 88256
rect 353300 88204 353352 88256
rect 292212 88136 292264 88188
rect 428464 88136 428516 88188
rect 105544 88068 105596 88120
rect 215484 88068 215536 88120
rect 272984 88068 273036 88120
rect 420920 88068 420972 88120
rect 88984 88000 89036 88052
rect 208860 88000 208912 88052
rect 286784 88000 286836 88052
rect 506480 88000 506532 88052
rect 71688 87932 71740 87984
rect 199384 87932 199436 87984
rect 288072 87932 288124 87984
rect 511264 87932 511316 87984
rect 75184 87864 75236 87916
rect 212724 87864 212776 87916
rect 300308 87864 300360 87916
rect 525800 87864 525852 87916
rect 61476 87796 61528 87848
rect 210148 87796 210200 87848
rect 288256 87796 288308 87848
rect 515404 87796 515456 87848
rect 41328 87728 41380 87780
rect 205824 87728 205876 87780
rect 289544 87728 289596 87780
rect 518164 87728 518216 87780
rect 28908 87660 28960 87712
rect 196624 87660 196676 87712
rect 293592 87660 293644 87712
rect 543004 87660 543056 87712
rect 30288 87592 30340 87644
rect 204444 87592 204496 87644
rect 209044 87592 209096 87644
rect 233516 87592 233568 87644
rect 248236 87592 248288 87644
rect 287060 87592 287112 87644
rect 297916 87592 297968 87644
rect 569960 87592 570012 87644
rect 254952 87524 255004 87576
rect 316132 87524 316184 87576
rect 253756 87456 253808 87508
rect 314016 87456 314068 87508
rect 259092 86912 259144 86964
rect 342260 86912 342312 86964
rect 342904 86912 342956 86964
rect 425060 86912 425112 86964
rect 259184 86844 259236 86896
rect 346400 86844 346452 86896
rect 271236 86776 271288 86828
rect 365812 86776 365864 86828
rect 261944 86708 261996 86760
rect 357440 86708 357492 86760
rect 267556 86640 267608 86692
rect 392032 86640 392084 86692
rect 123484 86572 123536 86624
rect 219900 86572 219952 86624
rect 275836 86572 275888 86624
rect 441620 86572 441672 86624
rect 106924 86504 106976 86556
rect 210056 86504 210108 86556
rect 292304 86504 292356 86556
rect 536104 86504 536156 86556
rect 111156 86436 111208 86488
rect 218520 86436 218572 86488
rect 293684 86436 293736 86488
rect 547144 86436 547196 86488
rect 86224 86368 86276 86420
rect 214104 86368 214156 86420
rect 244096 86368 244148 86420
rect 258080 86368 258132 86420
rect 294972 86368 295024 86420
rect 556160 86368 556212 86420
rect 79416 86300 79468 86352
rect 213092 86300 213144 86352
rect 249432 86300 249484 86352
rect 291292 86300 291344 86352
rect 296352 86300 296404 86352
rect 560392 86300 560444 86352
rect 68284 86232 68336 86284
rect 211712 86232 211764 86284
rect 250904 86232 250956 86284
rect 295340 86232 295392 86284
rect 299112 86232 299164 86284
rect 582748 86232 582800 86284
rect 3148 85484 3200 85536
rect 152464 85484 152516 85536
rect 262036 85416 262088 85468
rect 360200 85416 360252 85468
rect 263140 85348 263192 85400
rect 364340 85348 364392 85400
rect 263232 85280 263284 85332
rect 367100 85280 367152 85332
rect 266176 85212 266228 85264
rect 382372 85212 382424 85264
rect 268844 85144 268896 85196
rect 402980 85144 403032 85196
rect 153108 85076 153160 85128
rect 225420 85076 225472 85128
rect 278412 85076 278464 85128
rect 452660 85076 452712 85128
rect 124128 85008 124180 85060
rect 221096 85008 221148 85060
rect 291016 85008 291068 85060
rect 528560 85008 528612 85060
rect 95056 84940 95108 84992
rect 216128 84940 216180 84992
rect 300124 84940 300176 84992
rect 565820 84940 565872 84992
rect 88248 84872 88300 84924
rect 214932 84872 214984 84924
rect 245292 84872 245344 84924
rect 262220 84872 262272 84924
rect 296444 84872 296496 84924
rect 564532 84872 564584 84924
rect 10968 84804 11020 84856
rect 201776 84804 201828 84856
rect 252284 84804 252336 84856
rect 299480 84804 299532 84856
rect 301504 84804 301556 84856
rect 572812 84804 572864 84856
rect 260472 83988 260524 84040
rect 327724 83988 327776 84040
rect 264704 83920 264756 83972
rect 374092 83920 374144 83972
rect 264796 83852 264848 83904
rect 378140 83852 378192 83904
rect 265900 83784 265952 83836
rect 385040 83784 385092 83836
rect 267280 83716 267332 83768
rect 391940 83716 391992 83768
rect 268568 83648 268620 83700
rect 396080 83648 396132 83700
rect 270316 83580 270368 83632
rect 409972 83580 410024 83632
rect 45376 83512 45428 83564
rect 207480 83512 207532 83564
rect 274364 83512 274416 83564
rect 432052 83512 432104 83564
rect 35164 83444 35216 83496
rect 204720 83444 204772 83496
rect 246580 83444 246632 83496
rect 260104 83444 260156 83496
rect 281264 83444 281316 83496
rect 470600 83444 470652 83496
rect 268660 82560 268712 82612
rect 398932 82560 398984 82612
rect 270408 82492 270460 82544
rect 409880 82492 409932 82544
rect 271696 82424 271748 82476
rect 414020 82424 414072 82476
rect 273076 82356 273128 82408
rect 423772 82356 423824 82408
rect 276940 82288 276992 82340
rect 445760 82288 445812 82340
rect 5448 82220 5500 82272
rect 200948 82220 201000 82272
rect 278504 82220 278556 82272
rect 456892 82220 456944 82272
rect 21456 82152 21508 82204
rect 203156 82152 203208 82204
rect 246672 82152 246724 82204
rect 271236 82152 271288 82204
rect 284116 82152 284168 82204
rect 485780 82152 485832 82204
rect 200764 82084 200816 82136
rect 226800 82084 226852 82136
rect 249524 82084 249576 82136
rect 278136 82084 278188 82136
rect 298008 82084 298060 82136
rect 571340 82084 571392 82136
rect 255044 81132 255096 81184
rect 318064 81132 318116 81184
rect 271788 81064 271840 81116
rect 416780 81064 416832 81116
rect 273168 80996 273220 81048
rect 427820 80996 427872 81048
rect 274456 80928 274508 80980
rect 434720 80928 434772 80980
rect 278596 80860 278648 80912
rect 459560 80860 459612 80912
rect 282736 80792 282788 80844
rect 477500 80792 477552 80844
rect 286876 80724 286928 80776
rect 503720 80724 503772 80776
rect 299204 80656 299256 80708
rect 574100 80656 574152 80708
rect 257896 79704 257948 79756
rect 331864 79704 331916 79756
rect 260564 79636 260616 79688
rect 347780 79636 347832 79688
rect 277032 79568 277084 79620
rect 448612 79568 448664 79620
rect 281356 79500 281408 79552
rect 472624 79500 472676 79552
rect 282552 79432 282604 79484
rect 481732 79432 481784 79484
rect 286600 79364 286652 79416
rect 506572 79364 506624 79416
rect 256056 79296 256108 79348
rect 276020 79296 276072 79348
rect 290832 79296 290884 79348
rect 530584 79296 530636 79348
rect 258908 78276 258960 78328
rect 340972 78276 341024 78328
rect 261852 78208 261904 78260
rect 357532 78208 357584 78260
rect 283840 78140 283892 78192
rect 490012 78140 490064 78192
rect 285404 78072 285456 78124
rect 492680 78072 492732 78124
rect 287888 78004 287940 78056
rect 510620 78004 510672 78056
rect 293776 77936 293828 77988
rect 542360 77936 542412 77988
rect 276664 76712 276716 76764
rect 411260 76712 411312 76764
rect 289268 76644 289320 76696
rect 517520 76644 517572 76696
rect 292396 76576 292448 76628
rect 535460 76576 535512 76628
rect 295064 76508 295116 76560
rect 548524 76508 548576 76560
rect 275284 75284 275336 75336
rect 429200 75284 429252 75336
rect 296536 75216 296588 75268
rect 560300 75216 560352 75268
rect 250996 75148 251048 75200
rect 298100 75148 298152 75200
rect 299296 75148 299348 75200
rect 578240 75148 578292 75200
rect 279976 73856 280028 73908
rect 467840 73856 467892 73908
rect 299388 73788 299440 73840
rect 582932 73788 582984 73840
rect 305644 73108 305696 73160
rect 579988 73108 580040 73160
rect 3424 71680 3476 71732
rect 157984 71680 158036 71732
rect 158076 71000 158128 71052
rect 226708 71000 226760 71052
rect 68928 69640 68980 69692
rect 210516 69640 210568 69692
rect 278320 69640 278372 69692
rect 454040 69640 454092 69692
rect 313924 60664 313976 60716
rect 580172 60664 580224 60716
rect 3056 59304 3108 59356
rect 146944 59304 146996 59356
rect 3424 45500 3476 45552
rect 151084 45500 151136 45552
rect 249616 39312 249668 39364
rect 284300 39312 284352 39364
rect 242532 37884 242584 37936
rect 248420 37884 248472 37936
rect 89076 35164 89128 35216
rect 214288 35164 214340 35216
rect 580264 33940 580316 33992
rect 582564 33940 582616 33992
rect 275928 33736 275980 33788
rect 440332 33736 440384 33788
rect 2872 33056 2924 33108
rect 156604 33056 156656 33108
rect 273904 32376 273956 32428
rect 404360 32376 404412 32428
rect 248052 31016 248104 31068
rect 280160 31016 280212 31068
rect 280988 31016 281040 31068
rect 474740 31016 474792 31068
rect 257620 29656 257672 29708
rect 336096 29656 336148 29708
rect 336004 29588 336056 29640
rect 436100 29588 436152 29640
rect 259000 28228 259052 28280
rect 342904 28228 342956 28280
rect 256332 26868 256384 26920
rect 329840 26868 329892 26920
rect 113088 25508 113140 25560
rect 218336 25508 218388 25560
rect 295156 25508 295208 25560
rect 556252 25508 556304 25560
rect 253480 24080 253532 24132
rect 311900 24080 311952 24132
rect 312636 24080 312688 24132
rect 393320 24080 393372 24132
rect 26148 22720 26200 22772
rect 35256 22720 35308 22772
rect 252376 22720 252428 22772
rect 300860 22720 300912 22772
rect 44088 21360 44140 21412
rect 200856 21360 200908 21412
rect 3424 20612 3476 20664
rect 144184 20612 144236 20664
rect 177856 19932 177908 19984
rect 229468 19932 229520 19984
rect 296260 19932 296312 19984
rect 564624 19932 564676 19984
rect 246764 18708 246816 18760
rect 257344 18708 257396 18760
rect 243912 18640 243964 18692
rect 255320 18640 255372 18692
rect 143448 18572 143500 18624
rect 224040 18572 224092 18624
rect 245384 18572 245436 18624
rect 260196 18572 260248 18624
rect 268476 18572 268528 18624
rect 375380 18572 375432 18624
rect 232596 17892 232648 17944
rect 236736 17892 236788 17944
rect 250444 17892 250496 17944
rect 251180 17892 251232 17944
rect 249064 17824 249116 17876
rect 253940 17824 253992 17876
rect 97356 17212 97408 17264
rect 215576 17212 215628 17264
rect 254768 17212 254820 17264
rect 322940 17212 322992 17264
rect 436744 17212 436796 17264
rect 443000 17212 443052 17264
rect 454684 17212 454736 17264
rect 471980 17212 472032 17264
rect 39396 15852 39448 15904
rect 206284 15852 206336 15904
rect 227628 15852 227680 15904
rect 232504 15852 232556 15904
rect 293500 15852 293552 15904
rect 546684 15852 546736 15904
rect 236644 15172 236696 15224
rect 239036 15172 239088 15224
rect 245108 14492 245160 14544
rect 258724 14492 258776 14544
rect 119896 14424 119948 14476
rect 219808 14424 219860 14476
rect 246856 14424 246908 14476
rect 267740 14424 267792 14476
rect 287980 14424 288032 14476
rect 514760 14424 514812 14476
rect 234068 13812 234120 13864
rect 235080 13812 235132 13864
rect 64788 13064 64840 13116
rect 198004 13064 198056 13116
rect 285496 13064 285548 13116
rect 500224 13064 500276 13116
rect 357532 11772 357584 11824
rect 358728 11772 358780 11824
rect 398932 11772 398984 11824
rect 400128 11772 400180 11824
rect 35808 11704 35860 11756
rect 206008 11704 206060 11756
rect 219348 11704 219400 11756
rect 236368 11704 236420 11756
rect 242624 11704 242676 11756
rect 252560 11704 252612 11756
rect 329104 11704 329156 11756
rect 422576 11704 422628 11756
rect 423772 11704 423824 11756
rect 424968 11704 425020 11756
rect 448612 11704 448664 11756
rect 449808 11704 449860 11756
rect 223488 10344 223540 10396
rect 233976 10344 234028 10396
rect 81348 10276 81400 10328
rect 212908 10276 212960 10328
rect 217968 10276 218020 10328
rect 228548 10276 228600 10328
rect 267004 10276 267056 10328
rect 291200 10276 291252 10328
rect 292028 10276 292080 10328
rect 539600 10276 539652 10328
rect 234160 9868 234212 9920
rect 237840 9868 237892 9920
rect 234804 9596 234856 9648
rect 237748 9596 237800 9648
rect 70216 8916 70268 8968
rect 211436 8916 211488 8968
rect 227536 8916 227588 8968
rect 235356 8916 235408 8968
rect 285128 8916 285180 8968
rect 497096 8916 497148 8968
rect 233424 8372 233476 8424
rect 239128 8372 239180 8424
rect 242716 8236 242768 8288
rect 245660 8236 245712 8288
rect 393964 8236 394016 8288
rect 401324 8236 401376 8288
rect 443644 8236 443696 8288
rect 450912 8236 450964 8288
rect 202696 7692 202748 7744
rect 233884 7692 233936 7744
rect 124680 7624 124732 7676
rect 210424 7624 210476 7676
rect 102232 7556 102284 7608
rect 217508 7556 217560 7608
rect 400864 7556 400916 7608
rect 408408 7556 408460 7608
rect 450544 7556 450596 7608
rect 465172 7556 465224 7608
rect 229836 7420 229888 7472
rect 235264 7420 235316 7472
rect 3424 6808 3476 6860
rect 129004 6808 129056 6860
rect 199108 6264 199160 6316
rect 229744 6264 229796 6316
rect 131764 6196 131816 6248
rect 222476 6196 222528 6248
rect 107016 6128 107068 6180
rect 215944 6128 215996 6180
rect 249248 6128 249300 6180
rect 287796 6128 287848 6180
rect 289360 6128 289412 6180
rect 521844 6128 521896 6180
rect 241336 5516 241388 5568
rect 241704 5516 241756 5568
rect 242808 5516 242860 5568
rect 246396 5516 246448 5568
rect 245200 5448 245252 5500
rect 251088 5448 251140 5500
rect 250720 4972 250772 5024
rect 297272 4972 297324 5024
rect 212172 4904 212224 4956
rect 231124 4904 231176 4956
rect 278044 4904 278096 4956
rect 372896 4904 372948 4956
rect 99840 4836 99892 4888
rect 214564 4836 214616 4888
rect 271144 4836 271196 4888
rect 390652 4836 390704 4888
rect 98736 4768 98788 4820
rect 217140 4768 217192 4820
rect 269764 4768 269816 4820
rect 278320 4768 278372 4820
rect 294788 4768 294840 4820
rect 553768 4768 553820 4820
rect 15936 4088 15988 4140
rect 17224 4088 17276 4140
rect 20628 4088 20680 4140
rect 21456 4088 21508 4140
rect 72608 4088 72660 4140
rect 76564 4088 76616 4140
rect 148968 4088 149020 4140
rect 149520 4088 149572 4140
rect 17040 4020 17092 4072
rect 21364 4020 21416 4072
rect 58440 4020 58492 4072
rect 65524 4020 65576 4072
rect 78588 4020 78640 4072
rect 93124 4020 93176 4072
rect 13544 3952 13596 4004
rect 18604 3952 18656 4004
rect 24216 3952 24268 4004
rect 6460 3612 6512 3664
rect 14556 3680 14608 3732
rect 11152 3612 11204 3664
rect 12256 3612 12308 3664
rect 2872 3544 2924 3596
rect 19432 3884 19484 3936
rect 25504 3748 25556 3800
rect 54944 3952 54996 4004
rect 61384 3952 61436 4004
rect 63224 3952 63276 4004
rect 87604 3952 87656 4004
rect 91652 3952 91704 4004
rect 105544 4020 105596 4072
rect 111616 4020 111668 4072
rect 115204 4020 115256 4072
rect 117596 4020 117648 4072
rect 241428 4156 241480 4208
rect 242900 4156 242952 4208
rect 154212 4088 154264 4140
rect 155224 4088 155276 4140
rect 155408 4088 155460 4140
rect 156696 4088 156748 4140
rect 160100 4088 160152 4140
rect 161388 4088 161440 4140
rect 161480 4088 161532 4140
rect 200764 4088 200816 4140
rect 219256 4088 219308 4140
rect 228456 4088 228508 4140
rect 172152 4020 172204 4072
rect 189724 4020 189776 4072
rect 191196 4020 191248 4072
rect 198648 4020 198700 4072
rect 203892 4020 203944 4072
rect 209780 4020 209832 4072
rect 222844 4020 222896 4072
rect 255964 4020 256016 4072
rect 265348 4088 265400 4140
rect 353944 4088 353996 4140
rect 355232 4088 355284 4140
rect 382924 4088 382976 4140
rect 384764 4088 384816 4140
rect 460204 4088 460256 4140
rect 462780 4088 462832 4140
rect 479524 4088 479576 4140
rect 480536 4088 480588 4140
rect 547144 4088 547196 4140
rect 549076 4088 549128 4140
rect 566556 4088 566608 4140
rect 568028 4088 568080 4140
rect 260840 4020 260892 4072
rect 263600 4020 263652 4072
rect 276020 4020 276072 4072
rect 280252 4020 280304 4072
rect 347044 4020 347096 4072
rect 362316 4020 362368 4072
rect 93952 3952 94004 4004
rect 108304 3952 108356 4004
rect 130568 3952 130620 4004
rect 134524 3952 134576 4004
rect 137652 3952 137704 4004
rect 142804 3952 142856 4004
rect 148324 3952 148376 4004
rect 152556 3952 152608 4004
rect 152648 3952 152700 4004
rect 225236 3952 225288 4004
rect 225328 3952 225380 4004
rect 228364 3952 228416 4004
rect 228732 3952 228784 4004
rect 236644 3952 236696 4004
rect 257344 3952 257396 4004
rect 268844 3952 268896 4004
rect 279516 3952 279568 4004
rect 287060 3952 287112 4004
rect 327724 3952 327776 4004
rect 351644 3952 351696 4004
rect 360844 3952 360896 4004
rect 369400 3952 369452 4004
rect 377404 3952 377456 4004
rect 387156 3952 387208 4004
rect 52552 3884 52604 3936
rect 88984 3884 89036 3936
rect 92756 3884 92808 3936
rect 97356 3884 97408 3936
rect 103336 3884 103388 3936
rect 184204 3884 184256 3936
rect 200028 3884 200080 3936
rect 207388 3884 207440 3936
rect 214472 3884 214524 3936
rect 231216 3884 231268 3936
rect 257068 3884 257120 3936
rect 269120 3884 269172 3936
rect 271328 3884 271380 3936
rect 281540 3884 281592 3936
rect 304264 3884 304316 3936
rect 371700 3884 371752 3936
rect 385684 3884 385736 3936
rect 447416 3884 447468 3936
rect 475476 3884 475528 3936
rect 487620 3884 487672 3936
rect 40684 3816 40736 3868
rect 60832 3816 60884 3868
rect 106924 3816 106976 3868
rect 140044 3816 140096 3868
rect 223856 3816 223908 3868
rect 225144 3816 225196 3868
rect 234804 3816 234856 3868
rect 260104 3816 260156 3868
rect 273628 3816 273680 3868
rect 278136 3816 278188 3868
rect 288992 3816 289044 3868
rect 29644 3748 29696 3800
rect 39580 3748 39632 3800
rect 58624 3748 58676 3800
rect 75000 3748 75052 3800
rect 124864 3748 124916 3800
rect 150624 3748 150676 3800
rect 152648 3748 152700 3800
rect 172152 3748 172204 3800
rect 182824 3748 182876 3800
rect 221556 3748 221608 3800
rect 234160 3748 234212 3800
rect 245200 3748 245252 3800
rect 252652 3748 252704 3800
rect 253204 3748 253256 3800
rect 292580 3816 292632 3868
rect 311164 3816 311216 3868
rect 383568 3816 383620 3868
rect 411904 3816 411956 3868
rect 491116 3816 491168 3868
rect 518164 3816 518216 3868
rect 520740 3816 520792 3868
rect 536104 3816 536156 3868
rect 538404 3816 538456 3868
rect 290188 3748 290240 3800
rect 291292 3748 291344 3800
rect 296076 3748 296128 3800
rect 299572 3748 299624 3800
rect 322204 3748 322256 3800
rect 415492 3748 415544 3800
rect 429844 3748 429896 3800
rect 463976 3748 464028 3800
rect 465724 3748 465776 3800
rect 498200 3748 498252 3800
rect 14740 3680 14792 3732
rect 43444 3680 43496 3732
rect 62028 3680 62080 3732
rect 71044 3680 71096 3732
rect 82084 3680 82136 3732
rect 191104 3680 191156 3732
rect 215668 3680 215720 3732
rect 232596 3680 232648 3732
rect 251088 3680 251140 3732
rect 262956 3680 263008 3732
rect 264888 3680 264940 3732
rect 374092 3680 374144 3732
rect 381544 3680 381596 3732
rect 397736 3680 397788 3732
rect 421564 3680 421616 3732
rect 427268 3680 427320 3732
rect 428464 3680 428516 3732
rect 534908 3680 534960 3732
rect 21824 3612 21876 3664
rect 39304 3612 39356 3664
rect 41880 3612 41932 3664
rect 207296 3612 207348 3664
rect 213368 3612 213420 3664
rect 231308 3612 231360 3664
rect 249984 3612 250036 3664
rect 260840 3612 260892 3664
rect 261760 3612 261812 3664
rect 266452 3612 266504 3664
rect 274548 3612 274600 3664
rect 433248 3612 433300 3664
rect 447784 3612 447836 3664
rect 458088 3612 458140 3664
rect 458824 3612 458876 3664
rect 538864 3612 538916 3664
rect 25320 3544 25372 3596
rect 26148 3544 26200 3596
rect 26516 3544 26568 3596
rect 27528 3544 27580 3596
rect 32404 3544 32456 3596
rect 33048 3544 33100 3596
rect 33600 3544 33652 3596
rect 34428 3544 34480 3596
rect 34796 3544 34848 3596
rect 35808 3544 35860 3596
rect 35992 3544 36044 3596
rect 37096 3544 37148 3596
rect 38384 3544 38436 3596
rect 39396 3544 39448 3596
rect 40684 3544 40736 3596
rect 41328 3544 41380 3596
rect 43076 3544 43128 3596
rect 44088 3544 44140 3596
rect 44272 3544 44324 3596
rect 45376 3544 45428 3596
rect 50160 3544 50212 3596
rect 50988 3544 51040 3596
rect 51356 3544 51408 3596
rect 54484 3544 54536 3596
rect 56048 3544 56100 3596
rect 56508 3544 56560 3596
rect 57244 3544 57296 3596
rect 57888 3544 57940 3596
rect 59636 3544 59688 3596
rect 61476 3544 61528 3596
rect 64328 3544 64380 3596
rect 64788 3544 64840 3596
rect 67916 3544 67968 3596
rect 68928 3544 68980 3596
rect 69112 3544 69164 3596
rect 70308 3544 70360 3596
rect 79692 3544 79744 3596
rect 80704 3544 80756 3596
rect 80888 3544 80940 3596
rect 81348 3544 81400 3596
rect 83280 3544 83332 3596
rect 84108 3544 84160 3596
rect 84476 3544 84528 3596
rect 86224 3544 86276 3596
rect 90364 3544 90416 3596
rect 91008 3544 91060 3596
rect 91560 3544 91612 3596
rect 93860 3544 93912 3596
rect 93952 3544 94004 3596
rect 95056 3544 95108 3596
rect 97448 3544 97500 3596
rect 98644 3544 98696 3596
rect 101036 3544 101088 3596
rect 102048 3544 102100 3596
rect 105728 3544 105780 3596
rect 106188 3544 106240 3596
rect 109316 3544 109368 3596
rect 111156 3544 111208 3596
rect 114008 3544 114060 3596
rect 114468 3544 114520 3596
rect 115204 3544 115256 3596
rect 116584 3544 116636 3596
rect 122288 3544 122340 3596
rect 122748 3544 122800 3596
rect 123484 3544 123536 3596
rect 124128 3544 124180 3596
rect 125876 3544 125928 3596
rect 126888 3544 126940 3596
rect 129372 3544 129424 3596
rect 130384 3544 130436 3596
rect 132960 3544 133012 3596
rect 133788 3544 133840 3596
rect 134156 3544 134208 3596
rect 135168 3544 135220 3596
rect 136456 3544 136508 3596
rect 137284 3544 137336 3596
rect 138848 3544 138900 3596
rect 139308 3544 139360 3596
rect 141240 3544 141292 3596
rect 142068 3544 142120 3596
rect 142436 3544 142488 3596
rect 143448 3544 143500 3596
rect 147128 3544 147180 3596
rect 147588 3544 147640 3596
rect 157800 3544 157852 3596
rect 158628 3544 158680 3596
rect 158904 3544 158956 3596
rect 160008 3544 160060 3596
rect 163688 3544 163740 3596
rect 164148 3544 164200 3596
rect 164884 3544 164936 3596
rect 165528 3544 165580 3596
rect 166080 3544 166132 3596
rect 166908 3544 166960 3596
rect 167184 3544 167236 3596
rect 169024 3544 169076 3596
rect 169576 3544 169628 3596
rect 170404 3544 170456 3596
rect 171968 3544 172020 3596
rect 173164 3544 173216 3596
rect 175464 3544 175516 3596
rect 176568 3544 176620 3596
rect 176660 3544 176712 3596
rect 177948 3544 178000 3596
rect 180248 3544 180300 3596
rect 180708 3544 180760 3596
rect 181444 3544 181496 3596
rect 182088 3544 182140 3596
rect 182548 3544 182600 3596
rect 183468 3544 183520 3596
rect 183744 3544 183796 3596
rect 184848 3544 184900 3596
rect 186136 3544 186188 3596
rect 186964 3544 187016 3596
rect 187332 3544 187384 3596
rect 188344 3544 188396 3596
rect 188528 3544 188580 3596
rect 188988 3544 189040 3596
rect 192024 3544 192076 3596
rect 193128 3544 193180 3596
rect 193220 3544 193272 3596
rect 195244 3544 195296 3596
rect 197176 3544 197228 3596
rect 197912 3544 197964 3596
rect 572 3476 624 3528
rect 1308 3476 1360 3528
rect 9956 3476 10008 3528
rect 10968 3476 11020 3528
rect 200396 3544 200448 3596
rect 205088 3544 205140 3596
rect 225328 3544 225380 3596
rect 226340 3544 226392 3596
rect 227628 3544 227680 3596
rect 1676 3408 1728 3460
rect 7656 3340 7708 3392
rect 200304 3476 200356 3528
rect 202144 3476 202196 3528
rect 208584 3476 208636 3528
rect 234068 3544 234120 3596
rect 252100 3544 252152 3596
rect 299388 3544 299440 3596
rect 299480 3544 299532 3596
rect 300768 3544 300820 3596
rect 307024 3544 307076 3596
rect 307944 3544 307996 3596
rect 309140 3544 309192 3596
rect 310244 3544 310296 3596
rect 312544 3544 312596 3596
rect 313832 3544 313884 3596
rect 314016 3544 314068 3596
rect 315028 3544 315080 3596
rect 316684 3544 316736 3596
rect 485228 3544 485280 3596
rect 232228 3476 232280 3528
rect 233148 3476 233200 3528
rect 238668 3476 238720 3528
rect 244096 3476 244148 3528
rect 246488 3476 246540 3528
rect 200212 3408 200264 3460
rect 206192 3408 206244 3460
rect 234896 3408 234948 3460
rect 238116 3408 238168 3460
rect 251272 3408 251324 3460
rect 254860 3408 254912 3460
rect 66720 3340 66772 3392
rect 68284 3340 68336 3392
rect 85672 3340 85724 3392
rect 89076 3340 89128 3392
rect 89168 3340 89220 3392
rect 91560 3340 91612 3392
rect 96252 3340 96304 3392
rect 97264 3340 97316 3392
rect 110512 3340 110564 3392
rect 112444 3340 112496 3392
rect 135260 3340 135312 3392
rect 137376 3340 137428 3392
rect 156604 3340 156656 3392
rect 158076 3340 158128 3392
rect 168380 3340 168432 3392
rect 169668 3340 169720 3392
rect 173164 3340 173216 3392
rect 174544 3340 174596 3392
rect 184940 3340 184992 3392
rect 187056 3340 187108 3392
rect 190828 3340 190880 3392
rect 192484 3340 192536 3392
rect 196808 3340 196860 3392
rect 197268 3340 197320 3392
rect 210976 3340 211028 3392
rect 213184 3340 213236 3392
rect 216864 3340 216916 3392
rect 217968 3340 218020 3392
rect 218060 3340 218112 3392
rect 219348 3340 219400 3392
rect 65524 3272 65576 3324
rect 72424 3272 72476 3324
rect 108120 3272 108172 3324
rect 111064 3272 111116 3324
rect 116400 3272 116452 3324
rect 123392 3272 123444 3324
rect 151820 3272 151872 3324
rect 166264 3272 166316 3324
rect 258724 3408 258776 3460
rect 260656 3408 260708 3460
rect 258264 3340 258316 3392
rect 263692 3340 263744 3392
rect 268384 3476 268436 3528
rect 270040 3476 270092 3528
rect 279792 3476 279844 3528
rect 461584 3476 461636 3528
rect 464344 3476 464396 3528
rect 466276 3476 466328 3528
rect 272432 3340 272484 3392
rect 317328 3408 317380 3460
rect 320824 3408 320876 3460
rect 285404 3340 285456 3392
rect 288440 3340 288492 3392
rect 293684 3340 293736 3392
rect 295340 3340 295392 3392
rect 299388 3340 299440 3392
rect 305552 3340 305604 3392
rect 323584 3340 323636 3392
rect 325608 3340 325660 3392
rect 331864 3340 331916 3392
rect 333888 3340 333940 3392
rect 340880 3340 340932 3392
rect 342168 3340 342220 3392
rect 364984 3340 365036 3392
rect 367008 3340 367060 3392
rect 378784 3340 378836 3392
rect 381176 3340 381228 3392
rect 389824 3340 389876 3392
rect 391848 3340 391900 3392
rect 396724 3340 396776 3392
rect 402520 3340 402572 3392
rect 407764 3340 407816 3392
rect 409604 3340 409656 3392
rect 414664 3340 414716 3392
rect 416688 3340 416740 3392
rect 440240 3340 440292 3392
rect 441528 3340 441580 3392
rect 281908 3272 281960 3324
rect 285772 3272 285824 3324
rect 291844 3272 291896 3324
rect 294880 3272 294932 3324
rect 318156 3272 318208 3324
rect 319720 3272 319772 3324
rect 330484 3272 330536 3324
rect 332692 3272 332744 3324
rect 336096 3272 336148 3324
rect 337476 3272 337528 3324
rect 376116 3272 376168 3324
rect 379980 3272 380032 3324
rect 407212 3272 407264 3324
rect 409972 3272 410024 3324
rect 453304 3408 453356 3460
rect 455696 3408 455748 3460
rect 457444 3408 457496 3460
rect 459192 3408 459244 3460
rect 461676 3340 461728 3392
rect 472624 3476 472676 3528
rect 474556 3476 474608 3528
rect 485044 3476 485096 3528
rect 486424 3476 486476 3528
rect 488816 3476 488868 3528
rect 489184 3544 489236 3596
rect 515036 3544 515088 3596
rect 515404 3544 515456 3596
rect 517152 3544 517204 3596
rect 522304 3544 522356 3596
rect 524236 3544 524288 3596
rect 540796 3544 540848 3596
rect 572720 3612 572772 3664
rect 530584 3476 530636 3528
rect 532516 3476 532568 3528
rect 540244 3476 540296 3528
rect 541992 3476 542044 3528
rect 548524 3476 548576 3528
rect 550272 3476 550324 3528
rect 552664 3476 552716 3528
rect 553400 3476 553452 3528
rect 559748 3476 559800 3528
rect 560484 3476 560536 3528
rect 563244 3544 563296 3596
rect 564532 3544 564584 3596
rect 577412 3544 577464 3596
rect 582748 3544 582800 3596
rect 565636 3476 565688 3528
rect 582196 3476 582248 3528
rect 582932 3476 582984 3528
rect 467196 3272 467248 3324
rect 469864 3272 469916 3324
rect 479340 3340 479392 3392
rect 547880 3408 547932 3460
rect 581000 3408 581052 3460
rect 582840 3408 582892 3460
rect 490564 3340 490616 3392
rect 492312 3340 492364 3392
rect 497464 3340 497516 3392
rect 499396 3340 499448 3392
rect 502984 3340 503036 3392
rect 505376 3340 505428 3392
rect 520924 3340 520976 3392
rect 523040 3340 523092 3392
rect 18236 3136 18288 3188
rect 22744 3136 22796 3188
rect 31300 3068 31352 3120
rect 204628 3204 204680 3256
rect 48964 3136 49016 3188
rect 53104 3136 53156 3188
rect 126980 3136 127032 3188
rect 221188 3204 221240 3256
rect 324964 3204 325016 3256
rect 326804 3204 326856 3256
rect 500316 3204 500368 3256
rect 502984 3204 503036 3256
rect 220452 3136 220504 3188
rect 226984 3136 227036 3188
rect 260196 3136 260248 3188
rect 264152 3136 264204 3188
rect 271236 3136 271288 3188
rect 274824 3136 274876 3188
rect 299664 3136 299716 3188
rect 302332 3136 302384 3188
rect 389456 3136 389508 3188
rect 392032 3136 392084 3188
rect 143540 3068 143592 3120
rect 148232 3068 148284 3120
rect 231032 3068 231084 3120
rect 238024 3068 238076 3120
rect 239312 3068 239364 3120
rect 240600 3068 240652 3120
rect 543004 3068 543056 3120
rect 545488 3068 545540 3120
rect 8760 3000 8812 3052
rect 15844 3000 15896 3052
rect 27712 3000 27764 3052
rect 35164 3000 35216 3052
rect 73804 3000 73856 3052
rect 75184 3000 75236 3052
rect 118792 3000 118844 3052
rect 119988 3000 120040 3052
rect 174268 3000 174320 3052
rect 181352 3000 181404 3052
rect 252376 3000 252428 3052
rect 258080 3000 258132 3052
rect 259460 3000 259512 3052
rect 262220 3000 262272 3052
rect 280804 3000 280856 3052
rect 283104 3000 283156 3052
rect 342996 3000 343048 3052
rect 344560 3000 344612 3052
rect 374644 3000 374696 3052
rect 377680 3000 377732 3052
rect 446404 3000 446456 3052
rect 452108 3000 452160 3052
rect 493324 3000 493376 3052
rect 495900 3000 495952 3052
rect 504364 3000 504416 3052
rect 510068 3000 510120 3052
rect 511264 3000 511316 3052
rect 513564 3000 513616 3052
rect 529204 3000 529256 3052
rect 531320 3000 531372 3052
rect 23020 2932 23072 2984
rect 28264 2932 28316 2984
rect 76196 2932 76248 2984
rect 79324 2932 79376 2984
rect 222752 2932 222804 2984
rect 223488 2932 223540 2984
rect 245660 2932 245712 2984
rect 247592 2932 247644 2984
rect 435364 2932 435416 2984
rect 437940 2932 437992 2984
rect 525156 2932 525208 2984
rect 527824 2932 527876 2984
rect 77392 2864 77444 2916
rect 79416 2864 79468 2916
rect 201500 2864 201552 2916
rect 209044 2864 209096 2916
rect 223948 2864 224000 2916
rect 224868 2864 224920 2916
rect 417516 2864 417568 2916
rect 420184 2864 420236 2916
rect 432604 2864 432656 2916
rect 434444 2864 434496 2916
rect 442356 2864 442408 2916
rect 445024 2864 445076 2916
rect 471244 2864 471296 2916
rect 473452 2864 473504 2916
rect 515036 2796 515088 2848
rect 515956 2796 516008 2848
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 89364 703582 89668 703610
rect 8128 702434 8156 703520
rect 8128 702406 8248 702434
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 3436 683262 3464 684247
rect 3424 683256 3476 683262
rect 3424 683198 3476 683204
rect 3422 671256 3478 671265
rect 3422 671191 3478 671200
rect 3330 580000 3386 580009
rect 3330 579935 3386 579944
rect 3344 579698 3372 579935
rect 3332 579692 3384 579698
rect 3332 579634 3384 579640
rect 3238 566944 3294 566953
rect 3238 566879 3294 566888
rect 3252 565894 3280 566879
rect 3240 565888 3292 565894
rect 3240 565830 3292 565836
rect 3330 553888 3386 553897
rect 3330 553823 3386 553832
rect 3344 553450 3372 553823
rect 3332 553444 3384 553450
rect 3332 553386 3384 553392
rect 2962 527912 3018 527921
rect 2962 527847 3018 527856
rect 2976 527202 3004 527847
rect 2964 527196 3016 527202
rect 2964 527138 3016 527144
rect 3054 501800 3110 501809
rect 3054 501735 3110 501744
rect 3068 501022 3096 501735
rect 3056 501016 3108 501022
rect 3056 500958 3108 500964
rect 3054 475688 3110 475697
rect 3054 475623 3110 475632
rect 3068 474774 3096 475623
rect 3056 474768 3108 474774
rect 3056 474710 3108 474716
rect 3146 449576 3202 449585
rect 3146 449511 3202 449520
rect 3160 448594 3188 449511
rect 3148 448588 3200 448594
rect 3148 448530 3200 448536
rect 2870 410544 2926 410553
rect 2870 410479 2926 410488
rect 2884 409902 2912 410479
rect 2872 409896 2924 409902
rect 2872 409838 2924 409844
rect 3146 358456 3202 358465
rect 3146 358391 3202 358400
rect 3160 357474 3188 358391
rect 3148 357468 3200 357474
rect 3148 357410 3200 357416
rect 3330 345400 3386 345409
rect 3330 345335 3386 345344
rect 3344 345098 3372 345335
rect 3332 345092 3384 345098
rect 3332 345034 3384 345040
rect 3330 319288 3386 319297
rect 3330 319223 3386 319232
rect 3344 318850 3372 319223
rect 3332 318844 3384 318850
rect 3332 318786 3384 318792
rect 3436 308446 3464 671191
rect 3514 658200 3570 658209
rect 3514 658135 3570 658144
rect 3528 656946 3556 658135
rect 3516 656940 3568 656946
rect 3516 656882 3568 656888
rect 3516 632120 3568 632126
rect 3514 632088 3516 632097
rect 3568 632088 3570 632097
rect 3514 632023 3570 632032
rect 3514 619168 3570 619177
rect 3514 619103 3570 619112
rect 3528 618322 3556 619103
rect 3516 618316 3568 618322
rect 3516 618258 3568 618264
rect 3514 606112 3570 606121
rect 3514 606047 3570 606056
rect 3528 605878 3556 606047
rect 3516 605872 3568 605878
rect 3516 605814 3568 605820
rect 3514 514856 3570 514865
rect 3514 514791 3516 514800
rect 3568 514791 3570 514800
rect 3516 514762 3568 514768
rect 3514 462632 3570 462641
rect 3514 462567 3570 462576
rect 3528 462398 3556 462567
rect 3516 462392 3568 462398
rect 3516 462334 3568 462340
rect 3514 423600 3570 423609
rect 3514 423535 3570 423544
rect 3528 422346 3556 423535
rect 3516 422340 3568 422346
rect 3516 422282 3568 422288
rect 3516 397520 3568 397526
rect 3514 397488 3516 397497
rect 3568 397488 3570 397497
rect 3514 397423 3570 397432
rect 3514 371376 3570 371385
rect 3514 371311 3570 371320
rect 3528 371278 3556 371311
rect 3516 371272 3568 371278
rect 3516 371214 3568 371220
rect 3424 308440 3476 308446
rect 3424 308382 3476 308388
rect 8220 307154 8248 702406
rect 24320 700398 24348 703520
rect 40512 700466 40540 703520
rect 72988 700534 73016 703520
rect 89180 703474 89208 703520
rect 89364 703474 89392 703582
rect 89180 703446 89392 703474
rect 72976 700528 73028 700534
rect 72976 700470 73028 700476
rect 40500 700460 40552 700466
rect 40500 700402 40552 700408
rect 41328 700460 41380 700466
rect 41328 700402 41380 700408
rect 24308 700392 24360 700398
rect 24308 700334 24360 700340
rect 8208 307148 8260 307154
rect 8208 307090 8260 307096
rect 3238 306232 3294 306241
rect 3238 306167 3294 306176
rect 3252 305046 3280 306167
rect 41340 305862 41368 700402
rect 89640 307222 89668 703582
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 299492 703582 299980 703610
rect 105464 699718 105492 703520
rect 137848 702434 137876 703520
rect 137848 702406 137968 702434
rect 105452 699712 105504 699718
rect 105452 699654 105504 699660
rect 106188 699712 106240 699718
rect 106188 699654 106240 699660
rect 89628 307216 89680 307222
rect 89628 307158 89680 307164
rect 41328 305856 41380 305862
rect 41328 305798 41380 305804
rect 3240 305040 3292 305046
rect 3240 304982 3292 304988
rect 106200 304502 106228 699654
rect 137940 326398 137968 702406
rect 154132 699718 154160 703520
rect 170324 700942 170352 703520
rect 170312 700936 170364 700942
rect 170312 700878 170364 700884
rect 171048 700936 171100 700942
rect 171048 700878 171100 700884
rect 154120 699712 154172 699718
rect 154120 699654 154172 699660
rect 155224 699712 155276 699718
rect 155224 699654 155276 699660
rect 137928 326392 137980 326398
rect 137928 326334 137980 326340
rect 155236 305930 155264 699654
rect 155224 305924 155276 305930
rect 155224 305866 155276 305872
rect 171060 304638 171088 700878
rect 198556 337408 198608 337414
rect 198556 337350 198608 337356
rect 171048 304632 171100 304638
rect 171048 304574 171100 304580
rect 106188 304496 106240 304502
rect 106188 304438 106240 304444
rect 129004 303748 129056 303754
rect 129004 303690 129056 303696
rect 14464 302320 14516 302326
rect 14464 302262 14516 302268
rect 3424 298852 3476 298858
rect 3424 298794 3476 298800
rect 3056 293956 3108 293962
rect 3056 293898 3108 293904
rect 3068 293185 3096 293898
rect 3054 293176 3110 293185
rect 3054 293111 3110 293120
rect 3148 255264 3200 255270
rect 3148 255206 3200 255212
rect 3160 254153 3188 255206
rect 3146 254144 3202 254153
rect 3146 254079 3202 254088
rect 3332 215280 3384 215286
rect 3332 215222 3384 215228
rect 3344 214985 3372 215222
rect 3330 214976 3386 214985
rect 3330 214911 3386 214920
rect 3056 202836 3108 202842
rect 3056 202778 3108 202784
rect 3068 201929 3096 202778
rect 3054 201920 3110 201929
rect 3054 201855 3110 201864
rect 3240 164212 3292 164218
rect 3240 164154 3292 164160
rect 3252 162897 3280 164154
rect 3238 162888 3294 162897
rect 3238 162823 3294 162832
rect 3436 136785 3464 298794
rect 3516 267708 3568 267714
rect 3516 267650 3568 267656
rect 3528 267209 3556 267650
rect 3514 267200 3570 267209
rect 3514 267135 3570 267144
rect 3516 241460 3568 241466
rect 3516 241402 3568 241408
rect 3528 241097 3556 241402
rect 3514 241088 3570 241097
rect 3514 241023 3570 241032
rect 3516 189032 3568 189038
rect 3516 188974 3568 188980
rect 3528 188873 3556 188974
rect 3514 188864 3570 188873
rect 3514 188799 3570 188808
rect 3516 150408 3568 150414
rect 3516 150350 3568 150356
rect 3528 149841 3556 150350
rect 3514 149832 3570 149841
rect 3514 149767 3570 149776
rect 3422 136776 3478 136785
rect 3422 136711 3478 136720
rect 3424 111784 3476 111790
rect 3424 111726 3476 111732
rect 3436 110673 3464 111726
rect 3422 110664 3478 110673
rect 3422 110599 3478 110608
rect 14476 97986 14504 302262
rect 90364 301164 90416 301170
rect 90364 301106 90416 301112
rect 88984 299804 89036 299810
rect 88984 299746 89036 299752
rect 88996 164218 89024 299746
rect 90376 267714 90404 301106
rect 90364 267708 90416 267714
rect 90364 267650 90416 267656
rect 88984 164212 89036 164218
rect 88984 164154 89036 164160
rect 106188 100020 106240 100026
rect 106188 99962 106240 99968
rect 93124 99748 93176 99754
rect 93124 99690 93176 99696
rect 87604 99680 87656 99686
rect 87604 99622 87656 99628
rect 72424 99544 72476 99550
rect 72424 99486 72476 99492
rect 53104 99476 53156 99482
rect 53104 99418 53156 99424
rect 39304 99408 39356 99414
rect 39304 99350 39356 99356
rect 21364 98660 21416 98666
rect 21364 98602 21416 98608
rect 3424 97980 3476 97986
rect 3424 97922 3476 97928
rect 14464 97980 14516 97986
rect 14464 97922 14516 97928
rect 3436 97617 3464 97922
rect 3422 97608 3478 97617
rect 3422 97543 3478 97552
rect 14556 97300 14608 97306
rect 14556 97242 14608 97248
rect 12256 95940 12308 95946
rect 12256 95882 12308 95888
rect 1306 94480 1362 94489
rect 1306 94415 1362 94424
rect 1320 3534 1348 94415
rect 4066 93120 4122 93129
rect 4066 93055 4122 93064
rect 3148 85536 3200 85542
rect 3148 85478 3200 85484
rect 3160 84697 3188 85478
rect 3146 84688 3202 84697
rect 3146 84623 3202 84632
rect 3424 71732 3476 71738
rect 3424 71674 3476 71680
rect 3436 71641 3464 71674
rect 3422 71632 3478 71641
rect 3422 71567 3478 71576
rect 3056 59356 3108 59362
rect 3056 59298 3108 59304
rect 3068 58585 3096 59298
rect 3054 58576 3110 58585
rect 3054 58511 3110 58520
rect 3424 45552 3476 45558
rect 3422 45520 3424 45529
rect 3476 45520 3478 45529
rect 3422 45455 3478 45464
rect 2872 33108 2924 33114
rect 2872 33050 2924 33056
rect 2884 32473 2912 33050
rect 2870 32464 2926 32473
rect 2870 32399 2926 32408
rect 3424 20664 3476 20670
rect 3424 20606 3476 20612
rect 3436 19417 3464 20606
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 3424 6860 3476 6866
rect 3424 6802 3476 6808
rect 3436 6497 3464 6802
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 2872 3596 2924 3602
rect 2872 3538 2924 3544
rect 572 3528 624 3534
rect 572 3470 624 3476
rect 1308 3528 1360 3534
rect 1308 3470 1360 3476
rect 584 480 612 3470
rect 1676 3460 1728 3466
rect 1676 3402 1728 3408
rect 1688 480 1716 3402
rect 2884 480 2912 3538
rect 4080 480 4108 93055
rect 10968 84856 11020 84862
rect 10968 84798 11020 84804
rect 5448 82272 5500 82278
rect 5448 82214 5500 82220
rect 5460 6914 5488 82214
rect 5276 6886 5488 6914
rect 5276 480 5304 6886
rect 6460 3664 6512 3670
rect 6460 3606 6512 3612
rect 6472 480 6500 3606
rect 10980 3534 11008 84798
rect 12268 16574 12296 95882
rect 12346 95840 12402 95849
rect 12346 95775 12402 95784
rect 12176 16546 12296 16574
rect 11152 3664 11204 3670
rect 11152 3606 11204 3612
rect 9956 3528 10008 3534
rect 9956 3470 10008 3476
rect 10968 3528 11020 3534
rect 10968 3470 11020 3476
rect 7656 3392 7708 3398
rect 7656 3334 7708 3340
rect 7668 480 7696 3334
rect 8760 3052 8812 3058
rect 8760 2994 8812 3000
rect 8772 480 8800 2994
rect 9968 480 9996 3470
rect 11164 480 11192 3606
rect 12176 3482 12204 16546
rect 12360 6914 12388 95775
rect 12268 6886 12388 6914
rect 12268 3670 12296 6886
rect 13544 4004 13596 4010
rect 13544 3946 13596 3952
rect 12256 3664 12308 3670
rect 12256 3606 12308 3612
rect 12176 3454 12388 3482
rect 12360 480 12388 3454
rect 13556 480 13584 3946
rect 14568 3738 14596 97242
rect 17222 97200 17278 97209
rect 17222 97135 17278 97144
rect 15844 93152 15896 93158
rect 15844 93094 15896 93100
rect 14556 3732 14608 3738
rect 14556 3674 14608 3680
rect 14740 3732 14792 3738
rect 14740 3674 14792 3680
rect 14752 480 14780 3674
rect 15856 3058 15884 93094
rect 17236 4146 17264 97135
rect 18604 89004 18656 89010
rect 18604 88946 18656 88952
rect 15936 4140 15988 4146
rect 15936 4082 15988 4088
rect 17224 4140 17276 4146
rect 17224 4082 17276 4088
rect 15844 3052 15896 3058
rect 15844 2994 15896 3000
rect 15948 480 15976 4082
rect 17040 4072 17092 4078
rect 17040 4014 17092 4020
rect 17052 480 17080 4014
rect 18616 4010 18644 88946
rect 20628 4140 20680 4146
rect 20628 4082 20680 4088
rect 18604 4004 18656 4010
rect 18604 3946 18656 3952
rect 19432 3936 19484 3942
rect 19432 3878 19484 3884
rect 18236 3188 18288 3194
rect 18236 3130 18288 3136
rect 18248 480 18276 3130
rect 19444 480 19472 3878
rect 20640 480 20668 4082
rect 21376 4078 21404 98602
rect 35254 97472 35310 97481
rect 35254 97407 35310 97416
rect 29642 97336 29698 97345
rect 29642 97271 29698 97280
rect 22742 95976 22798 95985
rect 22742 95911 22798 95920
rect 21456 82204 21508 82210
rect 21456 82146 21508 82152
rect 21468 4146 21496 82146
rect 21456 4140 21508 4146
rect 21456 4082 21508 4088
rect 21364 4072 21416 4078
rect 21364 4014 21416 4020
rect 21824 3664 21876 3670
rect 21824 3606 21876 3612
rect 21836 480 21864 3606
rect 22756 3194 22784 95911
rect 28262 94616 28318 94625
rect 28262 94551 28318 94560
rect 25504 93220 25556 93226
rect 25504 93162 25556 93168
rect 24216 4004 24268 4010
rect 24216 3946 24268 3952
rect 22744 3188 22796 3194
rect 22744 3130 22796 3136
rect 23020 2984 23072 2990
rect 23020 2926 23072 2932
rect 23032 480 23060 2926
rect 24228 480 24256 3946
rect 25516 3806 25544 93162
rect 27528 89072 27580 89078
rect 27528 89014 27580 89020
rect 26148 22772 26200 22778
rect 26148 22714 26200 22720
rect 25504 3800 25556 3806
rect 25504 3742 25556 3748
rect 26160 3602 26188 22714
rect 27540 3602 27568 89014
rect 25320 3596 25372 3602
rect 25320 3538 25372 3544
rect 26148 3596 26200 3602
rect 26148 3538 26200 3544
rect 26516 3596 26568 3602
rect 26516 3538 26568 3544
rect 27528 3596 27580 3602
rect 27528 3538 27580 3544
rect 25332 480 25360 3538
rect 26528 480 26556 3538
rect 27712 3052 27764 3058
rect 27712 2994 27764 3000
rect 27724 480 27752 2994
rect 28276 2990 28304 94551
rect 28908 87712 28960 87718
rect 28908 87654 28960 87660
rect 28264 2984 28316 2990
rect 28264 2926 28316 2932
rect 28920 480 28948 87654
rect 29656 3806 29684 97271
rect 33048 93288 33100 93294
rect 33048 93230 33100 93236
rect 30288 87644 30340 87650
rect 30288 87586 30340 87592
rect 30300 6914 30328 87586
rect 30116 6886 30328 6914
rect 29644 3800 29696 3806
rect 29644 3742 29696 3748
rect 30116 480 30144 6886
rect 33060 3602 33088 93230
rect 34428 91792 34480 91798
rect 34428 91734 34480 91740
rect 34440 3602 34468 91734
rect 35164 83496 35216 83502
rect 35164 83438 35216 83444
rect 32404 3596 32456 3602
rect 32404 3538 32456 3544
rect 33048 3596 33100 3602
rect 33048 3538 33100 3544
rect 33600 3596 33652 3602
rect 33600 3538 33652 3544
rect 34428 3596 34480 3602
rect 34428 3538 34480 3544
rect 34796 3596 34848 3602
rect 34796 3538 34848 3544
rect 31300 3120 31352 3126
rect 31300 3062 31352 3068
rect 31312 480 31340 3062
rect 32416 480 32444 3538
rect 33612 480 33640 3538
rect 34808 480 34836 3538
rect 35176 3058 35204 83438
rect 35268 22778 35296 97407
rect 37188 96008 37240 96014
rect 37188 95950 37240 95956
rect 37096 89140 37148 89146
rect 37096 89082 37148 89088
rect 35256 22772 35308 22778
rect 35256 22714 35308 22720
rect 37108 16574 37136 89082
rect 37016 16546 37136 16574
rect 35808 11756 35860 11762
rect 35808 11698 35860 11704
rect 35820 3602 35848 11698
rect 35808 3596 35860 3602
rect 35808 3538 35860 3544
rect 35992 3596 36044 3602
rect 35992 3538 36044 3544
rect 35164 3052 35216 3058
rect 35164 2994 35216 3000
rect 36004 480 36032 3538
rect 37016 3482 37044 16546
rect 37200 6914 37228 95950
rect 37108 6886 37228 6914
rect 37108 3602 37136 6886
rect 39316 3670 39344 99350
rect 43444 98728 43496 98734
rect 43444 98670 43496 98676
rect 40684 97368 40736 97374
rect 40684 97310 40736 97316
rect 39396 15904 39448 15910
rect 39396 15846 39448 15852
rect 39304 3664 39356 3670
rect 39304 3606 39356 3612
rect 39408 3602 39436 15846
rect 40696 3874 40724 97310
rect 41328 87780 41380 87786
rect 41328 87722 41380 87728
rect 40684 3868 40736 3874
rect 40684 3810 40736 3816
rect 39580 3800 39632 3806
rect 39580 3742 39632 3748
rect 37096 3596 37148 3602
rect 37096 3538 37148 3544
rect 38384 3596 38436 3602
rect 38384 3538 38436 3544
rect 39396 3596 39448 3602
rect 39396 3538 39448 3544
rect 37016 3454 37228 3482
rect 37200 480 37228 3454
rect 38396 480 38424 3538
rect 39592 480 39620 3742
rect 41340 3602 41368 87722
rect 43456 3738 43484 98670
rect 50988 94580 51040 94586
rect 50988 94522 51040 94528
rect 48228 94512 48280 94518
rect 48228 94454 48280 94460
rect 46848 91860 46900 91866
rect 46848 91802 46900 91808
rect 45468 90364 45520 90370
rect 45468 90306 45520 90312
rect 45376 83564 45428 83570
rect 45376 83506 45428 83512
rect 44088 21412 44140 21418
rect 44088 21354 44140 21360
rect 43444 3732 43496 3738
rect 43444 3674 43496 3680
rect 41880 3664 41932 3670
rect 41880 3606 41932 3612
rect 40684 3596 40736 3602
rect 40684 3538 40736 3544
rect 41328 3596 41380 3602
rect 41328 3538 41380 3544
rect 40696 480 40724 3538
rect 41892 480 41920 3606
rect 44100 3602 44128 21354
rect 45388 16574 45416 83506
rect 45296 16546 45416 16574
rect 43076 3596 43128 3602
rect 43076 3538 43128 3544
rect 44088 3596 44140 3602
rect 44088 3538 44140 3544
rect 44272 3596 44324 3602
rect 44272 3538 44324 3544
rect 43088 480 43116 3538
rect 44284 480 44312 3538
rect 45296 3482 45324 16546
rect 45480 6914 45508 90306
rect 46860 6914 46888 91802
rect 48240 6914 48268 94454
rect 45388 6886 45508 6914
rect 46676 6886 46888 6914
rect 47872 6886 48268 6914
rect 45388 3602 45416 6886
rect 45376 3596 45428 3602
rect 45376 3538 45428 3544
rect 45296 3454 45508 3482
rect 45480 480 45508 3454
rect 46676 480 46704 6886
rect 47872 480 47900 6886
rect 51000 3602 51028 94522
rect 52552 3936 52604 3942
rect 52552 3878 52604 3884
rect 50160 3596 50212 3602
rect 50160 3538 50212 3544
rect 50988 3596 51040 3602
rect 50988 3538 51040 3544
rect 51356 3596 51408 3602
rect 51356 3538 51408 3544
rect 48964 3188 49016 3194
rect 48964 3130 49016 3136
rect 48976 480 49004 3130
rect 50172 480 50200 3538
rect 51368 480 51396 3538
rect 52564 480 52592 3878
rect 53116 3194 53144 99418
rect 54484 98796 54536 98802
rect 54484 98738 54536 98744
rect 53748 94648 53800 94654
rect 53748 94590 53800 94596
rect 53104 3188 53156 3194
rect 53104 3130 53156 3136
rect 53760 480 53788 94590
rect 54496 3602 54524 98738
rect 58624 97504 58676 97510
rect 58624 97446 58676 97452
rect 56508 97436 56560 97442
rect 56508 97378 56560 97384
rect 54944 4004 54996 4010
rect 54944 3946 54996 3952
rect 54484 3596 54536 3602
rect 54484 3538 54536 3544
rect 54956 480 54984 3946
rect 56520 3602 56548 97378
rect 57888 90432 57940 90438
rect 57888 90374 57940 90380
rect 57900 3602 57928 90374
rect 58440 4072 58492 4078
rect 58440 4014 58492 4020
rect 56048 3596 56100 3602
rect 56048 3538 56100 3544
rect 56508 3596 56560 3602
rect 56508 3538 56560 3544
rect 57244 3596 57296 3602
rect 57244 3538 57296 3544
rect 57888 3596 57940 3602
rect 57888 3538 57940 3544
rect 56060 480 56088 3538
rect 57256 480 57284 3538
rect 58452 480 58480 4014
rect 58636 3806 58664 97446
rect 65524 93424 65576 93430
rect 65524 93366 65576 93372
rect 61384 93356 61436 93362
rect 61384 93298 61436 93304
rect 61396 4010 61424 93298
rect 61476 87848 61528 87854
rect 61476 87790 61528 87796
rect 61384 4004 61436 4010
rect 61384 3946 61436 3952
rect 60832 3868 60884 3874
rect 60832 3810 60884 3816
rect 58624 3800 58676 3806
rect 58624 3742 58676 3748
rect 59636 3596 59688 3602
rect 59636 3538 59688 3544
rect 59648 480 59676 3538
rect 60844 480 60872 3810
rect 61488 3602 61516 87790
rect 64788 13116 64840 13122
rect 64788 13058 64840 13064
rect 63224 4004 63276 4010
rect 63224 3946 63276 3952
rect 62028 3732 62080 3738
rect 62028 3674 62080 3680
rect 61476 3596 61528 3602
rect 61476 3538 61528 3544
rect 62040 480 62068 3674
rect 63236 480 63264 3946
rect 64800 3602 64828 13058
rect 65536 4078 65564 93366
rect 71044 91996 71096 92002
rect 71044 91938 71096 91944
rect 70308 91928 70360 91934
rect 70308 91870 70360 91876
rect 68284 86284 68336 86290
rect 68284 86226 68336 86232
rect 65524 4072 65576 4078
rect 65524 4014 65576 4020
rect 64328 3596 64380 3602
rect 64328 3538 64380 3544
rect 64788 3596 64840 3602
rect 64788 3538 64840 3544
rect 67916 3596 67968 3602
rect 67916 3538 67968 3544
rect 64340 480 64368 3538
rect 66720 3392 66772 3398
rect 66720 3334 66772 3340
rect 65524 3324 65576 3330
rect 65524 3266 65576 3272
rect 65536 480 65564 3266
rect 66732 480 66760 3334
rect 67928 480 67956 3538
rect 68296 3398 68324 86226
rect 68928 69692 68980 69698
rect 68928 69634 68980 69640
rect 68940 3602 68968 69634
rect 70216 8968 70268 8974
rect 70216 8910 70268 8916
rect 68928 3596 68980 3602
rect 68928 3538 68980 3544
rect 69112 3596 69164 3602
rect 69112 3538 69164 3544
rect 68284 3392 68336 3398
rect 68284 3334 68336 3340
rect 69124 480 69152 3538
rect 70228 3482 70256 8910
rect 70320 3602 70348 91870
rect 71056 3738 71084 91938
rect 71688 87984 71740 87990
rect 71688 87926 71740 87932
rect 71700 6914 71728 87926
rect 71516 6886 71728 6914
rect 71044 3732 71096 3738
rect 71044 3674 71096 3680
rect 70308 3596 70360 3602
rect 70308 3538 70360 3544
rect 70228 3454 70348 3482
rect 70320 480 70348 3454
rect 71516 480 71544 6886
rect 72436 3330 72464 99486
rect 84108 98864 84160 98870
rect 84108 98806 84160 98812
rect 79324 94716 79376 94722
rect 79324 94658 79376 94664
rect 76564 90500 76616 90506
rect 76564 90442 76616 90448
rect 75184 87916 75236 87922
rect 75184 87858 75236 87864
rect 72608 4140 72660 4146
rect 72608 4082 72660 4088
rect 72424 3324 72476 3330
rect 72424 3266 72476 3272
rect 72620 480 72648 4082
rect 75000 3800 75052 3806
rect 75000 3742 75052 3748
rect 73804 3052 73856 3058
rect 73804 2994 73856 3000
rect 73816 480 73844 2994
rect 75012 480 75040 3742
rect 75196 3058 75224 87858
rect 76576 4146 76604 90442
rect 76564 4140 76616 4146
rect 76564 4082 76616 4088
rect 78588 4072 78640 4078
rect 78588 4014 78640 4020
rect 75184 3052 75236 3058
rect 75184 2994 75236 3000
rect 76196 2984 76248 2990
rect 76196 2926 76248 2932
rect 76208 480 76236 2926
rect 77392 2916 77444 2922
rect 77392 2858 77444 2864
rect 77404 480 77432 2858
rect 78600 480 78628 4014
rect 79336 2990 79364 94658
rect 80704 90568 80756 90574
rect 80704 90510 80756 90516
rect 79416 86352 79468 86358
rect 79416 86294 79468 86300
rect 79324 2984 79376 2990
rect 79324 2926 79376 2932
rect 79428 2922 79456 86294
rect 80716 3602 80744 90510
rect 81348 10328 81400 10334
rect 81348 10270 81400 10276
rect 81360 3602 81388 10270
rect 82084 3732 82136 3738
rect 82084 3674 82136 3680
rect 79692 3596 79744 3602
rect 79692 3538 79744 3544
rect 80704 3596 80756 3602
rect 80704 3538 80756 3544
rect 80888 3596 80940 3602
rect 80888 3538 80940 3544
rect 81348 3596 81400 3602
rect 81348 3538 81400 3544
rect 79416 2916 79468 2922
rect 79416 2858 79468 2864
rect 79704 480 79732 3538
rect 80900 480 80928 3538
rect 82096 480 82124 3674
rect 84120 3602 84148 98806
rect 86868 90636 86920 90642
rect 86868 90578 86920 90584
rect 86224 86420 86276 86426
rect 86224 86362 86276 86368
rect 86236 3602 86264 86362
rect 83280 3596 83332 3602
rect 83280 3538 83332 3544
rect 84108 3596 84160 3602
rect 84108 3538 84160 3544
rect 84476 3596 84528 3602
rect 84476 3538 84528 3544
rect 86224 3596 86276 3602
rect 86224 3538 86276 3544
rect 83292 480 83320 3538
rect 84488 480 84516 3538
rect 85672 3392 85724 3398
rect 85672 3334 85724 3340
rect 85684 480 85712 3334
rect 86880 480 86908 90578
rect 87616 4010 87644 99622
rect 91008 99612 91060 99618
rect 91008 99554 91060 99560
rect 88984 88052 89036 88058
rect 88984 87994 89036 88000
rect 88248 84924 88300 84930
rect 88248 84866 88300 84872
rect 88260 6914 88288 84866
rect 87984 6886 88288 6914
rect 87604 4004 87656 4010
rect 87604 3946 87656 3952
rect 87984 480 88012 6886
rect 88996 3942 89024 87994
rect 89076 35216 89128 35222
rect 89076 35158 89128 35164
rect 88984 3936 89036 3942
rect 88984 3878 89036 3884
rect 89088 3398 89116 35158
rect 91020 3602 91048 99554
rect 93136 4078 93164 99690
rect 97264 97572 97316 97578
rect 97264 97514 97316 97520
rect 95148 90704 95200 90710
rect 95148 90646 95200 90652
rect 95056 84992 95108 84998
rect 95056 84934 95108 84940
rect 95068 16574 95096 84934
rect 94976 16546 95096 16574
rect 93124 4072 93176 4078
rect 93124 4014 93176 4020
rect 91652 4004 91704 4010
rect 91652 3946 91704 3952
rect 93952 4004 94004 4010
rect 93952 3946 94004 3952
rect 90364 3596 90416 3602
rect 90364 3538 90416 3544
rect 91008 3596 91060 3602
rect 91008 3538 91060 3544
rect 91560 3596 91612 3602
rect 91560 3538 91612 3544
rect 89076 3392 89128 3398
rect 89076 3334 89128 3340
rect 89168 3392 89220 3398
rect 89168 3334 89220 3340
rect 89180 480 89208 3334
rect 90376 480 90404 3538
rect 91572 3398 91600 3538
rect 91560 3392 91612 3398
rect 91560 3334 91612 3340
rect 91664 2122 91692 3946
rect 92756 3936 92808 3942
rect 92756 3878 92808 3884
rect 91572 2094 91692 2122
rect 91572 480 91600 2094
rect 92768 480 92796 3878
rect 93964 3754 93992 3946
rect 93872 3726 93992 3754
rect 93872 3602 93900 3726
rect 93860 3596 93912 3602
rect 93860 3538 93912 3544
rect 93952 3596 94004 3602
rect 93952 3538 94004 3544
rect 93964 480 93992 3538
rect 94976 3482 95004 16546
rect 95160 6914 95188 90646
rect 95068 6886 95188 6914
rect 95068 3602 95096 6886
rect 95056 3596 95108 3602
rect 95056 3538 95108 3544
rect 94976 3454 95188 3482
rect 95160 480 95188 3454
rect 97276 3398 97304 97514
rect 98644 92064 98696 92070
rect 98644 92006 98696 92012
rect 97356 17264 97408 17270
rect 97356 17206 97408 17212
rect 97368 3942 97396 17206
rect 97356 3936 97408 3942
rect 97356 3878 97408 3884
rect 98656 3602 98684 92006
rect 104808 89276 104860 89282
rect 104808 89218 104860 89224
rect 102048 89208 102100 89214
rect 102048 89150 102100 89156
rect 99840 4888 99892 4894
rect 99840 4830 99892 4836
rect 98736 4820 98788 4826
rect 98736 4762 98788 4768
rect 97448 3596 97500 3602
rect 97448 3538 97500 3544
rect 98644 3596 98696 3602
rect 98644 3538 98696 3544
rect 96252 3392 96304 3398
rect 96252 3334 96304 3340
rect 97264 3392 97316 3398
rect 97264 3334 97316 3340
rect 96264 480 96292 3334
rect 97460 480 97488 3538
rect 98748 2394 98776 4762
rect 98656 2366 98776 2394
rect 98656 480 98684 2366
rect 99852 480 99880 4830
rect 102060 3602 102088 89150
rect 102232 7608 102284 7614
rect 102232 7550 102284 7556
rect 101036 3596 101088 3602
rect 101036 3538 101088 3544
rect 102048 3596 102100 3602
rect 102048 3538 102100 3544
rect 101048 480 101076 3538
rect 102244 480 102272 7550
rect 104820 6914 104848 89218
rect 105544 88120 105596 88126
rect 105544 88062 105596 88068
rect 104544 6886 104848 6914
rect 103336 3936 103388 3942
rect 103336 3878 103388 3884
rect 103348 480 103376 3878
rect 104544 480 104572 6886
rect 105556 4078 105584 88062
rect 105544 4072 105596 4078
rect 105544 4014 105596 4020
rect 106200 3602 106228 99962
rect 124864 99952 124916 99958
rect 124864 99894 124916 99900
rect 108304 99884 108356 99890
rect 108304 99826 108356 99832
rect 106924 86556 106976 86562
rect 106924 86498 106976 86504
rect 106936 3874 106964 86498
rect 107016 6180 107068 6186
rect 107016 6122 107068 6128
rect 106924 3868 106976 3874
rect 106924 3810 106976 3816
rect 105728 3596 105780 3602
rect 105728 3538 105780 3544
rect 106188 3596 106240 3602
rect 106188 3538 106240 3544
rect 105740 480 105768 3538
rect 107028 3074 107056 6122
rect 108316 4010 108344 99826
rect 111064 99816 111116 99822
rect 111064 99758 111116 99764
rect 108304 4004 108356 4010
rect 108304 3946 108356 3952
rect 109316 3596 109368 3602
rect 109316 3538 109368 3544
rect 108120 3324 108172 3330
rect 108120 3266 108172 3272
rect 106936 3046 107056 3074
rect 106936 480 106964 3046
rect 108132 480 108160 3266
rect 109328 480 109356 3538
rect 110512 3392 110564 3398
rect 110512 3334 110564 3340
rect 110524 480 110552 3334
rect 111076 3330 111104 99758
rect 121368 97708 121420 97714
rect 121368 97650 121420 97656
rect 112444 97640 112496 97646
rect 112444 97582 112496 97588
rect 111156 86488 111208 86494
rect 111156 86430 111208 86436
rect 111168 3602 111196 86430
rect 111616 4072 111668 4078
rect 111616 4014 111668 4020
rect 111156 3596 111208 3602
rect 111156 3538 111208 3544
rect 111064 3324 111116 3330
rect 111064 3266 111116 3272
rect 111628 480 111656 4014
rect 112456 3398 112484 97582
rect 114468 94784 114520 94790
rect 114468 94726 114520 94732
rect 113088 25560 113140 25566
rect 113088 25502 113140 25508
rect 113100 6914 113128 25502
rect 112824 6886 113128 6914
rect 112444 3392 112496 3398
rect 112444 3334 112496 3340
rect 112824 480 112852 6886
rect 114480 3602 114508 94726
rect 116584 90772 116636 90778
rect 116584 90714 116636 90720
rect 115204 89344 115256 89350
rect 115204 89286 115256 89292
rect 115216 4078 115244 89286
rect 115204 4072 115256 4078
rect 115204 4014 115256 4020
rect 116596 3602 116624 90714
rect 119988 89412 120040 89418
rect 119988 89354 120040 89360
rect 119896 14476 119948 14482
rect 119896 14418 119948 14424
rect 117596 4072 117648 4078
rect 117596 4014 117648 4020
rect 114008 3596 114060 3602
rect 114008 3538 114060 3544
rect 114468 3596 114520 3602
rect 114468 3538 114520 3544
rect 115204 3596 115256 3602
rect 115204 3538 115256 3544
rect 116584 3596 116636 3602
rect 116584 3538 116636 3544
rect 114020 480 114048 3538
rect 115216 480 115244 3538
rect 116400 3324 116452 3330
rect 116400 3266 116452 3272
rect 116412 480 116440 3266
rect 117608 480 117636 4014
rect 118792 3052 118844 3058
rect 118792 2994 118844 3000
rect 118804 480 118832 2994
rect 119908 480 119936 14418
rect 120000 3058 120028 89354
rect 121380 6914 121408 97650
rect 122748 89480 122800 89486
rect 122748 89422 122800 89428
rect 121104 6886 121408 6914
rect 119988 3052 120040 3058
rect 119988 2994 120040 3000
rect 121104 480 121132 6886
rect 122760 3602 122788 89422
rect 123484 86624 123536 86630
rect 123484 86566 123536 86572
rect 123496 6914 123524 86566
rect 124128 85060 124180 85066
rect 124128 85002 124180 85008
rect 123404 6886 123524 6914
rect 122288 3596 122340 3602
rect 122288 3538 122340 3544
rect 122748 3596 122800 3602
rect 122748 3538 122800 3544
rect 122300 480 122328 3538
rect 123404 3330 123432 6886
rect 124140 3602 124168 85002
rect 124680 7676 124732 7682
rect 124680 7618 124732 7624
rect 123484 3596 123536 3602
rect 123484 3538 123536 3544
rect 124128 3596 124180 3602
rect 124128 3538 124180 3544
rect 123392 3324 123444 3330
rect 123392 3266 123444 3272
rect 123496 480 123524 3538
rect 124692 480 124720 7618
rect 124876 3806 124904 99894
rect 126888 96076 126940 96082
rect 126888 96018 126940 96024
rect 124864 3800 124916 3806
rect 124864 3742 124916 3748
rect 126900 3602 126928 96018
rect 128268 93492 128320 93498
rect 128268 93434 128320 93440
rect 128280 6914 128308 93434
rect 128188 6886 128308 6914
rect 125876 3596 125928 3602
rect 125876 3538 125928 3544
rect 126888 3596 126940 3602
rect 126888 3538 126940 3544
rect 125888 480 125916 3538
rect 126980 3188 127032 3194
rect 126980 3130 127032 3136
rect 126992 480 127020 3130
rect 128188 480 128216 6886
rect 129016 6866 129044 303690
rect 180064 302796 180116 302802
rect 180064 302738 180116 302744
rect 166264 302524 166316 302530
rect 166264 302466 166316 302472
rect 148324 302456 148376 302462
rect 148324 302398 148376 302404
rect 144184 301232 144236 301238
rect 144184 301174 144236 301180
rect 134524 99136 134576 99142
rect 134524 99078 134576 99084
rect 133788 99000 133840 99006
rect 133788 98942 133840 98948
rect 130384 98932 130436 98938
rect 130384 98874 130436 98880
rect 129004 6860 129056 6866
rect 129004 6802 129056 6808
rect 130396 3602 130424 98874
rect 131764 6248 131816 6254
rect 131764 6190 131816 6196
rect 130568 4004 130620 4010
rect 130568 3946 130620 3952
rect 129372 3596 129424 3602
rect 129372 3538 129424 3544
rect 130384 3596 130436 3602
rect 130384 3538 130436 3544
rect 129384 480 129412 3538
rect 130580 480 130608 3946
rect 131776 480 131804 6190
rect 133800 3602 133828 98942
rect 134536 4010 134564 99078
rect 137284 94852 137336 94858
rect 137284 94794 137336 94800
rect 135168 93560 135220 93566
rect 135168 93502 135220 93508
rect 134524 4004 134576 4010
rect 134524 3946 134576 3952
rect 135180 3602 135208 93502
rect 137296 3602 137324 94794
rect 142068 93628 142120 93634
rect 142068 93570 142120 93576
rect 139308 90908 139360 90914
rect 139308 90850 139360 90856
rect 137376 90840 137428 90846
rect 137376 90782 137428 90788
rect 132960 3596 133012 3602
rect 132960 3538 133012 3544
rect 133788 3596 133840 3602
rect 133788 3538 133840 3544
rect 134156 3596 134208 3602
rect 134156 3538 134208 3544
rect 135168 3596 135220 3602
rect 135168 3538 135220 3544
rect 136456 3596 136508 3602
rect 136456 3538 136508 3544
rect 137284 3596 137336 3602
rect 137284 3538 137336 3544
rect 132972 480 133000 3538
rect 134168 480 134196 3538
rect 135260 3392 135312 3398
rect 135260 3334 135312 3340
rect 135272 480 135300 3334
rect 136468 480 136496 3538
rect 137388 3398 137416 90782
rect 137652 4004 137704 4010
rect 137652 3946 137704 3952
rect 137376 3392 137428 3398
rect 137376 3334 137428 3340
rect 137664 480 137692 3946
rect 139320 3602 139348 90850
rect 140044 3868 140096 3874
rect 140044 3810 140096 3816
rect 138848 3596 138900 3602
rect 138848 3538 138900 3544
rect 139308 3596 139360 3602
rect 139308 3538 139360 3544
rect 138860 480 138888 3538
rect 140056 480 140084 3810
rect 142080 3602 142108 93570
rect 142804 92132 142856 92138
rect 142804 92074 142856 92080
rect 142816 4010 142844 92074
rect 144196 20670 144224 301174
rect 146944 299872 146996 299878
rect 146944 299814 146996 299820
rect 146208 94920 146260 94926
rect 146208 94862 146260 94868
rect 144828 92200 144880 92206
rect 144828 92142 144880 92148
rect 144184 20664 144236 20670
rect 144184 20606 144236 20612
rect 143448 18624 143500 18630
rect 143448 18566 143500 18572
rect 142804 4004 142856 4010
rect 142804 3946 142856 3952
rect 143460 3602 143488 18566
rect 144840 6914 144868 92142
rect 146220 6914 146248 94862
rect 146956 59362 146984 299814
rect 148336 150414 148364 302398
rect 152464 301368 152516 301374
rect 152464 301310 152516 301316
rect 151084 299940 151136 299946
rect 151084 299882 151136 299888
rect 148324 150408 148376 150414
rect 148324 150350 148376 150356
rect 148324 99068 148376 99074
rect 148324 99010 148376 99016
rect 147588 94988 147640 94994
rect 147588 94930 147640 94936
rect 146944 59356 146996 59362
rect 146944 59298 146996 59304
rect 144748 6886 144868 6914
rect 145944 6886 146248 6914
rect 141240 3596 141292 3602
rect 141240 3538 141292 3544
rect 142068 3596 142120 3602
rect 142068 3538 142120 3544
rect 142436 3596 142488 3602
rect 142436 3538 142488 3544
rect 143448 3596 143500 3602
rect 143448 3538 143500 3544
rect 141252 480 141280 3538
rect 142448 480 142476 3538
rect 143540 3120 143592 3126
rect 143540 3062 143592 3068
rect 143552 480 143580 3062
rect 144748 480 144776 6886
rect 145944 480 145972 6886
rect 147600 3602 147628 94930
rect 148336 12434 148364 99010
rect 148968 92268 149020 92274
rect 148968 92210 149020 92216
rect 148244 12406 148364 12434
rect 147128 3596 147180 3602
rect 147128 3538 147180 3544
rect 147588 3596 147640 3602
rect 147588 3538 147640 3544
rect 147140 480 147168 3538
rect 148244 3126 148272 12406
rect 148980 4146 149008 92210
rect 151096 45558 151124 299882
rect 152476 85542 152504 301310
rect 156604 301300 156656 301306
rect 156604 301242 156656 301248
rect 155224 300076 155276 300082
rect 155224 300018 155276 300024
rect 155236 189038 155264 300018
rect 155224 189032 155276 189038
rect 155224 188974 155276 188980
rect 152556 99204 152608 99210
rect 152556 99146 152608 99152
rect 152464 85536 152516 85542
rect 152464 85478 152516 85484
rect 151084 45552 151136 45558
rect 151084 45494 151136 45500
rect 148968 4140 149020 4146
rect 148968 4082 149020 4088
rect 149520 4140 149572 4146
rect 149520 4082 149572 4088
rect 148324 4004 148376 4010
rect 148324 3946 148376 3952
rect 148232 3120 148284 3126
rect 148232 3062 148284 3068
rect 148336 480 148364 3946
rect 149532 480 149560 4082
rect 152568 4010 152596 99146
rect 155224 95056 155276 95062
rect 155224 94998 155276 95004
rect 153108 85128 153160 85134
rect 153108 85070 153160 85076
rect 152556 4004 152608 4010
rect 152556 3946 152608 3952
rect 152648 4004 152700 4010
rect 152648 3946 152700 3952
rect 152660 3806 152688 3946
rect 150624 3800 150676 3806
rect 150624 3742 150676 3748
rect 152648 3800 152700 3806
rect 152648 3742 152700 3748
rect 150636 480 150664 3742
rect 151820 3324 151872 3330
rect 151820 3266 151872 3272
rect 151832 480 151860 3266
rect 153120 2774 153148 85070
rect 155236 4146 155264 94998
rect 156616 33114 156644 301242
rect 159364 300144 159416 300150
rect 159364 300086 159416 300092
rect 157984 300008 158036 300014
rect 157984 299950 158036 299956
rect 156696 92336 156748 92342
rect 156696 92278 156748 92284
rect 156604 33108 156656 33114
rect 156604 33050 156656 33056
rect 156708 4146 156736 92278
rect 157996 71738 158024 299950
rect 159376 111790 159404 300086
rect 160008 209092 160060 209098
rect 160008 209034 160060 209040
rect 160020 161474 160048 209034
rect 166276 202842 166304 302466
rect 174544 301436 174596 301442
rect 174544 301378 174596 301384
rect 170404 294024 170456 294030
rect 170404 293966 170456 293972
rect 169668 276072 169720 276078
rect 169668 276014 169720 276020
rect 166264 202836 166316 202842
rect 166264 202778 166316 202784
rect 169680 186289 169708 276014
rect 169666 186280 169722 186289
rect 169666 186215 169722 186224
rect 160020 161446 160600 161474
rect 160572 160698 160600 161446
rect 169208 160812 169260 160818
rect 169208 160754 169260 160760
rect 169220 160698 169248 160754
rect 160572 160670 160954 160698
rect 168958 160670 169248 160698
rect 165160 160540 165212 160546
rect 165160 160482 165212 160488
rect 165172 160426 165200 160482
rect 164910 160398 165200 160426
rect 162872 158710 162900 160004
rect 162860 158704 162912 158710
rect 162860 158646 162912 158652
rect 166920 158030 166948 160004
rect 166908 158024 166960 158030
rect 166908 157966 166960 157972
rect 160940 122874 160968 124100
rect 162872 122942 162900 124100
rect 162860 122936 162912 122942
rect 162860 122878 162912 122884
rect 160928 122868 160980 122874
rect 160928 122810 160980 122816
rect 164896 122670 164924 124100
rect 166920 122806 166948 124100
rect 166908 122800 166960 122806
rect 166908 122742 166960 122748
rect 164884 122664 164936 122670
rect 164884 122606 164936 122612
rect 168944 122602 168972 124100
rect 170416 122806 170444 293966
rect 173164 278792 173216 278798
rect 173164 278734 173216 278740
rect 171784 248464 171836 248470
rect 171784 248406 171836 248412
rect 170496 212560 170548 212566
rect 170496 212502 170548 212508
rect 170508 152153 170536 212502
rect 171692 184816 171744 184822
rect 171692 184758 171744 184764
rect 171704 184249 171732 184758
rect 171690 184240 171746 184249
rect 171690 184175 171746 184184
rect 171796 171057 171824 248406
rect 171876 193180 171928 193186
rect 171876 193122 171928 193128
rect 171782 171048 171838 171057
rect 171782 170983 171838 170992
rect 171888 169289 171916 193122
rect 172428 190188 172480 190194
rect 172428 190130 172480 190136
rect 172440 189961 172468 190130
rect 172426 189952 172482 189961
rect 172426 189887 172482 189896
rect 172060 189032 172112 189038
rect 172060 188974 172112 188980
rect 172072 188737 172100 188974
rect 172058 188728 172114 188737
rect 172058 188663 172114 188672
rect 173176 187678 173204 278734
rect 173256 244316 173308 244322
rect 173256 244258 173308 244264
rect 173268 193186 173296 244258
rect 174556 241466 174584 301378
rect 175924 291236 175976 291242
rect 175924 291178 175976 291184
rect 174544 241460 174596 241466
rect 174544 241402 174596 241408
rect 174544 218068 174596 218074
rect 174544 218010 174596 218016
rect 173348 197396 173400 197402
rect 173348 197338 173400 197344
rect 173256 193180 173308 193186
rect 173256 193122 173308 193128
rect 172152 187672 172204 187678
rect 172150 187640 172152 187649
rect 173164 187672 173216 187678
rect 172204 187640 172206 187649
rect 173164 187614 173216 187620
rect 172150 187575 172206 187584
rect 171968 185564 172020 185570
rect 171968 185506 172020 185512
rect 171874 169280 171930 169289
rect 171874 169215 171930 169224
rect 171980 166977 172008 185506
rect 172426 184920 172482 184929
rect 172426 184855 172428 184864
rect 172480 184855 172482 184864
rect 172428 184826 172480 184832
rect 172428 183524 172480 183530
rect 172428 183466 172480 183472
rect 172440 183025 172468 183466
rect 172426 183016 172482 183025
rect 172426 182951 172482 182960
rect 172060 182164 172112 182170
rect 172060 182106 172112 182112
rect 172072 181801 172100 182106
rect 172058 181792 172114 181801
rect 172058 181727 172114 181736
rect 172428 180804 172480 180810
rect 172428 180746 172480 180752
rect 172440 180577 172468 180746
rect 172426 180568 172482 180577
rect 172426 180503 172482 180512
rect 172428 179376 172480 179382
rect 172428 179318 172480 179324
rect 172440 179217 172468 179318
rect 172426 179208 172482 179217
rect 172426 179143 172482 179152
rect 172428 178016 172480 178022
rect 172426 177984 172428 177993
rect 172480 177984 172482 177993
rect 172336 177948 172388 177954
rect 172426 177919 172482 177928
rect 172336 177890 172388 177896
rect 172348 177449 172376 177890
rect 172334 177440 172390 177449
rect 172334 177375 172390 177384
rect 172244 176656 172296 176662
rect 172244 176598 172296 176604
rect 172256 176089 172284 176598
rect 172242 176080 172298 176089
rect 172242 176015 172298 176024
rect 172428 175228 172480 175234
rect 172428 175170 172480 175176
rect 172440 174865 172468 175170
rect 172426 174856 172482 174865
rect 172426 174791 172482 174800
rect 172428 173664 172480 173670
rect 172426 173632 172428 173641
rect 172480 173632 172482 173641
rect 172426 173567 172482 173576
rect 172428 172440 172480 172446
rect 172426 172408 172428 172417
rect 172480 172408 172482 172417
rect 172426 172343 172482 172352
rect 172244 171080 172296 171086
rect 172244 171022 172296 171028
rect 172256 170513 172284 171022
rect 172242 170504 172298 170513
rect 172242 170439 172298 170448
rect 172244 169040 172296 169046
rect 172244 168982 172296 168988
rect 171966 166968 172022 166977
rect 171966 166903 172022 166912
rect 171784 166320 171836 166326
rect 171784 166262 171836 166268
rect 171600 154556 171652 154562
rect 171600 154498 171652 154504
rect 171612 153785 171640 154498
rect 171692 153808 171744 153814
rect 171598 153776 171654 153785
rect 171692 153750 171744 153756
rect 171598 153711 171654 153720
rect 171704 153241 171732 153750
rect 171690 153232 171746 153241
rect 171600 153196 171652 153202
rect 171690 153167 171746 153176
rect 171600 153138 171652 153144
rect 171612 152697 171640 153138
rect 171598 152688 171654 152697
rect 171598 152623 171654 152632
rect 170494 152144 170550 152153
rect 170494 152079 170550 152088
rect 171692 151632 171744 151638
rect 171692 151574 171744 151580
rect 171704 150521 171732 151574
rect 171690 150512 171746 150521
rect 171690 150447 171746 150456
rect 171508 149796 171560 149802
rect 171508 149738 171560 149744
rect 171520 149433 171548 149738
rect 171506 149424 171562 149433
rect 171506 149359 171562 149368
rect 171692 148368 171744 148374
rect 171690 148336 171692 148345
rect 171744 148336 171746 148345
rect 171690 148271 171746 148280
rect 171508 148028 171560 148034
rect 171508 147970 171560 147976
rect 171520 147801 171548 147970
rect 171506 147792 171562 147801
rect 171506 147727 171562 147736
rect 171692 147552 171744 147558
rect 171692 147494 171744 147500
rect 171704 147257 171732 147494
rect 171690 147248 171746 147257
rect 171690 147183 171746 147192
rect 171692 146192 171744 146198
rect 171692 146134 171744 146140
rect 171704 145081 171732 146134
rect 171690 145072 171746 145081
rect 171690 145007 171746 145016
rect 171692 144900 171744 144906
rect 171692 144842 171744 144848
rect 171704 144537 171732 144842
rect 171690 144528 171746 144537
rect 171690 144463 171746 144472
rect 171796 144129 171824 166262
rect 172060 165572 172112 165578
rect 172060 165514 172112 165520
rect 172072 165209 172100 165514
rect 172058 165200 172114 165209
rect 172058 165135 172114 165144
rect 172256 163577 172284 168982
rect 172428 168360 172480 168366
rect 172428 168302 172480 168308
rect 172440 167929 172468 168302
rect 172426 167920 172482 167929
rect 172426 167855 172482 167864
rect 172428 164212 172480 164218
rect 172428 164154 172480 164160
rect 172440 164121 172468 164154
rect 172426 164112 172482 164121
rect 172426 164047 172482 164056
rect 172242 163568 172298 163577
rect 172242 163503 172298 163512
rect 172152 162852 172204 162858
rect 172152 162794 172204 162800
rect 172164 162353 172192 162794
rect 172150 162344 172206 162353
rect 172150 162279 172206 162288
rect 172428 161220 172480 161226
rect 172428 161162 172480 161168
rect 172440 160993 172468 161162
rect 172426 160984 172482 160993
rect 172426 160919 172482 160928
rect 171968 156664 172020 156670
rect 171968 156606 172020 156612
rect 171782 144120 171838 144129
rect 171782 144055 171838 144064
rect 171876 144084 171928 144090
rect 171876 144026 171928 144032
rect 171888 143041 171916 144026
rect 171980 143585 172008 156606
rect 172244 151768 172296 151774
rect 172244 151710 172296 151716
rect 172256 151065 172284 151710
rect 172428 151700 172480 151706
rect 172428 151642 172480 151648
rect 172440 151609 172468 151642
rect 172426 151600 172482 151609
rect 172426 151535 172482 151544
rect 172242 151056 172298 151065
rect 172242 150991 172298 151000
rect 172428 150408 172480 150414
rect 172428 150350 172480 150356
rect 172440 149977 172468 150350
rect 172426 149968 172482 149977
rect 172426 149903 172482 149912
rect 172428 148912 172480 148918
rect 172426 148880 172428 148889
rect 172480 148880 172482 148889
rect 172426 148815 172482 148824
rect 173360 148374 173388 197338
rect 173440 194608 173492 194614
rect 173440 194550 173492 194556
rect 173348 148368 173400 148374
rect 173348 148310 173400 148316
rect 173164 148300 173216 148306
rect 173164 148242 173216 148248
rect 172336 147620 172388 147626
rect 172336 147562 172388 147568
rect 172348 146713 172376 147562
rect 172334 146704 172390 146713
rect 172334 146639 172390 146648
rect 172428 146260 172480 146266
rect 172428 146202 172480 146208
rect 172440 146169 172468 146202
rect 172426 146160 172482 146169
rect 172426 146095 172482 146104
rect 172428 145784 172480 145790
rect 172428 145726 172480 145732
rect 172440 145625 172468 145726
rect 172426 145616 172482 145625
rect 172426 145551 172482 145560
rect 171966 143576 172022 143585
rect 171966 143511 172022 143520
rect 172428 143540 172480 143546
rect 172428 143482 172480 143488
rect 171874 143032 171930 143041
rect 171874 142967 171930 142976
rect 172440 142497 172468 143482
rect 172426 142488 172482 142497
rect 172426 142423 172482 142432
rect 172428 142112 172480 142118
rect 172428 142054 172480 142060
rect 172336 142044 172388 142050
rect 172336 141986 172388 141992
rect 171876 141840 171928 141846
rect 171876 141782 171928 141788
rect 171888 141409 171916 141782
rect 171874 141400 171930 141409
rect 171874 141335 171930 141344
rect 172348 140865 172376 141986
rect 172440 141953 172468 142054
rect 172426 141944 172482 141953
rect 172426 141879 172482 141888
rect 172334 140856 172390 140865
rect 172334 140791 172390 140800
rect 172428 140752 172480 140758
rect 172428 140694 172480 140700
rect 172152 140344 172204 140350
rect 172150 140312 172152 140321
rect 172204 140312 172206 140321
rect 172150 140247 172206 140256
rect 171324 140072 171376 140078
rect 171324 140014 171376 140020
rect 171336 135425 171364 140014
rect 172440 139777 172468 140694
rect 173176 140350 173204 148242
rect 173452 148034 173480 194550
rect 174556 154562 174584 218010
rect 174636 216708 174688 216714
rect 174636 216650 174688 216656
rect 174544 154556 174596 154562
rect 174544 154498 174596 154504
rect 174648 153814 174676 216650
rect 174728 213988 174780 213994
rect 174728 213930 174780 213936
rect 174636 153808 174688 153814
rect 174636 153750 174688 153756
rect 174740 153202 174768 213930
rect 175936 160818 175964 291178
rect 176016 287088 176068 287094
rect 176016 287030 176068 287036
rect 175924 160812 175976 160818
rect 175924 160754 175976 160760
rect 176028 158710 176056 287030
rect 178684 282940 178736 282946
rect 178684 282882 178736 282888
rect 177304 271924 177356 271930
rect 177304 271866 177356 271872
rect 176108 193248 176160 193254
rect 176108 193190 176160 193196
rect 176016 158704 176068 158710
rect 176016 158646 176068 158652
rect 174728 153196 174780 153202
rect 174728 153138 174780 153144
rect 175924 151836 175976 151842
rect 175924 151778 175976 151784
rect 174544 149116 174596 149122
rect 174544 149058 174596 149064
rect 173440 148028 173492 148034
rect 173440 147970 173492 147976
rect 173164 140344 173216 140350
rect 173164 140286 173216 140292
rect 172426 139768 172482 139777
rect 172426 139703 172482 139712
rect 172428 139392 172480 139398
rect 172428 139334 172480 139340
rect 172336 139324 172388 139330
rect 172336 139266 172388 139272
rect 172244 139256 172296 139262
rect 172242 139224 172244 139233
rect 172296 139224 172298 139233
rect 172242 139159 172298 139168
rect 172348 138145 172376 139266
rect 172440 138689 172468 139334
rect 172426 138680 172482 138689
rect 172426 138615 172482 138624
rect 172334 138136 172390 138145
rect 172334 138071 172390 138080
rect 172060 137964 172112 137970
rect 172060 137906 172112 137912
rect 171692 137896 171744 137902
rect 171692 137838 171744 137844
rect 171704 137057 171732 137838
rect 172072 137601 172100 137906
rect 172058 137592 172114 137601
rect 172058 137527 172114 137536
rect 171690 137048 171746 137057
rect 171690 136983 171746 136992
rect 172244 136604 172296 136610
rect 172244 136546 172296 136552
rect 171876 136264 171928 136270
rect 171876 136206 171928 136212
rect 171322 135416 171378 135425
rect 171322 135351 171378 135360
rect 171692 135176 171744 135182
rect 171692 135118 171744 135124
rect 171704 134337 171732 135118
rect 171888 134881 171916 136206
rect 172256 135969 172284 136546
rect 174556 136542 174584 149058
rect 175936 137902 175964 151778
rect 176120 147558 176148 193190
rect 177316 184822 177344 271866
rect 177396 229152 177448 229158
rect 177396 229094 177448 229100
rect 177304 184816 177356 184822
rect 177304 184758 177356 184764
rect 177304 175296 177356 175302
rect 177304 175238 177356 175244
rect 176108 147552 176160 147558
rect 176108 147494 176160 147500
rect 177316 144090 177344 175238
rect 177408 161226 177436 229094
rect 178696 190194 178724 282882
rect 180076 255270 180104 302738
rect 196624 300280 196676 300286
rect 196624 300222 196676 300228
rect 196636 293962 196664 300222
rect 198568 298897 198596 337350
rect 202800 304706 202828 703520
rect 218992 700330 219020 703520
rect 235184 700466 235212 703520
rect 252468 700664 252520 700670
rect 252468 700606 252520 700612
rect 246948 700596 247000 700602
rect 246948 700538 247000 700544
rect 235172 700460 235224 700466
rect 235172 700402 235224 700408
rect 242164 700460 242216 700466
rect 242164 700402 242216 700408
rect 244188 700460 244240 700466
rect 244188 700402 244240 700408
rect 218980 700324 219032 700330
rect 218980 700266 219032 700272
rect 222844 700324 222896 700330
rect 222844 700266 222896 700272
rect 241428 700324 241480 700330
rect 241428 700266 241480 700272
rect 217324 618316 217376 618322
rect 217324 618258 217376 618264
rect 215944 565888 215996 565894
rect 215944 565830 215996 565836
rect 214564 462392 214616 462398
rect 214564 462334 214616 462340
rect 213184 409896 213236 409902
rect 213184 409838 213236 409844
rect 213196 307358 213224 409838
rect 213184 307352 213236 307358
rect 213184 307294 213236 307300
rect 214576 306066 214604 462334
rect 215956 307426 215984 565830
rect 217336 307494 217364 618258
rect 220728 324352 220780 324358
rect 220728 324294 220780 324300
rect 220636 311908 220688 311914
rect 220636 311850 220688 311856
rect 217324 307488 217376 307494
rect 217324 307430 217376 307436
rect 215944 307420 215996 307426
rect 215944 307362 215996 307368
rect 214564 306060 214616 306066
rect 214564 306002 214616 306008
rect 202788 304700 202840 304706
rect 202788 304642 202840 304648
rect 202052 303680 202104 303686
rect 202052 303622 202104 303628
rect 199384 301572 199436 301578
rect 199384 301514 199436 301520
rect 198554 298888 198610 298897
rect 198554 298823 198610 298832
rect 197910 294536 197966 294545
rect 197910 294471 197966 294480
rect 197924 294030 197952 294471
rect 197912 294024 197964 294030
rect 197912 293966 197964 293972
rect 196624 293956 196676 293962
rect 196624 293898 196676 293904
rect 197542 292360 197598 292369
rect 197542 292295 197598 292304
rect 197556 291242 197584 292295
rect 197544 291236 197596 291242
rect 197544 291178 197596 291184
rect 198738 290184 198794 290193
rect 198738 290119 198794 290128
rect 197542 288144 197598 288153
rect 197542 288079 197598 288088
rect 197556 287094 197584 288079
rect 197544 287088 197596 287094
rect 197544 287030 197596 287036
rect 198094 285968 198150 285977
rect 198094 285903 198150 285912
rect 197358 283792 197414 283801
rect 197358 283727 197414 283736
rect 197372 282946 197400 283727
rect 197360 282940 197412 282946
rect 197360 282882 197412 282888
rect 197358 281616 197414 281625
rect 181444 281580 181496 281586
rect 197358 281551 197360 281560
rect 181444 281522 181496 281528
rect 197412 281551 197414 281560
rect 197360 281522 197412 281528
rect 180064 255264 180116 255270
rect 180064 255206 180116 255212
rect 180064 252612 180116 252618
rect 180064 252554 180116 252560
rect 178776 251252 178828 251258
rect 178776 251194 178828 251200
rect 178684 190188 178736 190194
rect 178684 190130 178736 190136
rect 178684 186380 178736 186386
rect 178684 186322 178736 186328
rect 177396 161220 177448 161226
rect 177396 161162 177448 161168
rect 177488 160132 177540 160138
rect 177488 160074 177540 160080
rect 177304 144084 177356 144090
rect 177304 144026 177356 144032
rect 177500 139262 177528 160074
rect 178696 145790 178724 186322
rect 178788 172446 178816 251194
rect 180076 173670 180104 252554
rect 180156 240168 180208 240174
rect 180156 240110 180208 240116
rect 180168 185570 180196 240110
rect 180248 201544 180300 201550
rect 180248 201486 180300 201492
rect 180156 185564 180208 185570
rect 180156 185506 180208 185512
rect 180064 173664 180116 173670
rect 180064 173606 180116 173612
rect 180156 173188 180208 173194
rect 180156 173130 180208 173136
rect 178776 172440 178828 172446
rect 178776 172382 178828 172388
rect 178776 166388 178828 166394
rect 178776 166330 178828 166336
rect 178684 145784 178736 145790
rect 178684 145726 178736 145732
rect 178788 141846 178816 166330
rect 180168 144906 180196 173130
rect 180260 149802 180288 201486
rect 181456 189038 181484 281522
rect 197726 279440 197782 279449
rect 197726 279375 197782 279384
rect 197740 278798 197768 279375
rect 197728 278792 197780 278798
rect 197728 278734 197780 278740
rect 197358 277400 197414 277409
rect 197358 277335 197414 277344
rect 197372 276078 197400 277335
rect 197360 276072 197412 276078
rect 197360 276014 197412 276020
rect 196624 274712 196676 274718
rect 196624 274654 196676 274660
rect 195244 270564 195296 270570
rect 195244 270506 195296 270512
rect 192484 268184 192536 268190
rect 192484 268126 192536 268132
rect 191104 266484 191156 266490
rect 191104 266426 191156 266432
rect 188436 263628 188488 263634
rect 188436 263570 188488 263576
rect 187056 262268 187108 262274
rect 187056 262210 187108 262216
rect 184296 259480 184348 259486
rect 184296 259422 184348 259428
rect 182824 256760 182876 256766
rect 182824 256702 182876 256708
rect 181536 255332 181588 255338
rect 181536 255274 181588 255280
rect 181444 189032 181496 189038
rect 181444 188974 181496 188980
rect 181444 182844 181496 182850
rect 181444 182786 181496 182792
rect 180248 149796 180300 149802
rect 180248 149738 180300 149744
rect 181456 146198 181484 182786
rect 181548 175234 181576 255274
rect 181628 205692 181680 205698
rect 181628 205634 181680 205640
rect 181536 175228 181588 175234
rect 181536 175170 181588 175176
rect 181640 151638 181668 205634
rect 182836 176662 182864 256702
rect 184204 225004 184256 225010
rect 184204 224946 184256 224952
rect 182916 209840 182968 209846
rect 182916 209782 182968 209788
rect 182824 176656 182876 176662
rect 182824 176598 182876 176604
rect 182824 154624 182876 154630
rect 182824 154566 182876 154572
rect 181628 151632 181680 151638
rect 181628 151574 181680 151580
rect 181536 147688 181588 147694
rect 181536 147630 181588 147636
rect 181444 146192 181496 146198
rect 181444 146134 181496 146140
rect 180156 144900 180208 144906
rect 180156 144842 180208 144848
rect 179420 143608 179472 143614
rect 179420 143550 179472 143556
rect 178776 141840 178828 141846
rect 178776 141782 178828 141788
rect 178040 140820 178092 140826
rect 178040 140762 178092 140768
rect 177488 139256 177540 139262
rect 177488 139198 177540 139204
rect 175924 137896 175976 137902
rect 175924 137838 175976 137844
rect 176016 136672 176068 136678
rect 176016 136614 176068 136620
rect 172428 136536 172480 136542
rect 172426 136504 172428 136513
rect 174544 136536 174596 136542
rect 172480 136504 172482 136513
rect 174544 136478 174596 136484
rect 172426 136439 172482 136448
rect 172242 135960 172298 135969
rect 172242 135895 172298 135904
rect 172520 135924 172572 135930
rect 172520 135866 172572 135872
rect 171874 134872 171930 134881
rect 171874 134807 171930 134816
rect 172532 134722 172560 135866
rect 172440 134694 172560 134722
rect 171690 134328 171746 134337
rect 171690 134263 171746 134272
rect 172060 134292 172112 134298
rect 172060 134234 172112 134240
rect 172072 133385 172100 134234
rect 172440 133929 172468 134694
rect 172520 134564 172572 134570
rect 172520 134506 172572 134512
rect 172426 133920 172482 133929
rect 172426 133855 172482 133864
rect 172058 133376 172114 133385
rect 172058 133311 172114 133320
rect 172426 132832 172482 132841
rect 172532 132818 172560 134506
rect 176028 134298 176056 136614
rect 178052 135182 178080 140762
rect 179432 136270 179460 143550
rect 181548 136610 181576 147630
rect 182836 137970 182864 154566
rect 182928 151706 182956 209782
rect 183008 189100 183060 189106
rect 183008 189042 183060 189048
rect 182916 151700 182968 151706
rect 182916 151642 182968 151648
rect 183020 146266 183048 189042
rect 183008 146260 183060 146266
rect 183008 146202 183060 146208
rect 182824 137964 182876 137970
rect 182824 137906 182876 137912
rect 181536 136604 181588 136610
rect 181536 136546 181588 136552
rect 179420 136264 179472 136270
rect 179420 136206 179472 136212
rect 178040 135176 178092 135182
rect 178040 135118 178092 135124
rect 176016 134292 176068 134298
rect 176016 134234 176068 134240
rect 172482 132790 172560 132818
rect 172426 132767 172482 132776
rect 171140 132524 171192 132530
rect 171140 132466 171192 132472
rect 171152 132297 171180 132466
rect 171138 132288 171194 132297
rect 171138 132223 171194 132232
rect 172426 131744 172482 131753
rect 172426 131679 172482 131688
rect 171506 131200 171562 131209
rect 171506 131135 171562 131144
rect 171520 129742 171548 131135
rect 172440 131102 172468 131679
rect 172428 131096 172480 131102
rect 172428 131038 172480 131044
rect 171874 130656 171930 130665
rect 171874 130591 171930 130600
rect 171888 129810 171916 130591
rect 172426 130112 172482 130121
rect 172426 130047 172428 130056
rect 172480 130047 172482 130056
rect 175280 130076 175332 130082
rect 172428 130018 172480 130024
rect 175280 130018 175332 130024
rect 171876 129804 171928 129810
rect 171876 129746 171928 129752
rect 171508 129736 171560 129742
rect 171508 129678 171560 129684
rect 171874 129568 171930 129577
rect 171874 129503 171930 129512
rect 171506 129024 171562 129033
rect 171506 128959 171562 128968
rect 171520 128518 171548 128959
rect 171888 128586 171916 129503
rect 171876 128580 171928 128586
rect 171876 128522 171928 128528
rect 174452 128580 174504 128586
rect 174452 128522 174504 128528
rect 171508 128512 171560 128518
rect 173164 128512 173216 128518
rect 171508 128454 171560 128460
rect 171782 128480 171838 128489
rect 173164 128454 173216 128460
rect 171782 128415 171838 128424
rect 171690 127936 171746 127945
rect 171690 127871 171746 127880
rect 171704 127022 171732 127871
rect 171692 127016 171744 127022
rect 171692 126958 171744 126964
rect 171322 124672 171378 124681
rect 171322 124607 171324 124616
rect 171376 124607 171378 124616
rect 171324 124578 171376 124584
rect 170404 122800 170456 122806
rect 170404 122742 170456 122748
rect 168932 122596 168984 122602
rect 168932 122538 168984 122544
rect 171796 118658 171824 128415
rect 172426 127392 172482 127401
rect 172426 127327 172482 127336
rect 172440 127090 172468 127327
rect 172428 127084 172480 127090
rect 172428 127026 172480 127032
rect 172058 126848 172114 126857
rect 172058 126783 172114 126792
rect 172072 125662 172100 126783
rect 172334 126304 172390 126313
rect 172334 126239 172390 126248
rect 172348 125798 172376 126239
rect 172336 125792 172388 125798
rect 172336 125734 172388 125740
rect 172426 125760 172482 125769
rect 172426 125695 172428 125704
rect 172480 125695 172482 125704
rect 172428 125666 172480 125672
rect 172060 125656 172112 125662
rect 172060 125598 172112 125604
rect 172426 125216 172482 125225
rect 172426 125151 172428 125160
rect 172480 125151 172482 125160
rect 172428 125122 172480 125128
rect 171966 124264 172022 124273
rect 171966 124199 171968 124208
rect 172020 124199 172022 124208
rect 171968 124170 172020 124176
rect 173176 121446 173204 128454
rect 174464 127634 174492 128522
rect 174452 127628 174504 127634
rect 174452 127570 174504 127576
rect 175292 125594 175320 130018
rect 176660 129804 176712 129810
rect 176660 129746 176712 129752
rect 176672 126954 176700 129746
rect 182824 127084 182876 127090
rect 182824 127026 182876 127032
rect 176660 126948 176712 126954
rect 176660 126890 176712 126896
rect 180064 125792 180116 125798
rect 180064 125734 180116 125740
rect 178684 125724 178736 125730
rect 178684 125666 178736 125672
rect 175280 125588 175332 125594
rect 175280 125530 175332 125536
rect 177304 125180 177356 125186
rect 177304 125122 177356 125128
rect 175924 124636 175976 124642
rect 175924 124578 175976 124584
rect 174544 124228 174596 124234
rect 174544 124170 174596 124176
rect 173164 121440 173216 121446
rect 173164 121382 173216 121388
rect 171784 118652 171836 118658
rect 171784 118594 171836 118600
rect 159364 111784 159416 111790
rect 159364 111726 159416 111732
rect 174556 102134 174584 124170
rect 175936 103494 175964 124578
rect 177316 106282 177344 125122
rect 178696 107642 178724 125666
rect 180076 110430 180104 125734
rect 181444 125656 181496 125662
rect 181444 125598 181496 125604
rect 181456 111790 181484 125598
rect 182836 114510 182864 127026
rect 184216 122806 184244 224946
rect 184308 177954 184336 259422
rect 186964 227792 187016 227798
rect 186964 227734 187016 227740
rect 184296 177948 184348 177954
rect 184296 177890 184348 177896
rect 184296 173936 184348 173942
rect 184296 173878 184348 173884
rect 184308 143546 184336 173878
rect 184296 143540 184348 143546
rect 184296 143482 184348 143488
rect 184204 122800 184256 122806
rect 184204 122742 184256 122748
rect 186976 122738 187004 227734
rect 187068 178022 187096 262210
rect 188344 222216 188396 222222
rect 188344 222158 188396 222164
rect 187056 178016 187108 178022
rect 187056 177958 187108 177964
rect 188356 122942 188384 222158
rect 188448 179382 188476 263570
rect 191116 180810 191144 266426
rect 191196 241528 191248 241534
rect 191196 241470 191248 241476
rect 191104 180804 191156 180810
rect 191104 180746 191156 180752
rect 188436 179376 188488 179382
rect 188436 179318 188488 179324
rect 188528 178084 188580 178090
rect 188528 178026 188580 178032
rect 188540 156670 188568 178026
rect 191208 168366 191236 241470
rect 191288 191684 191340 191690
rect 191288 191626 191340 191632
rect 191196 168360 191248 168366
rect 191196 168302 191248 168308
rect 188528 156664 188580 156670
rect 188528 156606 188580 156612
rect 191104 155984 191156 155990
rect 191104 155926 191156 155932
rect 191116 139330 191144 155926
rect 191300 151774 191328 191626
rect 192496 182170 192524 268126
rect 192576 237448 192628 237454
rect 192576 237390 192628 237396
rect 192484 182164 192536 182170
rect 192484 182106 192536 182112
rect 192484 179444 192536 179450
rect 192484 179386 192536 179392
rect 192496 166326 192524 179386
rect 192484 166320 192536 166326
rect 192484 166262 192536 166268
rect 192588 165578 192616 237390
rect 193864 233844 193916 233850
rect 193864 233786 193916 233792
rect 193876 169046 193904 233786
rect 193956 198756 194008 198762
rect 193956 198698 194008 198704
rect 193864 169040 193916 169046
rect 193864 168982 193916 168988
rect 192576 165572 192628 165578
rect 192576 165514 192628 165520
rect 192484 164552 192536 164558
rect 192484 164494 192536 164500
rect 191288 151768 191340 151774
rect 191288 151710 191340 151716
rect 192496 142050 192524 164494
rect 192576 158840 192628 158846
rect 192576 158782 192628 158788
rect 192484 142044 192536 142050
rect 192484 141986 192536 141992
rect 192588 139398 192616 158782
rect 193968 150414 193996 198698
rect 195256 183530 195284 270506
rect 195336 236156 195388 236162
rect 195336 236098 195388 236104
rect 195244 183524 195296 183530
rect 195244 183466 195296 183472
rect 195348 164218 195376 236098
rect 195428 185224 195480 185230
rect 195428 185166 195480 185172
rect 195336 164212 195388 164218
rect 195336 164154 195388 164160
rect 195244 158024 195296 158030
rect 195244 157966 195296 157972
rect 193956 150408 194008 150414
rect 193956 150350 194008 150356
rect 192576 139392 192628 139398
rect 192576 139334 192628 139340
rect 191104 139324 191156 139330
rect 191104 139266 191156 139272
rect 191104 127016 191156 127022
rect 191104 126958 191156 126964
rect 188344 122936 188396 122942
rect 188344 122878 188396 122884
rect 186964 122732 187016 122738
rect 186964 122674 187016 122680
rect 191116 116686 191144 126958
rect 191104 116680 191156 116686
rect 191104 116622 191156 116628
rect 182824 114504 182876 114510
rect 182824 114446 182876 114452
rect 181444 111784 181496 111790
rect 181444 111726 181496 111732
rect 180064 110424 180116 110430
rect 180064 110366 180116 110372
rect 178684 107636 178736 107642
rect 178684 107578 178736 107584
rect 177304 106276 177356 106282
rect 177304 106218 177356 106224
rect 175924 103488 175976 103494
rect 175924 103430 175976 103436
rect 174544 102128 174596 102134
rect 174544 102070 174596 102076
rect 195256 100094 195284 157966
rect 195440 148918 195468 185166
rect 196636 184890 196664 274654
rect 197542 273048 197598 273057
rect 197542 272983 197598 272992
rect 197556 271930 197584 272983
rect 197544 271924 197596 271930
rect 197544 271866 197596 271872
rect 197726 270872 197782 270881
rect 197726 270807 197782 270816
rect 197740 270570 197768 270807
rect 197728 270564 197780 270570
rect 197728 270506 197780 270512
rect 197818 268696 197874 268705
rect 197818 268631 197874 268640
rect 197832 268190 197860 268631
rect 197820 268184 197872 268190
rect 197820 268126 197872 268132
rect 197358 266520 197414 266529
rect 197358 266455 197360 266464
rect 197412 266455 197414 266464
rect 197360 266426 197412 266432
rect 197358 264480 197414 264489
rect 197358 264415 197414 264424
rect 197372 263634 197400 264415
rect 197360 263628 197412 263634
rect 197360 263570 197412 263576
rect 197358 262304 197414 262313
rect 197358 262239 197360 262248
rect 197412 262239 197414 262248
rect 197360 262210 197412 262216
rect 197726 260128 197782 260137
rect 197726 260063 197782 260072
rect 197740 259486 197768 260063
rect 197728 259480 197780 259486
rect 197728 259422 197780 259428
rect 197542 257952 197598 257961
rect 197542 257887 197598 257896
rect 197556 256766 197584 257887
rect 197544 256760 197596 256766
rect 197544 256702 197596 256708
rect 197910 255776 197966 255785
rect 197910 255711 197966 255720
rect 197924 255338 197952 255711
rect 197912 255332 197964 255338
rect 197912 255274 197964 255280
rect 197542 253736 197598 253745
rect 197542 253671 197598 253680
rect 197556 252618 197584 253671
rect 197544 252612 197596 252618
rect 197544 252554 197596 252560
rect 197358 251560 197414 251569
rect 197358 251495 197414 251504
rect 197372 251258 197400 251495
rect 197360 251252 197412 251258
rect 197360 251194 197412 251200
rect 197634 249384 197690 249393
rect 197634 249319 197690 249328
rect 197648 248470 197676 249319
rect 197636 248464 197688 248470
rect 197636 248406 197688 248412
rect 198002 247208 198058 247217
rect 198002 247143 198058 247152
rect 197358 245032 197414 245041
rect 197358 244967 197414 244976
rect 197372 244322 197400 244967
rect 197360 244316 197412 244322
rect 197360 244258 197412 244264
rect 197910 242856 197966 242865
rect 197910 242791 197966 242800
rect 197924 241534 197952 242791
rect 197912 241528 197964 241534
rect 197912 241470 197964 241476
rect 197726 240816 197782 240825
rect 197726 240751 197782 240760
rect 197740 240174 197768 240751
rect 197728 240168 197780 240174
rect 197728 240110 197780 240116
rect 197542 238640 197598 238649
rect 197542 238575 197598 238584
rect 197556 237454 197584 238575
rect 197544 237448 197596 237454
rect 197544 237390 197596 237396
rect 197726 236464 197782 236473
rect 197726 236399 197782 236408
rect 197740 236162 197768 236399
rect 197728 236156 197780 236162
rect 197728 236098 197780 236104
rect 197726 234288 197782 234297
rect 197726 234223 197782 234232
rect 197740 233850 197768 234223
rect 197728 233844 197780 233850
rect 197728 233786 197780 233792
rect 196716 231940 196768 231946
rect 196716 231882 196768 231888
rect 196624 184884 196676 184890
rect 196624 184826 196676 184832
rect 196624 162852 196676 162858
rect 196624 162794 196676 162800
rect 195428 148912 195480 148918
rect 195428 148854 195480 148860
rect 195336 146260 195388 146266
rect 195336 146202 195388 146208
rect 195348 140758 195376 146202
rect 196636 142118 196664 162794
rect 196728 162790 196756 231882
rect 197634 230072 197690 230081
rect 197634 230007 197690 230016
rect 197648 229158 197676 230007
rect 197636 229152 197688 229158
rect 197636 229094 197688 229100
rect 197358 227896 197414 227905
rect 197358 227831 197414 227840
rect 197372 227798 197400 227831
rect 197360 227792 197412 227798
rect 197360 227734 197412 227740
rect 197358 225720 197414 225729
rect 197358 225655 197414 225664
rect 197372 225010 197400 225655
rect 197360 225004 197412 225010
rect 197360 224946 197412 224952
rect 197358 223544 197414 223553
rect 197358 223479 197414 223488
rect 197372 222222 197400 223479
rect 197360 222216 197412 222222
rect 197360 222158 197412 222164
rect 197542 219192 197598 219201
rect 197542 219127 197598 219136
rect 197556 218074 197584 219127
rect 197544 218068 197596 218074
rect 197544 218010 197596 218016
rect 197358 217152 197414 217161
rect 197358 217087 197414 217096
rect 197372 216714 197400 217087
rect 197360 216708 197412 216714
rect 197360 216650 197412 216656
rect 197542 214976 197598 214985
rect 197542 214911 197598 214920
rect 197556 213994 197584 214911
rect 197544 213988 197596 213994
rect 197544 213930 197596 213936
rect 197358 212800 197414 212809
rect 197358 212735 197414 212744
rect 197372 212566 197400 212735
rect 197360 212560 197412 212566
rect 197360 212502 197412 212508
rect 197358 210624 197414 210633
rect 197358 210559 197414 210568
rect 197372 209846 197400 210559
rect 197360 209840 197412 209846
rect 197360 209782 197412 209788
rect 197358 206408 197414 206417
rect 197358 206343 197414 206352
rect 197372 205698 197400 206343
rect 197360 205692 197412 205698
rect 197360 205634 197412 205640
rect 197358 202056 197414 202065
rect 197358 201991 197414 202000
rect 197372 201550 197400 201991
rect 197360 201544 197412 201550
rect 197360 201486 197412 201492
rect 197358 197704 197414 197713
rect 197358 197639 197414 197648
rect 197372 197402 197400 197639
rect 197360 197396 197412 197402
rect 197360 197338 197412 197344
rect 197634 195528 197690 195537
rect 197634 195463 197690 195472
rect 197648 194614 197676 195463
rect 197636 194608 197688 194614
rect 197636 194550 197688 194556
rect 197358 193488 197414 193497
rect 197358 193423 197414 193432
rect 197372 193254 197400 193423
rect 197360 193248 197412 193254
rect 197360 193190 197412 193196
rect 197358 189136 197414 189145
rect 197358 189071 197360 189080
rect 197412 189071 197414 189080
rect 197360 189042 197412 189048
rect 197358 186960 197414 186969
rect 197358 186895 197414 186904
rect 197372 186386 197400 186895
rect 197360 186380 197412 186386
rect 197360 186322 197412 186328
rect 197358 184784 197414 184793
rect 197358 184719 197414 184728
rect 196808 184204 196860 184210
rect 196808 184146 196860 184152
rect 196716 162784 196768 162790
rect 196716 162726 196768 162732
rect 196820 147626 196848 184146
rect 197372 182850 197400 184719
rect 197360 182844 197412 182850
rect 197360 182786 197412 182792
rect 197358 178392 197414 178401
rect 197358 178327 197414 178336
rect 197372 178090 197400 178327
rect 197360 178084 197412 178090
rect 197360 178026 197412 178032
rect 197634 176216 197690 176225
rect 197634 176151 197690 176160
rect 197648 175302 197676 176151
rect 197636 175296 197688 175302
rect 197636 175238 197688 175244
rect 197358 174040 197414 174049
rect 197358 173975 197414 173984
rect 197372 173942 197400 173975
rect 197360 173936 197412 173942
rect 197360 173878 197412 173884
rect 198016 171086 198044 247143
rect 198108 209098 198136 285903
rect 198646 275224 198702 275233
rect 198646 275159 198702 275168
rect 198660 274718 198688 275159
rect 198648 274712 198700 274718
rect 198648 274654 198700 274660
rect 198370 232112 198426 232121
rect 198370 232047 198426 232056
rect 198384 231946 198412 232047
rect 198372 231940 198424 231946
rect 198372 231882 198424 231888
rect 198096 209092 198148 209098
rect 198096 209034 198148 209040
rect 198186 208448 198242 208457
rect 198186 208383 198242 208392
rect 198094 199880 198150 199889
rect 198094 199815 198150 199824
rect 198108 185230 198136 199815
rect 198200 191690 198228 208383
rect 198278 204232 198334 204241
rect 198278 204167 198334 204176
rect 198292 198762 198320 204167
rect 198280 198756 198332 198762
rect 198280 198698 198332 198704
rect 198188 191684 198240 191690
rect 198188 191626 198240 191632
rect 198370 191312 198426 191321
rect 198370 191247 198426 191256
rect 198096 185224 198148 185230
rect 198096 185166 198148 185172
rect 198384 184210 198412 191247
rect 198372 184204 198424 184210
rect 198372 184146 198424 184152
rect 198094 182744 198150 182753
rect 198094 182679 198150 182688
rect 198108 173194 198136 182679
rect 198370 180568 198426 180577
rect 198370 180503 198426 180512
rect 198384 179450 198412 180503
rect 198372 179444 198424 179450
rect 198372 179386 198424 179392
rect 198096 173188 198148 173194
rect 198096 173130 198148 173136
rect 198186 171864 198242 171873
rect 198186 171799 198242 171808
rect 198004 171080 198056 171086
rect 198004 171022 198056 171028
rect 197726 169824 197782 169833
rect 197726 169759 197782 169768
rect 197542 167648 197598 167657
rect 197542 167583 197598 167592
rect 197556 164558 197584 167583
rect 197740 166394 197768 169759
rect 197728 166388 197780 166394
rect 197728 166330 197780 166336
rect 198094 165472 198150 165481
rect 198094 165407 198150 165416
rect 197544 164552 197596 164558
rect 197544 164494 197596 164500
rect 198002 163296 198058 163305
rect 198002 163231 198058 163240
rect 197542 161120 197598 161129
rect 197542 161055 197598 161064
rect 197556 160138 197584 161055
rect 197544 160132 197596 160138
rect 197544 160074 197596 160080
rect 197358 159080 197414 159089
rect 197358 159015 197414 159024
rect 197372 158846 197400 159015
rect 197360 158840 197412 158846
rect 197360 158782 197412 158788
rect 197818 156904 197874 156913
rect 197818 156839 197874 156848
rect 197832 155990 197860 156839
rect 197820 155984 197872 155990
rect 197820 155926 197872 155932
rect 197358 154728 197414 154737
rect 197358 154663 197414 154672
rect 197372 154630 197400 154663
rect 197360 154624 197412 154630
rect 197360 154566 197412 154572
rect 197358 152552 197414 152561
rect 197358 152487 197414 152496
rect 197372 151842 197400 152487
rect 197360 151836 197412 151842
rect 197360 151778 197412 151784
rect 197358 150376 197414 150385
rect 197358 150311 197414 150320
rect 197372 149122 197400 150311
rect 197360 149116 197412 149122
rect 197360 149058 197412 149064
rect 197358 148200 197414 148209
rect 197358 148135 197414 148144
rect 197372 147694 197400 148135
rect 197360 147688 197412 147694
rect 197360 147630 197412 147636
rect 196808 147620 196860 147626
rect 196808 147562 196860 147568
rect 198016 146266 198044 163231
rect 198108 148374 198136 165407
rect 198200 162858 198228 171799
rect 198188 162852 198240 162858
rect 198188 162794 198240 162800
rect 198752 160750 198780 290119
rect 198830 221368 198886 221377
rect 198830 221303 198886 221312
rect 198740 160744 198792 160750
rect 198740 160686 198792 160692
rect 198096 148368 198148 148374
rect 198096 148310 198148 148316
rect 198004 146260 198056 146266
rect 198004 146202 198056 146208
rect 198094 146160 198150 146169
rect 198094 146095 198150 146104
rect 197358 143984 197414 143993
rect 197358 143919 197414 143928
rect 197372 143614 197400 143919
rect 197360 143608 197412 143614
rect 197360 143550 197412 143556
rect 196624 142112 196676 142118
rect 196624 142054 196676 142060
rect 197542 141808 197598 141817
rect 197542 141743 197598 141752
rect 197556 140826 197584 141743
rect 197544 140820 197596 140826
rect 197544 140762 197596 140768
rect 195336 140752 195388 140758
rect 195336 140694 195388 140700
rect 198108 140078 198136 146095
rect 198096 140072 198148 140078
rect 198096 140014 198148 140020
rect 197726 139632 197782 139641
rect 197726 139567 197782 139576
rect 197358 137456 197414 137465
rect 197358 137391 197414 137400
rect 197372 136678 197400 137391
rect 197360 136672 197412 136678
rect 197360 136614 197412 136620
rect 197740 135930 197768 139567
rect 197728 135924 197780 135930
rect 197728 135866 197780 135872
rect 197358 135416 197414 135425
rect 197358 135351 197414 135360
rect 197372 134570 197400 135351
rect 197360 134564 197412 134570
rect 197360 134506 197412 134512
rect 197358 133240 197414 133249
rect 197358 133175 197414 133184
rect 197372 132530 197400 133175
rect 197360 132524 197412 132530
rect 197360 132466 197412 132472
rect 197360 131096 197412 131102
rect 197358 131064 197360 131073
rect 197412 131064 197414 131073
rect 197358 130999 197414 131008
rect 197360 129736 197412 129742
rect 197360 129678 197412 129684
rect 197372 128897 197400 129678
rect 197358 128888 197414 128897
rect 197358 128823 197414 128832
rect 198004 127628 198056 127634
rect 198004 127570 198056 127576
rect 197544 125588 197596 125594
rect 197544 125530 197596 125536
rect 197556 124545 197584 125530
rect 197542 124536 197598 124545
rect 197542 124471 197598 124480
rect 198016 122505 198044 127570
rect 198464 126948 198516 126954
rect 198464 126890 198516 126896
rect 198476 126721 198504 126890
rect 198462 126712 198518 126721
rect 198462 126647 198518 126656
rect 198844 122874 198872 221303
rect 199396 215286 199424 301514
rect 200396 300960 200448 300966
rect 200396 300902 200448 300908
rect 200408 299948 200436 300902
rect 201224 300892 201276 300898
rect 201224 300834 201276 300840
rect 201236 299948 201264 300834
rect 202064 299948 202092 303622
rect 209872 303136 209924 303142
rect 209872 303078 209924 303084
rect 209044 302864 209096 302870
rect 209044 302806 209096 302812
rect 204720 302660 204772 302666
rect 204720 302602 204772 302608
rect 202972 301028 203024 301034
rect 202972 300970 203024 300976
rect 202984 299948 203012 300970
rect 203800 300212 203852 300218
rect 203800 300154 203852 300160
rect 203812 299948 203840 300154
rect 204732 299948 204760 302602
rect 207296 302592 207348 302598
rect 207296 302534 207348 302540
rect 206468 301504 206520 301510
rect 206468 301446 206520 301452
rect 206480 299948 206508 301446
rect 207308 299948 207336 302534
rect 209056 299948 209084 302806
rect 209884 299948 209912 303078
rect 211620 302932 211672 302938
rect 211620 302874 211672 302880
rect 210792 301096 210844 301102
rect 210792 301038 210844 301044
rect 210804 299948 210832 301038
rect 211632 299948 211660 302874
rect 212540 302728 212592 302734
rect 212540 302670 212592 302676
rect 212552 299948 212580 302670
rect 215116 302388 215168 302394
rect 215116 302330 215168 302336
rect 213368 300348 213420 300354
rect 213368 300290 213420 300296
rect 213380 299948 213408 300290
rect 215128 299948 215156 302330
rect 216036 301640 216088 301646
rect 216036 301582 216088 301588
rect 216048 299948 216076 301582
rect 219348 300348 219400 300354
rect 219348 300290 219400 300296
rect 219440 300348 219492 300354
rect 219440 300290 219492 300296
rect 218888 299736 218940 299742
rect 218638 299684 218888 299690
rect 218638 299678 218940 299684
rect 218638 299662 218928 299678
rect 219360 299674 219388 300290
rect 219452 299948 219480 300290
rect 220648 299962 220676 311850
rect 220740 300354 220768 324294
rect 222856 306134 222884 700266
rect 238668 696992 238720 696998
rect 238668 696934 238720 696940
rect 238576 683188 238628 683194
rect 238576 683130 238628 683136
rect 237288 670744 237340 670750
rect 237288 670686 237340 670692
rect 235908 643136 235960 643142
rect 235908 643078 235960 643084
rect 234528 616888 234580 616894
rect 234528 616830 234580 616836
rect 233148 590708 233200 590714
rect 233148 590650 233200 590656
rect 231768 563100 231820 563106
rect 231768 563042 231820 563048
rect 230388 536852 230440 536858
rect 230388 536794 230440 536800
rect 229008 510672 229060 510678
rect 229008 510614 229060 510620
rect 227628 484424 227680 484430
rect 227628 484366 227680 484372
rect 227536 456816 227588 456822
rect 227536 456758 227588 456764
rect 224868 430636 224920 430642
rect 224868 430578 224920 430584
rect 224776 404388 224828 404394
rect 224776 404330 224828 404336
rect 222936 307080 222988 307086
rect 222936 307022 222988 307028
rect 222844 306128 222896 306134
rect 222844 306070 222896 306076
rect 222108 305720 222160 305726
rect 222108 305662 222160 305668
rect 221188 305652 221240 305658
rect 221188 305594 221240 305600
rect 220728 300348 220780 300354
rect 220728 300290 220780 300296
rect 220386 299934 220676 299962
rect 221200 299948 221228 305594
rect 222120 299948 222148 305662
rect 222948 299948 222976 307022
rect 224788 302122 224816 404330
rect 223856 302116 223908 302122
rect 223856 302058 223908 302064
rect 224776 302116 224828 302122
rect 224776 302058 224828 302064
rect 223868 299948 223896 302058
rect 224880 299962 224908 430578
rect 226248 418192 226300 418198
rect 226248 418134 226300 418140
rect 226260 306374 226288 418134
rect 225984 306346 226288 306374
rect 225984 299962 226012 306346
rect 227548 300354 227576 456758
rect 226432 300348 226484 300354
rect 226432 300290 226484 300296
rect 227536 300348 227588 300354
rect 227536 300290 227588 300296
rect 224710 299934 224908 299962
rect 225630 299934 226012 299962
rect 226444 299948 226472 300290
rect 227640 299962 227668 484366
rect 228916 470620 228968 470626
rect 228916 470562 228968 470568
rect 228928 302122 228956 470562
rect 228180 302116 228232 302122
rect 228180 302058 228232 302064
rect 228916 302116 228968 302122
rect 228916 302058 228968 302064
rect 227378 299934 227668 299962
rect 228192 299948 228220 302058
rect 229020 299948 229048 510614
rect 230400 299962 230428 536794
rect 231676 524476 231728 524482
rect 231676 524418 231728 524424
rect 231688 302122 231716 524418
rect 230756 302116 230808 302122
rect 230756 302058 230808 302064
rect 231676 302116 231728 302122
rect 231676 302058 231728 302064
rect 229954 299934 230428 299962
rect 230768 299948 230796 302058
rect 231780 299962 231808 563042
rect 233160 306374 233188 590650
rect 234436 576904 234488 576910
rect 234436 576846 234488 576852
rect 232976 306346 233188 306374
rect 232976 299962 233004 306346
rect 234448 302122 234476 576846
rect 233424 302116 233476 302122
rect 233424 302058 233476 302064
rect 234436 302116 234488 302122
rect 234436 302058 234488 302064
rect 231702 299934 231808 299962
rect 232530 299934 233004 299962
rect 233436 299948 233464 302058
rect 234540 299962 234568 616830
rect 235920 302122 235948 643078
rect 237196 630692 237248 630698
rect 237196 630634 237248 630640
rect 237208 302122 237236 630634
rect 235172 302116 235224 302122
rect 235172 302058 235224 302064
rect 235908 302116 235960 302122
rect 235908 302058 235960 302064
rect 236000 302116 236052 302122
rect 236000 302058 236052 302064
rect 237196 302116 237248 302122
rect 237196 302058 237248 302064
rect 234278 299934 234568 299962
rect 235184 299948 235212 302058
rect 236012 299948 236040 302058
rect 237300 300098 237328 670686
rect 237748 303000 237800 303006
rect 237748 302942 237800 302948
rect 237208 300070 237328 300098
rect 237208 299962 237236 300070
rect 236854 299934 237236 299962
rect 237760 299948 237788 302942
rect 238588 299948 238616 683130
rect 238680 303006 238708 696934
rect 240324 305788 240376 305794
rect 240324 305730 240376 305736
rect 239496 304292 239548 304298
rect 239496 304234 239548 304240
rect 238668 303000 238720 303006
rect 238668 302942 238720 302948
rect 239508 299948 239536 304234
rect 240336 299948 240364 305730
rect 241440 299962 241468 700266
rect 242176 304842 242204 700402
rect 242164 304836 242216 304842
rect 242164 304778 242216 304784
rect 242072 304360 242124 304366
rect 242072 304302 242124 304308
rect 241270 299934 241468 299962
rect 242084 299948 242112 304302
rect 242992 303544 243044 303550
rect 242992 303486 243044 303492
rect 243004 299948 243032 303486
rect 244200 299962 244228 700402
rect 245476 309800 245528 309806
rect 245476 309742 245528 309748
rect 244740 304428 244792 304434
rect 244740 304370 244792 304376
rect 243846 299934 244228 299962
rect 244752 299948 244780 304370
rect 245488 299962 245516 309742
rect 246960 306374 246988 700538
rect 249064 698964 249116 698970
rect 249064 698906 249116 698912
rect 246776 306346 246988 306374
rect 246776 299962 246804 306346
rect 248420 305992 248472 305998
rect 248420 305934 248472 305940
rect 247316 304564 247368 304570
rect 247316 304506 247368 304512
rect 245488 299934 245594 299962
rect 246422 299934 246804 299962
rect 247328 299948 247356 304506
rect 248432 302274 248460 305934
rect 249076 303550 249104 698906
rect 250996 607912 251048 607918
rect 250996 607854 251048 607860
rect 249432 307284 249484 307290
rect 249432 307226 249484 307232
rect 249064 303544 249116 303550
rect 249064 303486 249116 303492
rect 248340 302246 248460 302274
rect 248340 299962 248368 302246
rect 249444 299962 249472 307226
rect 249892 304768 249944 304774
rect 249892 304710 249944 304716
rect 248170 299934 248368 299962
rect 249090 299934 249472 299962
rect 249904 299948 249932 304710
rect 251008 299962 251036 607854
rect 251824 304700 251876 304706
rect 251824 304642 251876 304648
rect 251640 303000 251692 303006
rect 251640 302942 251692 302948
rect 250838 299934 251036 299962
rect 251652 299948 251680 302942
rect 251836 302258 251864 304642
rect 252480 303006 252508 700606
rect 258080 700528 258132 700534
rect 258080 700470 258132 700476
rect 253204 357468 253256 357474
rect 253204 357410 253256 357416
rect 253216 307562 253244 357410
rect 255320 326392 255372 326398
rect 255320 326334 255372 326340
rect 255332 325694 255360 326334
rect 258092 325694 258120 700470
rect 260104 700392 260156 700398
rect 260104 700334 260156 700340
rect 255332 325666 255544 325694
rect 258092 325666 258304 325694
rect 253204 307556 253256 307562
rect 253204 307498 253256 307504
rect 254308 306128 254360 306134
rect 254308 306070 254360 306076
rect 252560 304836 252612 304842
rect 252560 304778 252612 304784
rect 252468 303000 252520 303006
rect 252468 302942 252520 302948
rect 251824 302252 251876 302258
rect 251824 302194 251876 302200
rect 252572 299948 252600 304778
rect 253388 302252 253440 302258
rect 253388 302194 253440 302200
rect 253400 299948 253428 302194
rect 254320 299948 254348 306070
rect 255136 304632 255188 304638
rect 255136 304574 255188 304580
rect 255148 299948 255176 304574
rect 255516 299962 255544 325666
rect 256240 307216 256292 307222
rect 256240 307158 256292 307164
rect 256252 303346 256280 307158
rect 258080 307148 258132 307154
rect 258080 307090 258132 307096
rect 256884 305924 256936 305930
rect 256884 305866 256936 305872
rect 256240 303340 256292 303346
rect 256240 303282 256292 303288
rect 255516 299934 255990 299962
rect 256896 299948 256924 305866
rect 257712 304496 257764 304502
rect 257712 304438 257764 304444
rect 257724 299948 257752 304438
rect 258092 303074 258120 307090
rect 258080 303068 258132 303074
rect 258080 303010 258132 303016
rect 258276 299962 258304 325666
rect 259460 303340 259512 303346
rect 259460 303282 259512 303288
rect 258276 299934 258658 299962
rect 259472 299948 259500 303282
rect 260116 303006 260144 700334
rect 267660 697610 267688 703520
rect 283852 700670 283880 703520
rect 283840 700664 283892 700670
rect 283840 700606 283892 700612
rect 266360 697604 266412 697610
rect 266360 697546 266412 697552
rect 267648 697604 267700 697610
rect 267648 697546 267700 697552
rect 262220 683256 262272 683262
rect 262220 683198 262272 683204
rect 262232 325694 262260 683198
rect 263692 656940 263744 656946
rect 263692 656882 263744 656888
rect 262232 325666 262536 325694
rect 260380 305856 260432 305862
rect 260380 305798 260432 305804
rect 260104 303000 260156 303006
rect 260104 302942 260156 302948
rect 260392 299948 260420 305798
rect 261208 303068 261260 303074
rect 261208 303010 261260 303016
rect 261220 299948 261248 303010
rect 262128 303000 262180 303006
rect 262128 302942 262180 302948
rect 262140 299948 262168 302942
rect 262508 299962 262536 325666
rect 263232 308440 263284 308446
rect 263232 308382 263284 308388
rect 263244 303006 263272 308382
rect 263232 303000 263284 303006
rect 263232 302942 263284 302948
rect 263704 299962 263732 656882
rect 264980 632120 265032 632126
rect 264980 632062 265032 632068
rect 264992 325694 265020 632062
rect 266372 607918 266400 697546
rect 266360 607912 266412 607918
rect 266360 607854 266412 607860
rect 266360 605872 266412 605878
rect 266360 605814 266412 605820
rect 264992 325666 265112 325694
rect 264704 303000 264756 303006
rect 264704 302942 264756 302948
rect 262508 299934 262982 299962
rect 263704 299934 263902 299962
rect 264716 299948 264744 302942
rect 265084 299962 265112 325666
rect 266372 299962 266400 605814
rect 267740 579692 267792 579698
rect 267740 579634 267792 579640
rect 267280 307488 267332 307494
rect 267280 307430 267332 307436
rect 265084 299934 265558 299962
rect 266372 299934 266478 299962
rect 267292 299948 267320 307430
rect 267752 306374 267780 579634
rect 267832 553444 267884 553450
rect 267832 553386 267884 553392
rect 267844 325694 267872 553386
rect 270500 527196 270552 527202
rect 270500 527138 270552 527144
rect 269764 514820 269816 514826
rect 269764 514762 269816 514768
rect 267844 325666 268608 325694
rect 267752 306346 267872 306374
rect 267844 299962 267872 306346
rect 268580 299962 268608 325666
rect 269776 303006 269804 514762
rect 269948 307420 270000 307426
rect 269948 307362 270000 307368
rect 269764 303000 269816 303006
rect 269764 302942 269816 302948
rect 267844 299934 268226 299962
rect 268580 299934 269054 299962
rect 269960 299948 269988 307362
rect 270512 299962 270540 527138
rect 270592 501016 270644 501022
rect 270592 500958 270644 500964
rect 270604 325694 270632 500958
rect 273260 474768 273312 474774
rect 273260 474710 273312 474716
rect 270604 325666 271368 325694
rect 271340 299962 271368 325666
rect 272524 303000 272576 303006
rect 272524 302942 272576 302948
rect 270512 299934 270802 299962
rect 271340 299934 271722 299962
rect 272536 299948 272564 302942
rect 273272 299962 273300 474710
rect 273352 448588 273404 448594
rect 273352 448530 273404 448536
rect 273364 325694 273392 448530
rect 276020 422340 276072 422346
rect 276020 422282 276072 422288
rect 273364 325666 273944 325694
rect 273916 299962 273944 325666
rect 275100 306060 275152 306066
rect 275100 306002 275152 306008
rect 273272 299934 273378 299962
rect 273916 299934 274298 299962
rect 275112 299948 275140 306002
rect 276032 299948 276060 422282
rect 276112 397520 276164 397526
rect 276112 397462 276164 397468
rect 276124 325694 276152 397462
rect 277400 371272 277452 371278
rect 277400 371214 277452 371220
rect 277412 325694 277440 371214
rect 278780 345092 278832 345098
rect 278780 345034 278832 345040
rect 278792 325694 278820 345034
rect 276124 325666 276520 325694
rect 277412 325666 278176 325694
rect 278792 325666 279096 325694
rect 276492 299962 276520 325666
rect 277768 307352 277820 307358
rect 277768 307294 277820 307300
rect 276492 299934 276874 299962
rect 277780 299948 277808 307294
rect 278148 299962 278176 325666
rect 279068 299962 279096 325666
rect 280896 318844 280948 318850
rect 280896 318786 280948 318792
rect 280344 307556 280396 307562
rect 280344 307498 280396 307504
rect 278148 299934 278622 299962
rect 279068 299934 279542 299962
rect 280356 299948 280384 307498
rect 280908 299962 280936 318786
rect 282828 305040 282880 305046
rect 282828 304982 282880 304988
rect 282840 302274 282868 304982
rect 299492 304774 299520 703582
rect 299952 703474 299980 703582
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429212 703582 429700 703610
rect 300136 703474 300164 703520
rect 299952 703446 300164 703474
rect 332520 703050 332548 703520
rect 331220 703044 331272 703050
rect 331220 702986 331272 702992
rect 332508 703044 332560 703050
rect 332508 702986 332560 702992
rect 300768 337476 300820 337482
rect 300768 337418 300820 337424
rect 299480 304768 299532 304774
rect 299480 304710 299532 304716
rect 297732 303748 297784 303754
rect 297732 303690 297784 303696
rect 285588 302796 285640 302802
rect 285588 302738 285640 302744
rect 282840 302246 282960 302274
rect 282092 300280 282144 300286
rect 282092 300222 282144 300228
rect 280908 299934 281290 299962
rect 282104 299948 282132 300222
rect 282932 299948 282960 302246
rect 284668 301436 284720 301442
rect 284668 301378 284720 301384
rect 283840 301164 283892 301170
rect 283840 301106 283892 301112
rect 283852 299948 283880 301106
rect 284680 299948 284708 301378
rect 285600 299948 285628 302738
rect 288164 302524 288216 302530
rect 288164 302466 288216 302472
rect 285680 302252 285732 302258
rect 285680 302194 285732 302200
rect 219348 299668 219400 299674
rect 219348 299610 219400 299616
rect 208308 299600 208360 299606
rect 205574 299538 205680 299554
rect 208242 299548 208308 299554
rect 208242 299542 208360 299548
rect 205574 299532 205692 299538
rect 205574 299526 205640 299532
rect 208242 299526 208348 299542
rect 205640 299474 205692 299480
rect 216772 299464 216824 299470
rect 214314 299402 214696 299418
rect 216772 299406 216824 299412
rect 217414 299432 217470 299441
rect 214314 299396 214708 299402
rect 214314 299390 214656 299396
rect 214656 299338 214708 299344
rect 216784 299334 216812 299406
rect 217414 299367 217470 299376
rect 217966 299432 218022 299441
rect 217966 299367 217968 299376
rect 217428 299334 217456 299367
rect 218020 299367 218022 299376
rect 217968 299338 218020 299344
rect 285692 299334 285720 302194
rect 286416 301572 286468 301578
rect 286416 301514 286468 301520
rect 286428 299948 286456 301514
rect 287152 300076 287204 300082
rect 287152 300018 287204 300024
rect 287164 299962 287192 300018
rect 287164 299934 287362 299962
rect 288176 299948 288204 302466
rect 290832 302456 290884 302462
rect 290832 302398 290884 302404
rect 289912 302252 289964 302258
rect 289912 302194 289964 302200
rect 289924 299948 289952 302194
rect 290844 299948 290872 302398
rect 293408 302320 293460 302326
rect 293408 302262 293460 302268
rect 292488 301368 292540 301374
rect 292488 301310 292540 301316
rect 291660 300144 291712 300150
rect 291660 300086 291712 300092
rect 291672 299948 291700 300086
rect 292500 299948 292528 301310
rect 293420 299948 293448 302262
rect 296904 301300 296956 301306
rect 296904 301242 296956 301248
rect 293960 300008 294012 300014
rect 294012 299956 294262 299962
rect 293960 299950 294262 299956
rect 293972 299934 294262 299950
rect 294800 299946 295182 299962
rect 296916 299948 296944 301242
rect 297744 299948 297772 303690
rect 300780 302802 300808 337418
rect 331232 305998 331260 702986
rect 348804 699718 348832 703520
rect 364996 699718 365024 703520
rect 397472 699718 397500 703520
rect 413664 700602 413692 703520
rect 413652 700596 413704 700602
rect 413652 700538 413704 700544
rect 347044 699712 347096 699718
rect 347044 699654 347096 699660
rect 348792 699712 348844 699718
rect 348792 699654 348844 699660
rect 359464 699712 359516 699718
rect 359464 699654 359516 699660
rect 364984 699712 365036 699718
rect 364984 699654 365036 699660
rect 396724 699712 396776 699718
rect 396724 699654 396776 699660
rect 397460 699712 397512 699718
rect 397460 699654 397512 699660
rect 347056 307290 347084 699654
rect 347044 307284 347096 307290
rect 347044 307226 347096 307232
rect 331220 305992 331272 305998
rect 331220 305934 331272 305940
rect 359476 304570 359504 699654
rect 371882 369744 371938 369753
rect 371882 369679 371938 369688
rect 371606 369200 371662 369209
rect 371606 369135 371662 369144
rect 371620 368966 371648 369135
rect 371608 368960 371660 368966
rect 371608 368902 371660 368908
rect 371698 368112 371754 368121
rect 371698 368047 371754 368056
rect 371606 367568 371662 367577
rect 371606 367503 371662 367512
rect 371620 367198 371648 367503
rect 371608 367192 371660 367198
rect 371608 367134 371660 367140
rect 371712 367130 371740 368047
rect 371700 367124 371752 367130
rect 371700 367066 371752 367072
rect 371238 367024 371294 367033
rect 371238 366959 371294 366968
rect 371252 365838 371280 366959
rect 371514 366480 371570 366489
rect 371514 366415 371570 366424
rect 371240 365832 371292 365838
rect 371240 365774 371292 365780
rect 371528 365770 371556 366415
rect 371606 365936 371662 365945
rect 371606 365871 371608 365880
rect 371660 365871 371662 365880
rect 371608 365842 371660 365848
rect 371516 365764 371568 365770
rect 371516 365706 371568 365712
rect 371238 365392 371294 365401
rect 371238 365327 371294 365336
rect 371252 364682 371280 365327
rect 371606 364848 371662 364857
rect 371606 364783 371662 364792
rect 371240 364676 371292 364682
rect 371240 364618 371292 364624
rect 371620 364410 371648 364783
rect 371608 364404 371660 364410
rect 371608 364346 371660 364352
rect 371698 364304 371754 364313
rect 371698 364239 371754 364248
rect 371606 363760 371662 363769
rect 371606 363695 371662 363704
rect 371620 363118 371648 363695
rect 371608 363112 371660 363118
rect 371608 363054 371660 363060
rect 371712 362982 371740 364239
rect 371700 362976 371752 362982
rect 371700 362918 371752 362924
rect 371698 362672 371754 362681
rect 371698 362607 371754 362616
rect 371606 362128 371662 362137
rect 371606 362063 371662 362072
rect 371620 361690 371648 362063
rect 371608 361684 371660 361690
rect 371608 361626 371660 361632
rect 371712 361622 371740 362607
rect 371700 361616 371752 361622
rect 371606 361584 371662 361593
rect 371700 361558 371752 361564
rect 371606 361519 371608 361528
rect 371660 361519 371662 361528
rect 371608 361490 371660 361496
rect 371422 361040 371478 361049
rect 371422 360975 371478 360984
rect 371436 360398 371464 360975
rect 371606 360496 371662 360505
rect 371606 360431 371608 360440
rect 371660 360431 371662 360440
rect 371608 360402 371660 360408
rect 371424 360392 371476 360398
rect 371424 360334 371476 360340
rect 371896 359582 371924 369679
rect 374184 368960 374236 368966
rect 374184 368902 374236 368908
rect 372066 368656 372122 368665
rect 372066 368591 372122 368600
rect 371884 359576 371936 359582
rect 371884 359518 371936 359524
rect 372080 359514 372108 368591
rect 372526 363216 372582 363225
rect 372582 363174 372660 363202
rect 372526 363151 372582 363160
rect 372342 360088 372398 360097
rect 372342 360023 372398 360032
rect 372158 359544 372214 359553
rect 372068 359508 372120 359514
rect 372158 359479 372214 359488
rect 372068 359450 372120 359456
rect 371974 359000 372030 359009
rect 371974 358935 372030 358944
rect 371698 358456 371754 358465
rect 371698 358391 371754 358400
rect 371606 357912 371662 357921
rect 371606 357847 371662 357856
rect 371620 357474 371648 357847
rect 371712 357542 371740 358391
rect 371700 357536 371752 357542
rect 371700 357478 371752 357484
rect 371608 357468 371660 357474
rect 371608 357410 371660 357416
rect 371606 357368 371662 357377
rect 371606 357303 371662 357312
rect 371514 356824 371570 356833
rect 371514 356759 371570 356768
rect 371238 356280 371294 356289
rect 371238 356215 371294 356224
rect 371252 356182 371280 356215
rect 371240 356176 371292 356182
rect 371240 356118 371292 356124
rect 371528 356114 371556 356759
rect 371620 356250 371648 357303
rect 371608 356244 371660 356250
rect 371608 356186 371660 356192
rect 371516 356108 371568 356114
rect 371516 356050 371568 356056
rect 371606 355736 371662 355745
rect 371606 355671 371662 355680
rect 371514 355192 371570 355201
rect 371514 355127 371570 355136
rect 371528 354822 371556 355127
rect 371516 354816 371568 354822
rect 371516 354758 371568 354764
rect 371620 354754 371648 355671
rect 371608 354748 371660 354754
rect 371608 354690 371660 354696
rect 371330 354648 371386 354657
rect 371330 354583 371386 354592
rect 371344 353394 371372 354583
rect 371698 354104 371754 354113
rect 371698 354039 371754 354048
rect 371514 353560 371570 353569
rect 371514 353495 371570 353504
rect 371332 353388 371384 353394
rect 371332 353330 371384 353336
rect 369306 350568 369362 350577
rect 369306 350503 369362 350512
rect 369320 345014 369348 350503
rect 370318 348800 370374 348809
rect 370318 348735 370374 348744
rect 369398 347440 369454 347449
rect 369398 347375 369454 347384
rect 369136 344986 369348 345014
rect 360212 340054 360962 340082
rect 359464 304564 359516 304570
rect 359464 304506 359516 304512
rect 311164 302932 311216 302938
rect 311164 302874 311216 302880
rect 309784 302864 309836 302870
rect 309784 302806 309836 302812
rect 299480 302796 299532 302802
rect 299480 302738 299532 302744
rect 300768 302796 300820 302802
rect 300768 302738 300820 302744
rect 298652 301232 298704 301238
rect 298652 301174 298704 301180
rect 298664 299948 298692 301174
rect 299492 299948 299520 302738
rect 301504 301640 301556 301646
rect 301504 301582 301556 301588
rect 294788 299940 295182 299946
rect 294840 299934 295182 299940
rect 294788 299882 294840 299888
rect 295708 299872 295760 299878
rect 288728 299810 289110 299826
rect 295760 299820 296010 299826
rect 295708 299814 296010 299820
rect 288716 299804 289110 299810
rect 288768 299798 289110 299804
rect 295720 299798 296010 299814
rect 288716 299746 288768 299752
rect 216772 299328 216824 299334
rect 217416 299328 217468 299334
rect 217230 299296 217286 299305
rect 216772 299270 216824 299276
rect 216890 299254 217230 299282
rect 217692 299328 217744 299334
rect 217416 299270 217468 299276
rect 217690 299296 217692 299305
rect 218060 299328 218112 299334
rect 217744 299296 217746 299305
rect 217230 299231 217286 299240
rect 217810 299276 218060 299282
rect 217810 299270 218112 299276
rect 285680 299328 285732 299334
rect 285680 299270 285732 299276
rect 217810 299254 218100 299270
rect 217690 299231 217746 299240
rect 199844 298308 199896 298314
rect 199844 298250 199896 298256
rect 199856 296721 199884 298250
rect 199842 296712 199898 296721
rect 199842 296647 199898 296656
rect 301516 245614 301544 301582
rect 307024 301504 307076 301510
rect 307024 301446 307076 301452
rect 305644 300212 305696 300218
rect 305644 300154 305696 300160
rect 302790 298480 302846 298489
rect 302790 298415 302846 298424
rect 302804 298382 302832 298415
rect 302792 298376 302844 298382
rect 302792 298318 302844 298324
rect 302976 296812 303028 296818
rect 302976 296754 303028 296760
rect 302884 296744 302936 296750
rect 302884 296686 302936 296692
rect 302792 295384 302844 295390
rect 302790 295352 302792 295361
rect 302844 295352 302846 295361
rect 302790 295287 302846 295296
rect 302238 292224 302294 292233
rect 302238 292159 302294 292168
rect 302252 291514 302280 292159
rect 302240 291508 302292 291514
rect 302240 291450 302292 291456
rect 302698 289096 302754 289105
rect 302698 289031 302754 289040
rect 302712 288454 302740 289031
rect 302700 288448 302752 288454
rect 302700 288390 302752 288396
rect 302790 285968 302846 285977
rect 302790 285903 302846 285912
rect 302804 285734 302832 285903
rect 302792 285728 302844 285734
rect 302792 285670 302844 285676
rect 302514 282840 302570 282849
rect 302514 282775 302570 282784
rect 302528 281586 302556 282775
rect 302516 281580 302568 281586
rect 302516 281522 302568 281528
rect 302790 279712 302846 279721
rect 302790 279647 302846 279656
rect 302804 278798 302832 279647
rect 302792 278792 302844 278798
rect 302792 278734 302844 278740
rect 302790 276584 302846 276593
rect 302790 276519 302846 276528
rect 302804 276078 302832 276519
rect 302792 276072 302844 276078
rect 302792 276014 302844 276020
rect 302896 270337 302924 296686
rect 302988 273465 303016 296754
rect 304264 291508 304316 291514
rect 304264 291450 304316 291456
rect 302974 273456 303030 273465
rect 302974 273391 303030 273400
rect 302882 270328 302938 270337
rect 302882 270263 302938 270272
rect 303252 268388 303304 268394
rect 303252 268330 303304 268336
rect 303264 267209 303292 268330
rect 303250 267200 303306 267209
rect 303250 267135 303306 267144
rect 302792 264920 302844 264926
rect 302792 264862 302844 264868
rect 302804 264081 302832 264862
rect 302790 264072 302846 264081
rect 302790 264007 302846 264016
rect 302792 262200 302844 262206
rect 302792 262142 302844 262148
rect 302804 260953 302832 262142
rect 302790 260944 302846 260953
rect 302790 260879 302846 260888
rect 302790 257816 302846 257825
rect 302790 257751 302846 257760
rect 302804 256766 302832 257751
rect 302792 256760 302844 256766
rect 302792 256702 302844 256708
rect 302330 254688 302386 254697
rect 302330 254623 302386 254632
rect 302344 253978 302372 254623
rect 302332 253972 302384 253978
rect 302332 253914 302384 253920
rect 302974 251560 303030 251569
rect 302974 251495 303030 251504
rect 302792 248464 302844 248470
rect 302790 248432 302792 248441
rect 302844 248432 302846 248441
rect 302790 248367 302846 248376
rect 301504 245608 301556 245614
rect 301504 245550 301556 245556
rect 302882 245304 302938 245313
rect 302882 245239 302938 245248
rect 302698 229664 302754 229673
rect 302698 229599 302754 229608
rect 302712 229094 302740 229599
rect 302712 229066 302832 229094
rect 302698 226536 302754 226545
rect 302698 226471 302754 226480
rect 302712 224330 302740 226471
rect 302804 224398 302832 229066
rect 302896 225622 302924 245239
rect 302988 239426 303016 251495
rect 303066 242176 303122 242185
rect 303066 242111 303122 242120
rect 302976 239420 303028 239426
rect 302976 239362 303028 239368
rect 302974 235920 303030 235929
rect 302974 235855 303030 235864
rect 302884 225616 302936 225622
rect 302884 225558 302936 225564
rect 302792 224392 302844 224398
rect 302792 224334 302844 224340
rect 302700 224324 302752 224330
rect 302700 224266 302752 224272
rect 302988 224262 303016 235855
rect 303080 231130 303108 242111
rect 303158 239048 303214 239057
rect 303158 238983 303214 238992
rect 303068 231124 303120 231130
rect 303068 231066 303120 231072
rect 303172 229770 303200 238983
rect 303250 232792 303306 232801
rect 303250 232727 303306 232736
rect 303160 229764 303212 229770
rect 303160 229706 303212 229712
rect 303264 227050 303292 232727
rect 303252 227044 303304 227050
rect 303252 226986 303304 226992
rect 302976 224256 303028 224262
rect 302976 224198 303028 224204
rect 302792 223576 302844 223582
rect 302792 223518 302844 223524
rect 302804 223417 302832 223518
rect 302790 223408 302846 223417
rect 302790 223343 302846 223352
rect 302792 220788 302844 220794
rect 302792 220730 302844 220736
rect 302804 220289 302832 220730
rect 302790 220280 302846 220289
rect 302790 220215 302846 220224
rect 302516 218000 302568 218006
rect 302516 217942 302568 217948
rect 302528 217161 302556 217942
rect 302514 217152 302570 217161
rect 302514 217087 302570 217096
rect 199384 215280 199436 215286
rect 199384 215222 199436 215228
rect 302792 215280 302844 215286
rect 302792 215222 302844 215228
rect 302804 214033 302832 215222
rect 302790 214024 302846 214033
rect 302790 213959 302846 213968
rect 302792 211132 302844 211138
rect 302792 211074 302844 211080
rect 302804 210905 302832 211074
rect 302790 210896 302846 210905
rect 302790 210831 302846 210840
rect 302330 207768 302386 207777
rect 302330 207703 302386 207712
rect 302344 207058 302372 207703
rect 302332 207052 302384 207058
rect 302332 206994 302384 207000
rect 302698 204640 302754 204649
rect 302698 204575 302754 204584
rect 302712 204338 302740 204575
rect 302700 204332 302752 204338
rect 302700 204274 302752 204280
rect 302792 201544 302844 201550
rect 302790 201512 302792 201521
rect 302844 201512 302846 201521
rect 302790 201447 302846 201456
rect 302790 198384 302846 198393
rect 302790 198319 302846 198328
rect 302804 197402 302832 198319
rect 302792 197396 302844 197402
rect 302792 197338 302844 197344
rect 302884 196036 302936 196042
rect 302884 195978 302936 195984
rect 302332 195968 302384 195974
rect 302332 195910 302384 195916
rect 302344 195265 302372 195910
rect 302330 195256 302386 195265
rect 302330 195191 302386 195200
rect 301504 193860 301556 193866
rect 301504 193802 301556 193808
rect 198832 122868 198884 122874
rect 198832 122810 198884 122816
rect 198002 122496 198058 122505
rect 198002 122431 198058 122440
rect 197544 121440 197596 121446
rect 197544 121382 197596 121388
rect 197556 120329 197584 121382
rect 197542 120320 197598 120329
rect 197542 120255 197598 120264
rect 197912 118652 197964 118658
rect 197912 118594 197964 118600
rect 197924 118153 197952 118594
rect 197910 118144 197966 118153
rect 197910 118079 197966 118088
rect 198372 116680 198424 116686
rect 198372 116622 198424 116628
rect 198384 115977 198412 116622
rect 198370 115968 198426 115977
rect 198370 115903 198426 115912
rect 197360 114504 197412 114510
rect 197360 114446 197412 114452
rect 197372 113801 197400 114446
rect 197358 113792 197414 113801
rect 197358 113727 197414 113736
rect 197360 111784 197412 111790
rect 197358 111752 197360 111761
rect 197412 111752 197414 111761
rect 197358 111687 197414 111696
rect 197360 110424 197412 110430
rect 197360 110366 197412 110372
rect 197372 109585 197400 110366
rect 197358 109576 197414 109585
rect 197358 109511 197414 109520
rect 198556 107636 198608 107642
rect 198556 107578 198608 107584
rect 198568 107409 198596 107578
rect 198554 107400 198610 107409
rect 198554 107335 198610 107344
rect 197544 106276 197596 106282
rect 197544 106218 197596 106224
rect 197556 105233 197584 106218
rect 197542 105224 197598 105233
rect 197542 105159 197598 105168
rect 197912 103488 197964 103494
rect 197912 103430 197964 103436
rect 197924 103057 197952 103430
rect 197910 103048 197966 103057
rect 197910 102983 197966 102992
rect 197544 102128 197596 102134
rect 197544 102070 197596 102076
rect 197556 101017 197584 102070
rect 301516 101386 301544 193802
rect 302792 193180 302844 193186
rect 302792 193122 302844 193128
rect 302804 192137 302832 193122
rect 302790 192128 302846 192137
rect 302790 192063 302846 192072
rect 302792 189032 302844 189038
rect 302790 189000 302792 189009
rect 302844 189000 302846 189009
rect 302790 188935 302846 188944
rect 302700 186312 302752 186318
rect 302700 186254 302752 186260
rect 302712 185881 302740 186254
rect 302698 185872 302754 185881
rect 302698 185807 302754 185816
rect 302792 180124 302844 180130
rect 302792 180066 302844 180072
rect 302804 179625 302832 180066
rect 302790 179616 302846 179625
rect 302790 179551 302846 179560
rect 302790 176488 302846 176497
rect 302790 176423 302846 176432
rect 302804 175982 302832 176423
rect 302792 175976 302844 175982
rect 302792 175918 302844 175924
rect 302896 173369 302924 195978
rect 302976 195288 303028 195294
rect 302976 195230 303028 195236
rect 302988 182753 303016 195230
rect 304276 194546 304304 291450
rect 304264 194540 304316 194546
rect 304264 194482 304316 194488
rect 302974 182744 303030 182753
rect 302974 182679 303030 182688
rect 302882 173360 302938 173369
rect 302882 173295 302938 173304
rect 302792 170400 302844 170406
rect 302792 170342 302844 170348
rect 302804 170241 302832 170342
rect 302790 170232 302846 170241
rect 302790 170167 302846 170176
rect 303066 167104 303122 167113
rect 303066 167039 303122 167048
rect 302882 163976 302938 163985
rect 302882 163911 302938 163920
rect 302514 160848 302570 160857
rect 302514 160783 302570 160792
rect 302528 153202 302556 160783
rect 302790 157720 302846 157729
rect 302790 157655 302846 157664
rect 302606 154592 302662 154601
rect 302606 154527 302662 154536
rect 302516 153196 302568 153202
rect 302516 153138 302568 153144
rect 302620 153134 302648 154527
rect 302608 153128 302660 153134
rect 302608 153070 302660 153076
rect 302804 153066 302832 157655
rect 302896 155922 302924 163911
rect 303080 161430 303108 167039
rect 303068 161424 303120 161430
rect 303068 161366 303120 161372
rect 302884 155916 302936 155922
rect 302884 155858 302936 155864
rect 302792 153060 302844 153066
rect 302792 153002 302844 153008
rect 302700 151768 302752 151774
rect 302700 151710 302752 151716
rect 302712 151473 302740 151710
rect 302698 151464 302754 151473
rect 302698 151399 302754 151408
rect 302332 149048 302384 149054
rect 302332 148990 302384 148996
rect 302344 148345 302372 148990
rect 302330 148336 302386 148345
rect 302330 148271 302386 148280
rect 302792 146260 302844 146266
rect 302792 146202 302844 146208
rect 302804 145217 302832 146202
rect 302790 145208 302846 145217
rect 302790 145143 302846 145152
rect 302792 142112 302844 142118
rect 302790 142080 302792 142089
rect 302844 142080 302846 142089
rect 302790 142015 302846 142024
rect 302700 139392 302752 139398
rect 302700 139334 302752 139340
rect 302712 138961 302740 139334
rect 302698 138952 302754 138961
rect 302698 138887 302754 138896
rect 302882 135824 302938 135833
rect 302882 135759 302938 135768
rect 302606 129568 302662 129577
rect 302606 129503 302662 129512
rect 302620 125254 302648 129503
rect 302790 126440 302846 126449
rect 302790 126375 302846 126384
rect 302608 125248 302660 125254
rect 302608 125190 302660 125196
rect 302804 125118 302832 126375
rect 302792 125112 302844 125118
rect 302792 125054 302844 125060
rect 302896 125050 302924 135759
rect 302974 132696 303030 132705
rect 302974 132631 303030 132640
rect 302988 125186 303016 132631
rect 302976 125180 303028 125186
rect 302976 125122 303028 125128
rect 302884 125044 302936 125050
rect 302884 124986 302936 124992
rect 302792 124160 302844 124166
rect 302792 124102 302844 124108
rect 302804 123321 302832 124102
rect 302976 123616 303028 123622
rect 302976 123558 303028 123564
rect 302884 123480 302936 123486
rect 302884 123422 302936 123428
rect 302790 123312 302846 123321
rect 302790 123247 302846 123256
rect 302516 121440 302568 121446
rect 302516 121382 302568 121388
rect 302528 120193 302556 121382
rect 302514 120184 302570 120193
rect 302514 120119 302570 120128
rect 302792 117292 302844 117298
rect 302792 117234 302844 117240
rect 302804 117065 302832 117234
rect 302790 117056 302846 117065
rect 302790 116991 302846 117000
rect 302792 111784 302844 111790
rect 302792 111726 302844 111732
rect 302804 110809 302832 111726
rect 302790 110800 302846 110809
rect 302790 110735 302846 110744
rect 302792 108996 302844 109002
rect 302792 108938 302844 108944
rect 302804 107681 302832 108938
rect 302790 107672 302846 107681
rect 302790 107607 302846 107616
rect 302896 104553 302924 123422
rect 302988 113937 303016 123558
rect 302974 113928 303030 113937
rect 302974 113863 303030 113872
rect 302882 104544 302938 104553
rect 302882 104479 302938 104488
rect 302792 102808 302844 102814
rect 302792 102750 302844 102756
rect 302804 101561 302832 102750
rect 302790 101552 302846 101561
rect 302790 101487 302846 101496
rect 300216 101380 300268 101386
rect 300216 101322 300268 101328
rect 301504 101380 301556 101386
rect 301504 101322 301556 101328
rect 197542 101008 197598 101017
rect 197542 100943 197598 100952
rect 300228 100722 300256 101322
rect 299874 100694 300256 100722
rect 258106 100298 258212 100314
rect 258106 100292 258224 100298
rect 258106 100286 258172 100292
rect 258172 100234 258224 100240
rect 255780 100224 255832 100230
rect 255622 100172 255780 100178
rect 255622 100166 255832 100172
rect 255622 100150 255820 100166
rect 260682 100162 260788 100178
rect 260682 100156 260800 100162
rect 260682 100150 260748 100156
rect 260748 100098 260800 100104
rect 195244 100088 195296 100094
rect 299572 100088 299624 100094
rect 195244 100030 195296 100036
rect 180708 99340 180760 99346
rect 180708 99282 180760 99288
rect 174544 99272 174596 99278
rect 174544 99214 174596 99220
rect 173808 97776 173860 97782
rect 173808 97718 173860 97724
rect 161388 96416 161440 96422
rect 161388 96358 161440 96364
rect 158628 95124 158680 95130
rect 158628 95066 158680 95072
rect 157984 71732 158036 71738
rect 157984 71674 158036 71680
rect 158076 71052 158128 71058
rect 158076 70994 158128 71000
rect 154212 4140 154264 4146
rect 154212 4082 154264 4088
rect 155224 4140 155276 4146
rect 155224 4082 155276 4088
rect 155408 4140 155460 4146
rect 155408 4082 155460 4088
rect 156696 4140 156748 4146
rect 156696 4082 156748 4088
rect 153028 2746 153148 2774
rect 153028 480 153056 2746
rect 154224 480 154252 4082
rect 155420 480 155448 4082
rect 157800 3596 157852 3602
rect 157800 3538 157852 3544
rect 156604 3392 156656 3398
rect 156604 3334 156656 3340
rect 156616 480 156644 3334
rect 157812 480 157840 3538
rect 158088 3398 158116 70994
rect 158640 3602 158668 95066
rect 160008 92404 160060 92410
rect 160008 92346 160060 92352
rect 160020 3602 160048 92346
rect 161400 4146 161428 96358
rect 169668 96348 169720 96354
rect 169668 96290 169720 96296
rect 165528 96280 165580 96286
rect 165528 96222 165580 96228
rect 162768 95192 162820 95198
rect 162768 95134 162820 95140
rect 162780 6914 162808 95134
rect 164148 92472 164200 92478
rect 164148 92414 164200 92420
rect 162504 6886 162808 6914
rect 160100 4140 160152 4146
rect 160100 4082 160152 4088
rect 161388 4140 161440 4146
rect 161388 4082 161440 4088
rect 161480 4140 161532 4146
rect 161480 4082 161532 4088
rect 158628 3596 158680 3602
rect 158628 3538 158680 3544
rect 158904 3596 158956 3602
rect 158904 3538 158956 3544
rect 160008 3596 160060 3602
rect 160008 3538 160060 3544
rect 158076 3392 158128 3398
rect 158076 3334 158128 3340
rect 158916 480 158944 3538
rect 160112 480 160140 4082
rect 161492 4026 161520 4082
rect 161308 3998 161520 4026
rect 161308 480 161336 3998
rect 162504 480 162532 6886
rect 164160 3602 164188 92414
rect 165540 3602 165568 96222
rect 166264 96144 166316 96150
rect 166264 96086 166316 96092
rect 163688 3596 163740 3602
rect 163688 3538 163740 3544
rect 164148 3596 164200 3602
rect 164148 3538 164200 3544
rect 164884 3596 164936 3602
rect 164884 3538 164936 3544
rect 165528 3596 165580 3602
rect 165528 3538 165580 3544
rect 166080 3596 166132 3602
rect 166080 3538 166132 3544
rect 163700 480 163728 3538
rect 164896 480 164924 3538
rect 166092 480 166120 3538
rect 166276 3330 166304 96086
rect 166908 93696 166960 93702
rect 166908 93638 166960 93644
rect 166920 3602 166948 93638
rect 169024 90976 169076 90982
rect 169024 90918 169076 90924
rect 169036 3602 169064 90918
rect 166908 3596 166960 3602
rect 166908 3538 166960 3544
rect 167184 3596 167236 3602
rect 167184 3538 167236 3544
rect 169024 3596 169076 3602
rect 169024 3538 169076 3544
rect 169576 3596 169628 3602
rect 169576 3538 169628 3544
rect 166264 3324 166316 3330
rect 166264 3266 166316 3272
rect 167196 480 167224 3538
rect 168380 3392 168432 3398
rect 168380 3334 168432 3340
rect 168392 480 168420 3334
rect 169588 480 169616 3538
rect 169680 3398 169708 96290
rect 173164 96212 173216 96218
rect 173164 96154 173216 96160
rect 170404 93764 170456 93770
rect 170404 93706 170456 93712
rect 170416 3602 170444 93706
rect 171048 91724 171100 91730
rect 171048 91666 171100 91672
rect 171060 6914 171088 91666
rect 170784 6886 171088 6914
rect 170404 3596 170456 3602
rect 170404 3538 170456 3544
rect 169668 3392 169720 3398
rect 169668 3334 169720 3340
rect 170784 480 170812 6886
rect 172152 4072 172204 4078
rect 172152 4014 172204 4020
rect 172164 3806 172192 4014
rect 172152 3800 172204 3806
rect 172152 3742 172204 3748
rect 173176 3602 173204 96154
rect 173820 96014 173848 97718
rect 173808 96008 173860 96014
rect 173808 95950 173860 95956
rect 171968 3596 172020 3602
rect 171968 3538 172020 3544
rect 173164 3596 173216 3602
rect 173164 3538 173216 3544
rect 171980 480 172008 3538
rect 174556 3398 174584 99214
rect 176568 96552 176620 96558
rect 176568 96494 176620 96500
rect 176580 3602 176608 96494
rect 179328 95872 179380 95878
rect 179328 95814 179380 95820
rect 177948 94444 178000 94450
rect 177948 94386 178000 94392
rect 177856 19984 177908 19990
rect 177856 19926 177908 19932
rect 175464 3596 175516 3602
rect 175464 3538 175516 3544
rect 176568 3596 176620 3602
rect 176568 3538 176620 3544
rect 176660 3596 176712 3602
rect 176660 3538 176712 3544
rect 173164 3392 173216 3398
rect 173164 3334 173216 3340
rect 174544 3392 174596 3398
rect 174544 3334 174596 3340
rect 173176 480 173204 3334
rect 174268 3052 174320 3058
rect 174268 2994 174320 3000
rect 174280 480 174308 2994
rect 175476 480 175504 3538
rect 176672 480 176700 3538
rect 177868 480 177896 19926
rect 177960 3602 177988 94386
rect 179340 6914 179368 95814
rect 179064 6886 179368 6914
rect 177948 3596 178000 3602
rect 177948 3538 178000 3544
rect 179064 480 179092 6886
rect 180720 3602 180748 99282
rect 195888 98592 195940 98598
rect 195888 98534 195940 98540
rect 188988 98048 189040 98054
rect 188988 97990 189040 97996
rect 184204 97912 184256 97918
rect 184204 97854 184256 97860
rect 182824 97844 182876 97850
rect 182824 97786 182876 97792
rect 181444 93832 181496 93838
rect 181444 93774 181496 93780
rect 181456 6914 181484 93774
rect 182088 91656 182140 91662
rect 182088 91598 182140 91604
rect 181364 6886 181484 6914
rect 180248 3596 180300 3602
rect 180248 3538 180300 3544
rect 180708 3596 180760 3602
rect 180708 3538 180760 3544
rect 180260 480 180288 3538
rect 181364 3058 181392 6886
rect 182100 3602 182128 91598
rect 182836 3806 182864 97786
rect 183468 96008 183520 96014
rect 183468 95950 183520 95956
rect 182824 3800 182876 3806
rect 182824 3742 182876 3748
rect 183480 3602 183508 95950
rect 184216 3942 184244 97854
rect 186964 96484 187016 96490
rect 186964 96426 187016 96432
rect 184848 93084 184900 93090
rect 184848 93026 184900 93032
rect 184204 3936 184256 3942
rect 184204 3878 184256 3884
rect 184860 3602 184888 93026
rect 186976 3602 187004 96426
rect 188344 93016 188396 93022
rect 188344 92958 188396 92964
rect 187056 91044 187108 91050
rect 187056 90986 187108 90992
rect 181444 3596 181496 3602
rect 181444 3538 181496 3544
rect 182088 3596 182140 3602
rect 182088 3538 182140 3544
rect 182548 3596 182600 3602
rect 182548 3538 182600 3544
rect 183468 3596 183520 3602
rect 183468 3538 183520 3544
rect 183744 3596 183796 3602
rect 183744 3538 183796 3544
rect 184848 3596 184900 3602
rect 184848 3538 184900 3544
rect 186136 3596 186188 3602
rect 186136 3538 186188 3544
rect 186964 3596 187016 3602
rect 186964 3538 187016 3544
rect 181352 3052 181404 3058
rect 181352 2994 181404 3000
rect 181456 480 181484 3538
rect 182560 480 182588 3538
rect 183756 480 183784 3538
rect 184940 3392 184992 3398
rect 184940 3334 184992 3340
rect 184952 480 184980 3334
rect 186148 480 186176 3538
rect 187068 3398 187096 90986
rect 188356 3602 188384 92958
rect 189000 3602 189028 97990
rect 191104 97980 191156 97986
rect 191104 97922 191156 97928
rect 189724 4072 189776 4078
rect 189724 4014 189776 4020
rect 187332 3596 187384 3602
rect 187332 3538 187384 3544
rect 188344 3596 188396 3602
rect 188344 3538 188396 3544
rect 188528 3596 188580 3602
rect 188528 3538 188580 3544
rect 188988 3596 189040 3602
rect 188988 3538 189040 3544
rect 187056 3392 187108 3398
rect 187056 3334 187108 3340
rect 187344 480 187372 3538
rect 188540 480 188568 3538
rect 189736 480 189764 4014
rect 191116 3738 191144 97922
rect 192576 97232 192628 97238
rect 192576 97174 192628 97180
rect 191196 96620 191248 96626
rect 191196 96562 191248 96568
rect 191208 4078 191236 96562
rect 192484 94376 192536 94382
rect 192484 94318 192536 94324
rect 191196 4072 191248 4078
rect 191196 4014 191248 4020
rect 191104 3732 191156 3738
rect 191104 3674 191156 3680
rect 192024 3596 192076 3602
rect 192024 3538 192076 3544
rect 190828 3392 190880 3398
rect 190828 3334 190880 3340
rect 190840 480 190868 3334
rect 192036 480 192064 3538
rect 192496 3398 192524 94318
rect 192588 93294 192616 97174
rect 195244 95804 195296 95810
rect 195244 95746 195296 95752
rect 192576 93288 192628 93294
rect 192576 93230 192628 93236
rect 194508 93288 194560 93294
rect 194508 93230 194560 93236
rect 193128 90296 193180 90302
rect 193128 90238 193180 90244
rect 193140 3602 193168 90238
rect 194520 6914 194548 93230
rect 194428 6886 194548 6914
rect 193128 3596 193180 3602
rect 193128 3538 193180 3544
rect 193220 3596 193272 3602
rect 193220 3538 193272 3544
rect 192484 3392 192536 3398
rect 192484 3334 192536 3340
rect 193232 480 193260 3538
rect 194428 480 194456 6886
rect 195256 3602 195284 95746
rect 195900 6914 195928 98534
rect 198648 98524 198700 98530
rect 198648 98466 198700 98472
rect 196622 97608 196678 97617
rect 196622 97543 196678 97552
rect 196636 87718 196664 97543
rect 198004 97096 198056 97102
rect 198004 97038 198056 97044
rect 197268 95736 197320 95742
rect 197268 95678 197320 95684
rect 197176 92948 197228 92954
rect 197176 92890 197228 92896
rect 196624 87712 196676 87718
rect 196624 87654 196676 87660
rect 195624 6886 195928 6914
rect 195244 3596 195296 3602
rect 195244 3538 195296 3544
rect 195624 480 195652 6886
rect 197188 3602 197216 92890
rect 197176 3596 197228 3602
rect 197176 3538 197228 3544
rect 197280 3398 197308 95678
rect 198016 13122 198044 97038
rect 198004 13116 198056 13122
rect 198004 13058 198056 13064
rect 198660 4078 198688 98466
rect 199474 97880 199530 97889
rect 199474 97815 199530 97824
rect 199384 97164 199436 97170
rect 199384 97106 199436 97112
rect 199396 87990 199424 97106
rect 199488 93129 199516 97815
rect 200132 94489 200160 100028
rect 200224 100014 200330 100042
rect 200118 94480 200174 94489
rect 200118 94415 200174 94424
rect 200028 94308 200080 94314
rect 200028 94250 200080 94256
rect 199474 93120 199530 93129
rect 199474 93055 199530 93064
rect 199384 87984 199436 87990
rect 199384 87926 199436 87932
rect 199108 6316 199160 6322
rect 199108 6258 199160 6264
rect 198648 4072 198700 4078
rect 198648 4014 198700 4020
rect 197912 3596 197964 3602
rect 197912 3538 197964 3544
rect 196808 3392 196860 3398
rect 196808 3334 196860 3340
rect 197268 3392 197320 3398
rect 197268 3334 197320 3340
rect 196820 480 196848 3334
rect 197924 480 197952 3538
rect 199120 480 199148 6258
rect 200040 3942 200068 94250
rect 200028 3936 200080 3942
rect 200028 3878 200080 3884
rect 200224 3466 200252 100014
rect 200396 96960 200448 96966
rect 200396 96902 200448 96908
rect 200408 3602 200436 96902
rect 200500 93226 200528 100028
rect 200684 97889 200712 100028
rect 200882 100014 200988 100042
rect 200670 97880 200726 97889
rect 200670 97815 200726 97824
rect 200856 96824 200908 96830
rect 200856 96766 200908 96772
rect 200488 93220 200540 93226
rect 200488 93162 200540 93168
rect 200764 82136 200816 82142
rect 200764 82078 200816 82084
rect 200776 4146 200804 82078
rect 200868 21418 200896 96766
rect 200960 82278 200988 100014
rect 201052 97306 201080 100028
rect 201144 100014 201342 100042
rect 201040 97300 201092 97306
rect 201040 97242 201092 97248
rect 201144 96966 201172 100014
rect 201132 96960 201184 96966
rect 201132 96902 201184 96908
rect 201512 93158 201540 100028
rect 201710 100014 201816 100042
rect 201592 96960 201644 96966
rect 201592 96902 201644 96908
rect 201500 93152 201552 93158
rect 201500 93094 201552 93100
rect 201604 89010 201632 96902
rect 201592 89004 201644 89010
rect 201592 88946 201644 88952
rect 201788 84862 201816 100014
rect 201880 95849 201908 100028
rect 202064 95946 202092 100028
rect 202156 100014 202354 100042
rect 202156 96966 202184 100014
rect 202524 98734 202552 100028
rect 202512 98728 202564 98734
rect 202512 98670 202564 98676
rect 202708 97209 202736 100028
rect 202892 98666 202920 100028
rect 202880 98660 202932 98666
rect 202880 98602 202932 98608
rect 202694 97200 202750 97209
rect 202694 97135 202750 97144
rect 202144 96960 202196 96966
rect 202144 96902 202196 96908
rect 203076 95985 203104 100028
rect 203352 97345 203380 100028
rect 203444 100014 203550 100042
rect 203338 97336 203394 97345
rect 203338 97271 203394 97280
rect 203062 95976 203118 95985
rect 202052 95940 202104 95946
rect 202052 95882 202104 95888
rect 202144 95940 202196 95946
rect 203062 95911 203118 95920
rect 202144 95882 202196 95888
rect 201866 95840 201922 95849
rect 201866 95775 201922 95784
rect 201776 84856 201828 84862
rect 201776 84798 201828 84804
rect 200948 82272 201000 82278
rect 200948 82214 201000 82220
rect 200856 21412 200908 21418
rect 200856 21354 200908 21360
rect 200764 4140 200816 4146
rect 200764 4082 200816 4088
rect 200396 3596 200448 3602
rect 200396 3538 200448 3544
rect 202156 3534 202184 95882
rect 203444 84194 203472 100014
rect 203720 99414 203748 100028
rect 203708 99408 203760 99414
rect 203708 99350 203760 99356
rect 203524 97028 203576 97034
rect 203524 96970 203576 96976
rect 203536 91866 203564 96970
rect 203904 94625 203932 100028
rect 204088 97374 204116 100028
rect 204364 97481 204392 100028
rect 204350 97472 204406 97481
rect 204350 97407 204406 97416
rect 204076 97368 204128 97374
rect 204076 97310 204128 97316
rect 204444 96892 204496 96898
rect 204444 96834 204496 96840
rect 203890 94616 203946 94625
rect 203890 94551 203946 94560
rect 203524 91860 203576 91866
rect 203524 91802 203576 91808
rect 204456 87650 204484 96834
rect 204548 89078 204576 100028
rect 204628 96960 204680 96966
rect 204628 96902 204680 96908
rect 204536 89072 204588 89078
rect 204536 89014 204588 89020
rect 204444 87644 204496 87650
rect 204444 87586 204496 87592
rect 203168 84166 203472 84194
rect 203168 82210 203196 84166
rect 203156 82204 203208 82210
rect 203156 82146 203208 82152
rect 202696 7744 202748 7750
rect 202696 7686 202748 7692
rect 200304 3528 200356 3534
rect 200304 3470 200356 3476
rect 202144 3528 202196 3534
rect 202144 3470 202196 3476
rect 200212 3460 200264 3466
rect 200212 3402 200264 3408
rect 200316 480 200344 3470
rect 201500 2916 201552 2922
rect 201500 2858 201552 2864
rect 201512 480 201540 2858
rect 202708 480 202736 7686
rect 203892 4072 203944 4078
rect 203892 4014 203944 4020
rect 203904 480 203932 4014
rect 204640 3262 204668 96902
rect 204732 83502 204760 100028
rect 204916 97617 204944 100028
rect 205008 100014 205114 100042
rect 205192 100014 205390 100042
rect 204902 97608 204958 97617
rect 204902 97543 204958 97552
rect 204904 97232 204956 97238
rect 204904 97174 204956 97180
rect 204916 96082 204944 97174
rect 205008 96898 205036 100014
rect 205192 96966 205220 100014
rect 205560 97306 205588 100028
rect 205548 97300 205600 97306
rect 205548 97242 205600 97248
rect 205180 96960 205232 96966
rect 205180 96902 205232 96908
rect 204996 96892 205048 96898
rect 204996 96834 205048 96840
rect 204904 96076 204956 96082
rect 204904 96018 204956 96024
rect 205640 94716 205692 94722
rect 205640 94658 205692 94664
rect 205652 94246 205680 94658
rect 205640 94240 205692 94246
rect 205640 94182 205692 94188
rect 205744 91798 205772 100028
rect 205942 100014 206048 100042
rect 205824 94172 205876 94178
rect 205824 94114 205876 94120
rect 205732 91792 205784 91798
rect 205732 91734 205784 91740
rect 205836 87786 205864 94114
rect 205824 87780 205876 87786
rect 205824 87722 205876 87728
rect 204720 83496 204772 83502
rect 204720 83438 204772 83444
rect 206020 11762 206048 100014
rect 206112 97782 206140 100028
rect 206204 100014 206402 100042
rect 206480 100014 206586 100042
rect 206100 97776 206152 97782
rect 206100 97718 206152 97724
rect 206204 89146 206232 100014
rect 206192 89140 206244 89146
rect 206192 89082 206244 89088
rect 206480 84194 206508 100014
rect 206756 97510 206784 100028
rect 206848 100014 206954 100042
rect 207138 100014 207336 100042
rect 206744 97504 206796 97510
rect 206744 97446 206796 97452
rect 206848 94178 206876 100014
rect 206836 94172 206888 94178
rect 206836 94114 206888 94120
rect 206296 84166 206508 84194
rect 206296 15910 206324 84166
rect 206284 15904 206336 15910
rect 206284 15846 206336 15852
rect 206008 11756 206060 11762
rect 206008 11698 206060 11704
rect 207308 3670 207336 100014
rect 207400 96830 207428 100028
rect 207492 100014 207598 100042
rect 207676 100014 207782 100042
rect 207388 96824 207440 96830
rect 207388 96766 207440 96772
rect 207492 90370 207520 100014
rect 207480 90364 207532 90370
rect 207480 90306 207532 90312
rect 207676 84194 207704 100014
rect 207756 97776 207808 97782
rect 207756 97718 207808 97724
rect 207768 97646 207796 97718
rect 207756 97640 207808 97646
rect 207756 97582 207808 97588
rect 207952 97034 207980 100028
rect 207940 97028 207992 97034
rect 207940 96970 207992 96976
rect 208136 94518 208164 100028
rect 208412 99482 208440 100028
rect 208400 99476 208452 99482
rect 208400 99418 208452 99424
rect 208596 94654 208624 100028
rect 208780 98802 208808 100028
rect 208872 100014 208978 100042
rect 208768 98796 208820 98802
rect 208768 98738 208820 98744
rect 208584 94648 208636 94654
rect 208584 94590 208636 94596
rect 208124 94512 208176 94518
rect 208124 94454 208176 94460
rect 208872 88058 208900 100014
rect 209148 94722 209176 100028
rect 209240 100014 209438 100042
rect 209136 94716 209188 94722
rect 209136 94658 209188 94664
rect 209240 93362 209268 100014
rect 209608 97442 209636 100028
rect 209596 97436 209648 97442
rect 209596 97378 209648 97384
rect 209412 97368 209464 97374
rect 209412 97310 209464 97316
rect 209424 96422 209452 97310
rect 209792 96642 209820 100028
rect 209990 100014 210096 100042
rect 209700 96614 209820 96642
rect 209412 96416 209464 96422
rect 209412 96358 209464 96364
rect 209228 93356 209280 93362
rect 209228 93298 209280 93304
rect 209700 90438 209728 96614
rect 209964 94580 210016 94586
rect 209964 94522 210016 94528
rect 209688 90432 209740 90438
rect 209688 90374 209740 90380
rect 209976 89714 210004 94522
rect 210068 93430 210096 100014
rect 210056 93424 210108 93430
rect 210056 93366 210108 93372
rect 210160 93378 210188 100028
rect 210344 94586 210372 100028
rect 210424 97436 210476 97442
rect 210424 97378 210476 97384
rect 210332 94580 210384 94586
rect 210332 94522 210384 94528
rect 210160 93350 210372 93378
rect 210344 89714 210372 93350
rect 209976 89686 210096 89714
rect 208860 88052 208912 88058
rect 208860 87994 208912 88000
rect 209044 87644 209096 87650
rect 209044 87586 209096 87592
rect 207492 84166 207704 84194
rect 207492 83570 207520 84166
rect 207480 83564 207532 83570
rect 207480 83506 207532 83512
rect 207388 3936 207440 3942
rect 207388 3878 207440 3884
rect 207296 3664 207348 3670
rect 207296 3606 207348 3612
rect 205088 3596 205140 3602
rect 205088 3538 205140 3544
rect 204628 3256 204680 3262
rect 204628 3198 204680 3204
rect 205100 480 205128 3538
rect 206192 3460 206244 3466
rect 206192 3402 206244 3408
rect 206204 480 206232 3402
rect 207400 480 207428 3878
rect 208584 3528 208636 3534
rect 208584 3470 208636 3476
rect 208596 480 208624 3470
rect 209056 2922 209084 87586
rect 210068 86562 210096 89686
rect 210160 89686 210372 89714
rect 210160 87854 210188 89686
rect 210148 87848 210200 87854
rect 210148 87790 210200 87796
rect 210056 86556 210108 86562
rect 210056 86498 210108 86504
rect 210436 7682 210464 97378
rect 210516 96688 210568 96694
rect 210516 96630 210568 96636
rect 210528 69698 210556 96630
rect 210620 92002 210648 100028
rect 210804 99686 210832 100028
rect 210792 99680 210844 99686
rect 210792 99622 210844 99628
rect 210988 97102 211016 100028
rect 211172 99550 211200 100028
rect 211370 100014 211476 100042
rect 211160 99544 211212 99550
rect 211160 99486 211212 99492
rect 211448 99374 211476 100014
rect 211448 99346 211568 99374
rect 211160 97300 211212 97306
rect 211160 97242 211212 97248
rect 210976 97096 211028 97102
rect 210976 97038 211028 97044
rect 211172 95742 211200 97242
rect 211160 95736 211212 95742
rect 211160 95678 211212 95684
rect 211436 94580 211488 94586
rect 211436 94522 211488 94528
rect 210608 91996 210660 92002
rect 210608 91938 210660 91944
rect 210516 69692 210568 69698
rect 210516 69634 210568 69640
rect 211448 8974 211476 94522
rect 211540 89714 211568 99346
rect 211632 96694 211660 100028
rect 211620 96688 211672 96694
rect 211620 96630 211672 96636
rect 211816 91934 211844 100028
rect 211908 100014 212014 100042
rect 211908 94586 211936 100014
rect 212184 97170 212212 100028
rect 212276 100014 212382 100042
rect 212658 100014 212764 100042
rect 212172 97164 212224 97170
rect 212172 97106 212224 97112
rect 211896 94580 211948 94586
rect 211896 94522 211948 94528
rect 211804 91928 211856 91934
rect 211804 91870 211856 91876
rect 212276 90506 212304 100014
rect 212540 98048 212592 98054
rect 212540 97990 212592 97996
rect 212552 97170 212580 97990
rect 212540 97164 212592 97170
rect 212540 97106 212592 97112
rect 212264 90500 212316 90506
rect 212264 90442 212316 90448
rect 211540 89686 211752 89714
rect 211724 86290 211752 89686
rect 212736 87922 212764 100014
rect 212828 99958 212856 100028
rect 212816 99952 212868 99958
rect 212816 99894 212868 99900
rect 212908 94580 212960 94586
rect 212908 94522 212960 94528
rect 212724 87916 212776 87922
rect 212724 87858 212776 87864
rect 211712 86284 211764 86290
rect 211712 86226 211764 86232
rect 212920 10334 212948 94522
rect 213012 94246 213040 100028
rect 213104 100014 213210 100042
rect 213000 94240 213052 94246
rect 213000 94182 213052 94188
rect 213104 86358 213132 100014
rect 213380 99754 213408 100028
rect 213472 100014 213670 100042
rect 213748 100014 213854 100042
rect 213368 99748 213420 99754
rect 213368 99690 213420 99696
rect 213184 96076 213236 96082
rect 213184 96018 213236 96024
rect 213092 86352 213144 86358
rect 213092 86294 213144 86300
rect 212908 10328 212960 10334
rect 212908 10270 212960 10276
rect 211436 8968 211488 8974
rect 211436 8910 211488 8916
rect 210424 7676 210476 7682
rect 210424 7618 210476 7624
rect 212172 4956 212224 4962
rect 212172 4898 212224 4904
rect 209780 4072 209832 4078
rect 209780 4014 209832 4020
rect 209044 2916 209096 2922
rect 209044 2858 209096 2864
rect 209792 480 209820 4014
rect 210976 3392 211028 3398
rect 210976 3334 211028 3340
rect 210988 480 211016 3334
rect 212184 480 212212 4898
rect 213196 3398 213224 96018
rect 213472 90574 213500 100014
rect 213748 94586 213776 100014
rect 214024 97986 214052 100028
rect 214208 98870 214236 100028
rect 214300 100014 214406 100042
rect 214484 100014 214682 100042
rect 214760 100014 214866 100042
rect 214944 100014 215050 100042
rect 214196 98864 214248 98870
rect 214196 98806 214248 98812
rect 214012 97980 214064 97986
rect 214012 97922 214064 97928
rect 213736 94580 213788 94586
rect 213736 94522 213788 94528
rect 213460 90568 213512 90574
rect 213460 90510 213512 90516
rect 214300 89714 214328 100014
rect 214484 89714 214512 100014
rect 214564 97028 214616 97034
rect 214564 96970 214616 96976
rect 214116 89686 214328 89714
rect 214392 89686 214512 89714
rect 214116 86426 214144 89686
rect 214104 86420 214156 86426
rect 214104 86362 214156 86368
rect 214392 84194 214420 89686
rect 214300 84166 214420 84194
rect 214300 35222 214328 84166
rect 214288 35216 214340 35222
rect 214288 35158 214340 35164
rect 214576 4894 214604 96970
rect 214760 90642 214788 100014
rect 214748 90636 214800 90642
rect 214748 90578 214800 90584
rect 214944 84930 214972 100014
rect 215220 99890 215248 100028
rect 215208 99884 215260 99890
rect 215208 99826 215260 99832
rect 215404 99618 215432 100028
rect 215496 100014 215694 100042
rect 215772 100014 215878 100042
rect 215956 100014 216062 100042
rect 216140 100014 216246 100042
rect 215392 99612 215444 99618
rect 215392 99554 215444 99560
rect 215496 88126 215524 100014
rect 215772 97016 215800 100014
rect 215588 96988 215800 97016
rect 215484 88120 215536 88126
rect 215484 88062 215536 88068
rect 214932 84924 214984 84930
rect 214932 84866 214984 84872
rect 215588 17270 215616 96988
rect 215956 96914 215984 100014
rect 215772 96886 215984 96914
rect 215772 90710 215800 96886
rect 215944 96756 215996 96762
rect 215944 96698 215996 96704
rect 215760 90704 215812 90710
rect 215760 90646 215812 90652
rect 215576 17264 215628 17270
rect 215576 17206 215628 17212
rect 215956 6186 215984 96698
rect 216140 84998 216168 100014
rect 216416 97578 216444 100028
rect 216404 97572 216456 97578
rect 216404 97514 216456 97520
rect 216692 92070 216720 100028
rect 216772 97572 216824 97578
rect 216772 97514 216824 97520
rect 216784 96558 216812 97514
rect 216876 96830 216904 100028
rect 217060 97034 217088 100028
rect 217152 100014 217258 100042
rect 217442 100014 217548 100042
rect 217048 97028 217100 97034
rect 217048 96970 217100 96976
rect 217152 96914 217180 100014
rect 216968 96886 217180 96914
rect 216864 96824 216916 96830
rect 216864 96766 216916 96772
rect 216772 96552 216824 96558
rect 216772 96494 216824 96500
rect 216680 92064 216732 92070
rect 216680 92006 216732 92012
rect 216968 89214 216996 96886
rect 217140 96824 217192 96830
rect 217140 96766 217192 96772
rect 216956 89208 217008 89214
rect 216956 89150 217008 89156
rect 216128 84992 216180 84998
rect 216128 84934 216180 84940
rect 215944 6180 215996 6186
rect 215944 6122 215996 6128
rect 214564 4888 214616 4894
rect 214564 4830 214616 4836
rect 217152 4826 217180 96766
rect 217520 7614 217548 100014
rect 217704 97918 217732 100028
rect 217796 100014 217902 100042
rect 217980 100026 218086 100042
rect 217968 100020 218086 100026
rect 217692 97912 217744 97918
rect 217692 97854 217744 97860
rect 217796 89282 217824 100014
rect 218020 100014 218086 100020
rect 217968 99962 218020 99968
rect 218060 97640 218112 97646
rect 218060 97582 218112 97588
rect 218072 96286 218100 97582
rect 218152 97504 218204 97510
rect 218152 97446 218204 97452
rect 218060 96280 218112 96286
rect 218060 96222 218112 96228
rect 218164 95878 218192 97446
rect 218256 96762 218284 100028
rect 218440 99822 218468 100028
rect 218532 100014 218730 100042
rect 218428 99816 218480 99822
rect 218428 99758 218480 99764
rect 218336 96960 218388 96966
rect 218336 96902 218388 96908
rect 218244 96756 218296 96762
rect 218244 96698 218296 96704
rect 218152 95872 218204 95878
rect 218152 95814 218204 95820
rect 217784 89276 217836 89282
rect 217784 89218 217836 89224
rect 218348 25566 218376 96902
rect 218532 86494 218560 100014
rect 218900 97782 218928 100028
rect 218992 100014 219098 100042
rect 219176 100014 219282 100042
rect 218888 97776 218940 97782
rect 218888 97718 218940 97724
rect 218992 89350 219020 100014
rect 219176 96966 219204 100014
rect 219164 96960 219216 96966
rect 219164 96902 219216 96908
rect 219452 94790 219480 100028
rect 219624 96892 219676 96898
rect 219624 96834 219676 96840
rect 219440 94784 219492 94790
rect 219440 94726 219492 94732
rect 219636 89418 219664 96834
rect 219728 90778 219756 100028
rect 219808 96960 219860 96966
rect 219808 96902 219860 96908
rect 219716 90772 219768 90778
rect 219716 90714 219768 90720
rect 219624 89412 219676 89418
rect 219624 89354 219676 89360
rect 218980 89344 219032 89350
rect 218980 89286 219032 89292
rect 218520 86488 218572 86494
rect 218520 86430 218572 86436
rect 218336 25560 218388 25566
rect 218336 25502 218388 25508
rect 219820 14482 219848 96902
rect 219912 86630 219940 100028
rect 220096 97850 220124 100028
rect 220188 100014 220294 100042
rect 220372 100014 220478 100042
rect 220084 97844 220136 97850
rect 220084 97786 220136 97792
rect 220188 96898 220216 100014
rect 220372 96966 220400 100014
rect 220648 97714 220676 100028
rect 220938 100014 221044 100042
rect 220636 97708 220688 97714
rect 220636 97650 220688 97656
rect 220636 97096 220688 97102
rect 220636 97038 220688 97044
rect 220360 96960 220412 96966
rect 220360 96902 220412 96908
rect 220176 96892 220228 96898
rect 220176 96834 220228 96840
rect 220648 96354 220676 97038
rect 220636 96348 220688 96354
rect 220636 96290 220688 96296
rect 221016 89486 221044 100014
rect 221004 89480 221056 89486
rect 221004 89422 221056 89428
rect 219900 86624 219952 86630
rect 219900 86566 219952 86572
rect 221108 85066 221136 100028
rect 221292 97442 221320 100028
rect 221280 97436 221332 97442
rect 221280 97378 221332 97384
rect 221476 97238 221504 100028
rect 221568 100014 221674 100042
rect 221752 100014 221950 100042
rect 221464 97232 221516 97238
rect 221464 97174 221516 97180
rect 221568 96948 221596 100014
rect 221200 96920 221596 96948
rect 221096 85060 221148 85066
rect 221096 85002 221148 85008
rect 219808 14476 219860 14482
rect 219808 14418 219860 14424
rect 219348 11756 219400 11762
rect 219348 11698 219400 11704
rect 217968 10328 218020 10334
rect 217968 10270 218020 10276
rect 217508 7608 217560 7614
rect 217508 7550 217560 7556
rect 217140 4820 217192 4826
rect 217140 4762 217192 4768
rect 214472 3936 214524 3942
rect 214472 3878 214524 3884
rect 213368 3664 213420 3670
rect 213368 3606 213420 3612
rect 213184 3392 213236 3398
rect 213184 3334 213236 3340
rect 213380 480 213408 3606
rect 214484 480 214512 3878
rect 215668 3732 215720 3738
rect 215668 3674 215720 3680
rect 215680 480 215708 3674
rect 217980 3398 218008 10270
rect 219256 4140 219308 4146
rect 219256 4082 219308 4088
rect 216864 3392 216916 3398
rect 216864 3334 216916 3340
rect 217968 3392 218020 3398
rect 217968 3334 218020 3340
rect 218060 3392 218112 3398
rect 218060 3334 218112 3340
rect 216876 480 216904 3334
rect 218072 480 218100 3334
rect 219268 480 219296 4082
rect 219360 3398 219388 11698
rect 219348 3392 219400 3398
rect 219348 3334 219400 3340
rect 221200 3262 221228 96920
rect 221752 93498 221780 100014
rect 222120 98938 222148 100028
rect 222304 99142 222332 100028
rect 222292 99136 222344 99142
rect 222292 99078 222344 99084
rect 222108 98932 222160 98938
rect 222108 98874 222160 98880
rect 222384 96892 222436 96898
rect 222384 96834 222436 96840
rect 221740 93492 221792 93498
rect 221740 93434 221792 93440
rect 222396 92138 222424 96834
rect 222384 92132 222436 92138
rect 222384 92074 222436 92080
rect 222488 6254 222516 100028
rect 222672 99006 222700 100028
rect 222764 100014 222962 100042
rect 223040 100014 223146 100042
rect 222660 99000 222712 99006
rect 222660 98942 222712 98948
rect 222568 96960 222620 96966
rect 222568 96902 222620 96908
rect 222580 90846 222608 96902
rect 222764 93566 222792 100014
rect 223040 96966 223068 100014
rect 223028 96960 223080 96966
rect 223028 96902 223080 96908
rect 223316 94858 223344 100028
rect 223408 100014 223514 100042
rect 223698 100014 223804 100042
rect 223408 96898 223436 100014
rect 223580 97028 223632 97034
rect 223580 96970 223632 96976
rect 223396 96892 223448 96898
rect 223396 96834 223448 96840
rect 223592 94994 223620 96970
rect 223580 94988 223632 94994
rect 223580 94930 223632 94936
rect 223304 94852 223356 94858
rect 223304 94794 223356 94800
rect 222752 93560 222804 93566
rect 222752 93502 222804 93508
rect 222844 91792 222896 91798
rect 222844 91734 222896 91740
rect 222568 90840 222620 90846
rect 222568 90782 222620 90788
rect 222476 6248 222528 6254
rect 222476 6190 222528 6196
rect 222856 4078 222884 91734
rect 223776 90914 223804 100014
rect 223868 100014 223974 100042
rect 223764 90908 223816 90914
rect 223764 90850 223816 90856
rect 223488 10396 223540 10402
rect 223488 10338 223540 10344
rect 222844 4072 222896 4078
rect 222844 4014 222896 4020
rect 221556 3800 221608 3806
rect 221556 3742 221608 3748
rect 221188 3256 221240 3262
rect 221188 3198 221240 3204
rect 220452 3188 220504 3194
rect 220452 3130 220504 3136
rect 220464 480 220492 3130
rect 221568 480 221596 3742
rect 223500 2990 223528 10338
rect 223868 3874 223896 100014
rect 224144 93634 224172 100028
rect 224236 100014 224342 100042
rect 224132 93628 224184 93634
rect 224132 93570 224184 93576
rect 224236 84194 224264 100014
rect 224512 99074 224540 100028
rect 224604 100014 224710 100042
rect 224500 99068 224552 99074
rect 224500 99010 224552 99016
rect 224604 92206 224632 100014
rect 224868 97436 224920 97442
rect 224868 97378 224920 97384
rect 224592 92200 224644 92206
rect 224592 92142 224644 92148
rect 224052 84166 224264 84194
rect 224052 18630 224080 84166
rect 224040 18624 224092 18630
rect 224040 18566 224092 18572
rect 223856 3868 223908 3874
rect 223856 3810 223908 3816
rect 222752 2984 222804 2990
rect 222752 2926 222804 2932
rect 223488 2984 223540 2990
rect 223488 2926 223540 2932
rect 222764 480 222792 2926
rect 224880 2922 224908 97378
rect 224972 94926 225000 100028
rect 225156 97034 225184 100028
rect 225340 99210 225368 100028
rect 225328 99204 225380 99210
rect 225328 99146 225380 99152
rect 225144 97028 225196 97034
rect 225144 96970 225196 96976
rect 225236 96960 225288 96966
rect 225236 96902 225288 96908
rect 224960 94920 225012 94926
rect 224960 94862 225012 94868
rect 225248 4010 225276 96902
rect 225420 96892 225472 96898
rect 225420 96834 225472 96840
rect 225432 85134 225460 96834
rect 225524 92274 225552 100028
rect 225616 100014 225722 100042
rect 225616 96966 225644 100014
rect 225604 96960 225656 96966
rect 225604 96902 225656 96908
rect 225984 96150 226012 100028
rect 226076 100014 226182 100042
rect 226076 96898 226104 100014
rect 226064 96892 226116 96898
rect 226064 96834 226116 96840
rect 225972 96144 226024 96150
rect 225972 96086 226024 96092
rect 226352 95062 226380 100028
rect 226550 100014 226656 100042
rect 226628 96966 226656 100014
rect 226616 96960 226668 96966
rect 226616 96902 226668 96908
rect 226340 95056 226392 95062
rect 226340 94998 226392 95004
rect 225512 92268 225564 92274
rect 225512 92210 225564 92216
rect 225420 85128 225472 85134
rect 225420 85070 225472 85076
rect 226720 71058 226748 100028
rect 226892 96960 226944 96966
rect 226892 96902 226944 96908
rect 226800 96892 226852 96898
rect 226800 96834 226852 96840
rect 226812 82142 226840 96834
rect 226904 92342 226932 96902
rect 226996 95130 227024 100028
rect 227088 100014 227194 100042
rect 226984 95124 227036 95130
rect 226984 95066 227036 95072
rect 226984 94512 227036 94518
rect 226984 94454 227036 94460
rect 226892 92336 226944 92342
rect 226892 92278 226944 92284
rect 226800 82136 226852 82142
rect 226800 82078 226852 82084
rect 226708 71052 226760 71058
rect 226708 70994 226760 71000
rect 225236 4004 225288 4010
rect 225236 3946 225288 3952
rect 225328 4004 225380 4010
rect 225328 3946 225380 3952
rect 225144 3868 225196 3874
rect 225144 3810 225196 3816
rect 223948 2916 224000 2922
rect 223948 2858 224000 2864
rect 224868 2916 224920 2922
rect 224868 2858 224920 2864
rect 223960 480 223988 2858
rect 225156 480 225184 3810
rect 225340 3602 225368 3946
rect 225328 3596 225380 3602
rect 225328 3538 225380 3544
rect 226340 3596 226392 3602
rect 226340 3538 226392 3544
rect 226352 480 226380 3538
rect 226996 3194 227024 94454
rect 227088 92410 227116 100014
rect 227364 97374 227392 100028
rect 227456 100014 227562 100042
rect 227352 97368 227404 97374
rect 227352 97310 227404 97316
rect 227456 96898 227484 100014
rect 227444 96892 227496 96898
rect 227444 96834 227496 96840
rect 227732 95198 227760 100028
rect 227904 96892 227956 96898
rect 227904 96834 227956 96840
rect 227720 95192 227772 95198
rect 227720 95134 227772 95140
rect 227916 93770 227944 96834
rect 227904 93764 227956 93770
rect 227904 93706 227956 93712
rect 228008 92478 228036 100028
rect 228192 97646 228220 100028
rect 228284 100014 228390 100042
rect 228468 100014 228574 100042
rect 228180 97640 228232 97646
rect 228180 97582 228232 97588
rect 228088 96960 228140 96966
rect 228088 96902 228140 96908
rect 227996 92472 228048 92478
rect 227996 92414 228048 92420
rect 227076 92404 227128 92410
rect 227076 92346 227128 92352
rect 228100 90982 228128 96902
rect 228284 93702 228312 100014
rect 228468 96966 228496 100014
rect 228548 97368 228600 97374
rect 228548 97310 228600 97316
rect 228456 96960 228508 96966
rect 228456 96902 228508 96908
rect 228364 94580 228416 94586
rect 228364 94522 228416 94528
rect 228272 93696 228324 93702
rect 228272 93638 228324 93644
rect 228088 90976 228140 90982
rect 228088 90918 228140 90924
rect 227628 15904 227680 15910
rect 227628 15846 227680 15852
rect 227536 8968 227588 8974
rect 227536 8910 227588 8916
rect 226984 3188 227036 3194
rect 226984 3130 227036 3136
rect 227548 480 227576 8910
rect 227640 3602 227668 15846
rect 228376 4010 228404 94522
rect 228456 93152 228508 93158
rect 228456 93094 228508 93100
rect 228468 4146 228496 93094
rect 228560 10334 228588 97310
rect 228744 97102 228772 100028
rect 228836 100014 229034 100042
rect 228732 97096 228784 97102
rect 228732 97038 228784 97044
rect 228836 96898 228864 100014
rect 228824 96892 228876 96898
rect 228824 96834 228876 96840
rect 229204 91730 229232 100028
rect 229388 96218 229416 100028
rect 229572 99278 229600 100028
rect 229664 100014 229770 100042
rect 229560 99272 229612 99278
rect 229560 99214 229612 99220
rect 229468 96960 229520 96966
rect 229468 96902 229520 96908
rect 229376 96212 229428 96218
rect 229376 96154 229428 96160
rect 229192 91724 229244 91730
rect 229192 91666 229244 91672
rect 229480 19990 229508 96902
rect 229664 93838 229692 100014
rect 230032 97578 230060 100028
rect 230020 97572 230072 97578
rect 230020 97514 230072 97520
rect 229744 96824 229796 96830
rect 229744 96766 229796 96772
rect 229652 93832 229704 93838
rect 229652 93774 229704 93780
rect 229468 19984 229520 19990
rect 229468 19926 229520 19932
rect 228548 10328 228600 10334
rect 228548 10270 228600 10276
rect 229756 6322 229784 96766
rect 230216 94450 230244 100028
rect 230308 100014 230414 100042
rect 230308 96966 230336 100014
rect 230584 97510 230612 100028
rect 230768 99346 230796 100028
rect 230756 99340 230808 99346
rect 230756 99282 230808 99288
rect 230572 97504 230624 97510
rect 230572 97446 230624 97452
rect 230296 96960 230348 96966
rect 230296 96902 230348 96908
rect 230848 96960 230900 96966
rect 230848 96902 230900 96908
rect 230204 94444 230256 94450
rect 230204 94386 230256 94392
rect 230860 91050 230888 96902
rect 230952 91662 230980 100028
rect 231032 96892 231084 96898
rect 231032 96834 231084 96840
rect 231044 93090 231072 96834
rect 231124 96756 231176 96762
rect 231124 96698 231176 96704
rect 231032 93084 231084 93090
rect 231032 93026 231084 93032
rect 230940 91656 230992 91662
rect 230940 91598 230992 91604
rect 230848 91044 230900 91050
rect 230848 90986 230900 90992
rect 229836 7472 229888 7478
rect 229836 7414 229888 7420
rect 229744 6316 229796 6322
rect 229744 6258 229796 6264
rect 228456 4140 228508 4146
rect 228456 4082 228508 4088
rect 228364 4004 228416 4010
rect 228364 3946 228416 3952
rect 228732 4004 228784 4010
rect 228732 3946 228784 3952
rect 227628 3596 227680 3602
rect 227628 3538 227680 3544
rect 228744 480 228772 3946
rect 229848 480 229876 7414
rect 231136 4962 231164 96698
rect 231228 96014 231256 100028
rect 231320 100014 231426 100042
rect 231504 100014 231610 100042
rect 231320 96898 231348 100014
rect 231504 96966 231532 100014
rect 231492 96960 231544 96966
rect 231492 96902 231544 96908
rect 231308 96892 231360 96898
rect 231308 96834 231360 96840
rect 231780 96490 231808 100028
rect 231768 96484 231820 96490
rect 231768 96426 231820 96432
rect 231216 96008 231268 96014
rect 231216 95950 231268 95956
rect 231216 95872 231268 95878
rect 231216 95814 231268 95820
rect 231124 4956 231176 4962
rect 231124 4898 231176 4904
rect 231228 3942 231256 95814
rect 231964 93022 231992 100028
rect 232240 97170 232268 100028
rect 232332 100014 232438 100042
rect 232228 97164 232280 97170
rect 232228 97106 232280 97112
rect 232332 97050 232360 100014
rect 232056 97022 232360 97050
rect 232056 96626 232084 97022
rect 232044 96620 232096 96626
rect 232044 96562 232096 96568
rect 232608 94382 232636 100028
rect 232700 100014 232806 100042
rect 232596 94376 232648 94382
rect 232596 94318 232648 94324
rect 232700 94194 232728 100014
rect 232780 97096 232832 97102
rect 232780 97038 232832 97044
rect 232148 94166 232728 94194
rect 231952 93016 232004 93022
rect 231952 92958 232004 92964
rect 231308 91112 231360 91118
rect 231308 91054 231360 91060
rect 231216 3936 231268 3942
rect 231216 3878 231268 3884
rect 231320 3670 231348 91054
rect 232148 90302 232176 94166
rect 232136 90296 232188 90302
rect 232136 90238 232188 90244
rect 232792 84194 232820 97038
rect 232976 95810 233004 100028
rect 233266 100014 233372 100042
rect 233344 96898 233372 100014
rect 233436 98598 233464 100028
rect 233424 98592 233476 98598
rect 233424 98534 233476 98540
rect 233620 97306 233648 100028
rect 233712 100014 233818 100042
rect 233608 97300 233660 97306
rect 233608 97242 233660 97248
rect 233516 97028 233568 97034
rect 233516 96970 233568 96976
rect 233332 96892 233384 96898
rect 233332 96834 233384 96840
rect 232964 95804 233016 95810
rect 232964 95746 233016 95752
rect 233148 95328 233200 95334
rect 233148 95270 233200 95276
rect 232516 84166 232820 84194
rect 232516 15910 232544 84166
rect 232596 17944 232648 17950
rect 232596 17886 232648 17892
rect 232504 15904 232556 15910
rect 232504 15846 232556 15852
rect 232608 3738 232636 17886
rect 232596 3732 232648 3738
rect 232596 3674 232648 3680
rect 231308 3664 231360 3670
rect 231308 3606 231360 3612
rect 233160 3534 233188 95270
rect 233528 87650 233556 96970
rect 233712 92954 233740 100014
rect 233884 96960 233936 96966
rect 233884 96902 233936 96908
rect 233700 92948 233752 92954
rect 233700 92890 233752 92896
rect 233516 87644 233568 87650
rect 233516 87586 233568 87592
rect 233424 8424 233476 8430
rect 233424 8366 233476 8372
rect 232228 3528 232280 3534
rect 232228 3470 232280 3476
rect 233148 3528 233200 3534
rect 233148 3470 233200 3476
rect 231032 3120 231084 3126
rect 231032 3062 231084 3068
rect 231044 480 231072 3062
rect 232240 480 232268 3470
rect 233436 480 233464 8366
rect 233896 7750 233924 96902
rect 233988 96830 234016 100028
rect 234068 96892 234120 96898
rect 234068 96834 234120 96840
rect 233976 96824 234028 96830
rect 233976 96766 234028 96772
rect 233976 96688 234028 96694
rect 233976 96630 234028 96636
rect 233988 10402 234016 96630
rect 234080 93294 234108 96834
rect 234264 95946 234292 100028
rect 234356 100014 234462 100042
rect 234356 97034 234384 100014
rect 234344 97028 234396 97034
rect 234344 96970 234396 96976
rect 234632 96966 234660 100028
rect 234816 98530 234844 100028
rect 234908 100014 235014 100042
rect 235092 100014 235290 100042
rect 235368 100014 235474 100042
rect 235552 100014 235658 100042
rect 235736 100014 235842 100042
rect 234804 98524 234856 98530
rect 234804 98466 234856 98472
rect 234908 97050 234936 100014
rect 234816 97022 234936 97050
rect 234620 96960 234672 96966
rect 234620 96902 234672 96908
rect 234252 95940 234304 95946
rect 234252 95882 234304 95888
rect 234816 94586 234844 97022
rect 235092 96914 235120 100014
rect 234908 96886 235120 96914
rect 234804 94580 234856 94586
rect 234804 94522 234856 94528
rect 234068 93288 234120 93294
rect 234068 93230 234120 93236
rect 234528 92540 234580 92546
rect 234528 92482 234580 92488
rect 234068 13864 234120 13870
rect 234068 13806 234120 13812
rect 233976 10396 234028 10402
rect 233976 10338 234028 10344
rect 233884 7744 233936 7750
rect 233884 7686 233936 7692
rect 234080 3602 234108 13806
rect 234160 9920 234212 9926
rect 234160 9862 234212 9868
rect 234172 3806 234200 9862
rect 234160 3800 234212 3806
rect 234160 3742 234212 3748
rect 234068 3596 234120 3602
rect 234068 3538 234120 3544
rect 234540 3482 234568 92482
rect 234804 9648 234856 9654
rect 234804 9590 234856 9596
rect 234816 3874 234844 9590
rect 234804 3868 234856 3874
rect 234804 3810 234856 3816
rect 234540 3454 234660 3482
rect 234908 3466 234936 96886
rect 235080 96824 235132 96830
rect 235080 96766 235132 96772
rect 235092 13870 235120 96766
rect 235368 95690 235396 100014
rect 235552 96830 235580 100014
rect 235632 97232 235684 97238
rect 235632 97174 235684 97180
rect 235540 96824 235592 96830
rect 235540 96766 235592 96772
rect 235184 95662 235396 95690
rect 235184 94314 235212 95662
rect 235644 95554 235672 97174
rect 235276 95526 235672 95554
rect 235172 94308 235224 94314
rect 235172 94250 235224 94256
rect 235080 13864 235132 13870
rect 235080 13806 235132 13812
rect 235276 7478 235304 95526
rect 235356 95464 235408 95470
rect 235356 95406 235408 95412
rect 235368 8974 235396 95406
rect 235736 91798 235764 100014
rect 235816 97504 235868 97510
rect 235816 97446 235868 97452
rect 235828 95470 235856 97446
rect 236012 96082 236040 100028
rect 236104 100014 236302 100042
rect 236380 100014 236486 100042
rect 236104 96762 236132 100014
rect 236380 96914 236408 100014
rect 236196 96886 236408 96914
rect 236092 96756 236144 96762
rect 236092 96698 236144 96704
rect 236000 96076 236052 96082
rect 236000 96018 236052 96024
rect 235816 95464 235868 95470
rect 235816 95406 235868 95412
rect 235908 93900 235960 93906
rect 235908 93842 235960 93848
rect 235724 91792 235776 91798
rect 235724 91734 235776 91740
rect 235356 8968 235408 8974
rect 235356 8910 235408 8916
rect 235264 7472 235316 7478
rect 235264 7414 235316 7420
rect 235920 6914 235948 93842
rect 236196 91118 236224 96886
rect 236368 96824 236420 96830
rect 236368 96766 236420 96772
rect 236184 91112 236236 91118
rect 236184 91054 236236 91060
rect 236380 11762 236408 96766
rect 236656 95878 236684 100028
rect 236748 100014 236854 100042
rect 236644 95872 236696 95878
rect 236644 95814 236696 95820
rect 236748 17950 236776 100014
rect 237024 97374 237052 100028
rect 237116 100014 237314 100042
rect 237498 100014 237604 100042
rect 237012 97368 237064 97374
rect 237012 97310 237064 97316
rect 237116 96830 237144 100014
rect 237380 96892 237432 96898
rect 237380 96834 237432 96840
rect 237104 96824 237156 96830
rect 237104 96766 237156 96772
rect 237392 95316 237420 96834
rect 237300 95288 237420 95316
rect 236736 17944 236788 17950
rect 236736 17886 236788 17892
rect 236644 15224 236696 15230
rect 236644 15166 236696 15172
rect 236368 11756 236420 11762
rect 236368 11698 236420 11704
rect 235828 6886 235948 6914
rect 234632 480 234660 3454
rect 234896 3460 234948 3466
rect 234896 3402 234948 3408
rect 235828 480 235856 6886
rect 236656 4010 236684 15166
rect 237300 6914 237328 95288
rect 237576 94586 237604 100014
rect 237564 94580 237616 94586
rect 237564 94522 237616 94528
rect 237668 94518 237696 100028
rect 237760 100014 237866 100042
rect 238050 100014 238156 100042
rect 237760 96778 237788 100014
rect 238024 97776 238076 97782
rect 238024 97718 238076 97724
rect 237760 96750 237880 96778
rect 237748 96008 237800 96014
rect 237748 95950 237800 95956
rect 237656 94512 237708 94518
rect 237656 94454 237708 94460
rect 237760 9654 237788 95950
rect 237852 9926 237880 96750
rect 237932 94580 237984 94586
rect 237932 94522 237984 94528
rect 237944 93158 237972 94522
rect 237932 93152 237984 93158
rect 237932 93094 237984 93100
rect 237840 9920 237892 9926
rect 237840 9862 237892 9868
rect 237748 9648 237800 9654
rect 237748 9590 237800 9596
rect 237024 6886 237328 6914
rect 236644 4004 236696 4010
rect 236644 3946 236696 3952
rect 237024 480 237052 6886
rect 238036 3126 238064 97718
rect 238128 96694 238156 100014
rect 238312 97442 238340 100028
rect 238404 100014 238510 100042
rect 238300 97436 238352 97442
rect 238300 97378 238352 97384
rect 238116 96688 238168 96694
rect 238116 96630 238168 96636
rect 238404 96014 238432 100014
rect 238680 97102 238708 100028
rect 238864 97510 238892 100028
rect 238852 97504 238904 97510
rect 238852 97446 238904 97452
rect 238668 97096 238720 97102
rect 238668 97038 238720 97044
rect 238392 96008 238444 96014
rect 238392 95950 238444 95956
rect 238668 93152 238720 93158
rect 238668 93094 238720 93100
rect 238680 3534 238708 93094
rect 239048 15230 239076 100028
rect 239324 97238 239352 100028
rect 239508 97782 239536 100028
rect 239496 97776 239548 97782
rect 239496 97718 239548 97724
rect 239312 97232 239364 97238
rect 239312 97174 239364 97180
rect 239692 95334 239720 100028
rect 239784 100014 239890 100042
rect 239968 100014 240074 100042
rect 239680 95328 239732 95334
rect 239680 95270 239732 95276
rect 239784 95146 239812 100014
rect 239140 95118 239812 95146
rect 239036 15224 239088 15230
rect 239036 15166 239088 15172
rect 239140 8430 239168 95118
rect 239968 92546 239996 100014
rect 240140 96960 240192 96966
rect 240140 96902 240192 96908
rect 239956 92540 240008 92546
rect 239956 92482 240008 92488
rect 239128 8424 239180 8430
rect 239128 8366 239180 8372
rect 238668 3528 238720 3534
rect 238668 3470 238720 3476
rect 238116 3460 238168 3466
rect 238116 3402 238168 3408
rect 238024 3120 238076 3126
rect 238024 3062 238076 3068
rect 238128 480 238156 3402
rect 239312 3120 239364 3126
rect 239312 3062 239364 3068
rect 239324 480 239352 3062
rect 240152 490 240180 96902
rect 240244 93906 240272 100028
rect 240520 96898 240548 100028
rect 240508 96892 240560 96898
rect 240508 96834 240560 96840
rect 240704 94654 240732 100028
rect 240796 100014 240902 100042
rect 240692 94648 240744 94654
rect 240692 94590 240744 94596
rect 240232 93900 240284 93906
rect 240232 93842 240284 93848
rect 240796 84194 240824 100014
rect 241072 96966 241100 100028
rect 241270 100014 241376 100042
rect 241060 96960 241112 96966
rect 241060 96902 241112 96908
rect 240612 84166 240824 84194
rect 240612 3126 240640 84166
rect 241348 5574 241376 100014
rect 241532 96914 241560 100028
rect 241440 96886 241560 96914
rect 241336 5568 241388 5574
rect 241336 5510 241388 5516
rect 241440 4214 241468 96886
rect 241716 93158 241744 100028
rect 241900 96966 241928 100028
rect 242084 97034 242112 100028
rect 242072 97028 242124 97034
rect 242072 96970 242124 96976
rect 241888 96960 241940 96966
rect 241888 96902 241940 96908
rect 242268 96898 242296 100028
rect 242440 96960 242492 96966
rect 242440 96902 242492 96908
rect 242256 96892 242308 96898
rect 242256 96834 242308 96840
rect 241704 93152 241756 93158
rect 241704 93094 241756 93100
rect 242452 89078 242480 96902
rect 242440 89072 242492 89078
rect 242440 89014 242492 89020
rect 242544 37942 242572 100028
rect 242728 97374 242756 100028
rect 242716 97368 242768 97374
rect 242716 97310 242768 97316
rect 242912 97102 242940 100028
rect 242900 97096 242952 97102
rect 242900 97038 242952 97044
rect 242808 97028 242860 97034
rect 242808 96970 242860 96976
rect 242624 96960 242676 96966
rect 242624 96902 242676 96908
rect 242532 37936 242584 37942
rect 242532 37878 242584 37884
rect 242636 11762 242664 96902
rect 242716 96892 242768 96898
rect 242716 96834 242768 96840
rect 242624 11756 242676 11762
rect 242624 11698 242676 11704
rect 242728 8294 242756 96834
rect 242716 8288 242768 8294
rect 242716 8230 242768 8236
rect 242820 5574 242848 96970
rect 243096 96898 243124 100028
rect 243280 96966 243308 100028
rect 243556 97170 243584 100028
rect 243754 100014 243860 100042
rect 243544 97164 243596 97170
rect 243544 97106 243596 97112
rect 243268 96960 243320 96966
rect 243268 96902 243320 96908
rect 243084 96892 243136 96898
rect 243084 96834 243136 96840
rect 243832 93854 243860 100014
rect 243924 96082 243952 100028
rect 244016 100014 244122 100042
rect 243912 96076 243964 96082
rect 243912 96018 243964 96024
rect 243832 93826 243952 93854
rect 243924 18698 243952 93826
rect 244016 91866 244044 100014
rect 244292 96966 244320 100028
rect 244280 96960 244332 96966
rect 244280 96902 244332 96908
rect 244096 96892 244148 96898
rect 244096 96834 244148 96840
rect 244004 91860 244056 91866
rect 244004 91802 244056 91808
rect 244108 86426 244136 96834
rect 244568 96830 244596 100028
rect 244752 96898 244780 100028
rect 244950 100014 245056 100042
rect 245134 100014 245240 100042
rect 245318 100014 245516 100042
rect 245028 96914 245056 100014
rect 245212 97050 245240 100014
rect 245212 97022 245424 97050
rect 245292 96960 245344 96966
rect 244740 96892 244792 96898
rect 245028 96886 245240 96914
rect 245292 96902 245344 96908
rect 244740 96834 244792 96840
rect 244556 96824 244608 96830
rect 244556 96766 244608 96772
rect 245108 96824 245160 96830
rect 245108 96766 245160 96772
rect 244096 86420 244148 86426
rect 244096 86362 244148 86368
rect 243912 18692 243964 18698
rect 243912 18634 243964 18640
rect 245120 14550 245148 96766
rect 245108 14544 245160 14550
rect 245108 14486 245160 14492
rect 241704 5568 241756 5574
rect 241704 5510 241756 5516
rect 242808 5568 242860 5574
rect 242808 5510 242860 5516
rect 241428 4208 241480 4214
rect 241428 4150 241480 4156
rect 240600 3120 240652 3126
rect 240600 3062 240652 3068
rect 240336 598 240548 626
rect 240336 490 240364 598
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240152 462 240364 490
rect 240520 480 240548 598
rect 241716 480 241744 5510
rect 245212 5506 245240 96886
rect 245304 84930 245332 96902
rect 245292 84924 245344 84930
rect 245292 84866 245344 84872
rect 245396 18630 245424 97022
rect 245488 93158 245516 100014
rect 245580 97714 245608 100028
rect 245568 97708 245620 97714
rect 245568 97650 245620 97656
rect 245568 96892 245620 96898
rect 245568 96834 245620 96840
rect 245476 93152 245528 93158
rect 245476 93094 245528 93100
rect 245580 91798 245608 96834
rect 245764 96762 245792 100028
rect 245752 96756 245804 96762
rect 245752 96698 245804 96704
rect 245948 96694 245976 100028
rect 246146 100014 246252 100042
rect 245936 96688 245988 96694
rect 245936 96630 245988 96636
rect 245568 91792 245620 91798
rect 245568 91734 245620 91740
rect 246224 90438 246252 100014
rect 246316 96014 246344 100028
rect 246500 100014 246606 100042
rect 246684 100014 246790 100042
rect 246868 100014 246974 100042
rect 246304 96008 246356 96014
rect 246304 95950 246356 95956
rect 246212 90432 246264 90438
rect 246212 90374 246264 90380
rect 245384 18624 245436 18630
rect 245384 18566 245436 18572
rect 245660 8288 245712 8294
rect 245660 8230 245712 8236
rect 245200 5500 245252 5506
rect 245200 5442 245252 5448
rect 242900 4208 242952 4214
rect 242900 4150 242952 4156
rect 242912 480 242940 4150
rect 245200 3800 245252 3806
rect 245200 3742 245252 3748
rect 244096 3528 244148 3534
rect 244096 3470 244148 3476
rect 244108 480 244136 3470
rect 245212 480 245240 3742
rect 245672 2990 245700 8230
rect 246396 5568 246448 5574
rect 246396 5510 246448 5516
rect 245660 2984 245712 2990
rect 245660 2926 245712 2932
rect 246408 480 246436 5510
rect 246500 3534 246528 100014
rect 246684 96914 246712 100014
rect 246592 96886 246712 96914
rect 246592 83502 246620 96886
rect 246868 96812 246896 100014
rect 247144 96898 247172 100028
rect 247328 97578 247356 100028
rect 247316 97572 247368 97578
rect 247316 97514 247368 97520
rect 247604 97306 247632 100028
rect 247592 97300 247644 97306
rect 247592 97242 247644 97248
rect 247788 96966 247816 100028
rect 247986 100014 248092 100042
rect 247960 97028 248012 97034
rect 247960 96970 248012 96976
rect 247776 96960 247828 96966
rect 247776 96902 247828 96908
rect 247132 96892 247184 96898
rect 247132 96834 247184 96840
rect 246684 96784 246896 96812
rect 246580 83496 246632 83502
rect 246580 83438 246632 83444
rect 246684 82210 246712 96784
rect 246764 96688 246816 96694
rect 246764 96630 246816 96636
rect 246856 96688 246908 96694
rect 246856 96630 246908 96636
rect 246672 82204 246724 82210
rect 246672 82146 246724 82152
rect 246776 18766 246804 96630
rect 246764 18760 246816 18766
rect 246764 18702 246816 18708
rect 246868 14482 246896 96630
rect 247972 95946 248000 96970
rect 247960 95940 248012 95946
rect 247960 95882 248012 95888
rect 248064 31074 248092 100014
rect 248156 97034 248184 100028
rect 248340 97034 248368 100028
rect 248144 97028 248196 97034
rect 248144 96970 248196 96976
rect 248328 97028 248380 97034
rect 248328 96970 248380 96976
rect 248236 96960 248288 96966
rect 248236 96902 248288 96908
rect 248144 96892 248196 96898
rect 248144 96834 248196 96840
rect 248156 90370 248184 96834
rect 248144 90364 248196 90370
rect 248144 90306 248196 90312
rect 248248 87650 248276 96902
rect 248616 96830 248644 100028
rect 248604 96824 248656 96830
rect 248604 96766 248656 96772
rect 248800 94518 248828 100028
rect 248984 96966 249012 100028
rect 249182 100014 249288 100042
rect 249366 100014 249564 100042
rect 249064 97164 249116 97170
rect 249064 97106 249116 97112
rect 248972 96960 249024 96966
rect 248972 96902 249024 96908
rect 248788 94512 248840 94518
rect 248788 94454 248840 94460
rect 248236 87644 248288 87650
rect 248236 87586 248288 87592
rect 248420 37936 248472 37942
rect 248420 37878 248472 37884
rect 248052 31068 248104 31074
rect 248052 31010 248104 31016
rect 246856 14476 246908 14482
rect 246856 14418 246908 14424
rect 246488 3528 246540 3534
rect 246488 3470 246540 3476
rect 247592 2984 247644 2990
rect 247592 2926 247644 2932
rect 247604 480 247632 2926
rect 248432 490 248460 37878
rect 249076 17882 249104 97106
rect 249064 17876 249116 17882
rect 249064 17818 249116 17824
rect 249260 6186 249288 100014
rect 249340 96960 249392 96966
rect 249340 96902 249392 96908
rect 249432 96960 249484 96966
rect 249432 96902 249484 96908
rect 249352 89010 249380 96902
rect 249340 89004 249392 89010
rect 249340 88946 249392 88952
rect 249444 86358 249472 96902
rect 249432 86352 249484 86358
rect 249432 86294 249484 86300
rect 249536 82142 249564 100014
rect 249628 96966 249656 100028
rect 249812 97442 249840 100028
rect 249800 97436 249852 97442
rect 249800 97378 249852 97384
rect 249996 96966 250024 100028
rect 249616 96960 249668 96966
rect 249616 96902 249668 96908
rect 249984 96960 250036 96966
rect 249984 96902 250036 96908
rect 249616 96824 249668 96830
rect 249616 96766 249668 96772
rect 249524 82136 249576 82142
rect 249524 82078 249576 82084
rect 249628 39370 249656 96766
rect 250180 96762 250208 100028
rect 250364 97170 250392 100028
rect 250352 97164 250404 97170
rect 250352 97106 250404 97112
rect 250444 97096 250496 97102
rect 250444 97038 250496 97044
rect 250168 96756 250220 96762
rect 250168 96698 250220 96704
rect 249616 39364 249668 39370
rect 249616 39306 249668 39312
rect 250456 17950 250484 97038
rect 250548 95810 250576 100028
rect 250732 100014 250838 100042
rect 250536 95804 250588 95810
rect 250536 95746 250588 95752
rect 250444 17944 250496 17950
rect 250444 17886 250496 17892
rect 249248 6180 249300 6186
rect 249248 6122 249300 6128
rect 250732 5030 250760 100014
rect 250812 96960 250864 96966
rect 250812 96902 250864 96908
rect 250824 90030 250852 96902
rect 250904 96756 250956 96762
rect 250904 96698 250956 96704
rect 250812 90024 250864 90030
rect 250812 89966 250864 89972
rect 250916 86290 250944 96698
rect 250904 86284 250956 86290
rect 250904 86226 250956 86232
rect 251008 75206 251036 100028
rect 251192 96626 251220 100028
rect 251376 96898 251404 100028
rect 251364 96892 251416 96898
rect 251364 96834 251416 96840
rect 251560 96830 251588 100028
rect 251548 96824 251600 96830
rect 251548 96766 251600 96772
rect 251180 96620 251232 96626
rect 251180 96562 251232 96568
rect 251836 95878 251864 100028
rect 252020 96966 252048 100028
rect 252112 100014 252218 100042
rect 252008 96960 252060 96966
rect 252008 96902 252060 96908
rect 251824 95872 251876 95878
rect 251824 95814 251876 95820
rect 251272 94648 251324 94654
rect 251272 94590 251324 94596
rect 250996 75200 251048 75206
rect 250996 75142 251048 75148
rect 251180 17944 251232 17950
rect 251180 17886 251232 17892
rect 251088 5500 251140 5506
rect 251088 5442 251140 5448
rect 250720 5024 250772 5030
rect 250720 4966 250772 4972
rect 251100 3738 251128 5442
rect 251088 3732 251140 3738
rect 251088 3674 251140 3680
rect 249984 3664 250036 3670
rect 249984 3606 250036 3612
rect 248616 598 248828 626
rect 248616 490 248644 598
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248432 462 248644 490
rect 248800 480 248828 598
rect 249996 480 250024 3606
rect 251192 480 251220 17886
rect 251284 3466 251312 94590
rect 252112 3602 252140 100014
rect 252388 97646 252416 100028
rect 252376 97640 252428 97646
rect 252376 97582 252428 97588
rect 252192 96960 252244 96966
rect 252192 96902 252244 96908
rect 252204 92274 252232 96902
rect 252284 96892 252336 96898
rect 252284 96834 252336 96840
rect 252192 92268 252244 92274
rect 252192 92210 252244 92216
rect 252296 84862 252324 96834
rect 252572 96830 252600 100028
rect 252848 96898 252876 100028
rect 253032 99210 253060 100028
rect 253020 99204 253072 99210
rect 253020 99146 253072 99152
rect 253216 96966 253244 100028
rect 253414 100014 253520 100042
rect 253296 97708 253348 97714
rect 253296 97650 253348 97656
rect 253204 96960 253256 96966
rect 253204 96902 253256 96908
rect 252836 96892 252888 96898
rect 252836 96834 252888 96840
rect 252376 96824 252428 96830
rect 252376 96766 252428 96772
rect 252560 96824 252612 96830
rect 252560 96766 252612 96772
rect 252284 84856 252336 84862
rect 252284 84798 252336 84804
rect 252388 22778 252416 96766
rect 253308 90506 253336 97650
rect 253296 90500 253348 90506
rect 253296 90442 253348 90448
rect 253204 90024 253256 90030
rect 253204 89966 253256 89972
rect 252652 89072 252704 89078
rect 252652 89014 252704 89020
rect 252376 22772 252428 22778
rect 252376 22714 252428 22720
rect 252560 11756 252612 11762
rect 252560 11698 252612 11704
rect 252100 3596 252152 3602
rect 252100 3538 252152 3544
rect 252572 3482 252600 11698
rect 252664 3806 252692 89014
rect 253216 3806 253244 89966
rect 253492 24138 253520 100014
rect 253584 99142 253612 100028
rect 253768 100014 253874 100042
rect 253572 99136 253624 99142
rect 253572 99078 253624 99084
rect 253664 96960 253716 96966
rect 253664 96902 253716 96908
rect 253572 96892 253624 96898
rect 253572 96834 253624 96840
rect 253584 90234 253612 96834
rect 253572 90228 253624 90234
rect 253572 90170 253624 90176
rect 253676 88942 253704 96902
rect 253664 88936 253716 88942
rect 253664 88878 253716 88884
rect 253768 87514 253796 100014
rect 254044 96830 254072 100028
rect 254228 96966 254256 100028
rect 254216 96960 254268 96966
rect 254216 96902 254268 96908
rect 253848 96824 253900 96830
rect 253848 96766 253900 96772
rect 254032 96824 254084 96830
rect 254032 96766 254084 96772
rect 253860 92954 253888 96766
rect 254412 94450 254440 100028
rect 254610 100014 254808 100042
rect 254886 100014 254992 100042
rect 255070 100014 255176 100042
rect 254780 97050 254808 100014
rect 254964 98394 254992 100014
rect 254952 98388 255004 98394
rect 254952 98330 255004 98336
rect 254780 97022 255084 97050
rect 254860 96960 254912 96966
rect 254860 96902 254912 96908
rect 254768 96892 254820 96898
rect 254768 96834 254820 96840
rect 254400 94444 254452 94450
rect 254400 94386 254452 94392
rect 253848 92948 253900 92954
rect 253848 92890 253900 92896
rect 253756 87508 253808 87514
rect 253756 87450 253808 87456
rect 253480 24132 253532 24138
rect 253480 24074 253532 24080
rect 253940 17876 253992 17882
rect 253940 17818 253992 17824
rect 253952 16574 253980 17818
rect 254780 17270 254808 96834
rect 254768 17264 254820 17270
rect 254768 17206 254820 17212
rect 253952 16546 254256 16574
rect 252652 3800 252704 3806
rect 252652 3742 252704 3748
rect 253204 3800 253256 3806
rect 253204 3742 253256 3748
rect 251272 3460 251324 3466
rect 252572 3454 253520 3482
rect 251272 3402 251324 3408
rect 252376 3052 252428 3058
rect 252376 2994 252428 3000
rect 252388 480 252416 2994
rect 253492 480 253520 3454
rect 254228 490 254256 16546
rect 254872 3466 254900 96902
rect 254952 96824 255004 96830
rect 254952 96766 255004 96772
rect 254964 87582 254992 96766
rect 254952 87576 255004 87582
rect 254952 87518 255004 87524
rect 255056 81190 255084 97022
rect 255148 90302 255176 100014
rect 255240 96898 255268 100028
rect 255228 96892 255280 96898
rect 255228 96834 255280 96840
rect 255424 95198 255452 100028
rect 255884 99074 255912 100028
rect 255872 99068 255924 99074
rect 255872 99010 255924 99016
rect 255964 97572 256016 97578
rect 255964 97514 256016 97520
rect 255412 95192 255464 95198
rect 255412 95134 255464 95140
rect 255976 93854 256004 97514
rect 256068 95130 256096 100028
rect 256056 95124 256108 95130
rect 256056 95066 256108 95072
rect 255976 93826 256096 93854
rect 255964 93152 256016 93158
rect 255964 93094 256016 93100
rect 255136 90296 255188 90302
rect 255136 90238 255188 90244
rect 255044 81184 255096 81190
rect 255044 81126 255096 81132
rect 255320 18692 255372 18698
rect 255320 18634 255372 18640
rect 255332 16574 255360 18634
rect 255332 16546 255912 16574
rect 254860 3460 254912 3466
rect 254860 3402 254912 3408
rect 254504 598 254716 626
rect 254504 490 254532 598
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254228 462 254532 490
rect 254688 480 254716 598
rect 255884 480 255912 16546
rect 255976 4078 256004 93094
rect 256068 79354 256096 93826
rect 256252 89690 256280 100028
rect 256344 100014 256450 100042
rect 256528 100014 256634 100042
rect 256240 89684 256292 89690
rect 256240 89626 256292 89632
rect 256056 79348 256108 79354
rect 256056 79290 256108 79296
rect 256344 26926 256372 100014
rect 256528 93022 256556 100014
rect 256896 96966 256924 100028
rect 256884 96960 256936 96966
rect 256884 96902 256936 96908
rect 257080 96898 257108 100028
rect 257264 97986 257292 100028
rect 257252 97980 257304 97986
rect 257252 97922 257304 97928
rect 257068 96892 257120 96898
rect 257068 96834 257120 96840
rect 257448 96830 257476 100028
rect 257436 96824 257488 96830
rect 257436 96766 257488 96772
rect 256516 93016 256568 93022
rect 256516 92958 256568 92964
rect 257632 29714 257660 100028
rect 257922 100014 258028 100042
rect 257712 96960 257764 96966
rect 257712 96902 257764 96908
rect 257724 91730 257752 96902
rect 257896 96892 257948 96898
rect 257896 96834 257948 96840
rect 257804 96824 257856 96830
rect 257804 96766 257856 96772
rect 257712 91724 257764 91730
rect 257712 91666 257764 91672
rect 257816 88330 257844 96766
rect 257804 88324 257856 88330
rect 257804 88266 257856 88272
rect 257908 79762 257936 96834
rect 258000 93090 258028 100014
rect 258276 96966 258304 100028
rect 258264 96960 258316 96966
rect 258264 96902 258316 96908
rect 258460 95062 258488 100028
rect 258644 96830 258672 100028
rect 258934 100014 259040 100042
rect 258908 96960 258960 96966
rect 258908 96902 258960 96908
rect 258632 96824 258684 96830
rect 258632 96766 258684 96772
rect 258448 95056 258500 95062
rect 258448 94998 258500 95004
rect 257988 93084 258040 93090
rect 257988 93026 258040 93032
rect 258080 86420 258132 86426
rect 258080 86362 258132 86368
rect 257896 79756 257948 79762
rect 257896 79698 257948 79704
rect 257620 29708 257672 29714
rect 257620 29650 257672 29656
rect 256332 26920 256384 26926
rect 256332 26862 256384 26868
rect 257344 18760 257396 18766
rect 257344 18702 257396 18708
rect 255964 4072 256016 4078
rect 255964 4014 256016 4020
rect 257356 4010 257384 18702
rect 257344 4004 257396 4010
rect 257344 3946 257396 3952
rect 257068 3936 257120 3942
rect 257068 3878 257120 3884
rect 257080 480 257108 3878
rect 258092 3058 258120 86362
rect 258920 78334 258948 96902
rect 258908 78328 258960 78334
rect 258908 78270 258960 78276
rect 259012 28286 259040 100014
rect 259104 96966 259132 100028
rect 259196 100014 259302 100042
rect 259092 96960 259144 96966
rect 259092 96902 259144 96908
rect 259092 96824 259144 96830
rect 259092 96766 259144 96772
rect 259104 86970 259132 96766
rect 259092 86964 259144 86970
rect 259092 86906 259144 86912
rect 259196 86902 259224 100014
rect 259472 97102 259500 100028
rect 259460 97096 259512 97102
rect 259460 97038 259512 97044
rect 259368 96960 259420 96966
rect 259368 96902 259420 96908
rect 259380 93838 259408 96902
rect 259656 96830 259684 100028
rect 259946 100014 260052 100042
rect 259644 96824 259696 96830
rect 259644 96766 259696 96772
rect 260024 93854 260052 100014
rect 260116 96966 260144 100028
rect 260104 96960 260156 96966
rect 260104 96902 260156 96908
rect 260300 96898 260328 100028
rect 260392 100014 260498 100042
rect 260288 96892 260340 96898
rect 260288 96834 260340 96840
rect 259368 93832 259420 93838
rect 260024 93826 260328 93854
rect 259368 93774 259420 93780
rect 259184 86896 259236 86902
rect 259184 86838 259236 86844
rect 260104 83496 260156 83502
rect 260104 83438 260156 83444
rect 259000 28280 259052 28286
rect 259000 28222 259052 28228
rect 258724 14544 258776 14550
rect 258724 14486 258776 14492
rect 258736 3466 258764 14486
rect 260116 3874 260144 83438
rect 260196 18624 260248 18630
rect 260196 18566 260248 18572
rect 260104 3868 260156 3874
rect 260104 3810 260156 3816
rect 258724 3460 258776 3466
rect 258724 3402 258776 3408
rect 258264 3392 258316 3398
rect 258264 3334 258316 3340
rect 258080 3052 258132 3058
rect 258080 2994 258132 3000
rect 258276 480 258304 3334
rect 260208 3194 260236 18566
rect 260300 3505 260328 93826
rect 260392 88262 260420 100014
rect 260852 97578 260880 100028
rect 260840 97572 260892 97578
rect 260840 97514 260892 97520
rect 260564 97096 260616 97102
rect 260564 97038 260616 97044
rect 260472 96960 260524 96966
rect 260472 96902 260524 96908
rect 260380 88256 260432 88262
rect 260380 88198 260432 88204
rect 260484 84046 260512 96902
rect 260472 84040 260524 84046
rect 260472 83982 260524 83988
rect 260576 79694 260604 97038
rect 260748 96892 260800 96898
rect 260748 96834 260800 96840
rect 260656 96824 260708 96830
rect 260656 96766 260708 96772
rect 260564 79688 260616 79694
rect 260564 79630 260616 79636
rect 260668 16574 260696 96766
rect 260760 93770 260788 96834
rect 261128 96830 261156 100028
rect 261116 96824 261168 96830
rect 261116 96766 261168 96772
rect 261312 96762 261340 100028
rect 261496 97986 261524 100028
rect 261484 97980 261536 97986
rect 261484 97922 261536 97928
rect 261680 96966 261708 100028
rect 261864 97102 261892 100028
rect 261956 100014 262154 100042
rect 261852 97096 261904 97102
rect 261852 97038 261904 97044
rect 261668 96960 261720 96966
rect 261956 96948 261984 100014
rect 262128 97096 262180 97102
rect 262128 97038 262180 97044
rect 261668 96902 261720 96908
rect 261772 96920 261984 96948
rect 262036 96960 262088 96966
rect 261300 96756 261352 96762
rect 261300 96698 261352 96704
rect 260748 93764 260800 93770
rect 260748 93706 260800 93712
rect 261772 93702 261800 96920
rect 262036 96902 262088 96908
rect 261944 96824 261996 96830
rect 261944 96766 261996 96772
rect 261852 96756 261904 96762
rect 261852 96698 261904 96704
rect 261760 93696 261812 93702
rect 261760 93638 261812 93644
rect 261864 78266 261892 96698
rect 261956 86766 261984 96766
rect 261944 86760 261996 86766
rect 261944 86702 261996 86708
rect 262048 85474 262076 96902
rect 262140 96490 262168 97038
rect 262324 96830 262352 100028
rect 262508 97714 262536 100028
rect 262496 97708 262548 97714
rect 262496 97650 262548 97656
rect 262312 96824 262364 96830
rect 262312 96766 262364 96772
rect 262128 96484 262180 96490
rect 262128 96426 262180 96432
rect 262692 94994 262720 100028
rect 262890 100014 263088 100042
rect 263060 96948 263088 100014
rect 263152 99006 263180 100028
rect 263140 99000 263192 99006
rect 263140 98942 263192 98948
rect 263060 96920 263272 96948
rect 263140 96824 263192 96830
rect 263140 96766 263192 96772
rect 262680 94988 262732 94994
rect 262680 94930 262732 94936
rect 262036 85468 262088 85474
rect 262036 85410 262088 85416
rect 263152 85406 263180 96766
rect 263140 85400 263192 85406
rect 263140 85342 263192 85348
rect 263244 85338 263272 96920
rect 263336 92478 263364 100028
rect 263520 94314 263548 100028
rect 263704 97374 263732 100028
rect 263784 97640 263836 97646
rect 263784 97582 263836 97588
rect 263600 97368 263652 97374
rect 263600 97310 263652 97316
rect 263692 97368 263744 97374
rect 263692 97310 263744 97316
rect 263508 94308 263560 94314
rect 263508 94250 263560 94256
rect 263324 92472 263376 92478
rect 263324 92414 263376 92420
rect 263232 85332 263284 85338
rect 263232 85274 263284 85280
rect 262220 84924 262272 84930
rect 262220 84866 262272 84872
rect 261852 78260 261904 78266
rect 261852 78202 261904 78208
rect 260668 16546 260788 16574
rect 260286 3496 260342 3505
rect 260286 3431 260342 3440
rect 260656 3460 260708 3466
rect 260656 3402 260708 3408
rect 260196 3188 260248 3194
rect 260196 3130 260248 3136
rect 259460 3052 259512 3058
rect 259460 2994 259512 3000
rect 259472 480 259500 2994
rect 260668 480 260696 3402
rect 260760 3369 260788 16546
rect 260840 4072 260892 4078
rect 260840 4014 260892 4020
rect 260852 3670 260880 4014
rect 260840 3664 260892 3670
rect 260840 3606 260892 3612
rect 261760 3664 261812 3670
rect 261760 3606 261812 3612
rect 260746 3360 260802 3369
rect 260746 3295 260802 3304
rect 261772 480 261800 3606
rect 262232 3058 262260 84866
rect 263612 4078 263640 97310
rect 263796 94382 263824 97582
rect 263888 96898 263916 100028
rect 264164 96966 264192 100028
rect 264348 97782 264376 100028
rect 264546 100014 264652 100042
rect 264730 100014 264836 100042
rect 264914 100026 265020 100042
rect 264914 100020 265032 100026
rect 264914 100014 264980 100020
rect 264336 97776 264388 97782
rect 264336 97718 264388 97724
rect 264152 96960 264204 96966
rect 264152 96902 264204 96908
rect 263876 96892 263928 96898
rect 263876 96834 263928 96840
rect 263784 94376 263836 94382
rect 263784 94318 263836 94324
rect 264624 92410 264652 100014
rect 264704 96960 264756 96966
rect 264704 96902 264756 96908
rect 264612 92404 264664 92410
rect 264612 92346 264664 92352
rect 263692 91860 263744 91866
rect 263692 91802 263744 91808
rect 263600 4072 263652 4078
rect 263600 4014 263652 4020
rect 262956 3732 263008 3738
rect 262956 3674 263008 3680
rect 262220 3052 262272 3058
rect 262220 2994 262272 3000
rect 262968 480 262996 3674
rect 263704 3398 263732 91802
rect 264716 83978 264744 96902
rect 264704 83972 264756 83978
rect 264704 83914 264756 83920
rect 264808 83910 264836 100014
rect 264980 99962 265032 99968
rect 264888 96892 264940 96898
rect 264888 96834 264940 96840
rect 264796 83904 264848 83910
rect 264796 83846 264848 83852
rect 264900 3738 264928 96834
rect 265176 96830 265204 100028
rect 265360 96898 265388 100028
rect 265544 99278 265572 100028
rect 265532 99272 265584 99278
rect 265532 99214 265584 99220
rect 265728 96966 265756 100028
rect 265716 96960 265768 96966
rect 265716 96902 265768 96908
rect 265348 96892 265400 96898
rect 265348 96834 265400 96840
rect 265164 96824 265216 96830
rect 265164 96766 265216 96772
rect 265912 83842 265940 100028
rect 266096 100014 266202 100042
rect 265992 96960 266044 96966
rect 265992 96902 266044 96908
rect 266004 92206 266032 96902
rect 265992 92200 266044 92206
rect 265992 92142 266044 92148
rect 266096 89622 266124 100014
rect 266372 96966 266400 100028
rect 266360 96960 266412 96966
rect 266360 96902 266412 96908
rect 266176 96892 266228 96898
rect 266176 96834 266228 96840
rect 266084 89616 266136 89622
rect 266084 89558 266136 89564
rect 266188 85270 266216 96834
rect 266556 96830 266584 100028
rect 266740 97510 266768 100028
rect 266728 97504 266780 97510
rect 266728 97446 266780 97452
rect 266924 96898 266952 100028
rect 267214 100014 267320 100042
rect 267004 97436 267056 97442
rect 267004 97378 267056 97384
rect 266912 96892 266964 96898
rect 266912 96834 266964 96840
rect 266268 96824 266320 96830
rect 266268 96766 266320 96772
rect 266544 96824 266596 96830
rect 266544 96766 266596 96772
rect 266280 93634 266308 96766
rect 266268 93628 266320 93634
rect 266268 93570 266320 93576
rect 266452 91792 266504 91798
rect 266452 91734 266504 91740
rect 266360 90500 266412 90506
rect 266360 90442 266412 90448
rect 266176 85264 266228 85270
rect 266176 85206 266228 85212
rect 265900 83836 265952 83842
rect 265900 83778 265952 83784
rect 265348 4140 265400 4146
rect 265348 4082 265400 4088
rect 264888 3732 264940 3738
rect 264888 3674 264940 3680
rect 263692 3392 263744 3398
rect 263692 3334 263744 3340
rect 264152 3188 264204 3194
rect 264152 3130 264204 3136
rect 264164 480 264192 3130
rect 265360 480 265388 4082
rect 266372 3482 266400 90442
rect 266464 3670 266492 91734
rect 267016 10334 267044 97378
rect 267292 83774 267320 100014
rect 267384 97238 267412 100028
rect 267476 100014 267582 100042
rect 267372 97232 267424 97238
rect 267372 97174 267424 97180
rect 267372 96960 267424 96966
rect 267372 96902 267424 96908
rect 267384 92138 267412 96902
rect 267372 92132 267424 92138
rect 267372 92074 267424 92080
rect 267476 91050 267504 100014
rect 267648 96892 267700 96898
rect 267648 96834 267700 96840
rect 267556 96824 267608 96830
rect 267556 96766 267608 96772
rect 267464 91044 267516 91050
rect 267464 90986 267516 90992
rect 267568 86698 267596 96766
rect 267660 92070 267688 96834
rect 267752 96762 267780 100028
rect 267740 96756 267792 96762
rect 267740 96698 267792 96704
rect 267936 96694 267964 100028
rect 268212 96966 268240 100028
rect 268410 100014 268516 100042
rect 268384 97776 268436 97782
rect 268384 97718 268436 97724
rect 268200 96960 268252 96966
rect 268200 96902 268252 96908
rect 267924 96688 267976 96694
rect 267924 96630 267976 96636
rect 268396 93854 268424 97718
rect 268488 96914 268516 100014
rect 268580 97850 268608 100028
rect 268568 97844 268620 97850
rect 268568 97786 268620 97792
rect 268488 96886 268700 96914
rect 268568 96756 268620 96762
rect 268568 96698 268620 96704
rect 268396 93826 268516 93854
rect 267648 92064 267700 92070
rect 267648 92006 267700 92012
rect 268384 90432 268436 90438
rect 268384 90374 268436 90380
rect 267556 86692 267608 86698
rect 267556 86634 267608 86640
rect 267280 83768 267332 83774
rect 267280 83710 267332 83716
rect 267740 14476 267792 14482
rect 267740 14418 267792 14424
rect 267004 10328 267056 10334
rect 267004 10270 267056 10276
rect 266452 3664 266504 3670
rect 266452 3606 266504 3612
rect 266372 3454 266584 3482
rect 266556 480 266584 3454
rect 267752 480 267780 14418
rect 268396 3534 268424 90374
rect 268488 18630 268516 93826
rect 268580 83706 268608 96698
rect 268568 83700 268620 83706
rect 268568 83642 268620 83648
rect 268672 82618 268700 96886
rect 268764 90982 268792 100028
rect 268856 100014 268962 100042
rect 268752 90976 268804 90982
rect 268752 90918 268804 90924
rect 268856 85202 268884 100014
rect 268936 96960 268988 96966
rect 268936 96902 268988 96908
rect 268948 93566 268976 96902
rect 269224 96762 269252 100028
rect 269408 96966 269436 100028
rect 269396 96960 269448 96966
rect 269396 96902 269448 96908
rect 269592 96830 269620 100028
rect 269776 97782 269804 100028
rect 269974 100014 270080 100042
rect 270158 100014 270356 100042
rect 269764 97776 269816 97782
rect 269764 97718 269816 97724
rect 269764 97300 269816 97306
rect 269764 97242 269816 97248
rect 269580 96824 269632 96830
rect 269580 96766 269632 96772
rect 269212 96756 269264 96762
rect 269212 96698 269264 96704
rect 269028 96688 269080 96694
rect 269028 96630 269080 96636
rect 268936 93560 268988 93566
rect 268936 93502 268988 93508
rect 269040 92342 269068 96630
rect 269120 96076 269172 96082
rect 269120 96018 269172 96024
rect 269028 92336 269080 92342
rect 269028 92278 269080 92284
rect 268844 85196 268896 85202
rect 268844 85138 268896 85144
rect 268660 82612 268712 82618
rect 268660 82554 268712 82560
rect 268476 18624 268528 18630
rect 268476 18566 268528 18572
rect 268844 4004 268896 4010
rect 268844 3946 268896 3952
rect 268384 3528 268436 3534
rect 268384 3470 268436 3476
rect 268856 480 268884 3946
rect 269132 3942 269160 96018
rect 269776 4826 269804 97242
rect 269948 96960 270000 96966
rect 269948 96902 270000 96908
rect 269960 92002 269988 96902
rect 270052 96642 270080 100014
rect 270328 96914 270356 100014
rect 270420 97646 270448 100028
rect 270604 99958 270632 100028
rect 270592 99952 270644 99958
rect 270592 99894 270644 99900
rect 270408 97640 270460 97646
rect 270408 97582 270460 97588
rect 270328 96886 270448 96914
rect 270316 96824 270368 96830
rect 270316 96766 270368 96772
rect 270052 96614 270264 96642
rect 269948 91996 270000 92002
rect 269948 91938 270000 91944
rect 270236 90914 270264 96614
rect 270224 90908 270276 90914
rect 270224 90850 270276 90856
rect 270328 83638 270356 96766
rect 270316 83632 270368 83638
rect 270316 83574 270368 83580
rect 270420 82550 270448 96886
rect 270788 96830 270816 100028
rect 270972 96898 271000 100028
rect 271156 99890 271184 100028
rect 271144 99884 271196 99890
rect 271144 99826 271196 99832
rect 271236 97708 271288 97714
rect 271236 97650 271288 97656
rect 271144 97504 271196 97510
rect 271144 97446 271196 97452
rect 270960 96892 271012 96898
rect 270960 96834 271012 96840
rect 270776 96824 270828 96830
rect 270776 96766 270828 96772
rect 270408 82544 270460 82550
rect 270408 82486 270460 82492
rect 271156 4894 271184 97446
rect 271248 86834 271276 97650
rect 271432 96966 271460 100028
rect 271512 97572 271564 97578
rect 271512 97514 271564 97520
rect 271420 96960 271472 96966
rect 271420 96902 271472 96908
rect 271524 96558 271552 97514
rect 271616 97510 271644 100028
rect 271708 100014 271814 100042
rect 271604 97504 271656 97510
rect 271604 97446 271656 97452
rect 271708 96914 271736 100014
rect 271616 96886 271736 96914
rect 271788 96960 271840 96966
rect 271788 96902 271840 96908
rect 271512 96552 271564 96558
rect 271512 96494 271564 96500
rect 271616 90846 271644 96886
rect 271696 96824 271748 96830
rect 271696 96766 271748 96772
rect 271604 90840 271656 90846
rect 271604 90782 271656 90788
rect 271236 86828 271288 86834
rect 271236 86770 271288 86776
rect 271708 82482 271736 96766
rect 271696 82476 271748 82482
rect 271696 82418 271748 82424
rect 271236 82204 271288 82210
rect 271236 82146 271288 82152
rect 271144 4888 271196 4894
rect 271144 4830 271196 4836
rect 269764 4820 269816 4826
rect 269764 4762 269816 4768
rect 269120 3936 269172 3942
rect 269120 3878 269172 3884
rect 270040 3528 270092 3534
rect 270040 3470 270092 3476
rect 270052 480 270080 3470
rect 271248 3194 271276 82146
rect 271800 81122 271828 96902
rect 271984 96898 272012 100028
rect 272168 97442 272196 100028
rect 272444 99822 272472 100028
rect 272432 99816 272484 99822
rect 272432 99758 272484 99764
rect 272156 97436 272208 97442
rect 272156 97378 272208 97384
rect 272628 96966 272656 100028
rect 272812 97306 272840 100028
rect 272904 100014 273010 100042
rect 272800 97300 272852 97306
rect 272800 97242 272852 97248
rect 272616 96960 272668 96966
rect 272616 96902 272668 96908
rect 271972 96892 272024 96898
rect 271972 96834 272024 96840
rect 272904 91934 272932 100014
rect 273076 96960 273128 96966
rect 273076 96902 273128 96908
rect 272984 96892 273036 96898
rect 272984 96834 273036 96840
rect 272892 91928 272944 91934
rect 272892 91870 272944 91876
rect 272996 88126 273024 96834
rect 272984 88120 273036 88126
rect 272984 88062 273036 88068
rect 273088 82414 273116 96902
rect 273076 82408 273128 82414
rect 273076 82350 273128 82356
rect 271788 81116 271840 81122
rect 271788 81058 271840 81064
rect 273180 81054 273208 100028
rect 273456 97102 273484 100028
rect 273640 99754 273668 100028
rect 273628 99748 273680 99754
rect 273628 99690 273680 99696
rect 273444 97096 273496 97102
rect 273444 97038 273496 97044
rect 273824 96966 273852 100028
rect 273812 96960 273864 96966
rect 273812 96902 273864 96908
rect 274008 96898 274036 100028
rect 274206 100014 274312 100042
rect 273996 96892 274048 96898
rect 273996 96834 274048 96840
rect 273904 96756 273956 96762
rect 273904 96698 273956 96704
rect 273168 81048 273220 81054
rect 273168 80990 273220 80996
rect 273916 32434 273944 96698
rect 274284 90778 274312 100014
rect 274364 96960 274416 96966
rect 274364 96902 274416 96908
rect 274272 90772 274324 90778
rect 274272 90714 274324 90720
rect 274376 83570 274404 96902
rect 274364 83564 274416 83570
rect 274364 83506 274416 83512
rect 274468 80986 274496 100028
rect 274652 97918 274680 100028
rect 274836 99686 274864 100028
rect 274824 99680 274876 99686
rect 274824 99622 274876 99628
rect 274640 97912 274692 97918
rect 274640 97854 274692 97860
rect 274548 96892 274600 96898
rect 274548 96834 274600 96840
rect 274456 80980 274508 80986
rect 274456 80922 274508 80928
rect 273904 32428 273956 32434
rect 273904 32370 273956 32376
rect 271328 3936 271380 3942
rect 271328 3878 271380 3884
rect 271236 3188 271288 3194
rect 271236 3130 271288 3136
rect 271340 1986 271368 3878
rect 273628 3868 273680 3874
rect 273628 3810 273680 3816
rect 272432 3392 272484 3398
rect 272432 3334 272484 3340
rect 271248 1958 271368 1986
rect 271248 480 271276 1958
rect 272444 480 272472 3334
rect 273640 480 273668 3810
rect 274560 3670 274588 96834
rect 275020 96830 275048 100028
rect 275008 96824 275060 96830
rect 275008 96766 275060 96772
rect 275204 96762 275232 100028
rect 275480 99618 275508 100028
rect 275678 100014 275784 100042
rect 275468 99612 275520 99618
rect 275468 99554 275520 99560
rect 275376 97436 275428 97442
rect 275376 97378 275428 97384
rect 275388 97102 275416 97378
rect 275284 97096 275336 97102
rect 275284 97038 275336 97044
rect 275376 97096 275428 97102
rect 275376 97038 275428 97044
rect 275192 96756 275244 96762
rect 275192 96698 275244 96704
rect 275296 75342 275324 97038
rect 275756 96914 275784 100014
rect 275848 97578 275876 100028
rect 276032 99550 276060 100028
rect 276020 99544 276072 99550
rect 276020 99486 276072 99492
rect 275836 97572 275888 97578
rect 275836 97514 275888 97520
rect 276112 97504 276164 97510
rect 276112 97446 276164 97452
rect 275756 96886 275876 96914
rect 276124 96898 276152 97446
rect 275744 96824 275796 96830
rect 275744 96766 275796 96772
rect 275756 89554 275784 96766
rect 275744 89548 275796 89554
rect 275744 89490 275796 89496
rect 275848 86630 275876 96886
rect 276112 96892 276164 96898
rect 276112 96834 276164 96840
rect 276216 96830 276244 100028
rect 276204 96824 276256 96830
rect 276204 96766 276256 96772
rect 275928 96756 275980 96762
rect 275928 96698 275980 96704
rect 275836 86624 275888 86630
rect 275836 86566 275888 86572
rect 275284 75336 275336 75342
rect 275284 75278 275336 75284
rect 275940 33794 275968 96698
rect 276492 94926 276520 100028
rect 276572 97640 276624 97646
rect 276572 97582 276624 97588
rect 276480 94920 276532 94926
rect 276480 94862 276532 94868
rect 276584 93854 276612 97582
rect 276676 96762 276704 100028
rect 276874 100014 276980 100042
rect 276952 96914 276980 100014
rect 277044 97510 277072 100028
rect 277136 100014 277242 100042
rect 277032 97504 277084 97510
rect 277032 97446 277084 97452
rect 276952 96886 277072 96914
rect 276940 96824 276992 96830
rect 276940 96766 276992 96772
rect 276664 96756 276716 96762
rect 276664 96698 276716 96704
rect 276584 93826 276704 93854
rect 276020 79348 276072 79354
rect 276020 79290 276072 79296
rect 275928 33788 275980 33794
rect 275928 33730 275980 33736
rect 276032 16574 276060 79290
rect 276676 76770 276704 93826
rect 276952 82346 276980 96766
rect 276940 82340 276992 82346
rect 276940 82282 276992 82288
rect 277044 79626 277072 96886
rect 277136 90710 277164 100014
rect 277504 96830 277532 100028
rect 277584 97980 277636 97986
rect 277584 97922 277636 97928
rect 277596 96966 277624 97922
rect 277688 96966 277716 100028
rect 277584 96960 277636 96966
rect 277584 96902 277636 96908
rect 277676 96960 277728 96966
rect 277676 96902 277728 96908
rect 277492 96824 277544 96830
rect 277492 96766 277544 96772
rect 277308 96756 277360 96762
rect 277308 96698 277360 96704
rect 277320 93498 277348 96698
rect 277872 94790 277900 100028
rect 278070 100014 278176 100042
rect 278044 97368 278096 97374
rect 278044 97310 278096 97316
rect 277860 94784 277912 94790
rect 277860 94726 277912 94732
rect 277308 93492 277360 93498
rect 277308 93434 277360 93440
rect 277124 90704 277176 90710
rect 277124 90646 277176 90652
rect 277032 79620 277084 79626
rect 277032 79562 277084 79568
rect 276664 76764 276716 76770
rect 276664 76706 276716 76712
rect 276032 16546 276704 16574
rect 276020 4072 276072 4078
rect 276020 4014 276072 4020
rect 274548 3664 274600 3670
rect 274548 3606 274600 3612
rect 274824 3188 274876 3194
rect 274824 3130 274876 3136
rect 274836 480 274864 3130
rect 276032 480 276060 4014
rect 276676 490 276704 16546
rect 278056 4962 278084 97310
rect 278148 97050 278176 100014
rect 278240 97442 278268 100028
rect 278516 99482 278544 100028
rect 278608 100014 278714 100042
rect 278504 99476 278556 99482
rect 278504 99418 278556 99424
rect 278228 97436 278280 97442
rect 278228 97378 278280 97384
rect 278148 97022 278544 97050
rect 278320 96960 278372 96966
rect 278320 96902 278372 96908
rect 278136 82136 278188 82142
rect 278136 82078 278188 82084
rect 278044 4956 278096 4962
rect 278044 4898 278096 4904
rect 278148 3874 278176 82078
rect 278332 69698 278360 96902
rect 278412 96824 278464 96830
rect 278412 96766 278464 96772
rect 278424 85134 278452 96766
rect 278412 85128 278464 85134
rect 278412 85070 278464 85076
rect 278516 82278 278544 97022
rect 278504 82272 278556 82278
rect 278504 82214 278556 82220
rect 278608 80918 278636 100014
rect 278884 96966 278912 100028
rect 279068 98938 279096 100028
rect 279056 98932 279108 98938
rect 279056 98874 279108 98880
rect 278872 96960 278924 96966
rect 278872 96902 278924 96908
rect 279252 94858 279280 100028
rect 279528 97374 279556 100028
rect 279712 99414 279740 100028
rect 279700 99408 279752 99414
rect 279700 99350 279752 99356
rect 279516 97368 279568 97374
rect 279516 97310 279568 97316
rect 279792 96960 279844 96966
rect 279792 96902 279844 96908
rect 279240 94852 279292 94858
rect 279240 94794 279292 94800
rect 278596 80912 278648 80918
rect 278596 80854 278648 80860
rect 278320 69692 278372 69698
rect 278320 69634 278372 69640
rect 278320 4820 278372 4826
rect 278320 4762 278372 4768
rect 278136 3868 278188 3874
rect 278136 3810 278188 3816
rect 276952 598 277164 626
rect 276952 490 276980 598
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 276676 462 276980 490
rect 277136 480 277164 598
rect 278332 480 278360 4762
rect 279516 4004 279568 4010
rect 279516 3946 279568 3952
rect 279528 480 279556 3946
rect 279804 3534 279832 96902
rect 279896 93430 279924 100028
rect 279988 100014 280094 100042
rect 279884 93424 279936 93430
rect 279884 93366 279936 93372
rect 279988 73914 280016 100014
rect 280264 96694 280292 100028
rect 280448 96830 280476 100028
rect 280632 100014 280738 100042
rect 280922 100014 281028 100042
rect 280436 96824 280488 96830
rect 280436 96766 280488 96772
rect 280632 96762 280660 100014
rect 280712 97912 280764 97918
rect 280712 97854 280764 97860
rect 280724 97102 280752 97854
rect 280804 97776 280856 97782
rect 280804 97718 280856 97724
rect 280816 97306 280844 97718
rect 280804 97300 280856 97306
rect 280804 97242 280856 97248
rect 280896 97300 280948 97306
rect 280896 97242 280948 97248
rect 280712 97096 280764 97102
rect 280712 97038 280764 97044
rect 280804 97028 280856 97034
rect 280804 96970 280856 96976
rect 280620 96756 280672 96762
rect 280620 96698 280672 96704
rect 280252 96688 280304 96694
rect 280252 96630 280304 96636
rect 280252 90364 280304 90370
rect 280252 90306 280304 90312
rect 279976 73908 280028 73914
rect 279976 73850 280028 73856
rect 280160 31068 280212 31074
rect 280160 31010 280212 31016
rect 279792 3528 279844 3534
rect 279792 3470 279844 3476
rect 280172 3482 280200 31010
rect 280264 4078 280292 90306
rect 280252 4072 280304 4078
rect 280252 4014 280304 4020
rect 280172 3454 280752 3482
rect 280724 480 280752 3454
rect 280816 3058 280844 96970
rect 280908 93854 280936 97242
rect 281000 96948 281028 100014
rect 281092 97102 281120 100028
rect 281276 97306 281304 100028
rect 281368 100014 281474 100042
rect 281264 97300 281316 97306
rect 281264 97242 281316 97248
rect 281080 97096 281132 97102
rect 281080 97038 281132 97044
rect 281368 96948 281396 100014
rect 281448 97096 281500 97102
rect 281448 97038 281500 97044
rect 281000 96920 281120 96948
rect 280908 93826 281028 93854
rect 281000 31074 281028 93826
rect 281092 91866 281120 96920
rect 281184 96920 281396 96948
rect 281080 91860 281132 91866
rect 281080 91802 281132 91808
rect 281184 89486 281212 96920
rect 281264 96824 281316 96830
rect 281460 96812 281488 97038
rect 281736 97034 281764 100028
rect 281920 97481 281948 100028
rect 281906 97472 281962 97481
rect 281906 97407 281962 97416
rect 281724 97028 281776 97034
rect 281724 96970 281776 96976
rect 281264 96766 281316 96772
rect 281368 96784 281488 96812
rect 281172 89480 281224 89486
rect 281172 89422 281224 89428
rect 281276 83502 281304 96766
rect 281264 83496 281316 83502
rect 281264 83438 281316 83444
rect 281368 79558 281396 96784
rect 281448 96688 281500 96694
rect 281448 96630 281500 96636
rect 281460 90642 281488 96630
rect 282104 96218 282132 100028
rect 282288 96966 282316 100028
rect 282486 100014 282592 100042
rect 282762 100014 282868 100042
rect 282276 96960 282328 96966
rect 282276 96902 282328 96908
rect 282092 96212 282144 96218
rect 282092 96154 282144 96160
rect 281540 96008 281592 96014
rect 281540 95950 281592 95956
rect 281448 90636 281500 90642
rect 281448 90578 281500 90584
rect 281356 79552 281408 79558
rect 281356 79494 281408 79500
rect 280988 31068 281040 31074
rect 280988 31010 281040 31016
rect 281552 3942 281580 95950
rect 282564 79490 282592 100014
rect 282736 97028 282788 97034
rect 282736 96970 282788 96976
rect 282644 96960 282696 96966
rect 282644 96902 282696 96908
rect 282656 89418 282684 96902
rect 282644 89412 282696 89418
rect 282644 89354 282696 89360
rect 282748 80850 282776 96970
rect 282840 96082 282868 100014
rect 282932 99346 282960 100028
rect 282920 99340 282972 99346
rect 282920 99282 282972 99288
rect 283116 97034 283144 100028
rect 283104 97028 283156 97034
rect 283104 96970 283156 96976
rect 283300 96286 283328 100028
rect 283484 96966 283512 100028
rect 283774 100014 283880 100042
rect 283472 96960 283524 96966
rect 283472 96902 283524 96908
rect 283288 96280 283340 96286
rect 283288 96222 283340 96228
rect 282828 96076 282880 96082
rect 282828 96018 282880 96024
rect 282736 80844 282788 80850
rect 282736 80786 282788 80792
rect 282552 79484 282604 79490
rect 282552 79426 282604 79432
rect 283852 78198 283880 100014
rect 283944 97102 283972 100028
rect 284036 100014 284142 100042
rect 283932 97096 283984 97102
rect 283932 97038 283984 97044
rect 283932 96960 283984 96966
rect 283932 96902 283984 96908
rect 283944 90574 283972 96902
rect 283932 90568 283984 90574
rect 283932 90510 283984 90516
rect 284036 89350 284064 100014
rect 284208 97096 284260 97102
rect 284208 97038 284260 97044
rect 284116 97028 284168 97034
rect 284116 96970 284168 96976
rect 284024 89344 284076 89350
rect 284024 89286 284076 89292
rect 284128 82210 284156 96970
rect 284220 96422 284248 97038
rect 284312 97034 284340 100028
rect 284496 97209 284524 100028
rect 284482 97200 284538 97209
rect 284482 97135 284538 97144
rect 284300 97028 284352 97034
rect 284300 96970 284352 96976
rect 284772 96966 284800 100028
rect 284970 100014 285076 100042
rect 284760 96960 284812 96966
rect 284760 96902 284812 96908
rect 284208 96416 284260 96422
rect 284208 96358 284260 96364
rect 285048 93854 285076 100014
rect 285140 96354 285168 100028
rect 285232 100014 285338 100042
rect 285128 96348 285180 96354
rect 285128 96290 285180 96296
rect 285048 93826 285168 93854
rect 284116 82204 284168 82210
rect 284116 82146 284168 82152
rect 283840 78192 283892 78198
rect 283840 78134 283892 78140
rect 284300 39364 284352 39370
rect 284300 39306 284352 39312
rect 281540 3936 281592 3942
rect 281540 3878 281592 3884
rect 281908 3324 281960 3330
rect 281908 3266 281960 3272
rect 280804 3052 280856 3058
rect 280804 2994 280856 3000
rect 281920 480 281948 3266
rect 283104 3052 283156 3058
rect 283104 2994 283156 3000
rect 283116 480 283144 2994
rect 284312 480 284340 39306
rect 285140 8974 285168 93826
rect 285232 89214 285260 100014
rect 285404 97028 285456 97034
rect 285404 96970 285456 96976
rect 285312 96960 285364 96966
rect 285312 96902 285364 96908
rect 285324 89282 285352 96902
rect 285312 89276 285364 89282
rect 285312 89218 285364 89224
rect 285220 89208 285272 89214
rect 285220 89150 285272 89156
rect 285416 78130 285444 96970
rect 285404 78124 285456 78130
rect 285404 78066 285456 78072
rect 285508 13122 285536 100028
rect 285798 100014 285904 100042
rect 285876 96014 285904 100014
rect 285968 97034 285996 100028
rect 285956 97028 286008 97034
rect 285956 96970 286008 96976
rect 286152 96830 286180 100028
rect 286140 96824 286192 96830
rect 286140 96766 286192 96772
rect 285864 96008 285916 96014
rect 285864 95950 285916 95956
rect 285772 95940 285824 95946
rect 285772 95882 285824 95888
rect 285680 89004 285732 89010
rect 285680 88946 285732 88952
rect 285496 13116 285548 13122
rect 285496 13058 285548 13064
rect 285128 8968 285180 8974
rect 285128 8910 285180 8916
rect 285404 3392 285456 3398
rect 285404 3334 285456 3340
rect 285416 480 285444 3334
rect 285692 3210 285720 88946
rect 285784 3330 285812 95882
rect 286336 94654 286364 100028
rect 286520 96966 286548 100028
rect 286612 100014 286810 100042
rect 286508 96960 286560 96966
rect 286508 96902 286560 96908
rect 286324 94648 286376 94654
rect 286324 94590 286376 94596
rect 286612 79422 286640 100014
rect 286980 98802 287008 100028
rect 286968 98796 287020 98802
rect 286968 98738 287020 98744
rect 287164 97034 287192 100028
rect 286692 97028 286744 97034
rect 286692 96970 286744 96976
rect 287152 97028 287204 97034
rect 287152 96970 287204 96976
rect 286704 89146 286732 96970
rect 287348 96966 287376 100028
rect 287532 98734 287560 100028
rect 287520 98728 287572 98734
rect 287520 98670 287572 98676
rect 286784 96960 286836 96966
rect 286784 96902 286836 96908
rect 287336 96960 287388 96966
rect 287336 96902 287388 96908
rect 286692 89140 286744 89146
rect 286692 89082 286744 89088
rect 286796 88058 286824 96902
rect 287808 96898 287836 100028
rect 287888 96960 287940 96966
rect 287888 96902 287940 96908
rect 287796 96892 287848 96898
rect 287796 96834 287848 96840
rect 286876 96824 286928 96830
rect 286876 96766 286928 96772
rect 286784 88052 286836 88058
rect 286784 87994 286836 88000
rect 286888 80782 286916 96766
rect 287060 87644 287112 87650
rect 287060 87586 287112 87592
rect 286876 80776 286928 80782
rect 286876 80718 286928 80724
rect 286600 79416 286652 79422
rect 286600 79358 286652 79364
rect 287072 4010 287100 87586
rect 287900 78062 287928 96902
rect 287888 78056 287940 78062
rect 287888 77998 287940 78004
rect 287992 14482 288020 100028
rect 288072 96892 288124 96898
rect 288072 96834 288124 96840
rect 288084 87990 288112 96834
rect 288176 94722 288204 100028
rect 288268 100014 288374 100042
rect 288164 94716 288216 94722
rect 288164 94658 288216 94664
rect 288072 87984 288124 87990
rect 288072 87926 288124 87932
rect 288268 87854 288296 100014
rect 288348 97028 288400 97034
rect 288348 96970 288400 96976
rect 288360 90506 288388 96970
rect 288544 96694 288572 100028
rect 288532 96688 288584 96694
rect 288532 96630 288584 96636
rect 288820 94586 288848 100028
rect 289004 96966 289032 100028
rect 289202 100014 289308 100042
rect 288992 96960 289044 96966
rect 289280 96948 289308 100014
rect 289372 97306 289400 100028
rect 289464 100014 289570 100042
rect 289360 97300 289412 97306
rect 289360 97242 289412 97248
rect 289280 96920 289400 96948
rect 288992 96902 289044 96908
rect 289268 96688 289320 96694
rect 289268 96630 289320 96636
rect 288808 94580 288860 94586
rect 288808 94522 288860 94528
rect 288440 94512 288492 94518
rect 288440 94454 288492 94460
rect 288348 90500 288400 90506
rect 288348 90442 288400 90448
rect 288256 87848 288308 87854
rect 288256 87790 288308 87796
rect 287980 14476 288032 14482
rect 287980 14418 288032 14424
rect 287796 6180 287848 6186
rect 287796 6122 287848 6128
rect 287060 4004 287112 4010
rect 287060 3946 287112 3952
rect 285772 3324 285824 3330
rect 285772 3266 285824 3272
rect 285692 3182 286640 3210
rect 286612 480 286640 3182
rect 287808 480 287836 6122
rect 288452 3398 288480 94454
rect 289280 76702 289308 96630
rect 289268 76696 289320 76702
rect 289268 76638 289320 76644
rect 289372 6186 289400 96920
rect 289464 89078 289492 100014
rect 289728 97300 289780 97306
rect 289728 97242 289780 97248
rect 289544 96960 289596 96966
rect 289544 96902 289596 96908
rect 289452 89072 289504 89078
rect 289452 89014 289504 89020
rect 289556 87786 289584 96902
rect 289740 94518 289768 97242
rect 289832 96937 289860 100028
rect 290016 97617 290044 100028
rect 290002 97608 290058 97617
rect 290002 97543 290058 97552
rect 290200 96966 290228 100028
rect 290188 96960 290240 96966
rect 289818 96928 289874 96937
rect 290188 96902 290240 96908
rect 289818 96863 289874 96872
rect 290384 96762 290412 100028
rect 290568 98666 290596 100028
rect 290766 100014 290964 100042
rect 290556 98660 290608 98666
rect 290556 98602 290608 98608
rect 290832 96892 290884 96898
rect 290832 96834 290884 96840
rect 290372 96756 290424 96762
rect 290372 96698 290424 96704
rect 289728 94512 289780 94518
rect 289728 94454 289780 94460
rect 289544 87780 289596 87786
rect 289544 87722 289596 87728
rect 290844 79354 290872 96834
rect 290936 91798 290964 100014
rect 291028 96898 291056 100028
rect 291108 96960 291160 96966
rect 291108 96902 291160 96908
rect 291016 96892 291068 96898
rect 291016 96834 291068 96840
rect 291016 96756 291068 96762
rect 291016 96698 291068 96704
rect 290924 91792 290976 91798
rect 290924 91734 290976 91740
rect 291028 85066 291056 96698
rect 291120 93294 291148 96902
rect 291212 95946 291240 100028
rect 291396 96898 291424 100028
rect 291580 97034 291608 100028
rect 291672 100014 291778 100042
rect 291568 97028 291620 97034
rect 291568 96970 291620 96976
rect 291384 96892 291436 96898
rect 291384 96834 291436 96840
rect 291200 95940 291252 95946
rect 291200 95882 291252 95888
rect 291672 94761 291700 100014
rect 291844 97300 291896 97306
rect 291844 97242 291896 97248
rect 291752 97164 291804 97170
rect 291752 97106 291804 97112
rect 291658 94752 291714 94761
rect 291658 94687 291714 94696
rect 291764 93854 291792 97106
rect 291856 96830 291884 97242
rect 292040 96966 292068 100028
rect 292132 100014 292238 100042
rect 292028 96960 292080 96966
rect 291934 96928 291990 96937
rect 292028 96902 292080 96908
rect 291934 96863 291990 96872
rect 291844 96824 291896 96830
rect 291844 96766 291896 96772
rect 291764 93826 291884 93854
rect 291108 93288 291160 93294
rect 291108 93230 291160 93236
rect 291292 86352 291344 86358
rect 291292 86294 291344 86300
rect 291016 85060 291068 85066
rect 291016 85002 291068 85008
rect 290832 79348 290884 79354
rect 290832 79290 290884 79296
rect 291200 10328 291252 10334
rect 291200 10270 291252 10276
rect 289360 6180 289412 6186
rect 289360 6122 289412 6128
rect 288992 3868 289044 3874
rect 288992 3810 289044 3816
rect 288440 3392 288492 3398
rect 288440 3334 288492 3340
rect 289004 480 289032 3810
rect 290188 3800 290240 3806
rect 290188 3742 290240 3748
rect 290200 480 290228 3742
rect 291212 3482 291240 10270
rect 291304 3806 291332 86294
rect 291292 3800 291344 3806
rect 291292 3742 291344 3748
rect 291212 3454 291424 3482
rect 291396 480 291424 3454
rect 291856 3330 291884 93826
rect 291948 93362 291976 96863
rect 291936 93356 291988 93362
rect 291936 93298 291988 93304
rect 292132 84194 292160 100014
rect 292408 98870 292436 100028
rect 292396 98864 292448 98870
rect 292396 98806 292448 98812
rect 292396 97028 292448 97034
rect 292396 96970 292448 96976
rect 292304 96960 292356 96966
rect 292304 96902 292356 96908
rect 292212 96892 292264 96898
rect 292212 96834 292264 96840
rect 292224 88194 292252 96834
rect 292212 88188 292264 88194
rect 292212 88130 292264 88136
rect 292316 86562 292344 96902
rect 292304 86556 292356 86562
rect 292304 86498 292356 86504
rect 292040 84166 292160 84194
rect 292040 10334 292068 84166
rect 292408 76634 292436 96970
rect 292592 96898 292620 100028
rect 292776 97034 292804 100028
rect 293052 98841 293080 100028
rect 293038 98832 293094 98841
rect 293038 98767 293094 98776
rect 292764 97028 292816 97034
rect 292764 96970 292816 96976
rect 293236 96966 293264 100028
rect 293434 100014 293540 100042
rect 293224 96960 293276 96966
rect 293224 96902 293276 96908
rect 292580 96892 292632 96898
rect 292580 96834 292632 96840
rect 293408 96892 293460 96898
rect 293408 96834 293460 96840
rect 293420 90438 293448 96834
rect 293408 90432 293460 90438
rect 293408 90374 293460 90380
rect 292396 76628 292448 76634
rect 292396 76570 292448 76576
rect 293512 15910 293540 100014
rect 293604 97170 293632 100028
rect 293696 100014 293802 100042
rect 293592 97164 293644 97170
rect 293592 97106 293644 97112
rect 293592 96960 293644 96966
rect 293592 96902 293644 96908
rect 293604 87718 293632 96902
rect 293592 87712 293644 87718
rect 293592 87654 293644 87660
rect 293696 86494 293724 100014
rect 293868 97164 293920 97170
rect 293868 97106 293920 97112
rect 293776 97028 293828 97034
rect 293776 96970 293828 96976
rect 293684 86488 293736 86494
rect 293684 86430 293736 86436
rect 293788 77994 293816 96970
rect 293880 95742 293908 97106
rect 294064 97034 294092 100028
rect 294248 98705 294276 100028
rect 294234 98696 294290 98705
rect 294234 98631 294290 98640
rect 294052 97028 294104 97034
rect 294052 96970 294104 96976
rect 294432 96966 294460 100028
rect 294630 100014 294736 100042
rect 294420 96960 294472 96966
rect 294420 96902 294472 96908
rect 293868 95736 293920 95742
rect 293868 95678 293920 95684
rect 294708 93854 294736 100014
rect 294800 96898 294828 100028
rect 294984 100014 295090 100042
rect 295168 100014 295274 100042
rect 294880 96960 294932 96966
rect 294880 96902 294932 96908
rect 294788 96892 294840 96898
rect 294788 96834 294840 96840
rect 294708 93826 294828 93854
rect 293776 77988 293828 77994
rect 293776 77930 293828 77936
rect 293500 15904 293552 15910
rect 293500 15846 293552 15852
rect 292028 10328 292080 10334
rect 292028 10270 292080 10276
rect 294800 4826 294828 93826
rect 294892 89010 294920 96902
rect 294880 89004 294932 89010
rect 294880 88946 294932 88952
rect 294984 86426 295012 100014
rect 295064 97028 295116 97034
rect 295064 96970 295116 96976
rect 294972 86420 295024 86426
rect 294972 86362 295024 86368
rect 295076 76566 295104 96970
rect 295064 76560 295116 76566
rect 295064 76502 295116 76508
rect 295168 25566 295196 100014
rect 295444 96966 295472 100028
rect 295432 96960 295484 96966
rect 295432 96902 295484 96908
rect 295248 96892 295300 96898
rect 295248 96834 295300 96840
rect 295260 93158 295288 96834
rect 295628 96830 295656 100028
rect 295812 96898 295840 100028
rect 295800 96892 295852 96898
rect 295800 96834 295852 96840
rect 295616 96824 295668 96830
rect 295616 96766 295668 96772
rect 296088 94625 296116 100028
rect 296286 100014 296392 100042
rect 296260 97164 296312 97170
rect 296260 97106 296312 97112
rect 296074 94616 296130 94625
rect 296074 94551 296130 94560
rect 295248 93152 295300 93158
rect 295248 93094 295300 93100
rect 295340 86284 295392 86290
rect 295340 86226 295392 86232
rect 295156 25560 295208 25566
rect 295156 25502 295208 25508
rect 294788 4820 294840 4826
rect 294788 4762 294840 4768
rect 292580 3868 292632 3874
rect 292580 3810 292632 3816
rect 291844 3324 291896 3330
rect 291844 3266 291896 3272
rect 292592 480 292620 3810
rect 295352 3398 295380 86226
rect 296272 19990 296300 97106
rect 296364 96948 296392 100014
rect 296456 97170 296484 100028
rect 296444 97164 296496 97170
rect 296444 97106 296496 97112
rect 296364 96920 296484 96948
rect 296352 96824 296404 96830
rect 296352 96766 296404 96772
rect 296364 86358 296392 96766
rect 296352 86352 296404 86358
rect 296352 86294 296404 86300
rect 296456 84930 296484 96920
rect 296536 96892 296588 96898
rect 296536 96834 296588 96840
rect 296444 84924 296496 84930
rect 296444 84866 296496 84872
rect 296548 75274 296576 96834
rect 296640 93226 296668 100028
rect 296824 96937 296852 100028
rect 297114 100014 297220 100042
rect 296810 96928 296866 96937
rect 296810 96863 296866 96872
rect 296628 93220 296680 93226
rect 296628 93162 296680 93168
rect 297192 90370 297220 100014
rect 297284 96801 297312 100028
rect 297482 100014 297588 100042
rect 297666 100014 297772 100042
rect 297454 97200 297510 97209
rect 297454 97135 297510 97144
rect 297270 96792 297326 96801
rect 297270 96727 297326 96736
rect 297468 96150 297496 97135
rect 297560 96642 297588 100014
rect 297744 96948 297772 100014
rect 297836 98977 297864 100028
rect 297822 98968 297878 98977
rect 297822 98903 297878 98912
rect 297744 96920 298048 96948
rect 297560 96614 297956 96642
rect 297456 96144 297508 96150
rect 297456 96086 297508 96092
rect 297180 90364 297232 90370
rect 297180 90306 297232 90312
rect 297928 87650 297956 96614
rect 297916 87644 297968 87650
rect 297916 87586 297968 87592
rect 298020 82142 298048 96920
rect 298112 96898 298140 100028
rect 298100 96892 298152 96898
rect 298100 96834 298152 96840
rect 298296 96694 298324 100028
rect 298480 96966 298508 100028
rect 298678 100014 298784 100042
rect 298862 100014 299060 100042
rect 298756 97050 298784 100014
rect 299032 97152 299060 100014
rect 299124 97345 299152 100028
rect 299322 100014 299428 100042
rect 299624 100036 299690 100042
rect 299572 100030 299690 100036
rect 299110 97336 299166 97345
rect 299110 97271 299166 97280
rect 299032 97124 299336 97152
rect 298756 97022 299152 97050
rect 298376 96960 298428 96966
rect 298376 96902 298428 96908
rect 298468 96960 298520 96966
rect 298468 96902 298520 96908
rect 299020 96960 299072 96966
rect 299020 96902 299072 96908
rect 298284 96688 298336 96694
rect 298284 96630 298336 96636
rect 298388 95849 298416 96902
rect 298374 95840 298430 95849
rect 298374 95775 298430 95784
rect 299032 93129 299060 96902
rect 299018 93120 299074 93129
rect 299018 93055 299074 93064
rect 299124 86290 299152 97022
rect 299204 96688 299256 96694
rect 299204 96630 299256 96636
rect 299112 86284 299164 86290
rect 299112 86226 299164 86232
rect 298008 82136 298060 82142
rect 298008 82078 298060 82084
rect 299216 80714 299244 96630
rect 299204 80708 299256 80714
rect 299204 80650 299256 80656
rect 296536 75268 296588 75274
rect 296536 75210 296588 75216
rect 299308 75206 299336 97124
rect 298100 75200 298152 75206
rect 298100 75142 298152 75148
rect 299296 75200 299348 75206
rect 299296 75142 299348 75148
rect 296260 19984 296312 19990
rect 296260 19926 296312 19932
rect 297272 5024 297324 5030
rect 297272 4966 297324 4972
rect 296076 3800 296128 3806
rect 296076 3742 296128 3748
rect 293684 3392 293736 3398
rect 293684 3334 293736 3340
rect 295340 3392 295392 3398
rect 295340 3334 295392 3340
rect 293696 480 293724 3334
rect 294880 3324 294932 3330
rect 294880 3266 294932 3272
rect 294892 480 294920 3266
rect 296088 480 296116 3742
rect 297284 480 297312 4966
rect 298112 490 298140 75142
rect 299400 73846 299428 100014
rect 299492 97345 299520 100028
rect 299584 100014 299690 100030
rect 300306 97608 300362 97617
rect 300306 97543 300362 97552
rect 299478 97336 299534 97345
rect 299478 97271 299534 97280
rect 300122 96928 300178 96937
rect 300122 96863 300178 96872
rect 299572 95804 299624 95810
rect 299572 95746 299624 95752
rect 299480 84856 299532 84862
rect 299480 84798 299532 84804
rect 299388 73840 299440 73846
rect 299388 73782 299440 73788
rect 299492 3602 299520 84798
rect 299584 3806 299612 95746
rect 300136 84998 300164 96863
rect 300320 87922 300348 97543
rect 304356 97096 304408 97102
rect 304356 97038 304408 97044
rect 301504 96892 301556 96898
rect 301504 96834 301556 96840
rect 300766 96792 300822 96801
rect 300766 96727 300822 96736
rect 300780 94489 300808 96727
rect 300766 94480 300822 94489
rect 300766 94415 300822 94424
rect 300308 87916 300360 87922
rect 300308 87858 300360 87864
rect 300124 84992 300176 84998
rect 300124 84934 300176 84940
rect 301516 84862 301544 96834
rect 302332 96620 302384 96626
rect 302332 96562 302384 96568
rect 302240 95872 302292 95878
rect 302240 95814 302292 95820
rect 301504 84856 301556 84862
rect 301504 84798 301556 84804
rect 300860 22772 300912 22778
rect 300860 22714 300912 22720
rect 300872 16574 300900 22714
rect 300872 16546 301544 16574
rect 299572 3800 299624 3806
rect 299572 3742 299624 3748
rect 299388 3596 299440 3602
rect 299388 3538 299440 3544
rect 299480 3596 299532 3602
rect 299480 3538 299532 3544
rect 300768 3596 300820 3602
rect 300768 3538 300820 3544
rect 299400 3398 299428 3538
rect 299388 3392 299440 3398
rect 299388 3334 299440 3340
rect 299664 3188 299716 3194
rect 299664 3130 299716 3136
rect 298296 598 298508 626
rect 298296 490 298324 598
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298112 462 298324 490
rect 298480 480 298508 598
rect 299676 480 299704 3130
rect 300780 480 300808 3538
rect 301516 490 301544 16546
rect 302252 3074 302280 95814
rect 302344 3194 302372 96562
rect 304264 94308 304316 94314
rect 304264 94250 304316 94256
rect 303620 92268 303672 92274
rect 303620 92210 303672 92216
rect 303632 16574 303660 92210
rect 303632 16546 303936 16574
rect 302332 3188 302384 3194
rect 302332 3130 302384 3136
rect 302252 3046 303200 3074
rect 301792 598 302004 626
rect 301792 490 301820 598
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301516 462 301820 490
rect 301976 480 302004 598
rect 303172 480 303200 3046
rect 303908 490 303936 16546
rect 304276 3942 304304 94250
rect 304368 92274 304396 97038
rect 304356 92268 304408 92274
rect 304356 92210 304408 92216
rect 305656 73166 305684 300154
rect 307036 113150 307064 301446
rect 309796 156670 309824 302806
rect 311176 228410 311204 302874
rect 318064 302728 318116 302734
rect 318064 302670 318116 302676
rect 313924 302660 313976 302666
rect 313924 302602 313976 302608
rect 312544 298240 312596 298246
rect 312544 298182 312596 298188
rect 312556 233238 312584 298182
rect 312544 233232 312596 233238
rect 312544 233174 312596 233180
rect 311164 228404 311216 228410
rect 311164 228346 311216 228352
rect 309784 156664 309836 156670
rect 309784 156606 309836 156612
rect 307024 113144 307076 113150
rect 307024 113086 307076 113092
rect 311164 99272 311216 99278
rect 311164 99214 311216 99220
rect 309140 99204 309192 99210
rect 309140 99146 309192 99152
rect 306380 94376 306432 94382
rect 306380 94318 306432 94324
rect 305644 73160 305696 73166
rect 305644 73102 305696 73108
rect 304264 3936 304316 3942
rect 304264 3878 304316 3884
rect 305552 3392 305604 3398
rect 305552 3334 305604 3340
rect 304184 598 304396 626
rect 304184 490 304212 598
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 303908 462 304212 490
rect 304368 480 304396 598
rect 305564 480 305592 3334
rect 306392 490 306420 94318
rect 307024 92948 307076 92954
rect 307024 92890 307076 92896
rect 307036 3602 307064 92890
rect 309152 3602 309180 99146
rect 309232 90228 309284 90234
rect 309232 90170 309284 90176
rect 307024 3596 307076 3602
rect 307024 3538 307076 3544
rect 307944 3596 307996 3602
rect 307944 3538 307996 3544
rect 309140 3596 309192 3602
rect 309140 3538 309192 3544
rect 306576 598 306788 626
rect 306576 490 306604 598
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306392 462 306604 490
rect 306760 480 306788 598
rect 307956 480 307984 3538
rect 309244 3482 309272 90170
rect 310520 88936 310572 88942
rect 310520 88878 310572 88884
rect 310532 16574 310560 88878
rect 310532 16546 311112 16574
rect 310244 3596 310296 3602
rect 310244 3538 310296 3544
rect 309060 3454 309272 3482
rect 309060 480 309088 3454
rect 310256 480 310284 3538
rect 311084 3482 311112 16546
rect 311176 3874 311204 99214
rect 312544 99136 312596 99142
rect 312544 99078 312596 99084
rect 311900 24132 311952 24138
rect 311900 24074 311952 24080
rect 311912 16574 311940 24074
rect 311912 16546 312216 16574
rect 311164 3868 311216 3874
rect 311164 3810 311216 3816
rect 311084 3454 311480 3482
rect 311452 480 311480 3454
rect 312188 490 312216 16546
rect 312556 3602 312584 99078
rect 312636 97232 312688 97238
rect 312636 97174 312688 97180
rect 312648 24138 312676 97174
rect 313936 60722 313964 302602
rect 316684 302592 316736 302598
rect 316684 302534 316736 302540
rect 316696 100706 316724 302534
rect 318076 179382 318104 302670
rect 323584 298376 323636 298382
rect 323584 298318 323636 298324
rect 322204 295384 322256 295390
rect 322204 295326 322256 295332
rect 320824 288448 320876 288454
rect 320824 288390 320876 288396
rect 318064 179376 318116 179382
rect 318064 179318 318116 179324
rect 320836 122738 320864 288390
rect 322216 122806 322244 295326
rect 323596 267714 323624 298318
rect 359464 298308 359516 298314
rect 359464 298250 359516 298256
rect 327724 295928 327776 295934
rect 327724 295870 327776 295876
rect 324964 285728 325016 285734
rect 324964 285670 325016 285676
rect 323584 267708 323636 267714
rect 323584 267650 323636 267656
rect 324976 266218 325004 285670
rect 327736 268394 327764 295870
rect 352564 295860 352616 295866
rect 352564 295802 352616 295808
rect 327724 268388 327776 268394
rect 327724 268330 327776 268336
rect 324964 266212 325016 266218
rect 324964 266154 325016 266160
rect 352576 264926 352604 295802
rect 353944 281580 353996 281586
rect 353944 281522 353996 281528
rect 353956 266257 353984 281522
rect 356704 278792 356756 278798
rect 356704 278734 356756 278740
rect 353942 266248 353998 266257
rect 353942 266183 353998 266192
rect 356716 266121 356744 278734
rect 359476 266354 359504 298250
rect 360212 276078 360240 340054
rect 362880 337793 362908 340068
rect 364904 337793 364932 340068
rect 362866 337784 362922 337793
rect 362866 337719 362922 337728
rect 364890 337784 364946 337793
rect 364890 337719 364946 337728
rect 366928 337414 366956 340068
rect 368966 340054 369072 340082
rect 366916 337408 366968 337414
rect 366916 337350 366968 337356
rect 369044 335374 369072 340054
rect 369032 335368 369084 335374
rect 369032 335310 369084 335316
rect 369136 278662 369164 344986
rect 369412 340218 369440 347375
rect 369858 345808 369914 345817
rect 369858 345743 369914 345752
rect 369228 340190 369440 340218
rect 369124 278656 369176 278662
rect 369124 278598 369176 278604
rect 369136 277394 369164 278598
rect 369044 277366 369164 277394
rect 360200 276072 360252 276078
rect 360200 276014 360252 276020
rect 360660 276072 360712 276078
rect 360660 276014 360712 276020
rect 360672 268138 360700 276014
rect 369044 268802 369072 277366
rect 369228 275398 369256 340190
rect 369308 335368 369360 335374
rect 369308 335310 369360 335316
rect 369216 275392 369268 275398
rect 369216 275334 369268 275340
rect 369032 268796 369084 268802
rect 369032 268738 369084 268744
rect 369320 268546 369348 335310
rect 369490 297392 369546 297401
rect 369490 297327 369546 297336
rect 369398 296848 369454 296857
rect 369504 296818 369532 297327
rect 369398 296783 369454 296792
rect 369492 296812 369544 296818
rect 369412 296750 369440 296783
rect 369492 296754 369544 296760
rect 369400 296744 369452 296750
rect 369400 296686 369452 296692
rect 369398 296304 369454 296313
rect 369398 296239 369454 296248
rect 369412 296002 369440 296239
rect 369400 295996 369452 296002
rect 369400 295938 369452 295944
rect 369398 295896 369454 295905
rect 369398 295831 369400 295840
rect 369452 295831 369454 295840
rect 369400 295802 369452 295808
rect 369490 279032 369546 279041
rect 369490 278967 369546 278976
rect 369400 278656 369452 278662
rect 369398 278624 369400 278633
rect 369452 278624 369454 278633
rect 369398 278559 369454 278568
rect 369412 275398 369440 275429
rect 369400 275392 369452 275398
rect 369398 275360 369400 275369
rect 369452 275360 369454 275369
rect 369398 275295 369454 275304
rect 369044 268518 369348 268546
rect 369044 268138 369072 268518
rect 369124 268456 369176 268462
rect 369412 268410 369440 275295
rect 369124 268398 369176 268404
rect 360672 268124 360962 268138
rect 360672 268110 360976 268124
rect 359464 266348 359516 266354
rect 359464 266290 359516 266296
rect 356702 266112 356758 266121
rect 356702 266047 356758 266056
rect 360948 265742 360976 268110
rect 362880 266286 362908 268124
rect 362868 266280 362920 266286
rect 362868 266222 362920 266228
rect 362880 266121 362908 266222
rect 364904 266218 364932 268124
rect 366928 266354 366956 268124
rect 368492 268110 369072 268138
rect 366916 266348 366968 266354
rect 366916 266290 366968 266296
rect 364892 266212 364944 266218
rect 364892 266154 364944 266160
rect 364904 266121 364932 266154
rect 368492 266150 368520 268110
rect 368480 266144 368532 266150
rect 362866 266112 362922 266121
rect 362866 266047 362922 266056
rect 364890 266112 364946 266121
rect 368480 266086 368532 266092
rect 364890 266047 364946 266056
rect 360200 265736 360252 265742
rect 360200 265678 360252 265684
rect 360936 265736 360988 265742
rect 360936 265678 360988 265684
rect 352564 264920 352616 264926
rect 352564 264862 352616 264868
rect 359464 253972 359516 253978
rect 359464 253914 359516 253920
rect 359372 225208 359424 225214
rect 359372 225150 359424 225156
rect 359384 223582 359412 225150
rect 359476 224466 359504 253914
rect 359648 225344 359700 225350
rect 359648 225286 359700 225292
rect 359556 225140 359608 225146
rect 359556 225082 359608 225088
rect 359464 224460 359516 224466
rect 359464 224402 359516 224408
rect 359464 223916 359516 223922
rect 359464 223858 359516 223864
rect 359372 223576 359424 223582
rect 359372 223518 359424 223524
rect 359476 220794 359504 223858
rect 359464 220788 359516 220794
rect 359464 220730 359516 220736
rect 359568 211138 359596 225082
rect 359660 215286 359688 225286
rect 359740 223984 359792 223990
rect 359740 223926 359792 223932
rect 359752 218006 359780 223926
rect 359740 218000 359792 218006
rect 359740 217942 359792 217948
rect 359648 215280 359700 215286
rect 359648 215222 359700 215228
rect 359556 211132 359608 211138
rect 359556 211074 359608 211080
rect 360212 209774 360240 265678
rect 368492 265674 368520 266086
rect 368480 265668 368532 265674
rect 368480 265610 368532 265616
rect 360212 209746 360608 209774
rect 359464 207052 359516 207058
rect 359464 206994 359516 207000
rect 359476 197130 359504 206994
rect 359556 204332 359608 204338
rect 359556 204274 359608 204280
rect 359464 197124 359516 197130
rect 359464 197066 359516 197072
rect 359568 197062 359596 204274
rect 360108 201544 360160 201550
rect 360108 201486 360160 201492
rect 360120 197266 360148 201486
rect 360108 197260 360160 197266
rect 360108 197202 360160 197208
rect 359556 197056 359608 197062
rect 359556 196998 359608 197004
rect 360580 196058 360608 209746
rect 369136 206174 369164 268398
rect 369228 268382 369440 268410
rect 369228 206394 369256 268382
rect 369308 265668 369360 265674
rect 369308 265610 369360 265616
rect 369320 206514 369348 265610
rect 369400 224460 369452 224466
rect 369400 224402 369452 224408
rect 369412 222873 369440 224402
rect 369398 222864 369454 222873
rect 369398 222799 369454 222808
rect 369504 209774 369532 278967
rect 369872 274281 369900 345743
rect 370226 345536 370282 345545
rect 370226 345471 370282 345480
rect 370240 345014 370268 345471
rect 370056 344986 370268 345014
rect 369952 340604 370004 340610
rect 369952 340546 370004 340552
rect 369858 274272 369914 274281
rect 369858 274207 369914 274216
rect 369964 268977 369992 340546
rect 370056 273329 370084 344986
rect 370134 340640 370190 340649
rect 370134 340575 370136 340584
rect 370188 340575 370190 340584
rect 370136 340546 370188 340552
rect 370226 340232 370282 340241
rect 370226 340167 370282 340176
rect 370136 296132 370188 296138
rect 370136 296074 370188 296080
rect 370148 295633 370176 296074
rect 370134 295624 370190 295633
rect 370134 295559 370190 295568
rect 370042 273320 370098 273329
rect 370042 273255 370098 273264
rect 369950 268968 370006 268977
rect 369950 268903 370006 268912
rect 369584 231124 369636 231130
rect 369584 231066 369636 231072
rect 369596 220697 369624 231066
rect 369860 225616 369912 225622
rect 369860 225558 369912 225564
rect 369872 220794 369900 225558
rect 369952 224392 370004 224398
rect 369952 224334 370004 224340
rect 369860 220788 369912 220794
rect 369860 220730 369912 220736
rect 369872 220697 369900 220730
rect 369582 220688 369638 220697
rect 369582 220623 369638 220632
rect 369858 220688 369914 220697
rect 369858 220623 369914 220632
rect 369964 218521 369992 224334
rect 369950 218512 370006 218521
rect 369950 218447 370006 218456
rect 369504 209746 369624 209774
rect 369596 206553 369624 209746
rect 369688 208758 369716 208789
rect 369676 208752 369728 208758
rect 369674 208720 369676 208729
rect 369728 208720 369730 208729
rect 369674 208655 369730 208664
rect 369582 206544 369638 206553
rect 369308 206508 369360 206514
rect 369582 206479 369638 206488
rect 369308 206450 369360 206456
rect 369228 206366 369532 206394
rect 369216 206304 369268 206310
rect 369216 206246 369268 206252
rect 369124 206168 369176 206174
rect 369124 206110 369176 206116
rect 369228 196330 369256 206246
rect 369412 206174 369440 206205
rect 369400 206168 369452 206174
rect 369398 206136 369400 206145
rect 369452 206136 369454 206145
rect 369398 206071 369454 206080
rect 369412 200114 369440 206071
rect 369504 204105 369532 206366
rect 369490 204096 369546 204105
rect 369596 204066 369624 206479
rect 369490 204031 369546 204040
rect 369584 204060 369636 204066
rect 369584 204002 369636 204008
rect 369688 203946 369716 208655
rect 369766 207088 369822 207097
rect 369766 207023 369822 207032
rect 369780 206990 369808 207023
rect 369768 206984 369820 206990
rect 369768 206926 369820 206932
rect 369044 196302 369256 196330
rect 369320 200086 369440 200114
rect 369504 203918 369716 203946
rect 364522 196072 364578 196081
rect 360580 196030 360962 196058
rect 360580 180794 360608 196030
rect 362880 194585 362908 196044
rect 369044 196058 369072 196302
rect 364578 196044 364918 196058
rect 364578 196030 364932 196044
rect 364522 196007 364578 196016
rect 364904 194585 364932 196030
rect 362866 194576 362922 194585
rect 362866 194511 362922 194520
rect 364890 194576 364946 194585
rect 366928 194546 366956 196044
rect 368966 196030 369072 196058
rect 364890 194511 364946 194520
rect 366916 194540 366968 194546
rect 366916 194482 366968 194488
rect 360212 180766 360608 180794
rect 359464 152176 359516 152182
rect 359464 152118 359516 152124
rect 358912 152108 358964 152114
rect 358912 152050 358964 152056
rect 358924 146266 358952 152050
rect 358912 146260 358964 146266
rect 358912 146202 358964 146208
rect 359476 139398 359504 152118
rect 360108 152040 360160 152046
rect 360108 151982 360160 151988
rect 359556 151972 359608 151978
rect 359556 151914 359608 151920
rect 359568 142118 359596 151914
rect 360120 149054 360148 151982
rect 360108 149048 360160 149054
rect 360108 148990 360160 148996
rect 359556 142112 359608 142118
rect 359556 142054 359608 142060
rect 359464 139392 359516 139398
rect 359464 139334 359516 139340
rect 360212 132494 360240 180766
rect 360212 132466 360608 132494
rect 359464 124908 359516 124914
rect 359464 124850 359516 124856
rect 322204 122800 322256 122806
rect 322204 122742 322256 122748
rect 320824 122732 320876 122738
rect 320824 122674 320876 122680
rect 359476 109002 359504 124850
rect 360580 124794 360608 132466
rect 369044 124794 369072 196030
rect 369320 180794 369348 200086
rect 369504 196042 369532 203918
rect 369584 203856 369636 203862
rect 369584 203798 369636 203804
rect 369492 196036 369544 196042
rect 369492 195978 369544 195984
rect 369136 180766 369348 180794
rect 369136 167958 369164 180766
rect 369124 167952 369176 167958
rect 369124 167894 369176 167900
rect 369308 167000 369360 167006
rect 369308 166942 369360 166948
rect 369320 153202 369348 166942
rect 369400 158704 369452 158710
rect 369400 158646 369452 158652
rect 369308 153196 369360 153202
rect 369308 153138 369360 153144
rect 369306 152960 369362 152969
rect 369306 152895 369362 152904
rect 369320 152862 369348 152895
rect 369308 152856 369360 152862
rect 369308 152798 369360 152804
rect 369124 152176 369176 152182
rect 369124 152118 369176 152124
rect 369136 130914 369164 152118
rect 369216 152108 369268 152114
rect 369216 152050 369268 152056
rect 369228 132002 369256 152050
rect 369412 152046 369440 158646
rect 369400 152040 369452 152046
rect 369400 151982 369452 151988
rect 369412 132433 369440 151982
rect 369504 136649 369532 195978
rect 369596 155922 369624 203798
rect 369676 171148 369728 171154
rect 369676 171090 369728 171096
rect 369584 155916 369636 155922
rect 369584 155858 369636 155864
rect 369584 153196 369636 153202
rect 369584 153138 369636 153144
rect 369596 151978 369624 153138
rect 369688 152930 369716 171090
rect 369780 161430 369808 206926
rect 370056 201929 370084 273255
rect 370148 262206 370176 295559
rect 370240 268297 370268 340167
rect 370332 276865 370360 348735
rect 370410 347168 370466 347177
rect 370410 347103 370466 347112
rect 370318 276856 370374 276865
rect 370318 276791 370374 276800
rect 370332 274718 370360 276791
rect 370424 275233 370452 347103
rect 371528 345014 371556 353495
rect 371712 353326 371740 354039
rect 371988 354006 372016 358935
rect 371976 354000 372028 354006
rect 371976 353942 372028 353948
rect 371700 353320 371752 353326
rect 371700 353262 371752 353268
rect 371974 353016 372030 353025
rect 371974 352951 372030 352960
rect 371606 349344 371662 349353
rect 371606 349279 371608 349288
rect 371660 349279 371662 349288
rect 371608 349250 371660 349256
rect 371606 348256 371662 348265
rect 371606 348191 371608 348200
rect 371660 348191 371662 348200
rect 371608 348162 371660 348168
rect 371528 344986 371648 345014
rect 371422 344448 371478 344457
rect 371422 344383 371478 344392
rect 371330 342272 371386 342281
rect 371330 342207 371386 342216
rect 371240 295316 371292 295322
rect 371240 295258 371292 295264
rect 371252 294001 371280 295258
rect 371238 293992 371294 294001
rect 371238 293927 371294 293936
rect 371240 292460 371292 292466
rect 371240 292402 371292 292408
rect 371252 291825 371280 292402
rect 371238 291816 371294 291825
rect 371238 291751 371294 291760
rect 371240 290556 371292 290562
rect 371240 290498 371292 290504
rect 371252 290193 371280 290498
rect 371238 290184 371294 290193
rect 371238 290119 371294 290128
rect 371238 287056 371294 287065
rect 371238 286991 371294 287000
rect 371252 286346 371280 286991
rect 371240 286340 371292 286346
rect 371240 286282 371292 286288
rect 371238 281616 371294 281625
rect 371238 281551 371294 281560
rect 370410 275224 370466 275233
rect 370410 275159 370466 275168
rect 370320 274712 370372 274718
rect 370320 274654 370372 274660
rect 370594 274136 370650 274145
rect 370594 274071 370650 274080
rect 370226 268288 370282 268297
rect 370226 268223 370282 268232
rect 370136 262200 370188 262206
rect 370136 262142 370188 262148
rect 370504 256760 370556 256766
rect 370504 256702 370556 256708
rect 370228 249756 370280 249762
rect 370228 249698 370280 249704
rect 370240 248470 370268 249698
rect 370228 248464 370280 248470
rect 370228 248406 370280 248412
rect 370240 229094 370268 248406
rect 370320 239420 370372 239426
rect 370320 239362 370372 239368
rect 370148 229066 370268 229094
rect 370148 221474 370176 229066
rect 370228 224324 370280 224330
rect 370228 224266 370280 224272
rect 370136 221468 370188 221474
rect 370136 221410 370188 221416
rect 370148 221377 370176 221410
rect 370134 221368 370190 221377
rect 370134 221303 370190 221312
rect 370240 218006 370268 224266
rect 370332 221921 370360 239362
rect 370412 224256 370464 224262
rect 370412 224198 370464 224204
rect 370318 221912 370374 221921
rect 370318 221847 370374 221856
rect 370424 219201 370452 224198
rect 370516 223009 370544 256702
rect 370502 223000 370558 223009
rect 370502 222935 370558 222944
rect 370410 219192 370466 219201
rect 370410 219127 370466 219136
rect 370424 218754 370452 219127
rect 370412 218748 370464 218754
rect 370412 218690 370464 218696
rect 370228 218000 370280 218006
rect 370228 217942 370280 217948
rect 370240 217569 370268 217942
rect 370226 217560 370282 217569
rect 370226 217495 370282 217504
rect 370410 211712 370466 211721
rect 370410 211647 370466 211656
rect 370424 211206 370452 211647
rect 370412 211200 370464 211206
rect 370412 211142 370464 211148
rect 370318 209536 370374 209545
rect 370318 209471 370374 209480
rect 370134 208992 370190 209001
rect 370134 208927 370190 208936
rect 370042 201920 370098 201929
rect 370042 201855 370098 201864
rect 370056 201618 370084 201855
rect 370044 201612 370096 201618
rect 370044 201554 370096 201560
rect 370148 175982 370176 208927
rect 370226 202056 370282 202065
rect 370226 201991 370282 202000
rect 370136 175976 370188 175982
rect 370136 175918 370188 175924
rect 370044 168360 370096 168366
rect 370044 168302 370096 168308
rect 370056 167958 370084 168302
rect 370044 167952 370096 167958
rect 370044 167894 370096 167900
rect 369768 161424 369820 161430
rect 369768 161366 369820 161372
rect 370056 153066 370084 167894
rect 370240 164218 370268 201991
rect 370332 180130 370360 209471
rect 370424 193186 370452 211142
rect 370502 203144 370558 203153
rect 370502 203079 370558 203088
rect 370412 193180 370464 193186
rect 370412 193122 370464 193128
rect 370320 180124 370372 180130
rect 370320 180066 370372 180072
rect 370228 164212 370280 164218
rect 370228 164154 370280 164160
rect 370228 161424 370280 161430
rect 370228 161366 370280 161372
rect 370240 153270 370268 161366
rect 370228 153264 370280 153270
rect 370228 153206 370280 153212
rect 370136 153196 370188 153202
rect 370136 153138 370188 153144
rect 370044 153060 370096 153066
rect 370044 153002 370096 153008
rect 369676 152924 369728 152930
rect 369676 152866 369728 152872
rect 369584 151972 369636 151978
rect 369584 151914 369636 151920
rect 369490 136640 369546 136649
rect 369490 136575 369546 136584
rect 369398 132424 369454 132433
rect 369398 132359 369454 132368
rect 369306 132016 369362 132025
rect 369228 131974 369306 132002
rect 369306 131951 369362 131960
rect 369596 131481 369624 151914
rect 369688 151814 369716 152866
rect 369688 151786 369900 151814
rect 369872 133657 369900 151786
rect 370056 142154 370084 153002
rect 370148 151910 370176 153138
rect 370136 151904 370188 151910
rect 370136 151846 370188 151852
rect 369964 142126 370084 142154
rect 369964 134609 369992 142126
rect 369950 134600 370006 134609
rect 369950 134535 370006 134544
rect 369858 133648 369914 133657
rect 369858 133583 369914 133592
rect 370148 132841 370176 151846
rect 370240 135425 370268 153206
rect 370332 137601 370360 180066
rect 370516 167006 370544 203079
rect 370608 202065 370636 274071
rect 370686 268288 370742 268297
rect 370686 268223 370742 268232
rect 370594 202056 370650 202065
rect 370594 201991 370650 202000
rect 370700 196217 370728 268223
rect 371252 225078 371280 281551
rect 371344 270337 371372 342207
rect 371436 272513 371464 344383
rect 371514 342816 371570 342825
rect 371514 342751 371570 342760
rect 371422 272504 371478 272513
rect 371422 272439 371478 272448
rect 371528 270881 371556 342751
rect 371620 286550 371648 344986
rect 371882 344992 371938 345001
rect 371882 344927 371938 344936
rect 371790 341728 371846 341737
rect 371790 341663 371846 341672
rect 371698 295080 371754 295089
rect 371698 295015 371754 295024
rect 371712 294642 371740 295015
rect 371700 294636 371752 294642
rect 371700 294578 371752 294584
rect 371698 294536 371754 294545
rect 371698 294471 371754 294480
rect 371712 294030 371740 294471
rect 371700 294024 371752 294030
rect 371700 293966 371752 293972
rect 371700 293276 371752 293282
rect 371700 293218 371752 293224
rect 371712 292913 371740 293218
rect 371698 292904 371754 292913
rect 371698 292839 371754 292848
rect 371700 292392 371752 292398
rect 371698 292360 371700 292369
rect 371752 292360 371754 292369
rect 371698 292295 371754 292304
rect 371698 290728 371754 290737
rect 371698 290663 371754 290672
rect 371712 290494 371740 290663
rect 371700 290488 371752 290494
rect 371700 290430 371752 290436
rect 371698 289640 371754 289649
rect 371698 289575 371700 289584
rect 371752 289575 371754 289584
rect 371700 289546 371752 289552
rect 371700 289128 371752 289134
rect 371698 289096 371700 289105
rect 371752 289096 371754 289105
rect 371698 289031 371754 289040
rect 371698 288552 371754 288561
rect 371698 288487 371700 288496
rect 371752 288487 371754 288496
rect 371700 288458 371752 288464
rect 371700 288380 371752 288386
rect 371700 288322 371752 288328
rect 371712 288153 371740 288322
rect 371698 288144 371754 288153
rect 371698 288079 371754 288088
rect 371700 287700 371752 287706
rect 371700 287642 371752 287648
rect 371712 287609 371740 287642
rect 371698 287600 371754 287609
rect 371698 287535 371754 287544
rect 371700 287020 371752 287026
rect 371700 286962 371752 286968
rect 371608 286544 371660 286550
rect 371712 286521 371740 286962
rect 371608 286486 371660 286492
rect 371698 286512 371754 286521
rect 371698 286447 371754 286456
rect 371608 286408 371660 286414
rect 371608 286350 371660 286356
rect 371620 285977 371648 286350
rect 371606 285968 371662 285977
rect 371606 285903 371662 285912
rect 371700 285660 371752 285666
rect 371700 285602 371752 285608
rect 371608 285524 371660 285530
rect 371608 285466 371660 285472
rect 371620 285433 371648 285466
rect 371606 285424 371662 285433
rect 371606 285359 371662 285368
rect 371606 284880 371662 284889
rect 371606 284815 371662 284824
rect 371620 284374 371648 284815
rect 371608 284368 371660 284374
rect 371712 284345 371740 285602
rect 371608 284310 371660 284316
rect 371698 284336 371754 284345
rect 371698 284271 371754 284280
rect 371606 283792 371662 283801
rect 371606 283727 371662 283736
rect 371620 283626 371648 283727
rect 371700 283688 371752 283694
rect 371700 283630 371752 283636
rect 371608 283620 371660 283626
rect 371608 283562 371660 283568
rect 371712 283257 371740 283630
rect 371698 283248 371754 283257
rect 371698 283183 371754 283192
rect 371608 282736 371660 282742
rect 371606 282704 371608 282713
rect 371660 282704 371662 282713
rect 371606 282639 371662 282648
rect 371608 282192 371660 282198
rect 371606 282160 371608 282169
rect 371660 282160 371662 282169
rect 371606 282095 371662 282104
rect 371606 281072 371662 281081
rect 371606 281007 371662 281016
rect 371514 270872 371570 270881
rect 371514 270807 371570 270816
rect 371330 270328 371386 270337
rect 371386 270286 371556 270314
rect 371330 270263 371386 270272
rect 371422 270192 371478 270201
rect 371422 270127 371478 270136
rect 371436 269249 371464 270127
rect 371422 269240 371478 269249
rect 371422 269175 371478 269184
rect 371240 225072 371292 225078
rect 371240 225014 371292 225020
rect 371330 224632 371386 224641
rect 371330 224567 371386 224576
rect 371344 224330 371372 224567
rect 371332 224324 371384 224330
rect 371332 224266 371384 224272
rect 371330 223000 371386 223009
rect 371330 222935 371386 222944
rect 371238 222456 371294 222465
rect 371238 222391 371240 222400
rect 371292 222391 371294 222400
rect 371240 222362 371292 222368
rect 371344 222290 371372 222935
rect 371332 222284 371384 222290
rect 371332 222226 371384 222232
rect 371238 221912 371294 221921
rect 371238 221847 371294 221856
rect 371252 220930 371280 221847
rect 371240 220924 371292 220930
rect 371240 220866 371292 220872
rect 371240 220720 371292 220726
rect 371240 220662 371292 220668
rect 371056 218136 371108 218142
rect 371054 218104 371056 218113
rect 371108 218104 371110 218113
rect 371054 218039 371110 218048
rect 371252 209545 371280 220662
rect 371330 216472 371386 216481
rect 371330 216407 371386 216416
rect 371344 216034 371372 216407
rect 371332 216028 371384 216034
rect 371332 215970 371384 215976
rect 371330 213888 371386 213897
rect 371330 213823 371386 213832
rect 371344 213314 371372 213823
rect 371332 213308 371384 213314
rect 371332 213250 371384 213256
rect 371332 213172 371384 213178
rect 371332 213114 371384 213120
rect 371238 209536 371294 209545
rect 371238 209471 371294 209480
rect 371344 209001 371372 213114
rect 371330 208992 371386 209001
rect 371330 208927 371386 208936
rect 371238 203688 371294 203697
rect 371238 203623 371294 203632
rect 371252 202502 371280 203623
rect 371240 202496 371292 202502
rect 371240 202438 371292 202444
rect 371436 200114 371464 269175
rect 371344 200086 371464 200114
rect 371238 198792 371294 198801
rect 371238 198727 371294 198736
rect 371252 196738 371280 198727
rect 371344 197169 371372 200086
rect 371528 198257 371556 270286
rect 371620 225758 371648 281007
rect 371698 277400 371754 277409
rect 371698 277335 371700 277344
rect 371752 277335 371754 277344
rect 371700 277306 371752 277312
rect 371698 276312 371754 276321
rect 371698 276247 371754 276256
rect 371712 276146 371740 276247
rect 371700 276140 371752 276146
rect 371700 276082 371752 276088
rect 371698 273048 371754 273057
rect 371698 272983 371754 272992
rect 371608 225752 371660 225758
rect 371608 225694 371660 225700
rect 371608 225616 371660 225622
rect 371608 225558 371660 225564
rect 371620 225185 371648 225558
rect 371606 225176 371662 225185
rect 371606 225111 371662 225120
rect 371608 224256 371660 224262
rect 371608 224198 371660 224204
rect 371620 224097 371648 224198
rect 371606 224088 371662 224097
rect 371606 224023 371662 224032
rect 371606 223544 371662 223553
rect 371606 223479 371662 223488
rect 371620 222902 371648 223479
rect 371608 222896 371660 222902
rect 371608 222838 371660 222844
rect 371608 222352 371660 222358
rect 371608 222294 371660 222300
rect 371620 217190 371648 222294
rect 371608 217184 371660 217190
rect 371608 217126 371660 217132
rect 371608 217048 371660 217054
rect 371606 217016 371608 217025
rect 371660 217016 371662 217025
rect 371606 216951 371662 216960
rect 371606 216064 371662 216073
rect 371606 215999 371662 216008
rect 371620 215966 371648 215999
rect 371608 215960 371660 215966
rect 371608 215902 371660 215908
rect 371608 215280 371660 215286
rect 371608 215222 371660 215228
rect 371620 214985 371648 215222
rect 371606 214976 371662 214985
rect 371606 214911 371662 214920
rect 371606 214432 371662 214441
rect 371606 214367 371662 214376
rect 371620 213994 371648 214367
rect 371608 213988 371660 213994
rect 371608 213930 371660 213936
rect 371606 213344 371662 213353
rect 371606 213279 371662 213288
rect 371620 213246 371648 213279
rect 371608 213240 371660 213246
rect 371608 213182 371660 213188
rect 371608 211268 371660 211274
rect 371608 211210 371660 211216
rect 371620 211177 371648 211210
rect 371606 211168 371662 211177
rect 371606 211103 371662 211112
rect 371608 210656 371660 210662
rect 371606 210624 371608 210633
rect 371660 210624 371662 210633
rect 371606 210559 371662 210568
rect 371606 205864 371662 205873
rect 371606 205799 371608 205808
rect 371660 205799 371662 205808
rect 371608 205770 371660 205776
rect 371608 205352 371660 205358
rect 371606 205320 371608 205329
rect 371660 205320 371662 205329
rect 371606 205255 371662 205264
rect 371608 204808 371660 204814
rect 371606 204776 371608 204785
rect 371660 204776 371662 204785
rect 371606 204711 371662 204720
rect 371608 204264 371660 204270
rect 371606 204232 371608 204241
rect 371660 204232 371662 204241
rect 371606 204167 371662 204176
rect 371712 200977 371740 272983
rect 371804 269793 371832 341663
rect 371896 273057 371924 344927
rect 371988 286686 372016 352951
rect 372172 352646 372200 359479
rect 372160 352640 372212 352646
rect 372160 352582 372212 352588
rect 372356 352578 372384 360023
rect 372632 354674 372660 363174
rect 372896 359508 372948 359514
rect 372896 359450 372948 359456
rect 372632 354646 372752 354674
rect 372344 352572 372396 352578
rect 372344 352514 372396 352520
rect 372434 351928 372490 351937
rect 372434 351863 372490 351872
rect 372066 343904 372122 343913
rect 372066 343839 372122 343848
rect 371976 286680 372028 286686
rect 371976 286622 372028 286628
rect 371976 286544 372028 286550
rect 371976 286486 372028 286492
rect 371988 281625 372016 286486
rect 371974 281616 372030 281625
rect 371974 281551 372030 281560
rect 371974 279440 372030 279449
rect 371974 279375 372030 279384
rect 371988 279002 372016 279375
rect 371976 278996 372028 279002
rect 371976 278938 372028 278944
rect 371882 273048 371938 273057
rect 371882 272983 371938 272992
rect 371974 272504 372030 272513
rect 371974 272439 372030 272448
rect 371882 270872 371938 270881
rect 371882 270807 371938 270816
rect 371790 269784 371846 269793
rect 371790 269719 371846 269728
rect 371698 200968 371754 200977
rect 371698 200903 371754 200912
rect 371606 198928 371662 198937
rect 371606 198863 371662 198872
rect 371514 198248 371570 198257
rect 371514 198183 371570 198192
rect 371330 197160 371386 197169
rect 371330 197095 371386 197104
rect 371160 196710 371280 196738
rect 370686 196208 370742 196217
rect 370686 196143 370742 196152
rect 370596 175228 370648 175234
rect 370596 175170 370648 175176
rect 370608 170406 370636 175170
rect 370596 170400 370648 170406
rect 370596 170342 370648 170348
rect 370504 167000 370556 167006
rect 370504 166942 370556 166948
rect 370608 166818 370636 170342
rect 370424 166790 370636 166818
rect 370318 137592 370374 137601
rect 370318 137527 370374 137536
rect 370424 135969 370452 166790
rect 370504 164212 370556 164218
rect 370504 164154 370556 164160
rect 370596 164212 370648 164218
rect 370596 164154 370648 164160
rect 370410 135960 370466 135969
rect 370410 135895 370466 135904
rect 370226 135416 370282 135425
rect 370226 135351 370282 135360
rect 370134 132832 370190 132841
rect 370134 132767 370190 132776
rect 369582 131472 369638 131481
rect 369582 131407 369638 131416
rect 369306 130928 369362 130937
rect 369136 130886 369306 130914
rect 369306 130863 369362 130872
rect 370516 130121 370544 164154
rect 370608 153202 370636 164154
rect 370596 153196 370648 153202
rect 370596 153138 370648 153144
rect 370502 130112 370558 130121
rect 370502 130047 370558 130056
rect 369950 129840 370006 129849
rect 369950 129775 370006 129784
rect 369860 129600 369912 129606
rect 369860 129542 369912 129548
rect 369872 129169 369900 129542
rect 369858 129160 369914 129169
rect 369858 129095 369914 129104
rect 369398 126440 369454 126449
rect 369398 126375 369454 126384
rect 369306 124944 369362 124953
rect 369306 124879 369308 124888
rect 369360 124879 369362 124888
rect 369308 124850 369360 124856
rect 360580 124766 360962 124794
rect 368966 124766 369072 124794
rect 362788 124086 362894 124114
rect 364918 124086 365208 124114
rect 362788 124001 362816 124086
rect 365180 124001 365208 124086
rect 362774 123992 362830 124001
rect 362774 123927 362830 123936
rect 365166 123992 365222 124001
rect 365166 123927 365222 123936
rect 366928 122738 366956 124100
rect 369412 124098 369440 126375
rect 369872 125186 369900 129095
rect 369860 125180 369912 125186
rect 369860 125122 369912 125128
rect 369964 125050 369992 129775
rect 370240 129062 370268 129093
rect 370228 129056 370280 129062
rect 370226 129024 370228 129033
rect 370280 129024 370282 129033
rect 370226 128959 370282 128968
rect 370042 128616 370098 128625
rect 370042 128551 370098 128560
rect 370056 125118 370084 128551
rect 370134 125760 370190 125769
rect 370134 125695 370190 125704
rect 370044 125112 370096 125118
rect 370044 125054 370096 125060
rect 369952 125044 370004 125050
rect 369952 124986 370004 124992
rect 369858 124400 369914 124409
rect 369858 124335 369914 124344
rect 367652 124092 367704 124098
rect 367652 124034 367704 124040
rect 369400 124092 369452 124098
rect 369400 124034 369452 124040
rect 366916 122732 366968 122738
rect 366916 122674 366968 122680
rect 367664 117298 367692 124034
rect 367652 117292 367704 117298
rect 367652 117234 367704 117240
rect 359464 108996 359516 109002
rect 359464 108938 359516 108944
rect 369872 102814 369900 124335
rect 370148 118694 370176 125695
rect 370240 125254 370268 128959
rect 370318 127392 370374 127401
rect 370318 127327 370374 127336
rect 370228 125248 370280 125254
rect 370228 125190 370280 125196
rect 370226 124672 370282 124681
rect 370226 124607 370282 124616
rect 370240 123486 370268 124607
rect 370228 123480 370280 123486
rect 370228 123422 370280 123428
rect 370332 121446 370360 127327
rect 370410 126304 370466 126313
rect 370410 126239 370466 126248
rect 370424 123622 370452 126239
rect 370700 124273 370728 196143
rect 371160 195786 371188 196710
rect 371238 196616 371294 196625
rect 371238 196551 371294 196560
rect 371252 195974 371280 196551
rect 371240 195968 371292 195974
rect 371240 195910 371292 195916
rect 371160 195758 371280 195786
rect 370780 175976 370832 175982
rect 370780 175918 370832 175924
rect 370792 137057 370820 175918
rect 370872 155916 370924 155922
rect 370872 155858 370924 155864
rect 370884 153338 370912 155858
rect 370872 153332 370924 153338
rect 370872 153274 370924 153280
rect 370778 137048 370834 137057
rect 370778 136983 370834 136992
rect 370884 134881 370912 153274
rect 370870 134872 370926 134881
rect 370870 134807 370926 134816
rect 371252 126449 371280 195758
rect 371238 126440 371294 126449
rect 371238 126375 371294 126384
rect 371252 126070 371280 126375
rect 371240 126064 371292 126070
rect 371240 126006 371292 126012
rect 371240 125520 371292 125526
rect 371240 125462 371292 125468
rect 371252 124681 371280 125462
rect 371344 125225 371372 197095
rect 371424 154488 371476 154494
rect 371424 154430 371476 154436
rect 371436 153785 371464 154430
rect 371422 153776 371478 153785
rect 371422 153711 371478 153720
rect 371424 153128 371476 153134
rect 371424 153070 371476 153076
rect 371436 152697 371464 153070
rect 371422 152688 371478 152697
rect 371422 152623 371478 152632
rect 371424 151768 371476 151774
rect 371424 151710 371476 151716
rect 371436 151609 371464 151710
rect 371422 151600 371478 151609
rect 371422 151535 371478 151544
rect 371424 150952 371476 150958
rect 371424 150894 371476 150900
rect 371436 150521 371464 150894
rect 371422 150512 371478 150521
rect 371422 150447 371478 150456
rect 371424 150340 371476 150346
rect 371424 150282 371476 150288
rect 371436 149977 371464 150282
rect 371422 149968 371478 149977
rect 371422 149903 371478 149912
rect 371424 148980 371476 148986
rect 371424 148922 371476 148928
rect 371436 148889 371464 148922
rect 371422 148880 371478 148889
rect 371422 148815 371478 148824
rect 371424 147552 371476 147558
rect 371424 147494 371476 147500
rect 371436 147257 371464 147494
rect 371422 147248 371478 147257
rect 371422 147183 371478 147192
rect 371424 146192 371476 146198
rect 371422 146160 371424 146169
rect 371476 146160 371478 146169
rect 371422 146095 371478 146104
rect 371424 145920 371476 145926
rect 371424 145862 371476 145868
rect 371436 145081 371464 145862
rect 371422 145072 371478 145081
rect 371422 145007 371478 145016
rect 371424 144764 371476 144770
rect 371424 144706 371476 144712
rect 371436 144537 371464 144706
rect 371422 144528 371478 144537
rect 371422 144463 371478 144472
rect 371424 144288 371476 144294
rect 371424 144230 371476 144236
rect 371436 144129 371464 144230
rect 371422 144120 371478 144129
rect 371422 144055 371478 144064
rect 371424 143948 371476 143954
rect 371424 143890 371476 143896
rect 371436 143585 371464 143890
rect 371422 143576 371478 143585
rect 371422 143511 371478 143520
rect 371424 143472 371476 143478
rect 371424 143414 371476 143420
rect 371436 142497 371464 143414
rect 371422 142488 371478 142497
rect 371422 142423 371478 142432
rect 371424 141976 371476 141982
rect 371422 141944 371424 141953
rect 371476 141944 371478 141953
rect 371422 141879 371478 141888
rect 371424 140684 371476 140690
rect 371424 140626 371476 140632
rect 371436 139777 371464 140626
rect 371422 139768 371478 139777
rect 371422 139703 371478 139712
rect 371424 139392 371476 139398
rect 371424 139334 371476 139340
rect 371436 139233 371464 139334
rect 371422 139224 371478 139233
rect 371422 139159 371478 139168
rect 371424 138712 371476 138718
rect 371422 138680 371424 138689
rect 371476 138680 371478 138689
rect 371422 138615 371478 138624
rect 371528 126313 371556 198183
rect 371620 127945 371648 198863
rect 371712 129062 371740 200903
rect 371804 197713 371832 269719
rect 371896 198801 371924 270807
rect 371988 200433 372016 272439
rect 372080 271969 372108 343839
rect 372250 341184 372306 341193
rect 372250 341119 372306 341128
rect 372160 293480 372212 293486
rect 372158 293448 372160 293457
rect 372212 293448 372214 293457
rect 372158 293383 372214 293392
rect 372160 291984 372212 291990
rect 372160 291926 372212 291932
rect 372172 291281 372200 291926
rect 372158 291272 372214 291281
rect 372158 291207 372214 291216
rect 372160 286680 372212 286686
rect 372160 286622 372212 286628
rect 372172 281081 372200 286622
rect 372158 281072 372214 281081
rect 372158 281007 372214 281016
rect 372066 271960 372122 271969
rect 372066 271895 372122 271904
rect 372080 267734 372108 271895
rect 372264 270201 372292 341119
rect 372448 279993 372476 351863
rect 372526 346624 372582 346633
rect 372582 346582 372660 346610
rect 372526 346559 372582 346568
rect 372434 279984 372490 279993
rect 372434 279919 372490 279928
rect 372632 274786 372660 346582
rect 372724 291990 372752 354646
rect 372802 349888 372858 349897
rect 372802 349823 372858 349832
rect 372712 291984 372764 291990
rect 372712 291926 372764 291932
rect 372816 277953 372844 349823
rect 372908 296721 372936 359450
rect 374092 353320 374144 353326
rect 374092 353262 374144 353268
rect 374000 349308 374052 349314
rect 374000 349250 374052 349256
rect 373264 297492 373316 297498
rect 373264 297434 373316 297440
rect 373276 296818 373304 297434
rect 373264 296812 373316 296818
rect 373264 296754 373316 296760
rect 372894 296712 372950 296721
rect 372894 296647 372950 296656
rect 372908 296070 372936 296647
rect 372896 296064 372948 296070
rect 372896 296006 372948 296012
rect 372802 277944 372858 277953
rect 372802 277879 372858 277888
rect 372816 277394 372844 277879
rect 372724 277366 372844 277394
rect 372620 274780 372672 274786
rect 372620 274722 372672 274728
rect 372526 274680 372582 274689
rect 372632 274666 372660 274722
rect 372582 274638 372660 274666
rect 372526 274615 372582 274624
rect 372250 270192 372306 270201
rect 372250 270127 372306 270136
rect 372080 267706 372200 267734
rect 372068 220652 372120 220658
rect 372068 220594 372120 220600
rect 372080 219745 372108 220594
rect 372066 219736 372122 219745
rect 372066 219671 372122 219680
rect 372068 213784 372120 213790
rect 372068 213726 372120 213732
rect 372080 212809 372108 213726
rect 372066 212800 372122 212809
rect 372066 212735 372122 212744
rect 372068 202836 372120 202842
rect 372068 202778 372120 202784
rect 372080 202609 372108 202778
rect 372066 202600 372122 202609
rect 372066 202535 372122 202544
rect 371974 200424 372030 200433
rect 371974 200359 372030 200368
rect 371882 198792 371938 198801
rect 371882 198727 371938 198736
rect 371790 197704 371846 197713
rect 371790 197639 371846 197648
rect 371700 129056 371752 129062
rect 371700 128998 371752 129004
rect 371606 127936 371662 127945
rect 371606 127871 371662 127880
rect 371514 126304 371570 126313
rect 371514 126239 371570 126248
rect 371528 125934 371556 126239
rect 371516 125928 371568 125934
rect 371516 125870 371568 125876
rect 371330 125216 371386 125225
rect 371330 125151 371386 125160
rect 371238 124672 371294 124681
rect 371238 124607 371294 124616
rect 370686 124264 370742 124273
rect 370686 124199 370742 124208
rect 371620 124166 371648 127871
rect 371804 126002 371832 197639
rect 371988 156754 372016 200359
rect 372172 199889 372200 267706
rect 372620 227044 372672 227050
rect 372620 226986 372672 226992
rect 372344 225752 372396 225758
rect 372250 225720 372306 225729
rect 372344 225694 372396 225700
rect 372250 225655 372252 225664
rect 372304 225655 372306 225664
rect 372252 225626 372304 225632
rect 372356 222358 372384 225694
rect 372526 225040 372582 225049
rect 372526 224975 372528 224984
rect 372580 224975 372582 224984
rect 372528 224946 372580 224952
rect 372344 222352 372396 222358
rect 372344 222294 372396 222300
rect 372632 219434 372660 226986
rect 372620 219428 372672 219434
rect 372620 219370 372672 219376
rect 372632 218657 372660 219370
rect 372618 218648 372674 218657
rect 372618 218583 372674 218592
rect 372252 217184 372304 217190
rect 372252 217126 372304 217132
rect 372264 213178 372292 217126
rect 372342 215520 372398 215529
rect 372342 215455 372344 215464
rect 372396 215455 372398 215464
rect 372344 215426 372396 215432
rect 372724 214554 372752 277366
rect 373080 274780 373132 274786
rect 373080 274722 373132 274728
rect 372896 274712 372948 274718
rect 372896 274654 372948 274660
rect 372804 229764 372856 229770
rect 372804 229706 372856 229712
rect 372816 225282 372844 229706
rect 372804 225276 372856 225282
rect 372804 225218 372856 225224
rect 372804 225072 372856 225078
rect 372804 225014 372856 225020
rect 372816 220726 372844 225014
rect 372804 220720 372856 220726
rect 372804 220662 372856 220668
rect 372802 220280 372858 220289
rect 372802 220215 372858 220224
rect 372632 214526 372752 214554
rect 372252 213172 372304 213178
rect 372252 213114 372304 213120
rect 372250 212256 372306 212265
rect 372250 212191 372306 212200
rect 372264 211818 372292 212191
rect 372252 211812 372304 211818
rect 372252 211754 372304 211760
rect 372632 205834 372660 214526
rect 372724 210118 372752 210149
rect 372712 210112 372764 210118
rect 372710 210080 372712 210089
rect 372764 210080 372766 210089
rect 372710 210015 372766 210024
rect 372620 205828 372672 205834
rect 372620 205770 372672 205776
rect 372724 200114 372752 210015
rect 372632 200086 372752 200114
rect 372158 199880 372214 199889
rect 372158 199815 372214 199824
rect 372066 199336 372122 199345
rect 372066 199271 372122 199280
rect 372080 159361 372108 199271
rect 372172 198937 372200 199815
rect 372158 198928 372214 198937
rect 372158 198863 372214 198872
rect 372632 195294 372660 200086
rect 372620 195288 372672 195294
rect 372620 195230 372672 195236
rect 372620 160744 372672 160750
rect 372620 160686 372672 160692
rect 372066 159352 372122 159361
rect 372066 159287 372122 159296
rect 371988 156738 372108 156754
rect 371988 156732 372120 156738
rect 371988 156726 372068 156732
rect 372068 156674 372120 156680
rect 371976 154556 372028 154562
rect 371976 154498 372028 154504
rect 371988 153241 372016 154498
rect 371974 153232 372030 153241
rect 371884 153196 371936 153202
rect 371974 153167 372030 153176
rect 371884 153138 371936 153144
rect 371896 152153 371924 153138
rect 371882 152144 371938 152153
rect 371882 152079 371938 152088
rect 372080 151814 372108 156674
rect 372632 152182 372660 160686
rect 372620 152176 372672 152182
rect 372620 152118 372672 152124
rect 372816 151814 372844 220215
rect 372908 204814 372936 274654
rect 372988 225752 373040 225758
rect 372988 225694 373040 225700
rect 373000 225350 373028 225694
rect 372988 225344 373040 225350
rect 372988 225286 373040 225292
rect 372988 225004 373040 225010
rect 372988 224946 373040 224952
rect 373000 208758 373028 224946
rect 372988 208752 373040 208758
rect 372988 208694 373040 208700
rect 372896 204808 372948 204814
rect 372896 204750 372948 204756
rect 372908 164218 372936 204750
rect 373092 202842 373120 274722
rect 373276 225690 373304 296754
rect 373356 293956 373408 293962
rect 373356 293898 373408 293904
rect 373368 293486 373396 293898
rect 373356 293480 373408 293486
rect 373356 293422 373408 293428
rect 373368 249762 373396 293422
rect 374012 277370 374040 349250
rect 374104 282198 374132 353262
rect 374196 297430 374224 368902
rect 378140 367192 378192 367198
rect 378140 367134 378192 367140
rect 376944 365900 376996 365906
rect 376944 365842 376996 365848
rect 375564 364676 375616 364682
rect 375564 364618 375616 364624
rect 374276 362976 374328 362982
rect 374276 362918 374328 362924
rect 374184 297424 374236 297430
rect 374184 297366 374236 297372
rect 374196 296750 374224 297366
rect 374184 296744 374236 296750
rect 374184 296686 374236 296692
rect 374288 292482 374316 362918
rect 375380 361548 375432 361554
rect 375380 361490 375432 361496
rect 374460 360460 374512 360466
rect 374460 360402 374512 360408
rect 374368 348220 374420 348226
rect 374368 348162 374420 348168
rect 374196 292454 374316 292482
rect 374196 292398 374224 292454
rect 374184 292392 374236 292398
rect 374184 292334 374236 292340
rect 374092 282192 374144 282198
rect 374092 282134 374144 282140
rect 374092 278996 374144 279002
rect 374092 278938 374144 278944
rect 374000 277364 374052 277370
rect 374000 277306 374052 277312
rect 374012 276078 374040 277306
rect 374000 276072 374052 276078
rect 374000 276014 374052 276020
rect 373356 249756 373408 249762
rect 373356 249698 373408 249704
rect 373540 225752 373592 225758
rect 373540 225694 373592 225700
rect 373264 225684 373316 225690
rect 373264 225626 373316 225632
rect 373172 225276 373224 225282
rect 373172 225218 373224 225224
rect 373184 220726 373212 225218
rect 373172 220720 373224 220726
rect 373172 220662 373224 220668
rect 373552 215490 373580 225694
rect 374000 223848 374052 223854
rect 374000 223790 374052 223796
rect 374012 222358 374040 223790
rect 374000 222352 374052 222358
rect 374000 222294 374052 222300
rect 373540 215484 373592 215490
rect 373540 215426 373592 215432
rect 373172 211812 373224 211818
rect 373172 211754 373224 211760
rect 373080 202836 373132 202842
rect 373080 202778 373132 202784
rect 373184 195906 373212 211754
rect 374104 206990 374132 278938
rect 374196 231130 374224 292334
rect 374276 282192 374328 282198
rect 374276 282134 374328 282140
rect 374184 231124 374236 231130
rect 374184 231066 374236 231072
rect 374288 210118 374316 282134
rect 374380 276146 374408 348162
rect 374472 288522 374500 360402
rect 375392 289610 375420 361490
rect 375472 353388 375524 353394
rect 375472 353330 375524 353336
rect 375380 289604 375432 289610
rect 375380 289546 375432 289552
rect 374460 288516 374512 288522
rect 374460 288458 374512 288464
rect 374368 276140 374420 276146
rect 374368 276082 374420 276088
rect 374368 225208 374420 225214
rect 374368 225150 374420 225156
rect 374380 217054 374408 225150
rect 374472 223922 374500 288458
rect 374644 286408 374696 286414
rect 374644 286350 374696 286356
rect 374552 276072 374604 276078
rect 374552 276014 374604 276020
rect 374460 223916 374512 223922
rect 374460 223858 374512 223864
rect 374368 217048 374420 217054
rect 374368 216990 374420 216996
rect 374276 210112 374328 210118
rect 374276 210054 374328 210060
rect 374092 206984 374144 206990
rect 374092 206926 374144 206932
rect 373264 205828 373316 205834
rect 373264 205770 373316 205776
rect 373172 195900 373224 195906
rect 373172 195842 373224 195848
rect 372896 164212 372948 164218
rect 372896 164154 372948 164160
rect 371896 151786 372108 151814
rect 372632 151786 372844 151814
rect 371896 128625 371924 151786
rect 371976 151632 372028 151638
rect 371976 151574 372028 151580
rect 371988 151065 372016 151574
rect 371974 151056 372030 151065
rect 371974 150991 372030 151000
rect 371976 150408 372028 150414
rect 371976 150350 372028 150356
rect 371988 149433 372016 150350
rect 371974 149424 372030 149433
rect 371974 149359 372030 149368
rect 371976 149048 372028 149054
rect 371976 148990 372028 148996
rect 371988 147801 372016 148990
rect 372526 148336 372582 148345
rect 372632 148322 372660 151786
rect 372582 148294 372660 148322
rect 372526 148271 372582 148280
rect 371974 147792 372030 147801
rect 371974 147727 372030 147736
rect 371976 147620 372028 147626
rect 371976 147562 372028 147568
rect 371988 146713 372016 147562
rect 371974 146704 372030 146713
rect 371974 146639 372030 146648
rect 371976 146124 372028 146130
rect 371976 146066 372028 146072
rect 371988 145625 372016 146066
rect 371974 145616 372030 145625
rect 371974 145551 372030 145560
rect 371976 143540 372028 143546
rect 371976 143482 372028 143488
rect 371988 143041 372016 143482
rect 371974 143032 372030 143041
rect 371974 142967 372030 142976
rect 371976 142112 372028 142118
rect 371976 142054 372028 142060
rect 371988 141409 372016 142054
rect 372068 142044 372120 142050
rect 372068 141986 372120 141992
rect 371974 141400 372030 141409
rect 371974 141335 372030 141344
rect 372080 140865 372108 141986
rect 372066 140856 372122 140865
rect 372066 140791 372122 140800
rect 373184 140350 373212 195842
rect 373276 162178 373304 205770
rect 374000 204264 374052 204270
rect 374000 204206 374052 204212
rect 374012 202874 374040 204206
rect 373920 202846 374040 202874
rect 373356 202836 373408 202842
rect 373356 202778 373408 202784
rect 373264 162172 373316 162178
rect 373264 162114 373316 162120
rect 373276 153105 373304 162114
rect 373368 160750 373396 202778
rect 373356 160744 373408 160750
rect 373356 160686 373408 160692
rect 373920 158710 373948 202846
rect 374000 201612 374052 201618
rect 374000 201554 374052 201560
rect 373908 158704 373960 158710
rect 373908 158646 373960 158652
rect 373262 153096 373318 153105
rect 373262 153031 373318 153040
rect 371976 140344 372028 140350
rect 371974 140312 371976 140321
rect 373172 140344 373224 140350
rect 372028 140312 372030 140321
rect 373172 140286 373224 140292
rect 371974 140247 372030 140256
rect 371976 139052 372028 139058
rect 371976 138994 372028 139000
rect 371988 138145 372016 138994
rect 371974 138136 372030 138145
rect 371974 138071 372030 138080
rect 374012 129606 374040 201554
rect 374092 195968 374144 195974
rect 374092 195910 374144 195916
rect 374000 129600 374052 129606
rect 374000 129542 374052 129548
rect 371882 128616 371938 128625
rect 371882 128551 371938 128560
rect 371792 125996 371844 126002
rect 371792 125938 371844 125944
rect 371804 125769 371832 125938
rect 371790 125760 371846 125769
rect 371790 125695 371846 125704
rect 374104 125526 374132 195910
rect 374184 195288 374236 195294
rect 374184 195230 374236 195236
rect 374196 139058 374224 195230
rect 374380 145926 374408 216990
rect 374472 216034 374500 223858
rect 374460 216028 374512 216034
rect 374460 215970 374512 215976
rect 374564 205358 374592 276014
rect 374656 213314 374684 286350
rect 375380 285524 375432 285530
rect 375380 285466 375432 285472
rect 375104 276140 375156 276146
rect 375104 276082 375156 276088
rect 374920 222896 374972 222902
rect 374920 222838 374972 222844
rect 374644 213308 374696 213314
rect 374644 213250 374696 213256
rect 374736 211132 374788 211138
rect 374736 211074 374788 211080
rect 374748 210662 374776 211074
rect 374736 210656 374788 210662
rect 374736 210598 374788 210604
rect 374552 205352 374604 205358
rect 374552 205294 374604 205300
rect 374564 172514 374592 205294
rect 374644 202496 374696 202502
rect 374644 202438 374696 202444
rect 374552 172508 374604 172514
rect 374552 172450 374604 172456
rect 374564 171154 374592 172450
rect 374552 171148 374604 171154
rect 374552 171090 374604 171096
rect 374656 154630 374684 202438
rect 374748 186318 374776 210598
rect 374736 186312 374788 186318
rect 374736 186254 374788 186260
rect 374644 154624 374696 154630
rect 374644 154566 374696 154572
rect 374656 152114 374684 154566
rect 374644 152108 374696 152114
rect 374644 152050 374696 152056
rect 374932 151774 374960 222838
rect 375012 215484 375064 215490
rect 375012 215426 375064 215432
rect 374920 151768 374972 151774
rect 374920 151710 374972 151716
rect 374368 145920 374420 145926
rect 374368 145862 374420 145868
rect 375024 143954 375052 215426
rect 375116 204270 375144 276082
rect 375392 213246 375420 285466
rect 375484 282742 375512 353330
rect 375576 293962 375604 364618
rect 376760 357536 376812 357542
rect 376760 357478 376812 357484
rect 375656 356244 375708 356250
rect 375656 356186 375708 356192
rect 375564 293956 375616 293962
rect 375564 293898 375616 293904
rect 375564 289604 375616 289610
rect 375564 289546 375616 289552
rect 375472 282736 375524 282742
rect 375472 282678 375524 282684
rect 375380 213240 375432 213246
rect 375380 213182 375432 213188
rect 375484 211138 375512 282678
rect 375576 218006 375604 289546
rect 375668 285530 375696 356186
rect 376024 293276 376076 293282
rect 376024 293218 376076 293224
rect 375656 285524 375708 285530
rect 375656 285466 375708 285472
rect 375656 222420 375708 222426
rect 375656 222362 375708 222368
rect 375564 218000 375616 218006
rect 375564 217942 375616 217948
rect 375576 216714 375604 217942
rect 375564 216708 375616 216714
rect 375564 216650 375616 216656
rect 375564 215960 375616 215966
rect 375564 215902 375616 215908
rect 375472 211132 375524 211138
rect 375472 211074 375524 211080
rect 375104 204264 375156 204270
rect 375104 204206 375156 204212
rect 375288 186312 375340 186318
rect 375340 186260 375420 186266
rect 375288 186254 375420 186260
rect 375300 186238 375420 186254
rect 375392 180794 375420 186238
rect 375392 180766 375512 180794
rect 375012 143948 375064 143954
rect 375012 143890 375064 143896
rect 374184 139052 374236 139058
rect 374184 138994 374236 139000
rect 375484 138718 375512 180766
rect 375576 144294 375604 215902
rect 375668 150958 375696 222362
rect 376036 220794 376064 293218
rect 376772 287026 376800 357478
rect 376852 354816 376904 354822
rect 376852 354758 376904 354764
rect 376760 287020 376812 287026
rect 376760 286962 376812 286968
rect 376772 285734 376800 286962
rect 376760 285728 376812 285734
rect 376760 285670 376812 285676
rect 376864 283778 376892 354758
rect 376956 295322 376984 365842
rect 377036 361684 377088 361690
rect 377036 361626 377088 361632
rect 376944 295316 376996 295322
rect 376944 295258 376996 295264
rect 376944 294024 376996 294030
rect 376944 293966 376996 293972
rect 376772 283750 376892 283778
rect 376772 283694 376800 283750
rect 376760 283688 376812 283694
rect 376760 283630 376812 283636
rect 376024 220788 376076 220794
rect 376024 220730 376076 220736
rect 375932 218136 375984 218142
rect 375932 218078 375984 218084
rect 375840 209840 375892 209846
rect 375840 209782 375892 209788
rect 375746 208448 375802 208457
rect 375746 208383 375802 208392
rect 375760 175234 375788 208383
rect 375852 189038 375880 209782
rect 375840 189032 375892 189038
rect 375840 188974 375892 188980
rect 375748 175228 375800 175234
rect 375748 175170 375800 175176
rect 375656 150952 375708 150958
rect 375656 150894 375708 150900
rect 375944 146198 375972 218078
rect 376772 211274 376800 283630
rect 376956 222426 376984 293966
rect 377048 290562 377076 361626
rect 378152 296138 378180 367134
rect 383660 367124 383712 367130
rect 383660 367066 383712 367072
rect 382280 365832 382332 365838
rect 382280 365774 382332 365780
rect 378324 363112 378376 363118
rect 378324 363054 378376 363060
rect 378232 360392 378284 360398
rect 378232 360334 378284 360340
rect 378140 296132 378192 296138
rect 378140 296074 378192 296080
rect 377036 290556 377088 290562
rect 377036 290498 377088 290504
rect 376944 222420 376996 222426
rect 376944 222362 376996 222368
rect 377048 218142 377076 290498
rect 377404 284368 377456 284374
rect 377404 284310 377456 284316
rect 377036 218136 377088 218142
rect 377036 218078 377088 218084
rect 376944 216708 376996 216714
rect 376944 216650 376996 216656
rect 376852 212492 376904 212498
rect 376852 212434 376904 212440
rect 376760 211268 376812 211274
rect 376760 211210 376812 211216
rect 376772 209846 376800 211210
rect 376864 211206 376892 212434
rect 376852 211200 376904 211206
rect 376852 211142 376904 211148
rect 376760 209840 376812 209846
rect 376760 209782 376812 209788
rect 375932 146192 375984 146198
rect 375932 146134 375984 146140
rect 375564 144288 375616 144294
rect 375564 144230 375616 144236
rect 376772 139398 376800 209782
rect 376864 140690 376892 211142
rect 376956 146130 376984 216650
rect 377416 213790 377444 284310
rect 378152 222902 378180 296074
rect 378244 289134 378272 360334
rect 378336 292466 378364 363054
rect 380992 361616 381044 361622
rect 380992 361558 381044 361564
rect 379520 359576 379572 359582
rect 379520 359518 379572 359524
rect 378416 352640 378468 352646
rect 378416 352582 378468 352588
rect 378324 292460 378376 292466
rect 378324 292402 378376 292408
rect 378336 292058 378364 292402
rect 378324 292052 378376 292058
rect 378324 291994 378376 292000
rect 378232 289128 378284 289134
rect 378232 289070 378284 289076
rect 378244 287054 378272 289070
rect 378428 287706 378456 352582
rect 379532 297498 379560 359518
rect 380900 354748 380952 354754
rect 380900 354690 380952 354696
rect 379612 352572 379664 352578
rect 379612 352514 379664 352520
rect 379520 297492 379572 297498
rect 379520 297434 379572 297440
rect 379520 296064 379572 296070
rect 379520 296006 379572 296012
rect 378508 291984 378560 291990
rect 378508 291926 378560 291932
rect 378416 287700 378468 287706
rect 378416 287642 378468 287648
rect 378244 287026 378364 287054
rect 378336 225214 378364 287026
rect 378428 225758 378456 287642
rect 378416 225752 378468 225758
rect 378416 225694 378468 225700
rect 378324 225208 378376 225214
rect 378324 225150 378376 225156
rect 378324 223576 378376 223582
rect 378324 223518 378376 223524
rect 378140 222896 378192 222902
rect 378140 222838 378192 222844
rect 378336 222290 378364 223518
rect 378324 222284 378376 222290
rect 378324 222226 378376 222232
rect 378232 218272 378284 218278
rect 378232 218214 378284 218220
rect 378140 216028 378192 216034
rect 378140 215970 378192 215976
rect 377404 213784 377456 213790
rect 377404 213726 377456 213732
rect 377036 213308 377088 213314
rect 377036 213250 377088 213256
rect 377048 197062 377076 213250
rect 377036 197056 377088 197062
rect 377036 196998 377088 197004
rect 376944 146124 376996 146130
rect 376944 146066 376996 146072
rect 377048 141982 377076 196998
rect 378152 144770 378180 215970
rect 378244 147558 378272 218214
rect 378336 151638 378364 222226
rect 378520 218754 378548 291926
rect 379532 224330 379560 296006
rect 379624 288386 379652 352514
rect 379612 288380 379664 288386
rect 379612 288322 379664 288328
rect 379624 287094 379652 288322
rect 379612 287088 379664 287094
rect 379612 287030 379664 287036
rect 380912 283626 380940 354690
rect 381004 290494 381032 361558
rect 381084 356176 381136 356182
rect 381084 356118 381136 356124
rect 380992 290488 381044 290494
rect 380992 290430 381044 290436
rect 380900 283620 380952 283626
rect 380900 283562 380952 283568
rect 380912 282946 380940 283562
rect 380900 282940 380952 282946
rect 380900 282882 380952 282888
rect 379520 224324 379572 224330
rect 379520 224266 379572 224272
rect 378508 218748 378560 218754
rect 378508 218690 378560 218696
rect 378520 218278 378548 218690
rect 378508 218272 378560 218278
rect 378508 218214 378560 218220
rect 378416 214396 378468 214402
rect 378416 214338 378468 214344
rect 378428 213994 378456 214338
rect 378416 213988 378468 213994
rect 378416 213930 378468 213936
rect 378428 197130 378456 213930
rect 378416 197124 378468 197130
rect 378416 197066 378468 197072
rect 378324 151632 378376 151638
rect 378324 151574 378376 151580
rect 378232 147552 378284 147558
rect 378232 147494 378284 147500
rect 378140 144764 378192 144770
rect 378140 144706 378192 144712
rect 378428 143478 378456 197066
rect 379532 153134 379560 224266
rect 380900 220788 380952 220794
rect 380900 220730 380952 220736
rect 379520 153128 379572 153134
rect 379520 153070 379572 153076
rect 380912 148986 380940 220730
rect 381004 219434 381032 290430
rect 381096 285666 381124 356118
rect 382292 294642 382320 365774
rect 382372 364404 382424 364410
rect 382372 364346 382424 364352
rect 382280 294636 382332 294642
rect 382280 294578 382332 294584
rect 382292 292754 382320 294578
rect 382384 293282 382412 364346
rect 382556 357468 382608 357474
rect 382556 357410 382608 357416
rect 382372 293276 382424 293282
rect 382372 293218 382424 293224
rect 382292 292726 382504 292754
rect 382372 292052 382424 292058
rect 382372 291994 382424 292000
rect 381268 285728 381320 285734
rect 381268 285670 381320 285676
rect 381084 285660 381136 285666
rect 381084 285602 381136 285608
rect 381096 284442 381124 285602
rect 381084 284436 381136 284442
rect 381084 284378 381136 284384
rect 381176 282940 381228 282946
rect 381176 282882 381228 282888
rect 381084 225684 381136 225690
rect 381084 225626 381136 225632
rect 380992 219428 381044 219434
rect 380992 219370 381044 219376
rect 380900 148980 380952 148986
rect 380900 148922 380952 148928
rect 381004 147626 381032 219370
rect 381096 154494 381124 225626
rect 381188 212498 381216 282882
rect 381280 214402 381308 285670
rect 382280 284436 382332 284442
rect 382280 284378 382332 284384
rect 381268 214396 381320 214402
rect 381268 214338 381320 214344
rect 381176 212492 381228 212498
rect 381176 212434 381228 212440
rect 382292 211818 382320 284378
rect 382384 220726 382412 291994
rect 382476 223582 382504 292726
rect 382568 286414 382596 357410
rect 383672 296002 383700 367066
rect 385040 365764 385092 365770
rect 385040 365706 385092 365712
rect 383752 354000 383804 354006
rect 383752 353942 383804 353948
rect 383660 295996 383712 296002
rect 383660 295938 383712 295944
rect 382556 286408 382608 286414
rect 382556 286350 382608 286356
rect 383672 224262 383700 295938
rect 383764 286346 383792 353942
rect 385052 294030 385080 365706
rect 385224 356108 385276 356114
rect 385224 356050 385276 356056
rect 385132 297424 385184 297430
rect 385132 297366 385184 297372
rect 385040 294024 385092 294030
rect 385040 293966 385092 293972
rect 383752 286340 383804 286346
rect 383752 286282 383804 286288
rect 383764 225146 383792 286282
rect 385144 225622 385172 297366
rect 385236 284374 385264 356050
rect 396736 309806 396764 699654
rect 396724 309800 396776 309806
rect 396724 309742 396776 309748
rect 429212 304434 429240 703582
rect 429672 703474 429700 703582
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494072 703582 494652 703610
rect 429856 703474 429884 703520
rect 429672 703446 429884 703474
rect 462332 698970 462360 703520
rect 478524 700466 478552 703520
rect 478512 700460 478564 700466
rect 478512 700402 478564 700408
rect 479524 700392 479576 700398
rect 479524 700334 479576 700340
rect 462320 698964 462372 698970
rect 462320 698906 462372 698912
rect 445206 369472 445262 369481
rect 445206 369407 445262 369416
rect 445220 368558 445248 369407
rect 445208 368552 445260 368558
rect 445208 368494 445260 368500
rect 454040 368552 454092 368558
rect 454040 368494 454092 368500
rect 445666 368384 445722 368393
rect 445722 368342 445800 368370
rect 445666 368319 445722 368328
rect 445666 367160 445722 367169
rect 445666 367095 445668 367104
rect 445720 367095 445722 367104
rect 445668 367066 445720 367072
rect 445298 366072 445354 366081
rect 445298 366007 445354 366016
rect 445312 365770 445340 366007
rect 445300 365764 445352 365770
rect 445300 365706 445352 365712
rect 445666 364848 445722 364857
rect 445666 364783 445722 364792
rect 445680 364410 445708 364783
rect 445668 364404 445720 364410
rect 445668 364346 445720 364352
rect 444930 363760 444986 363769
rect 444930 363695 444986 363704
rect 444944 362982 444972 363695
rect 444932 362976 444984 362982
rect 444932 362918 444984 362924
rect 445206 362536 445262 362545
rect 445206 362471 445262 362480
rect 445220 361622 445248 362471
rect 445208 361616 445260 361622
rect 445208 361558 445260 361564
rect 445114 361448 445170 361457
rect 445114 361383 445170 361392
rect 445128 360806 445156 361383
rect 445116 360800 445168 360806
rect 445116 360742 445168 360748
rect 444564 360324 444616 360330
rect 444564 360266 444616 360272
rect 444576 360233 444604 360266
rect 444562 360224 444618 360233
rect 444562 360159 444618 360168
rect 444562 357912 444618 357921
rect 444562 357847 444618 357856
rect 444576 357474 444604 357847
rect 444564 357468 444616 357474
rect 444564 357410 444616 357416
rect 444378 356824 444434 356833
rect 444378 356759 444434 356768
rect 444392 356250 444420 356759
rect 444380 356244 444432 356250
rect 444380 356186 444432 356192
rect 444746 355600 444802 355609
rect 444746 355535 444802 355544
rect 444760 355094 444788 355535
rect 444748 355088 444800 355094
rect 444748 355030 444800 355036
rect 444746 353288 444802 353297
rect 444746 353223 444802 353232
rect 444760 352510 444788 353223
rect 444748 352504 444800 352510
rect 444748 352446 444800 352452
rect 444470 352200 444526 352209
rect 444470 352135 444526 352144
rect 444484 352034 444512 352135
rect 444472 352028 444524 352034
rect 444472 351970 444524 351976
rect 444378 350976 444434 350985
rect 444378 350911 444434 350920
rect 431972 340054 432952 340082
rect 434732 340054 434884 340082
rect 436112 340054 436908 340082
rect 438932 340054 438992 340082
rect 440956 340054 441292 340082
rect 429200 304428 429252 304434
rect 429200 304370 429252 304376
rect 385408 295316 385460 295322
rect 385408 295258 385460 295264
rect 385316 287088 385368 287094
rect 385316 287030 385368 287036
rect 385224 284368 385276 284374
rect 385224 284310 385276 284316
rect 385132 225616 385184 225622
rect 385132 225558 385184 225564
rect 383752 225140 383804 225146
rect 383752 225082 383804 225088
rect 383660 224256 383712 224262
rect 383660 224198 383712 224204
rect 382464 223576 382516 223582
rect 382464 223518 382516 223524
rect 382464 220924 382516 220930
rect 382464 220866 382516 220872
rect 382372 220720 382424 220726
rect 382372 220662 382424 220668
rect 382280 211812 382332 211818
rect 382280 211754 382332 211760
rect 382280 196784 382332 196790
rect 382280 196726 382332 196732
rect 381084 154488 381136 154494
rect 381084 154430 381136 154436
rect 380992 147620 381044 147626
rect 380992 147562 381044 147568
rect 378416 143472 378468 143478
rect 378416 143414 378468 143420
rect 382292 142050 382320 196726
rect 382384 149054 382412 220662
rect 382476 150346 382504 220866
rect 382556 213784 382608 213790
rect 382556 213726 382608 213732
rect 382568 197198 382596 213726
rect 382556 197192 382608 197198
rect 382556 197134 382608 197140
rect 382568 196790 382596 197134
rect 382556 196784 382608 196790
rect 382556 196726 382608 196732
rect 383672 153202 383700 224198
rect 383764 215218 383792 225082
rect 385040 221468 385092 221474
rect 385040 221410 385092 221416
rect 383752 215212 383804 215218
rect 383752 215154 383804 215160
rect 383752 213240 383804 213246
rect 383752 213182 383804 213188
rect 383764 197266 383792 213182
rect 383752 197260 383804 197266
rect 383752 197202 383804 197208
rect 383660 153196 383712 153202
rect 383660 153138 383712 153144
rect 382464 150340 382516 150346
rect 382464 150282 382516 150288
rect 382372 149048 382424 149054
rect 382372 148990 382424 148996
rect 383764 142118 383792 197202
rect 385052 150414 385080 221410
rect 385144 154562 385172 225558
rect 385328 223990 385356 287030
rect 385316 223984 385368 223990
rect 385316 223926 385368 223932
rect 385328 219434 385356 223926
rect 385420 220930 385448 295258
rect 431972 287054 432000 340054
rect 434732 297634 434760 340054
rect 436112 297702 436140 340054
rect 438964 337482 438992 340054
rect 438952 337476 439004 337482
rect 438952 337418 439004 337424
rect 441264 336802 441292 340054
rect 441252 336796 441304 336802
rect 441252 336738 441304 336744
rect 441620 336796 441672 336802
rect 441620 336738 441672 336744
rect 436100 297696 436152 297702
rect 436100 297638 436152 297644
rect 434720 297628 434772 297634
rect 434720 297570 434772 297576
rect 431972 287026 432552 287054
rect 432524 268682 432552 287026
rect 432524 268654 432952 268682
rect 432616 265742 432644 268654
rect 441632 268138 441660 336738
rect 443644 302388 443696 302394
rect 443644 302330 443696 302336
rect 442264 298172 442316 298178
rect 442264 298114 442316 298120
rect 441712 297628 441764 297634
rect 441712 297570 441764 297576
rect 434884 268110 435220 268138
rect 436908 268110 437244 268138
rect 440956 268124 441660 268138
rect 435192 266354 435220 268110
rect 437216 267734 437244 268110
rect 438918 268002 438946 268124
rect 440942 268110 441660 268124
rect 440942 268002 440970 268110
rect 438872 267974 438946 268002
rect 440896 267974 440970 268002
rect 437216 267706 437428 267734
rect 438872 267714 438900 267974
rect 435180 266348 435232 266354
rect 435180 266290 435232 266296
rect 437400 266286 437428 267706
rect 438860 267708 438912 267714
rect 438860 267650 438912 267656
rect 437388 266280 437440 266286
rect 437388 266222 437440 266228
rect 431960 265736 432012 265742
rect 431960 265678 432012 265684
rect 432604 265736 432656 265742
rect 432604 265678 432656 265684
rect 385408 220924 385460 220930
rect 385408 220866 385460 220872
rect 385236 219406 385356 219434
rect 385236 215966 385264 219406
rect 385224 215960 385276 215966
rect 385224 215902 385276 215908
rect 385224 215212 385276 215218
rect 385224 215154 385276 215160
rect 385132 154556 385184 154562
rect 385132 154498 385184 154504
rect 385040 150408 385092 150414
rect 385040 150350 385092 150356
rect 385236 143546 385264 215154
rect 431972 209774 432000 265678
rect 437400 226234 437428 266222
rect 440896 265674 440924 267974
rect 441724 267734 441752 297570
rect 442276 273222 442304 298114
rect 443000 297696 443052 297702
rect 443000 297638 443052 297644
rect 442264 273216 442316 273222
rect 442264 273158 442316 273164
rect 441632 267706 441752 267734
rect 441632 266354 441660 267706
rect 441620 266348 441672 266354
rect 441620 266290 441672 266296
rect 440884 265668 440936 265674
rect 440884 265610 440936 265616
rect 440896 226302 440924 265610
rect 440884 226296 440936 226302
rect 440884 226238 440936 226244
rect 437388 226228 437440 226234
rect 437388 226170 437440 226176
rect 431972 209746 432552 209774
rect 432524 196058 432552 209746
rect 441344 197328 441396 197334
rect 441344 197270 441396 197276
rect 441356 196058 441384 197270
rect 432524 196030 432952 196058
rect 434884 196030 435220 196058
rect 436908 196030 437244 196058
rect 438932 196030 438992 196058
rect 440956 196030 441384 196058
rect 432524 180794 432552 196030
rect 435192 193730 435220 196030
rect 436008 194540 436060 194546
rect 436008 194482 436060 194488
rect 436020 193730 436048 194482
rect 437216 194478 437244 196030
rect 437204 194472 437256 194478
rect 437204 194414 437256 194420
rect 438964 193866 438992 196030
rect 438952 193860 439004 193866
rect 438952 193802 439004 193808
rect 435180 193724 435232 193730
rect 435180 193666 435232 193672
rect 436008 193724 436060 193730
rect 436008 193666 436060 193672
rect 436020 181694 436048 193666
rect 441356 190454 441384 196030
rect 441632 194546 441660 266290
rect 443012 266286 443040 297638
rect 443000 266280 443052 266286
rect 443000 266222 443052 266228
rect 443000 226296 443052 226302
rect 443000 226238 443052 226244
rect 441712 226228 441764 226234
rect 441712 226170 441764 226176
rect 441620 194540 441672 194546
rect 441620 194482 441672 194488
rect 441724 194478 441752 226170
rect 441804 225072 441856 225078
rect 441802 225040 441804 225049
rect 441856 225040 441858 225049
rect 441802 224975 441858 224984
rect 441804 224256 441856 224262
rect 441802 224224 441804 224233
rect 441856 224224 441858 224233
rect 441802 224159 441858 224168
rect 443012 197334 443040 226238
rect 443656 219434 443684 302330
rect 444392 279682 444420 350911
rect 444470 349888 444526 349897
rect 444470 349823 444526 349832
rect 444380 279676 444432 279682
rect 444380 279618 444432 279624
rect 444484 277953 444512 349823
rect 445666 348664 445722 348673
rect 445666 348599 445722 348608
rect 445680 347818 445708 348599
rect 445668 347812 445720 347818
rect 445668 347754 445720 347760
rect 444654 347576 444710 347585
rect 444654 347511 444710 347520
rect 444668 346458 444696 347511
rect 444656 346452 444708 346458
rect 444656 346394 444708 346400
rect 445298 346352 445354 346361
rect 445298 346287 445354 346296
rect 445312 345166 445340 346287
rect 445666 345264 445722 345273
rect 445666 345199 445722 345208
rect 445300 345160 445352 345166
rect 445300 345102 445352 345108
rect 445680 345098 445708 345199
rect 445668 345092 445720 345098
rect 445668 345034 445720 345040
rect 445666 344040 445722 344049
rect 445666 343975 445722 343984
rect 445680 343738 445708 343975
rect 445668 343732 445720 343738
rect 445668 343674 445720 343680
rect 445022 342952 445078 342961
rect 445022 342887 445078 342896
rect 445036 342310 445064 342887
rect 445024 342304 445076 342310
rect 445024 342246 445076 342252
rect 444562 341728 444618 341737
rect 444562 341663 444618 341672
rect 444576 341290 444604 341663
rect 444564 341284 444616 341290
rect 444564 341226 444616 341232
rect 444562 340640 444618 340649
rect 444562 340575 444618 340584
rect 444576 340202 444604 340575
rect 444564 340196 444616 340202
rect 444564 340138 444616 340144
rect 445666 297528 445722 297537
rect 445666 297463 445722 297472
rect 445680 297090 445708 297463
rect 445668 297084 445720 297090
rect 445668 297026 445720 297032
rect 445666 296440 445722 296449
rect 445772 296426 445800 368342
rect 449900 367124 449952 367130
rect 449900 367066 449952 367072
rect 448612 362976 448664 362982
rect 448612 362918 448664 362924
rect 445850 359136 445906 359145
rect 445850 359071 445906 359080
rect 445722 296398 445800 296426
rect 445666 296375 445722 296384
rect 445772 296002 445800 296398
rect 445760 295996 445812 296002
rect 445760 295938 445812 295944
rect 445668 295316 445720 295322
rect 445668 295258 445720 295264
rect 445680 295225 445708 295258
rect 445666 295216 445722 295225
rect 445666 295151 445722 295160
rect 445668 294636 445720 294642
rect 445668 294578 445720 294584
rect 445680 294137 445708 294578
rect 445666 294128 445722 294137
rect 445666 294063 445722 294072
rect 445668 293276 445720 293282
rect 445668 293218 445720 293224
rect 445680 292913 445708 293218
rect 445666 292904 445722 292913
rect 445666 292839 445722 292848
rect 445666 291816 445722 291825
rect 445666 291751 445722 291760
rect 445680 291242 445708 291751
rect 445668 291236 445720 291242
rect 445668 291178 445720 291184
rect 445666 290592 445722 290601
rect 445722 290550 445800 290578
rect 445666 290527 445722 290536
rect 445772 290494 445800 290550
rect 445760 290488 445812 290494
rect 445760 290430 445812 290436
rect 445666 289504 445722 289513
rect 445666 289439 445722 289448
rect 445680 289202 445708 289439
rect 445668 289196 445720 289202
rect 445668 289138 445720 289144
rect 445666 288280 445722 288289
rect 445666 288215 445722 288224
rect 445484 287292 445536 287298
rect 445484 287234 445536 287240
rect 445496 287201 445524 287234
rect 445482 287192 445538 287201
rect 445680 287162 445708 288215
rect 445482 287127 445538 287136
rect 445668 287156 445720 287162
rect 445668 287098 445720 287104
rect 445668 286000 445720 286006
rect 445666 285968 445668 285977
rect 445720 285968 445722 285977
rect 445666 285903 445722 285912
rect 445390 284880 445446 284889
rect 445390 284815 445392 284824
rect 445444 284815 445446 284824
rect 445392 284786 445444 284792
rect 445666 283656 445722 283665
rect 445666 283591 445668 283600
rect 445720 283591 445722 283600
rect 445668 283562 445720 283568
rect 445668 281376 445720 281382
rect 445666 281344 445668 281353
rect 445720 281344 445722 281353
rect 445666 281279 445722 281288
rect 445024 280288 445076 280294
rect 445022 280256 445024 280265
rect 445076 280256 445078 280265
rect 445022 280191 445078 280200
rect 444656 279676 444708 279682
rect 444656 279618 444708 279624
rect 444668 279041 444696 279618
rect 444654 279032 444710 279041
rect 444654 278967 444710 278976
rect 444470 277944 444526 277953
rect 444470 277879 444526 277888
rect 443644 219428 443696 219434
rect 443644 219370 443696 219376
rect 444484 205873 444512 277879
rect 444564 268728 444616 268734
rect 444562 268696 444564 268705
rect 444616 268696 444618 268705
rect 444562 268631 444618 268640
rect 444564 225004 444616 225010
rect 444564 224946 444616 224952
rect 444576 223582 444604 224946
rect 444564 223576 444616 223582
rect 444564 223518 444616 223524
rect 444576 223145 444604 223518
rect 444562 223136 444618 223145
rect 444562 223071 444618 223080
rect 444564 210520 444616 210526
rect 444562 210488 444564 210497
rect 444616 210488 444618 210497
rect 444562 210423 444618 210432
rect 444668 209774 444696 278967
rect 445666 276720 445722 276729
rect 445666 276655 445668 276664
rect 445720 276655 445722 276664
rect 445668 276626 445720 276632
rect 445668 276004 445720 276010
rect 445668 275946 445720 275952
rect 445680 275641 445708 275946
rect 445666 275632 445722 275641
rect 445666 275567 445722 275576
rect 445668 274644 445720 274650
rect 445668 274586 445720 274592
rect 445680 274417 445708 274586
rect 445666 274408 445722 274417
rect 445666 274343 445722 274352
rect 445024 273964 445076 273970
rect 445024 273906 445076 273912
rect 445036 273329 445064 273906
rect 445022 273320 445078 273329
rect 445022 273255 445078 273264
rect 445668 272536 445720 272542
rect 445668 272478 445720 272484
rect 445680 272105 445708 272478
rect 445666 272096 445722 272105
rect 445666 272031 445722 272040
rect 445666 271008 445722 271017
rect 445666 270943 445722 270952
rect 445680 270570 445708 270943
rect 445668 270564 445720 270570
rect 445668 270506 445720 270512
rect 445392 269816 445444 269822
rect 445390 269784 445392 269793
rect 445444 269784 445446 269793
rect 445390 269719 445446 269728
rect 445668 222148 445720 222154
rect 445668 222090 445720 222096
rect 445680 222057 445708 222090
rect 445666 222048 445722 222057
rect 445666 221983 445722 221992
rect 445114 220824 445170 220833
rect 445114 220759 445170 220768
rect 445128 220114 445156 220759
rect 445116 220108 445168 220114
rect 445116 220050 445168 220056
rect 445666 219736 445722 219745
rect 445666 219671 445722 219680
rect 445680 219638 445708 219671
rect 445668 219632 445720 219638
rect 445668 219574 445720 219580
rect 445666 218512 445722 218521
rect 445772 218498 445800 290430
rect 445864 287298 445892 359071
rect 448520 357468 448572 357474
rect 448520 357410 448572 357416
rect 447140 356244 447192 356250
rect 447140 356186 447192 356192
rect 445942 354512 445998 354521
rect 445942 354447 445998 354456
rect 445852 287292 445904 287298
rect 445852 287234 445904 287240
rect 445956 287054 445984 354447
rect 446036 340196 446088 340202
rect 446036 340138 446088 340144
rect 445864 287026 445984 287054
rect 445864 282577 445892 287026
rect 445850 282568 445906 282577
rect 445850 282503 445906 282512
rect 445722 218470 445800 218498
rect 445666 218447 445722 218456
rect 445772 218074 445800 218470
rect 445760 218068 445812 218074
rect 445760 218010 445812 218016
rect 445666 217424 445722 217433
rect 445666 217359 445722 217368
rect 445680 217326 445708 217359
rect 445668 217320 445720 217326
rect 445668 217262 445720 217268
rect 445666 216200 445722 216209
rect 445666 216135 445668 216144
rect 445720 216135 445722 216144
rect 445668 216106 445720 216112
rect 445666 215112 445722 215121
rect 445666 215047 445722 215056
rect 445680 214062 445708 215047
rect 445668 214056 445720 214062
rect 445668 213998 445720 214004
rect 445668 213920 445720 213926
rect 445666 213888 445668 213897
rect 445720 213888 445722 213897
rect 445666 213823 445722 213832
rect 445300 212832 445352 212838
rect 445298 212800 445300 212809
rect 445352 212800 445354 212809
rect 445298 212735 445354 212744
rect 445668 211608 445720 211614
rect 445666 211576 445668 211585
rect 445720 211576 445722 211585
rect 445666 211511 445722 211520
rect 445864 211138 445892 282503
rect 446048 268734 446076 340138
rect 447152 284850 447180 356186
rect 447232 352028 447284 352034
rect 447232 351970 447284 351976
rect 447140 284844 447192 284850
rect 447140 284786 447192 284792
rect 447152 284374 447180 284786
rect 447140 284368 447192 284374
rect 447140 284310 447192 284316
rect 447244 280294 447272 351970
rect 447508 346452 447560 346458
rect 447508 346394 447560 346400
rect 447416 341284 447468 341290
rect 447416 341226 447468 341232
rect 447324 284368 447376 284374
rect 447324 284310 447376 284316
rect 447232 280288 447284 280294
rect 447232 280230 447284 280236
rect 447244 277394 447272 280230
rect 447152 277366 447272 277394
rect 446404 274644 446456 274650
rect 446404 274586 446456 274592
rect 446036 268728 446088 268734
rect 446036 268670 446088 268676
rect 446048 258074 446076 268670
rect 445956 258046 446076 258074
rect 445852 211132 445904 211138
rect 445852 211074 445904 211080
rect 444668 209746 444788 209774
rect 444760 206961 444788 209746
rect 445666 209264 445722 209273
rect 445666 209199 445668 209208
rect 445720 209199 445722 209208
rect 445668 209170 445720 209176
rect 445116 208208 445168 208214
rect 445114 208176 445116 208185
rect 445168 208176 445170 208185
rect 445114 208111 445170 208120
rect 444746 206952 444802 206961
rect 444746 206887 444802 206896
rect 444470 205864 444526 205873
rect 444470 205799 444526 205808
rect 443000 197328 443052 197334
rect 443000 197270 443052 197276
rect 441712 194472 441764 194478
rect 441712 194414 441764 194420
rect 443184 194472 443236 194478
rect 443184 194414 443236 194420
rect 441356 190426 441568 190454
rect 436008 181688 436060 181694
rect 436008 181630 436060 181636
rect 431972 180766 432552 180794
rect 385224 143540 385276 143546
rect 385224 143482 385276 143488
rect 383752 142112 383804 142118
rect 383752 142054 383804 142060
rect 382280 142044 382332 142050
rect 382280 141986 382332 141992
rect 377036 141976 377088 141982
rect 377036 141918 377088 141924
rect 376852 140684 376904 140690
rect 376852 140626 376904 140632
rect 376760 139392 376812 139398
rect 376760 139334 376812 139340
rect 375472 138712 375524 138718
rect 375472 138654 375524 138660
rect 431972 132494 432000 180766
rect 441540 154574 441568 190426
rect 441712 181688 441764 181694
rect 441712 181630 441764 181636
rect 441540 154546 441660 154574
rect 431972 132466 432552 132494
rect 375288 129600 375340 129606
rect 375288 129542 375340 129548
rect 375300 129130 375328 129542
rect 375288 129124 375340 129130
rect 375288 129066 375340 129072
rect 429200 129124 429252 129130
rect 429200 129066 429252 129072
rect 374092 125520 374144 125526
rect 374092 125462 374144 125468
rect 429212 125458 429240 129066
rect 430580 129056 430632 129062
rect 430580 128998 430632 129004
rect 429200 125452 429252 125458
rect 429200 125394 429252 125400
rect 430592 125390 430620 128998
rect 430580 125384 430632 125390
rect 430580 125326 430632 125332
rect 372528 125316 372580 125322
rect 372528 125258 372580 125264
rect 372540 125225 372568 125258
rect 372526 125216 372582 125225
rect 372526 125151 372582 125160
rect 372436 124908 372488 124914
rect 372436 124850 372488 124856
rect 372448 124273 372476 124850
rect 432524 124794 432552 132466
rect 441632 125594 441660 154546
rect 441356 125566 441660 125594
rect 441356 124794 441384 125566
rect 432524 124766 432952 124794
rect 440956 124766 441384 124794
rect 372434 124264 372490 124273
rect 372434 124199 372490 124208
rect 371608 124160 371660 124166
rect 371608 124102 371660 124108
rect 434884 124086 435220 124114
rect 436908 124098 437244 124114
rect 436908 124092 437256 124098
rect 436908 124086 437204 124092
rect 370412 123616 370464 123622
rect 370412 123558 370464 123564
rect 435192 122738 435220 124086
rect 437204 124034 437256 124040
rect 438918 123842 438946 124100
rect 438872 123814 438946 123842
rect 438872 122806 438900 123814
rect 438860 122800 438912 122806
rect 438860 122742 438912 122748
rect 441724 122738 441752 181630
rect 441804 153264 441856 153270
rect 441804 153206 441856 153212
rect 441816 149025 441844 153206
rect 441802 149016 441858 149025
rect 441802 148951 441858 148960
rect 441802 129840 441858 129849
rect 441802 129775 441858 129784
rect 441816 126070 441844 129775
rect 442998 129296 443054 129305
rect 442998 129231 443054 129240
rect 441894 126440 441950 126449
rect 441894 126375 441950 126384
rect 441804 126064 441856 126070
rect 441804 126006 441856 126012
rect 441804 125520 441856 125526
rect 441802 125488 441804 125497
rect 441856 125488 441858 125497
rect 441802 125423 441858 125432
rect 441908 125322 441936 126375
rect 443012 125934 443040 129231
rect 443000 125928 443052 125934
rect 443000 125870 443052 125876
rect 441896 125316 441948 125322
rect 441896 125258 441948 125264
rect 441802 124944 441858 124953
rect 441802 124879 441804 124888
rect 441856 124879 441858 124888
rect 441804 124850 441856 124856
rect 443196 124098 443224 194414
rect 444484 156738 444512 205799
rect 444472 156732 444524 156738
rect 444472 156674 444524 156680
rect 444380 153400 444432 153406
rect 444380 153342 444432 153348
rect 444392 147801 444420 153342
rect 444378 147792 444434 147801
rect 444378 147727 444434 147736
rect 444380 146600 444432 146606
rect 444378 146568 444380 146577
rect 444432 146568 444434 146577
rect 444378 146503 444434 146512
rect 444380 136332 444432 136338
rect 444380 136274 444432 136280
rect 444392 136241 444420 136274
rect 444378 136232 444434 136241
rect 444378 136167 444434 136176
rect 444484 133929 444512 156674
rect 444564 155916 444616 155922
rect 444564 155858 444616 155864
rect 444576 154630 444604 155858
rect 444564 154624 444616 154630
rect 444564 154566 444616 154572
rect 444576 140865 444604 154566
rect 444562 140856 444618 140865
rect 444562 140791 444618 140800
rect 444564 136332 444616 136338
rect 444564 136274 444616 136280
rect 444470 133920 444526 133929
rect 444470 133855 444526 133864
rect 444472 133204 444524 133210
rect 444472 133146 444524 133152
rect 444484 132705 444512 133146
rect 444470 132696 444526 132705
rect 444470 132631 444526 132640
rect 443642 128072 443698 128081
rect 443642 128007 443698 128016
rect 443656 127022 443684 128007
rect 443644 127016 443696 127022
rect 443644 126958 443696 126964
rect 443276 126268 443328 126274
rect 443276 126210 443328 126216
rect 443288 125769 443316 126210
rect 443656 126002 443684 126958
rect 443644 125996 443696 126002
rect 443644 125938 443696 125944
rect 443274 125760 443330 125769
rect 443274 125695 443330 125704
rect 444484 124166 444512 132631
rect 444576 125458 444604 136274
rect 444760 135017 444788 206887
rect 445300 205624 445352 205630
rect 445300 205566 445352 205572
rect 445312 204649 445340 205566
rect 445298 204640 445354 204649
rect 445298 204575 445354 204584
rect 445022 203552 445078 203561
rect 445022 203487 445078 203496
rect 445036 202910 445064 203487
rect 445024 202904 445076 202910
rect 445024 202846 445076 202852
rect 445666 202328 445722 202337
rect 445666 202263 445722 202272
rect 445680 201550 445708 202263
rect 445668 201544 445720 201550
rect 445668 201486 445720 201492
rect 445666 201240 445722 201249
rect 445666 201175 445722 201184
rect 445680 200802 445708 201175
rect 445668 200796 445720 200802
rect 445668 200738 445720 200744
rect 445956 200114 445984 258046
rect 446128 218068 446180 218074
rect 446128 218010 446180 218016
rect 446036 211132 446088 211138
rect 446036 211074 446088 211080
rect 446048 210526 446076 211074
rect 446036 210520 446088 210526
rect 446036 210462 446088 210468
rect 445864 200086 445984 200114
rect 445666 200016 445722 200025
rect 445666 199951 445722 199960
rect 445680 199442 445708 199951
rect 445668 199436 445720 199442
rect 445668 199378 445720 199384
rect 445666 198928 445722 198937
rect 445666 198863 445722 198872
rect 445680 198830 445708 198863
rect 445668 198824 445720 198830
rect 445720 198784 445800 198812
rect 445668 198766 445720 198772
rect 445390 197704 445446 197713
rect 445390 197639 445392 197648
rect 445444 197639 445446 197648
rect 445392 197610 445444 197616
rect 444932 154080 444984 154086
rect 444932 154022 444984 154028
rect 444944 153513 444972 154022
rect 444930 153504 444986 153513
rect 444930 153439 444986 153448
rect 445300 153264 445352 153270
rect 445300 153206 445352 153212
rect 444932 151768 444984 151774
rect 444932 151710 444984 151716
rect 444944 151201 444972 151710
rect 444930 151192 444986 151201
rect 444930 151127 444986 151136
rect 444932 150204 444984 150210
rect 444932 150146 444984 150152
rect 444944 150113 444972 150146
rect 444930 150104 444986 150113
rect 444930 150039 444986 150048
rect 445312 149054 445340 153206
rect 445668 153196 445720 153202
rect 445668 153138 445720 153144
rect 445680 152425 445708 153138
rect 445666 152416 445722 152425
rect 445666 152351 445722 152360
rect 445300 149048 445352 149054
rect 445300 148990 445352 148996
rect 445668 146260 445720 146266
rect 445668 146202 445720 146208
rect 445680 145489 445708 146202
rect 445666 145480 445722 145489
rect 445666 145415 445722 145424
rect 445300 144832 445352 144838
rect 445300 144774 445352 144780
rect 445312 144265 445340 144774
rect 445298 144256 445354 144265
rect 445298 144191 445354 144200
rect 445206 143168 445262 143177
rect 445206 143103 445262 143112
rect 445220 142254 445248 143103
rect 445208 142248 445260 142254
rect 445208 142190 445260 142196
rect 445116 141976 445168 141982
rect 445114 141944 445116 141953
rect 445168 141944 445170 141953
rect 445114 141879 445170 141888
rect 445116 140412 445168 140418
rect 445116 140354 445168 140360
rect 445128 139641 445156 140354
rect 445114 139632 445170 139641
rect 445114 139567 445170 139576
rect 444840 137964 444892 137970
rect 444840 137906 444892 137912
rect 444852 137329 444880 137906
rect 444838 137320 444894 137329
rect 444838 137255 444894 137264
rect 444746 135008 444802 135017
rect 444746 134943 444802 134952
rect 444564 125452 444616 125458
rect 444564 125394 444616 125400
rect 444760 125390 444788 134943
rect 445668 132456 445720 132462
rect 445668 132398 445720 132404
rect 445680 131617 445708 132398
rect 445666 131608 445722 131617
rect 445666 131543 445722 131552
rect 444840 130484 444892 130490
rect 444840 130426 444892 130432
rect 444852 130393 444880 130426
rect 444838 130384 444894 130393
rect 444838 130319 444894 130328
rect 444840 129736 444892 129742
rect 444840 129678 444892 129684
rect 444852 129305 444880 129678
rect 444838 129296 444894 129305
rect 444838 129231 444894 129240
rect 445666 126984 445722 126993
rect 445772 126970 445800 198784
rect 445864 196625 445892 200086
rect 445850 196616 445906 196625
rect 445850 196551 445906 196560
rect 445722 126942 445800 126970
rect 445666 126919 445722 126928
rect 444748 125384 444800 125390
rect 444748 125326 444800 125332
rect 445864 124914 445892 196551
rect 446048 161474 446076 210462
rect 446140 168434 446168 218010
rect 446416 201550 446444 274586
rect 447152 208214 447180 277366
rect 447232 270496 447284 270502
rect 447232 270438 447284 270444
rect 447244 269822 447272 270438
rect 447232 269816 447284 269822
rect 447232 269758 447284 269764
rect 447140 208208 447192 208214
rect 447140 208150 447192 208156
rect 446404 201544 446456 201550
rect 446404 201486 446456 201492
rect 446128 168428 446180 168434
rect 446128 168370 446180 168376
rect 445956 161446 446076 161474
rect 445956 160750 445984 161446
rect 445944 160744 445996 160750
rect 445944 160686 445996 160692
rect 445956 138553 445984 160686
rect 446140 146606 446168 168370
rect 446128 146600 446180 146606
rect 446128 146542 446180 146548
rect 445942 138544 445998 138553
rect 445942 138479 445998 138488
rect 447152 136338 447180 208150
rect 447244 197674 447272 269758
rect 447336 212838 447364 284310
rect 447428 270502 447456 341226
rect 447520 276010 447548 346394
rect 448532 286006 448560 357410
rect 448624 291242 448652 362918
rect 448704 352504 448756 352510
rect 448704 352446 448756 352452
rect 448612 291236 448664 291242
rect 448612 291178 448664 291184
rect 448520 286000 448572 286006
rect 448520 285942 448572 285948
rect 447508 276004 447560 276010
rect 447508 275946 447560 275952
rect 447520 275330 447548 275946
rect 447508 275324 447560 275330
rect 447508 275266 447560 275272
rect 447416 270496 447468 270502
rect 447416 270438 447468 270444
rect 448532 213926 448560 285942
rect 448716 281382 448744 352446
rect 449912 295322 449940 367066
rect 452752 364404 452804 364410
rect 452752 364346 452804 364352
rect 449992 360800 450044 360806
rect 449992 360742 450044 360748
rect 449900 295316 449952 295322
rect 449900 295258 449952 295264
rect 449912 294710 449940 295258
rect 449900 294704 449952 294710
rect 449900 294646 449952 294652
rect 448796 294636 448848 294642
rect 448796 294578 448848 294584
rect 448704 281376 448756 281382
rect 448704 281318 448756 281324
rect 448612 222148 448664 222154
rect 448612 222090 448664 222096
rect 448520 213920 448572 213926
rect 448520 213862 448572 213868
rect 447324 212832 447376 212838
rect 447324 212774 447376 212780
rect 447232 197668 447284 197674
rect 447232 197610 447284 197616
rect 447140 136332 447192 136338
rect 447140 136274 447192 136280
rect 447244 126274 447272 197610
rect 447336 155922 447364 212774
rect 448532 158710 448560 213862
rect 448624 175234 448652 222090
rect 448716 209234 448744 281318
rect 448808 222154 448836 294578
rect 450004 289202 450032 360742
rect 452660 360324 452712 360330
rect 452660 360266 452712 360272
rect 450084 355088 450136 355094
rect 450084 355030 450136 355036
rect 449992 289196 450044 289202
rect 449992 289138 450044 289144
rect 449992 287428 450044 287434
rect 449992 287370 450044 287376
rect 450004 287162 450032 287370
rect 449992 287156 450044 287162
rect 449992 287098 450044 287104
rect 449900 225004 449952 225010
rect 449900 224946 449952 224952
rect 448796 222148 448848 222154
rect 448796 222090 448848 222096
rect 448704 209228 448756 209234
rect 448704 209170 448756 209176
rect 448612 175228 448664 175234
rect 448612 175170 448664 175176
rect 448520 158704 448572 158710
rect 448520 158646 448572 158652
rect 447324 155916 447376 155922
rect 447324 155858 447376 155864
rect 448532 141982 448560 158646
rect 448624 150210 448652 175170
rect 448716 164286 448744 209170
rect 448704 164280 448756 164286
rect 448704 164222 448756 164228
rect 448612 150204 448664 150210
rect 448612 150146 448664 150152
rect 448520 141976 448572 141982
rect 448520 141918 448572 141924
rect 448716 137970 448744 164222
rect 449912 154086 449940 224946
rect 450004 216170 450032 287098
rect 450096 283626 450124 355030
rect 451280 343732 451332 343738
rect 451280 343674 451332 343680
rect 450176 297424 450228 297430
rect 450176 297366 450228 297372
rect 450188 297090 450216 297366
rect 450176 297084 450228 297090
rect 450176 297026 450228 297032
rect 450084 283620 450136 283626
rect 450084 283562 450136 283568
rect 449992 216164 450044 216170
rect 449992 216106 450044 216112
rect 450004 215354 450032 216106
rect 449992 215348 450044 215354
rect 449992 215290 450044 215296
rect 450096 211614 450124 283562
rect 450188 225010 450216 297026
rect 451292 272542 451320 343674
rect 452672 287434 452700 360266
rect 452764 293282 452792 364346
rect 452844 345160 452896 345166
rect 452844 345102 452896 345108
rect 452752 293276 452804 293282
rect 452752 293218 452804 293224
rect 452752 291236 452804 291242
rect 452752 291178 452804 291184
rect 452660 287428 452712 287434
rect 452660 287370 452712 287376
rect 452660 287292 452712 287298
rect 452660 287234 452712 287240
rect 451280 272536 451332 272542
rect 451280 272478 451332 272484
rect 451372 270564 451424 270570
rect 451372 270506 451424 270512
rect 450176 225004 450228 225010
rect 450176 224946 450228 224952
rect 450176 215348 450228 215354
rect 450176 215290 450228 215296
rect 450084 211608 450136 211614
rect 450084 211550 450136 211556
rect 450096 200114 450124 211550
rect 450004 200086 450124 200114
rect 450004 167074 450032 200086
rect 450188 172514 450216 215290
rect 451280 201544 451332 201550
rect 451280 201486 451332 201492
rect 450176 172508 450228 172514
rect 450176 172450 450228 172456
rect 449992 167068 450044 167074
rect 449992 167010 450044 167016
rect 449900 154080 449952 154086
rect 449900 154022 449952 154028
rect 450004 140418 450032 167010
rect 450188 161474 450216 172450
rect 450096 161446 450216 161474
rect 450096 144838 450124 161446
rect 450084 144832 450136 144838
rect 450084 144774 450136 144780
rect 449992 140412 450044 140418
rect 449992 140354 450044 140360
rect 448704 137964 448756 137970
rect 448704 137906 448756 137912
rect 451292 130490 451320 201486
rect 451384 198830 451412 270506
rect 452672 214062 452700 287234
rect 452764 219638 452792 291178
rect 452856 274650 452884 345102
rect 454052 297430 454080 368494
rect 456800 365764 456852 365770
rect 456800 365706 456852 365712
rect 454132 361616 454184 361622
rect 454132 361558 454184 361564
rect 454040 297424 454092 297430
rect 454040 297366 454092 297372
rect 454040 294704 454092 294710
rect 454040 294646 454092 294652
rect 452844 274644 452896 274650
rect 452844 274586 452896 274592
rect 453304 273964 453356 273970
rect 453304 273906 453356 273912
rect 452752 219632 452804 219638
rect 452752 219574 452804 219580
rect 452660 214056 452712 214062
rect 452660 213998 452712 214004
rect 452660 199436 452712 199442
rect 452660 199378 452712 199384
rect 451372 198824 451424 198830
rect 451372 198766 451424 198772
rect 451280 130484 451332 130490
rect 451280 130426 451332 130432
rect 452672 127022 452700 199378
rect 452764 153406 452792 219574
rect 452844 214056 452896 214062
rect 452844 213998 452896 214004
rect 452856 164218 452884 213998
rect 453316 200802 453344 273906
rect 454052 223582 454080 294646
rect 454144 290494 454172 361558
rect 454224 347812 454276 347818
rect 454224 347754 454276 347760
rect 454132 290488 454184 290494
rect 454132 290430 454184 290436
rect 454132 289196 454184 289202
rect 454132 289138 454184 289144
rect 454040 223576 454092 223582
rect 454040 223518 454092 223524
rect 453304 200796 453356 200802
rect 453304 200738 453356 200744
rect 452844 164212 452896 164218
rect 452844 164154 452896 164160
rect 452752 153400 452804 153406
rect 452752 153342 452804 153348
rect 452856 142254 452884 164154
rect 454052 151774 454080 223518
rect 454144 217326 454172 289138
rect 454236 276690 454264 347754
rect 456812 294642 456840 365706
rect 456892 345092 456944 345098
rect 456892 345034 456944 345040
rect 456800 294636 456852 294642
rect 456800 294578 456852 294584
rect 456800 293276 456852 293282
rect 456800 293218 456852 293224
rect 454224 276684 454276 276690
rect 454224 276626 454276 276632
rect 454132 217320 454184 217326
rect 454132 217262 454184 217268
rect 454144 162178 454172 217262
rect 454236 205630 454264 276626
rect 456812 220794 456840 293218
rect 456904 273970 456932 345034
rect 458180 342304 458232 342310
rect 458180 342246 458232 342252
rect 456892 273964 456944 273970
rect 456892 273906 456944 273912
rect 456892 272536 456944 272542
rect 456892 272478 456944 272484
rect 456800 220788 456852 220794
rect 456800 220730 456852 220736
rect 454224 205624 454276 205630
rect 454224 205566 454276 205572
rect 454224 204264 454276 204270
rect 454224 204206 454276 204212
rect 454236 202910 454264 204206
rect 454224 202904 454276 202910
rect 454224 202846 454276 202852
rect 454132 162172 454184 162178
rect 454132 162114 454184 162120
rect 454040 151768 454092 151774
rect 454040 151710 454092 151716
rect 454144 146266 454172 162114
rect 454236 159361 454264 202846
rect 456800 200796 456852 200802
rect 456800 200738 456852 200744
rect 454222 159352 454278 159361
rect 454222 159287 454278 159296
rect 454132 146260 454184 146266
rect 454132 146202 454184 146208
rect 452844 142248 452896 142254
rect 452844 142190 452896 142196
rect 454236 132462 454264 159287
rect 454224 132456 454276 132462
rect 454224 132398 454276 132404
rect 456812 129742 456840 200738
rect 456904 199442 456932 272478
rect 458192 270570 458220 342246
rect 479536 305794 479564 700334
rect 479524 305788 479576 305794
rect 479524 305730 479576 305736
rect 494072 304366 494100 703582
rect 494624 703474 494652 703582
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 494808 703474 494836 703520
rect 494624 703446 494836 703474
rect 527192 700398 527220 703520
rect 527180 700392 527232 700398
rect 527180 700334 527232 700340
rect 543476 700330 543504 703520
rect 559668 702434 559696 703520
rect 558932 702406 559696 702434
rect 543464 700324 543516 700330
rect 543464 700266 543516 700272
rect 494060 304360 494112 304366
rect 494060 304302 494112 304308
rect 558932 304298 558960 702406
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 580184 696998 580212 697167
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 580170 683904 580226 683913
rect 580170 683839 580226 683848
rect 580184 683194 580212 683839
rect 580172 683188 580224 683194
rect 580172 683130 580224 683136
rect 580172 670744 580224 670750
rect 580170 670712 580172 670721
rect 580224 670712 580226 670721
rect 580170 670647 580226 670656
rect 580170 644056 580226 644065
rect 580170 643991 580226 644000
rect 580184 643142 580212 643991
rect 580172 643136 580224 643142
rect 580172 643078 580224 643084
rect 580170 630864 580226 630873
rect 580170 630799 580226 630808
rect 580184 630698 580212 630799
rect 580172 630692 580224 630698
rect 580172 630634 580224 630640
rect 580170 617536 580226 617545
rect 580170 617471 580226 617480
rect 580184 616894 580212 617471
rect 580172 616888 580224 616894
rect 580172 616830 580224 616836
rect 579802 591016 579858 591025
rect 579802 590951 579858 590960
rect 579816 590714 579844 590951
rect 579804 590708 579856 590714
rect 579804 590650 579856 590656
rect 580170 577688 580226 577697
rect 580170 577623 580226 577632
rect 580184 576910 580212 577623
rect 580172 576904 580224 576910
rect 580172 576846 580224 576852
rect 579802 564360 579858 564369
rect 579802 564295 579858 564304
rect 579816 563106 579844 564295
rect 579804 563100 579856 563106
rect 579804 563042 579856 563048
rect 580170 537840 580226 537849
rect 580170 537775 580226 537784
rect 580184 536858 580212 537775
rect 580172 536852 580224 536858
rect 580172 536794 580224 536800
rect 580170 524512 580226 524521
rect 580170 524447 580172 524456
rect 580224 524447 580226 524456
rect 580172 524418 580224 524424
rect 580170 511320 580226 511329
rect 580170 511255 580226 511264
rect 580184 510678 580212 511255
rect 580172 510672 580224 510678
rect 580172 510614 580224 510620
rect 580170 484664 580226 484673
rect 580170 484599 580226 484608
rect 580184 484430 580212 484599
rect 580172 484424 580224 484430
rect 580172 484366 580224 484372
rect 579986 471472 580042 471481
rect 579986 471407 580042 471416
rect 580000 470626 580028 471407
rect 579988 470620 580040 470626
rect 579988 470562 580040 470568
rect 580170 458144 580226 458153
rect 580170 458079 580226 458088
rect 580184 456822 580212 458079
rect 580172 456816 580224 456822
rect 580172 456758 580224 456764
rect 580170 431624 580226 431633
rect 580170 431559 580226 431568
rect 580184 430642 580212 431559
rect 580172 430636 580224 430642
rect 580172 430578 580224 430584
rect 580170 418296 580226 418305
rect 580170 418231 580226 418240
rect 580184 418198 580212 418231
rect 580172 418192 580224 418198
rect 580172 418134 580224 418140
rect 580170 404968 580226 404977
rect 580170 404903 580226 404912
rect 580184 404394 580212 404903
rect 580172 404388 580224 404394
rect 580172 404330 580224 404336
rect 582378 378448 582434 378457
rect 582378 378383 582434 378392
rect 580170 325272 580226 325281
rect 580170 325207 580226 325216
rect 580184 324358 580212 325207
rect 580172 324352 580224 324358
rect 580172 324294 580224 324300
rect 580170 312080 580226 312089
rect 580170 312015 580226 312024
rect 580184 311914 580212 312015
rect 580172 311908 580224 311914
rect 580172 311850 580224 311856
rect 582392 305726 582420 378383
rect 582470 365120 582526 365129
rect 582470 365055 582526 365064
rect 582484 307086 582512 365055
rect 582562 351928 582618 351937
rect 582562 351863 582618 351872
rect 582472 307080 582524 307086
rect 582472 307022 582524 307028
rect 582380 305720 582432 305726
rect 582380 305662 582432 305668
rect 582576 305658 582604 351863
rect 582564 305652 582616 305658
rect 582564 305594 582616 305600
rect 558920 304292 558972 304298
rect 558920 304234 558972 304240
rect 582472 303680 582524 303686
rect 582472 303622 582524 303628
rect 548524 303136 548576 303142
rect 548524 303078 548576 303084
rect 458272 295996 458324 296002
rect 458272 295938 458324 295944
rect 458180 270564 458232 270570
rect 458180 270506 458232 270512
rect 458284 224262 458312 295938
rect 458364 275324 458416 275330
rect 458364 275266 458416 275272
rect 458272 224256 458324 224262
rect 458272 224198 458324 224204
rect 456984 220788 457036 220794
rect 456984 220730 457036 220736
rect 456996 220114 457024 220730
rect 456984 220108 457036 220114
rect 456984 220050 457036 220056
rect 456892 199436 456944 199442
rect 456892 199378 456944 199384
rect 456996 149054 457024 220050
rect 458180 205624 458232 205630
rect 458180 205566 458232 205572
rect 456984 149048 457036 149054
rect 456984 148990 457036 148996
rect 458192 133210 458220 205566
rect 458284 153202 458312 224198
rect 458376 204270 458404 275266
rect 458364 204264 458416 204270
rect 458364 204206 458416 204212
rect 458272 153196 458324 153202
rect 458272 153138 458324 153144
rect 548536 139398 548564 303078
rect 582380 300960 582432 300966
rect 582380 300902 582432 300908
rect 579896 299736 579948 299742
rect 579896 299678 579948 299684
rect 579908 298761 579936 299678
rect 580264 298784 580316 298790
rect 579894 298752 579950 298761
rect 580264 298726 580316 298732
rect 579894 298687 579950 298696
rect 579896 273216 579948 273222
rect 579896 273158 579948 273164
rect 579908 272241 579936 273158
rect 579894 272232 579950 272241
rect 579894 272167 579950 272176
rect 580276 258913 580304 298726
rect 580262 258904 580318 258913
rect 580262 258839 580318 258848
rect 580172 245608 580224 245614
rect 580170 245576 580172 245585
rect 580224 245576 580226 245585
rect 580170 245511 580226 245520
rect 579988 233232 580040 233238
rect 579988 233174 580040 233180
rect 580000 232393 580028 233174
rect 579986 232384 580042 232393
rect 579986 232319 580042 232328
rect 580264 228404 580316 228410
rect 580264 228346 580316 228352
rect 579896 219428 579948 219434
rect 579896 219370 579948 219376
rect 579908 219065 579936 219370
rect 579894 219056 579950 219065
rect 579894 218991 579950 219000
rect 580276 192545 580304 228346
rect 580262 192536 580318 192545
rect 580262 192471 580318 192480
rect 580172 179376 580224 179382
rect 580172 179318 580224 179324
rect 580184 179217 580212 179318
rect 580170 179208 580226 179217
rect 580170 179143 580226 179152
rect 579620 156664 579672 156670
rect 579620 156606 579672 156612
rect 579632 152697 579660 156606
rect 579618 152688 579674 152697
rect 579618 152623 579674 152632
rect 548524 139392 548576 139398
rect 580172 139392 580224 139398
rect 548524 139334 548576 139340
rect 580170 139360 580172 139369
rect 580224 139360 580226 139369
rect 580170 139295 580226 139304
rect 458180 133204 458232 133210
rect 458180 133146 458232 133152
rect 456800 129736 456852 129742
rect 456800 129678 456852 129684
rect 452660 127016 452712 127022
rect 452660 126958 452712 126964
rect 447232 126268 447284 126274
rect 447232 126210 447284 126216
rect 445852 124908 445904 124914
rect 445852 124850 445904 124856
rect 444472 124160 444524 124166
rect 444472 124102 444524 124108
rect 443184 124092 443236 124098
rect 443184 124034 443236 124040
rect 435180 122732 435232 122738
rect 435180 122674 435232 122680
rect 441712 122732 441764 122738
rect 441712 122674 441764 122680
rect 370320 121440 370372 121446
rect 370320 121382 370372 121388
rect 369964 118666 370176 118694
rect 369964 111790 369992 118666
rect 579804 113144 579856 113150
rect 579804 113086 579856 113092
rect 579816 112849 579844 113086
rect 579802 112840 579858 112849
rect 579802 112775 579858 112784
rect 369952 111784 370004 111790
rect 369952 111726 370004 111732
rect 369860 102808 369912 102814
rect 369860 102750 369912 102756
rect 316684 100700 316736 100706
rect 316684 100642 316736 100648
rect 580172 100700 580224 100706
rect 580172 100642 580224 100648
rect 339500 100292 339552 100298
rect 339500 100234 339552 100240
rect 323584 100224 323636 100230
rect 323584 100166 323636 100172
rect 316684 99340 316736 99346
rect 316684 99282 316736 99288
rect 316132 87576 316184 87582
rect 316132 87518 316184 87524
rect 314016 87508 314068 87514
rect 314016 87450 314068 87456
rect 313924 60716 313976 60722
rect 313924 60658 313976 60664
rect 312636 24132 312688 24138
rect 312636 24074 312688 24080
rect 314028 3602 314056 87450
rect 316144 16574 316172 87518
rect 316144 16546 316264 16574
rect 312544 3596 312596 3602
rect 312544 3538 312596 3544
rect 313832 3596 313884 3602
rect 313832 3538 313884 3544
rect 314016 3596 314068 3602
rect 314016 3538 314068 3544
rect 315028 3596 315080 3602
rect 315028 3538 315080 3544
rect 312464 598 312676 626
rect 312464 490 312492 598
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312188 462 312492 490
rect 312648 480 312676 598
rect 313844 480 313872 3538
rect 315040 480 315068 3538
rect 316236 480 316264 16546
rect 316696 3602 316724 99282
rect 320180 98184 320232 98190
rect 320180 98126 320232 98132
rect 317420 94444 317472 94450
rect 317420 94386 317472 94392
rect 317432 6914 317460 94386
rect 318064 81184 318116 81190
rect 318064 81126 318116 81132
rect 318076 16574 318104 81126
rect 320192 16574 320220 98126
rect 322204 97980 322256 97986
rect 322204 97922 322256 97928
rect 320824 95736 320876 95742
rect 320824 95678 320876 95684
rect 318076 16546 318196 16574
rect 320192 16546 320496 16574
rect 317432 6886 318104 6914
rect 316684 3596 316736 3602
rect 316684 3538 316736 3544
rect 317328 3460 317380 3466
rect 317328 3402 317380 3408
rect 317340 480 317368 3402
rect 318076 490 318104 6886
rect 318168 3330 318196 16546
rect 318156 3324 318208 3330
rect 318156 3266 318208 3272
rect 319720 3324 319772 3330
rect 319720 3266 319772 3272
rect 318352 598 318564 626
rect 318352 490 318380 598
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318076 462 318380 490
rect 318536 480 318564 598
rect 319732 480 319760 3266
rect 320468 490 320496 16546
rect 320836 3466 320864 95678
rect 321560 90296 321612 90302
rect 321560 90238 321612 90244
rect 321572 16574 321600 90238
rect 321572 16546 322152 16574
rect 320824 3460 320876 3466
rect 320824 3402 320876 3408
rect 320744 598 320956 626
rect 320744 490 320772 598
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320468 462 320772 490
rect 320928 480 320956 598
rect 322124 480 322152 16546
rect 322216 3806 322244 97922
rect 322940 17264 322992 17270
rect 322940 17206 322992 17212
rect 322204 3800 322256 3806
rect 322204 3742 322256 3748
rect 322952 490 322980 17206
rect 323596 3398 323624 100166
rect 324964 99068 325016 99074
rect 324964 99010 325016 99016
rect 324412 95192 324464 95198
rect 324412 95134 324464 95140
rect 323584 3392 323636 3398
rect 323584 3334 323636 3340
rect 323136 598 323348 626
rect 323136 490 323164 598
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 322952 462 323164 490
rect 323320 480 323348 598
rect 324424 480 324452 95134
rect 324976 3262 325004 99010
rect 333980 98116 334032 98122
rect 333980 98058 334032 98064
rect 329104 97912 329156 97918
rect 329104 97854 329156 97860
rect 327080 95124 327132 95130
rect 327080 95066 327132 95072
rect 327092 16574 327120 95066
rect 328460 89684 328512 89690
rect 328460 89626 328512 89632
rect 327724 84040 327776 84046
rect 327724 83982 327776 83988
rect 327092 16546 327672 16574
rect 327644 3482 327672 16546
rect 327736 4010 327764 83982
rect 328472 16574 328500 89626
rect 328472 16546 328776 16574
rect 327724 4004 327776 4010
rect 327724 3946 327776 3952
rect 327644 3454 328040 3482
rect 325608 3392 325660 3398
rect 325608 3334 325660 3340
rect 324964 3256 325016 3262
rect 324964 3198 325016 3204
rect 325620 480 325648 3334
rect 326804 3256 326856 3262
rect 326804 3198 326856 3204
rect 326816 480 326844 3198
rect 328012 480 328040 3454
rect 328748 490 328776 16546
rect 329116 11762 329144 97854
rect 331220 93016 331272 93022
rect 331220 92958 331272 92964
rect 330484 91724 330536 91730
rect 330484 91666 330536 91672
rect 329840 26920 329892 26926
rect 329840 26862 329892 26868
rect 329852 16574 329880 26862
rect 329852 16546 330432 16574
rect 329104 11756 329156 11762
rect 329104 11698 329156 11704
rect 329024 598 329236 626
rect 329024 490 329052 598
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 328748 462 329052 490
rect 329208 480 329236 598
rect 330404 480 330432 16546
rect 330496 3330 330524 91666
rect 330484 3324 330536 3330
rect 330484 3266 330536 3272
rect 331232 490 331260 92958
rect 331864 79756 331916 79762
rect 331864 79698 331916 79704
rect 331876 3398 331904 79698
rect 333992 16574 334020 98058
rect 336004 97844 336056 97850
rect 336004 97786 336056 97792
rect 335360 88324 335412 88330
rect 335360 88266 335412 88272
rect 335372 16574 335400 88266
rect 336016 29646 336044 97786
rect 338120 93084 338172 93090
rect 338120 93026 338172 93032
rect 336096 29708 336148 29714
rect 336096 29650 336148 29656
rect 336004 29640 336056 29646
rect 336004 29582 336056 29588
rect 333992 16546 334664 16574
rect 335372 16546 336044 16574
rect 331864 3392 331916 3398
rect 331864 3334 331916 3340
rect 333888 3392 333940 3398
rect 333888 3334 333940 3340
rect 332692 3324 332744 3330
rect 332692 3266 332744 3272
rect 331416 598 331628 626
rect 331416 490 331444 598
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331232 462 331444 490
rect 331600 480 331628 598
rect 332704 480 332732 3266
rect 333900 480 333928 3334
rect 334636 490 334664 16546
rect 336016 3210 336044 16546
rect 336108 3330 336136 29650
rect 338132 16574 338160 93026
rect 338132 16546 338712 16574
rect 336096 3324 336148 3330
rect 336096 3266 336148 3272
rect 337476 3324 337528 3330
rect 337476 3266 337528 3272
rect 336016 3182 336320 3210
rect 334912 598 335124 626
rect 334912 490 334940 598
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 334636 462 334940 490
rect 335096 480 335124 598
rect 336292 480 336320 3182
rect 337488 480 337516 3266
rect 338684 480 338712 16546
rect 339512 490 339540 100234
rect 353944 100156 353996 100162
rect 353944 100098 353996 100104
rect 342904 97776 342956 97782
rect 342904 97718 342956 97724
rect 340880 95056 340932 95062
rect 340880 94998 340932 95004
rect 340892 3398 340920 94998
rect 342916 86970 342944 97718
rect 347044 96484 347096 96490
rect 347044 96426 347096 96432
rect 345020 93832 345072 93838
rect 345020 93774 345072 93780
rect 342260 86964 342312 86970
rect 342260 86906 342312 86912
rect 342904 86964 342956 86970
rect 342904 86906 342956 86912
rect 340972 78328 341024 78334
rect 340972 78270 341024 78276
rect 340880 3392 340932 3398
rect 340880 3334 340932 3340
rect 339696 598 339908 626
rect 339696 490 339724 598
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339512 462 339724 490
rect 339880 480 339908 598
rect 340984 480 341012 78270
rect 342272 6914 342300 86906
rect 342904 28280 342956 28286
rect 342904 28222 342956 28228
rect 342916 16574 342944 28222
rect 345032 16574 345060 93774
rect 346400 86896 346452 86902
rect 346400 86838 346452 86844
rect 346412 16574 346440 86838
rect 342916 16546 343036 16574
rect 345032 16546 345336 16574
rect 346412 16546 346992 16574
rect 342272 6886 342944 6914
rect 342168 3392 342220 3398
rect 342168 3334 342220 3340
rect 342180 480 342208 3334
rect 342916 490 342944 6886
rect 343008 3058 343036 16546
rect 342996 3052 343048 3058
rect 342996 2994 343048 3000
rect 344560 3052 344612 3058
rect 344560 2994 344612 3000
rect 343192 598 343404 626
rect 343192 490 343220 598
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 342916 462 343220 490
rect 343376 480 343404 598
rect 344572 480 344600 2994
rect 345308 490 345336 16546
rect 345584 598 345796 626
rect 345584 490 345612 598
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345308 462 345612 490
rect 345768 480 345796 598
rect 346964 480 346992 16546
rect 347056 4078 347084 96426
rect 351920 93764 351972 93770
rect 351920 93706 351972 93712
rect 347780 79688 347832 79694
rect 347780 79630 347832 79636
rect 347792 16574 347820 79630
rect 351932 16574 351960 93706
rect 353300 88256 353352 88262
rect 353300 88198 353352 88204
rect 353312 16574 353340 88198
rect 347792 16546 348096 16574
rect 351932 16546 352880 16574
rect 353312 16546 353616 16574
rect 347044 4072 347096 4078
rect 347044 4014 347096 4020
rect 348068 480 348096 16546
rect 351644 4004 351696 4010
rect 351644 3946 351696 3952
rect 350446 3496 350502 3505
rect 350446 3431 350502 3440
rect 349250 3360 349306 3369
rect 349250 3295 349306 3304
rect 349264 480 349292 3295
rect 350460 480 350488 3431
rect 351656 480 351684 3946
rect 352852 480 352880 16546
rect 353588 490 353616 16546
rect 353956 4146 353984 100098
rect 376024 100020 376076 100026
rect 376024 99962 376076 99968
rect 360844 99000 360896 99006
rect 360844 98942 360896 98948
rect 358820 98048 358872 98054
rect 358820 97990 358872 97996
rect 356060 96552 356112 96558
rect 356060 96494 356112 96500
rect 356072 16574 356100 96494
rect 357440 86760 357492 86766
rect 357440 86702 357492 86708
rect 356072 16546 356376 16574
rect 353944 4140 353996 4146
rect 353944 4082 353996 4088
rect 355232 4140 355284 4146
rect 355232 4082 355284 4088
rect 353864 598 354076 626
rect 353864 490 353892 598
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 353588 462 353892 490
rect 354048 480 354076 598
rect 355244 480 355272 4082
rect 356348 480 356376 16546
rect 357452 6914 357480 86702
rect 357532 78260 357584 78266
rect 357532 78202 357584 78208
rect 357544 11830 357572 78202
rect 358832 16574 358860 97990
rect 360200 85468 360252 85474
rect 360200 85410 360252 85416
rect 360212 16574 360240 85410
rect 358832 16546 359504 16574
rect 360212 16546 360792 16574
rect 357532 11824 357584 11830
rect 357532 11766 357584 11772
rect 358728 11824 358780 11830
rect 358728 11766 358780 11772
rect 357452 6886 357572 6914
rect 357544 480 357572 6886
rect 358740 480 358768 11766
rect 359476 490 359504 16546
rect 360764 3482 360792 16546
rect 360856 4010 360884 98942
rect 364984 94988 365036 94994
rect 364984 94930 365036 94936
rect 362960 93696 363012 93702
rect 362960 93638 363012 93644
rect 362972 16574 363000 93638
rect 364340 85400 364392 85406
rect 364340 85342 364392 85348
rect 364352 16574 364380 85342
rect 362972 16546 363552 16574
rect 364352 16546 364656 16574
rect 362316 4072 362368 4078
rect 362316 4014 362368 4020
rect 360844 4004 360896 4010
rect 360844 3946 360896 3952
rect 360764 3454 361160 3482
rect 359752 598 359964 626
rect 359752 490 359780 598
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359476 462 359780 490
rect 359936 480 359964 598
rect 361132 480 361160 3454
rect 362328 480 362356 4014
rect 363524 480 363552 16546
rect 364628 480 364656 16546
rect 364996 3398 365024 94930
rect 369860 92472 369912 92478
rect 369860 92414 369912 92420
rect 365812 86828 365864 86834
rect 365812 86770 365864 86776
rect 364984 3392 365036 3398
rect 364984 3334 365036 3340
rect 365824 480 365852 86770
rect 367100 85332 367152 85338
rect 367100 85274 367152 85280
rect 367112 16574 367140 85274
rect 369872 16574 369900 92414
rect 374644 92404 374696 92410
rect 374644 92346 374696 92352
rect 374092 83972 374144 83978
rect 374092 83914 374144 83920
rect 374104 16574 374132 83914
rect 367112 16546 367784 16574
rect 369872 16546 370176 16574
rect 374104 16546 374592 16574
rect 367008 3392 367060 3398
rect 367008 3334 367060 3340
rect 367020 480 367048 3334
rect 367756 490 367784 16546
rect 369400 4004 369452 4010
rect 369400 3946 369452 3952
rect 368032 598 368244 626
rect 368032 490 368060 598
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 367756 462 368060 490
rect 368216 480 368244 598
rect 369412 480 369440 3946
rect 370148 490 370176 16546
rect 372896 4956 372948 4962
rect 372896 4898 372948 4904
rect 371700 3936 371752 3942
rect 371700 3878 371752 3884
rect 370424 598 370636 626
rect 370424 490 370452 598
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370148 462 370452 490
rect 370608 480 370636 598
rect 371712 480 371740 3878
rect 372908 480 372936 4898
rect 374092 3732 374144 3738
rect 374092 3674 374144 3680
rect 374104 480 374132 3674
rect 374564 2938 374592 16546
rect 374656 3058 374684 92346
rect 375380 18624 375432 18630
rect 375380 18566 375432 18572
rect 375392 6914 375420 18566
rect 376036 16574 376064 99962
rect 412640 99952 412692 99958
rect 412640 99894 412692 99900
rect 393964 97708 394016 97714
rect 393964 97650 394016 97656
rect 385684 94920 385736 94926
rect 385684 94862 385736 94868
rect 378784 93628 378836 93634
rect 378784 93570 378836 93576
rect 377404 89616 377456 89622
rect 377404 89558 377456 89564
rect 376036 16546 376156 16574
rect 375392 6886 376064 6914
rect 374644 3052 374696 3058
rect 374644 2994 374696 3000
rect 374564 2910 375328 2938
rect 375300 480 375328 2910
rect 376036 490 376064 6886
rect 376128 3330 376156 16546
rect 377416 4010 377444 89558
rect 378140 83904 378192 83910
rect 378140 83846 378192 83852
rect 378152 16574 378180 83846
rect 378152 16546 378456 16574
rect 377404 4004 377456 4010
rect 377404 3946 377456 3952
rect 376116 3324 376168 3330
rect 376116 3266 376168 3272
rect 377680 3052 377732 3058
rect 377680 2994 377732 3000
rect 376312 598 376524 626
rect 376312 490 376340 598
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376036 462 376340 490
rect 376496 480 376524 598
rect 377692 480 377720 2994
rect 378428 490 378456 16546
rect 378796 3398 378824 93570
rect 381544 92336 381596 92342
rect 381544 92278 381596 92284
rect 381556 3738 381584 92278
rect 382924 92200 382976 92206
rect 382924 92142 382976 92148
rect 382372 85264 382424 85270
rect 382372 85206 382424 85212
rect 381544 3732 381596 3738
rect 381544 3674 381596 3680
rect 378784 3392 378836 3398
rect 378784 3334 378836 3340
rect 381176 3392 381228 3398
rect 381176 3334 381228 3340
rect 379980 3324 380032 3330
rect 379980 3266 380032 3272
rect 378704 598 378916 626
rect 378704 490 378732 598
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378428 462 378732 490
rect 378888 480 378916 598
rect 379992 480 380020 3266
rect 381188 480 381216 3334
rect 382384 480 382412 85206
rect 382936 4146 382964 92142
rect 385040 83836 385092 83842
rect 385040 83778 385092 83784
rect 385052 16574 385080 83778
rect 385052 16546 385632 16574
rect 382924 4140 382976 4146
rect 382924 4082 382976 4088
rect 384764 4140 384816 4146
rect 384764 4082 384816 4088
rect 383568 3868 383620 3874
rect 383568 3810 383620 3816
rect 383580 480 383608 3810
rect 384776 480 384804 4082
rect 385604 3482 385632 16546
rect 385696 3942 385724 94862
rect 387800 92132 387852 92138
rect 387800 92074 387852 92080
rect 387156 4004 387208 4010
rect 387156 3946 387208 3952
rect 385684 3936 385736 3942
rect 385684 3878 385736 3884
rect 385604 3454 386000 3482
rect 385972 480 386000 3454
rect 387168 480 387196 3946
rect 387812 490 387840 92074
rect 389824 92064 389876 92070
rect 389824 92006 389876 92012
rect 389836 3398 389864 92006
rect 392032 86692 392084 86698
rect 392032 86634 392084 86640
rect 391940 83768 391992 83774
rect 391940 83710 391992 83716
rect 390652 4888 390704 4894
rect 390652 4830 390704 4836
rect 389824 3392 389876 3398
rect 389824 3334 389876 3340
rect 389456 3188 389508 3194
rect 389456 3130 389508 3136
rect 388088 598 388300 626
rect 388088 490 388116 598
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 387812 462 388116 490
rect 388272 480 388300 598
rect 389468 480 389496 3130
rect 390664 480 390692 4830
rect 391848 3392 391900 3398
rect 391848 3334 391900 3340
rect 391860 480 391888 3334
rect 391952 2530 391980 83710
rect 392044 3194 392072 86634
rect 393320 24132 393372 24138
rect 393320 24074 393372 24080
rect 393332 6914 393360 24074
rect 393976 8294 394004 97650
rect 400864 97640 400916 97646
rect 400864 97582 400916 97588
rect 398840 93560 398892 93566
rect 398840 93502 398892 93508
rect 394700 91044 394752 91050
rect 394700 90986 394752 90992
rect 394712 16574 394740 90986
rect 396724 90976 396776 90982
rect 396724 90918 396776 90924
rect 396080 83700 396132 83706
rect 396080 83642 396132 83648
rect 394712 16546 395384 16574
rect 393964 8288 394016 8294
rect 393964 8230 394016 8236
rect 393332 6886 394280 6914
rect 392032 3188 392084 3194
rect 392032 3130 392084 3136
rect 391952 2502 392624 2530
rect 392596 490 392624 2502
rect 392872 598 393084 626
rect 392872 490 392900 598
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 392596 462 392900 490
rect 393056 480 393084 598
rect 394252 480 394280 6886
rect 395356 480 395384 16546
rect 396092 490 396120 83642
rect 396736 3398 396764 90918
rect 398852 6914 398880 93502
rect 398932 82612 398984 82618
rect 398932 82554 398984 82560
rect 398944 11830 398972 82554
rect 398932 11824 398984 11830
rect 398932 11766 398984 11772
rect 400128 11824 400180 11830
rect 400128 11766 400180 11772
rect 398852 6886 398972 6914
rect 397736 3732 397788 3738
rect 397736 3674 397788 3680
rect 396724 3392 396776 3398
rect 396724 3334 396776 3340
rect 396368 598 396580 626
rect 396368 490 396396 598
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396092 462 396396 490
rect 396552 480 396580 598
rect 397748 480 397776 3674
rect 398944 480 398972 6886
rect 400140 480 400168 11766
rect 400876 7614 400904 97582
rect 411904 96416 411956 96422
rect 411904 96358 411956 96364
rect 405740 91996 405792 92002
rect 405740 91938 405792 91944
rect 402980 85196 403032 85202
rect 402980 85138 403032 85144
rect 402992 16574 403020 85138
rect 404360 32428 404412 32434
rect 404360 32370 404412 32376
rect 402992 16546 403664 16574
rect 401324 8288 401376 8294
rect 401324 8230 401376 8236
rect 400864 7608 400916 7614
rect 400864 7550 400916 7556
rect 401336 480 401364 8230
rect 402520 3392 402572 3398
rect 402520 3334 402572 3340
rect 402532 480 402560 3334
rect 403636 480 403664 16546
rect 404372 490 404400 32370
rect 405752 16574 405780 91938
rect 407764 90908 407816 90914
rect 407764 90850 407816 90856
rect 405752 16546 406056 16574
rect 404648 598 404860 626
rect 404648 490 404676 598
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404372 462 404676 490
rect 404832 480 404860 598
rect 406028 480 406056 16546
rect 407776 3398 407804 90850
rect 409972 83632 410024 83638
rect 409972 83574 410024 83580
rect 409880 82544 409932 82550
rect 409880 82486 409932 82492
rect 408408 7608 408460 7614
rect 408408 7550 408460 7556
rect 407764 3392 407816 3398
rect 407764 3334 407816 3340
rect 407212 3324 407264 3330
rect 407212 3266 407264 3272
rect 407224 480 407252 3266
rect 408420 480 408448 7550
rect 409604 3392 409656 3398
rect 409604 3334 409656 3340
rect 409616 480 409644 3334
rect 409892 3210 409920 82486
rect 409984 3330 410012 83574
rect 411260 76764 411312 76770
rect 411260 76706 411312 76712
rect 411272 16574 411300 76706
rect 411272 16546 411852 16574
rect 411824 3482 411852 16546
rect 411916 3874 411944 96358
rect 411904 3868 411956 3874
rect 411904 3810 411956 3816
rect 411824 3454 411944 3482
rect 409972 3324 410024 3330
rect 409972 3266 410024 3272
rect 409892 3182 410840 3210
rect 410812 480 410840 3182
rect 411916 480 411944 3454
rect 412652 490 412680 99894
rect 414664 99884 414716 99890
rect 414664 99826 414716 99832
rect 414020 82476 414072 82482
rect 414020 82418 414072 82424
rect 414032 16574 414060 82418
rect 414032 16546 414336 16574
rect 412928 598 413140 626
rect 412928 490 412956 598
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 412652 462 412956 490
rect 413112 480 413140 598
rect 414308 480 414336 16546
rect 414676 3398 414704 99826
rect 423680 99816 423732 99822
rect 423680 99758 423732 99764
rect 418160 92268 418212 92274
rect 418160 92210 418212 92216
rect 417424 90840 417476 90846
rect 417424 90782 417476 90788
rect 416780 81116 416832 81122
rect 416780 81058 416832 81064
rect 416792 6914 416820 81058
rect 417436 16574 417464 90782
rect 418172 16574 418200 92210
rect 421564 91928 421616 91934
rect 421564 91870 421616 91876
rect 420920 88120 420972 88126
rect 420920 88062 420972 88068
rect 417436 16546 417556 16574
rect 418172 16546 418568 16574
rect 416792 6886 417464 6914
rect 415492 3800 415544 3806
rect 415492 3742 415544 3748
rect 414664 3392 414716 3398
rect 414664 3334 414716 3340
rect 415504 480 415532 3742
rect 416688 3392 416740 3398
rect 416688 3334 416740 3340
rect 416700 480 416728 3334
rect 417436 490 417464 6886
rect 417528 2922 417556 16546
rect 417516 2916 417568 2922
rect 417516 2858 417568 2864
rect 417712 598 417924 626
rect 417712 490 417740 598
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417436 462 417740 490
rect 417896 480 417924 598
rect 418540 490 418568 16546
rect 420184 2916 420236 2922
rect 420184 2858 420236 2864
rect 418816 598 419028 626
rect 418816 490 418844 598
rect 417854 -960 417966 480
rect 418540 462 418844 490
rect 419000 480 419028 598
rect 420196 480 420224 2858
rect 420932 490 420960 88062
rect 421576 3738 421604 91870
rect 422576 11756 422628 11762
rect 422576 11698 422628 11704
rect 421564 3732 421616 3738
rect 421564 3674 421616 3680
rect 421208 598 421420 626
rect 421208 490 421236 598
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 420932 462 421236 490
rect 421392 480 421420 598
rect 422588 480 422616 11698
rect 423692 6914 423720 99758
rect 430580 99748 430632 99754
rect 430580 99690 430632 99696
rect 429844 94852 429896 94858
rect 429844 94794 429896 94800
rect 428464 88188 428516 88194
rect 428464 88130 428516 88136
rect 425060 86964 425112 86970
rect 425060 86906 425112 86912
rect 423772 82408 423824 82414
rect 423772 82350 423824 82356
rect 423784 11762 423812 82350
rect 425072 16574 425100 86906
rect 427820 81048 427872 81054
rect 427820 80990 427872 80996
rect 427832 16574 427860 80990
rect 425072 16546 425744 16574
rect 427832 16546 428412 16574
rect 423772 11756 423824 11762
rect 423772 11698 423824 11704
rect 424968 11756 425020 11762
rect 424968 11698 425020 11704
rect 423692 6886 423812 6914
rect 423784 480 423812 6886
rect 424980 480 425008 11698
rect 425716 490 425744 16546
rect 427268 3732 427320 3738
rect 427268 3674 427320 3680
rect 425992 598 426204 626
rect 425992 490 426020 598
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 425716 462 426020 490
rect 426176 480 426204 598
rect 427280 480 427308 3674
rect 428384 3482 428412 16546
rect 428476 3738 428504 88130
rect 429200 75336 429252 75342
rect 429200 75278 429252 75284
rect 428464 3732 428516 3738
rect 428464 3674 428516 3680
rect 428384 3454 428504 3482
rect 428476 480 428504 3454
rect 429212 490 429240 75278
rect 429856 3806 429884 94794
rect 430592 16574 430620 99690
rect 435364 99680 435416 99686
rect 435364 99622 435416 99628
rect 432604 90772 432656 90778
rect 432604 90714 432656 90720
rect 432052 83564 432104 83570
rect 432052 83506 432104 83512
rect 430592 16546 430896 16574
rect 429844 3800 429896 3806
rect 429844 3742 429896 3748
rect 429488 598 429700 626
rect 429488 490 429516 598
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429212 462 429516 490
rect 429672 480 429700 598
rect 430868 480 430896 16546
rect 432064 480 432092 83506
rect 432616 2922 432644 90714
rect 434720 80980 434772 80986
rect 434720 80922 434772 80928
rect 434732 16574 434760 80922
rect 434732 16546 435128 16574
rect 433248 3664 433300 3670
rect 433248 3606 433300 3612
rect 432604 2916 432656 2922
rect 432604 2858 432656 2864
rect 433260 480 433288 3606
rect 434444 2916 434496 2922
rect 434444 2858 434496 2864
rect 434456 480 434484 2858
rect 435100 490 435128 16546
rect 435376 2990 435404 99622
rect 440240 99612 440292 99618
rect 440240 99554 440292 99560
rect 436744 97572 436796 97578
rect 436744 97514 436796 97520
rect 436100 29640 436152 29646
rect 436100 29582 436152 29588
rect 436112 16574 436140 29582
rect 436756 17270 436784 97514
rect 438860 89548 438912 89554
rect 438860 89490 438912 89496
rect 436744 17264 436796 17270
rect 436744 17206 436796 17212
rect 438872 16574 438900 89490
rect 436112 16546 436784 16574
rect 438872 16546 439176 16574
rect 435364 2984 435416 2990
rect 435364 2926 435416 2932
rect 435376 598 435588 626
rect 435376 490 435404 598
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435100 462 435404 490
rect 435560 480 435588 598
rect 436756 480 436784 16546
rect 437940 2984 437992 2990
rect 437940 2926 437992 2932
rect 437952 480 437980 2926
rect 439148 480 439176 16546
rect 440252 3398 440280 99554
rect 442264 99544 442316 99550
rect 580184 99521 580212 100642
rect 442264 99486 442316 99492
rect 580170 99512 580226 99521
rect 441620 86624 441672 86630
rect 441620 86566 441672 86572
rect 440332 33788 440384 33794
rect 440332 33730 440384 33736
rect 440240 3392 440292 3398
rect 440240 3334 440292 3340
rect 440344 480 440372 33730
rect 441632 6914 441660 86566
rect 442276 16574 442304 99486
rect 457444 99476 457496 99482
rect 580170 99447 580226 99456
rect 457444 99418 457496 99424
rect 443644 97504 443696 97510
rect 443644 97446 443696 97452
rect 443000 17264 443052 17270
rect 443000 17206 443052 17212
rect 443012 16574 443040 17206
rect 442276 16546 442396 16574
rect 443012 16546 443408 16574
rect 441632 6886 442304 6914
rect 441528 3392 441580 3398
rect 441528 3334 441580 3340
rect 441540 480 441568 3334
rect 442276 2802 442304 6886
rect 442368 2922 442396 16546
rect 442356 2916 442408 2922
rect 442356 2858 442408 2864
rect 442276 2774 442672 2802
rect 442644 480 442672 2774
rect 443380 490 443408 16546
rect 443656 8294 443684 97446
rect 447784 97436 447836 97442
rect 447784 97378 447836 97384
rect 446404 90704 446456 90710
rect 446404 90646 446456 90652
rect 445760 82340 445812 82346
rect 445760 82282 445812 82288
rect 443644 8288 443696 8294
rect 443644 8230 443696 8236
rect 445024 2916 445076 2922
rect 445024 2858 445076 2864
rect 443656 598 443868 626
rect 443656 490 443684 598
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443380 462 443684 490
rect 443840 480 443868 598
rect 445036 480 445064 2858
rect 445772 490 445800 82282
rect 446416 3058 446444 90646
rect 447416 3936 447468 3942
rect 447416 3878 447468 3884
rect 446404 3052 446456 3058
rect 446404 2994 446456 3000
rect 446048 598 446260 626
rect 446048 490 446076 598
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 445772 462 446076 490
rect 446232 480 446260 598
rect 447428 480 447456 3878
rect 447796 3670 447824 97378
rect 450544 97368 450596 97374
rect 450544 97310 450596 97316
rect 448520 93492 448572 93498
rect 448520 93434 448572 93440
rect 448532 6914 448560 93434
rect 448612 79620 448664 79626
rect 448612 79562 448664 79568
rect 448624 11762 448652 79562
rect 448612 11756 448664 11762
rect 448612 11698 448664 11704
rect 449808 11756 449860 11762
rect 449808 11698 449860 11704
rect 448532 6886 448652 6914
rect 447784 3664 447836 3670
rect 447784 3606 447836 3612
rect 448624 480 448652 6886
rect 449820 480 449848 11698
rect 450556 7614 450584 97310
rect 454684 97300 454736 97306
rect 454684 97242 454736 97248
rect 453304 94784 453356 94790
rect 453304 94726 453356 94732
rect 452660 85128 452712 85134
rect 452660 85070 452712 85076
rect 452672 16574 452700 85070
rect 452672 16546 453252 16574
rect 450912 8288 450964 8294
rect 450912 8230 450964 8236
rect 450544 7608 450596 7614
rect 450544 7550 450596 7556
rect 450924 480 450952 8230
rect 453224 3346 453252 16546
rect 453316 3466 453344 94726
rect 454040 69692 454092 69698
rect 454040 69634 454092 69640
rect 453304 3460 453356 3466
rect 453304 3402 453356 3408
rect 453224 3318 453344 3346
rect 452108 3052 452160 3058
rect 452108 2994 452160 3000
rect 452120 480 452148 2994
rect 453316 480 453344 3318
rect 454052 490 454080 69634
rect 454696 17270 454724 97242
rect 456892 82272 456944 82278
rect 456892 82214 456944 82220
rect 454684 17264 454736 17270
rect 454684 17206 454736 17212
rect 455696 3460 455748 3466
rect 455696 3402 455748 3408
rect 454328 598 454540 626
rect 454328 490 454356 598
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454052 462 454356 490
rect 454512 480 454540 598
rect 455708 480 455736 3402
rect 456904 480 456932 82214
rect 457456 3466 457484 99418
rect 464344 99408 464396 99414
rect 464344 99350 464396 99356
rect 458822 98968 458878 98977
rect 458822 98903 458878 98912
rect 460204 98932 460256 98938
rect 458836 3670 458864 98903
rect 460204 98874 460256 98880
rect 459560 80912 459612 80918
rect 459560 80854 459612 80860
rect 459572 16574 459600 80854
rect 459572 16546 459968 16574
rect 458088 3664 458140 3670
rect 458088 3606 458140 3612
rect 458824 3664 458876 3670
rect 458824 3606 458876 3612
rect 457444 3460 457496 3466
rect 457444 3402 457496 3408
rect 458100 480 458128 3606
rect 459192 3460 459244 3466
rect 459192 3402 459244 3408
rect 459204 480 459232 3402
rect 459940 490 459968 16546
rect 460216 4146 460244 98874
rect 461582 97472 461638 97481
rect 461582 97407 461638 97416
rect 461596 16574 461624 97407
rect 461596 16546 461716 16574
rect 460204 4140 460256 4146
rect 460204 4082 460256 4088
rect 461584 3528 461636 3534
rect 461584 3470 461636 3476
rect 460216 598 460428 626
rect 460216 490 460244 598
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 459940 462 460244 490
rect 460400 480 460428 598
rect 461596 480 461624 3470
rect 461688 3398 461716 16546
rect 462780 4140 462832 4146
rect 462780 4082 462832 4088
rect 461676 3392 461728 3398
rect 461676 3334 461728 3340
rect 462792 480 462820 4082
rect 463976 3800 464028 3806
rect 463976 3742 464028 3748
rect 463988 480 464016 3742
rect 464356 3534 464384 99350
rect 485044 98864 485096 98870
rect 485044 98806 485096 98812
rect 543738 98832 543794 98841
rect 465724 96348 465776 96354
rect 465724 96290 465776 96296
rect 465172 7608 465224 7614
rect 465172 7550 465224 7556
rect 464344 3528 464396 3534
rect 464344 3470 464396 3476
rect 465184 480 465212 7550
rect 465736 3806 465764 96290
rect 475384 96280 475436 96286
rect 475384 96222 475436 96228
rect 466460 93424 466512 93430
rect 466460 93366 466512 93372
rect 466472 6914 466500 93366
rect 471244 91860 471296 91866
rect 471244 91802 471296 91808
rect 467104 90636 467156 90642
rect 467104 90578 467156 90584
rect 467116 16574 467144 90578
rect 470600 83496 470652 83502
rect 470600 83438 470652 83444
rect 467840 73908 467892 73914
rect 467840 73850 467892 73856
rect 467852 16574 467880 73850
rect 467116 16546 467236 16574
rect 467852 16546 468248 16574
rect 466472 6886 467144 6914
rect 465724 3800 465776 3806
rect 465724 3742 465776 3748
rect 466276 3528 466328 3534
rect 466276 3470 466328 3476
rect 466288 480 466316 3470
rect 467116 3210 467144 6886
rect 467208 3330 467236 16546
rect 467196 3324 467248 3330
rect 467196 3266 467248 3272
rect 467116 3182 467512 3210
rect 467484 480 467512 3182
rect 468220 490 468248 16546
rect 469864 3324 469916 3330
rect 469864 3266 469916 3272
rect 468496 598 468708 626
rect 468496 490 468524 598
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468220 462 468524 490
rect 468680 480 468708 598
rect 469876 480 469904 3266
rect 470612 490 470640 83438
rect 471256 2922 471284 91802
rect 472624 79552 472676 79558
rect 472624 79494 472676 79500
rect 471980 17264 472032 17270
rect 471980 17206 472032 17212
rect 471992 16574 472020 17206
rect 471992 16546 472296 16574
rect 471244 2916 471296 2922
rect 471244 2858 471296 2864
rect 470888 598 471100 626
rect 470888 490 470916 598
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 470612 462 470916 490
rect 471072 480 471100 598
rect 472268 480 472296 16546
rect 472636 3534 472664 79494
rect 474740 31068 474792 31074
rect 474740 31010 474792 31016
rect 474752 6914 474780 31010
rect 475396 16574 475424 96222
rect 479524 96212 479576 96218
rect 479524 96154 479576 96160
rect 476120 89480 476172 89486
rect 476120 89422 476172 89428
rect 476132 16574 476160 89422
rect 477500 80844 477552 80850
rect 477500 80786 477552 80792
rect 477512 16574 477540 80786
rect 475396 16546 475516 16574
rect 476132 16546 476528 16574
rect 477512 16546 478184 16574
rect 474752 6886 475424 6914
rect 472624 3528 472676 3534
rect 472624 3470 472676 3476
rect 474556 3528 474608 3534
rect 474556 3470 474608 3476
rect 475396 3482 475424 6886
rect 475488 3942 475516 16546
rect 475476 3936 475528 3942
rect 475476 3878 475528 3884
rect 473452 2916 473504 2922
rect 473452 2858 473504 2864
rect 473464 480 473492 2858
rect 474568 480 474596 3470
rect 475396 3454 475792 3482
rect 475764 480 475792 3454
rect 476500 490 476528 16546
rect 476776 598 476988 626
rect 476776 490 476804 598
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476500 462 476804 490
rect 476960 480 476988 598
rect 478156 480 478184 16546
rect 479536 4146 479564 96154
rect 483020 96076 483072 96082
rect 483020 96018 483072 96024
rect 481640 89412 481692 89418
rect 481640 89354 481692 89360
rect 481652 6914 481680 89354
rect 481732 79484 481784 79490
rect 481732 79426 481784 79432
rect 481744 16574 481772 79426
rect 483032 16574 483060 96018
rect 481744 16546 482416 16574
rect 483032 16546 484072 16574
rect 481652 6886 481772 6914
rect 479524 4140 479576 4146
rect 479524 4082 479576 4088
rect 480536 4140 480588 4146
rect 480536 4082 480588 4088
rect 479340 3392 479392 3398
rect 479340 3334 479392 3340
rect 479352 480 479380 3334
rect 480548 480 480576 4082
rect 481744 480 481772 6886
rect 482388 490 482416 16546
rect 482664 598 482876 626
rect 482664 490 482692 598
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482388 462 482692 490
rect 482848 480 482876 598
rect 484044 480 484072 16546
rect 485056 3534 485084 98806
rect 507860 98796 507912 98802
rect 543738 98767 543794 98776
rect 507860 98738 507912 98744
rect 494060 96144 494112 96150
rect 494060 96086 494112 96092
rect 489184 94716 489236 94722
rect 489184 94658 489236 94664
rect 486424 90568 486476 90574
rect 486424 90510 486476 90516
rect 485780 82204 485832 82210
rect 485780 82146 485832 82152
rect 485792 16574 485820 82146
rect 485792 16546 486372 16574
rect 485228 3596 485280 3602
rect 485228 3538 485280 3544
rect 485044 3528 485096 3534
rect 485044 3470 485096 3476
rect 485240 480 485268 3538
rect 486344 3346 486372 16546
rect 486436 3534 486464 90510
rect 487620 3936 487672 3942
rect 487620 3878 487672 3884
rect 486424 3528 486476 3534
rect 486424 3470 486476 3476
rect 486344 3318 486464 3346
rect 486436 480 486464 3318
rect 487632 480 487660 3878
rect 489196 3602 489224 94658
rect 490564 89344 490616 89350
rect 490564 89286 490616 89292
rect 490012 78192 490064 78198
rect 490012 78134 490064 78140
rect 490024 6914 490052 78134
rect 489932 6886 490052 6914
rect 489184 3596 489236 3602
rect 489184 3538 489236 3544
rect 488816 3528 488868 3534
rect 488816 3470 488868 3476
rect 488828 480 488856 3470
rect 489932 480 489960 6886
rect 490576 3398 490604 89286
rect 493324 89276 493376 89282
rect 493324 89218 493376 89224
rect 492680 78124 492732 78130
rect 492680 78066 492732 78072
rect 492692 16574 492720 78066
rect 492692 16546 493088 16574
rect 491116 3868 491168 3874
rect 491116 3810 491168 3816
rect 490564 3392 490616 3398
rect 490564 3334 490616 3340
rect 491128 480 491156 3810
rect 492312 3392 492364 3398
rect 492312 3334 492364 3340
rect 492324 480 492352 3334
rect 493060 490 493088 16546
rect 493336 3058 493364 89218
rect 494072 16574 494100 96086
rect 500960 96008 501012 96014
rect 500960 95950 501012 95956
rect 497464 89208 497516 89214
rect 497464 89150 497516 89156
rect 494072 16546 494744 16574
rect 493324 3052 493376 3058
rect 493324 2994 493376 3000
rect 493336 598 493548 626
rect 493336 490 493364 598
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493060 462 493364 490
rect 493520 480 493548 598
rect 494716 480 494744 16546
rect 497096 8968 497148 8974
rect 497096 8910 497148 8916
rect 495900 3052 495952 3058
rect 495900 2994 495952 3000
rect 495912 480 495940 2994
rect 497108 480 497136 8910
rect 497476 3398 497504 89150
rect 500224 89140 500276 89146
rect 500224 89082 500276 89088
rect 500236 16574 500264 89082
rect 500972 16574 501000 95950
rect 502984 94648 503036 94654
rect 502984 94590 503036 94596
rect 500236 16546 500356 16574
rect 500972 16546 501368 16574
rect 500224 13116 500276 13122
rect 500224 13058 500276 13064
rect 498200 3800 498252 3806
rect 498200 3742 498252 3748
rect 497464 3392 497516 3398
rect 497464 3334 497516 3340
rect 498212 480 498240 3742
rect 499396 3392 499448 3398
rect 499396 3334 499448 3340
rect 499408 480 499436 3334
rect 500236 3074 500264 13058
rect 500328 3262 500356 16546
rect 500316 3256 500368 3262
rect 500316 3198 500368 3204
rect 500236 3046 500632 3074
rect 500604 480 500632 3046
rect 501340 490 501368 16546
rect 502996 3398 503024 94590
rect 504364 90500 504416 90506
rect 504364 90442 504416 90448
rect 503720 80776 503772 80782
rect 503720 80718 503772 80724
rect 502984 3392 503036 3398
rect 502984 3334 503036 3340
rect 502984 3256 503036 3262
rect 502984 3198 503036 3204
rect 501616 598 501828 626
rect 501616 490 501644 598
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501340 462 501644 490
rect 501800 480 501828 598
rect 502996 480 503024 3198
rect 503732 490 503760 80718
rect 504376 3058 504404 90442
rect 506480 88052 506532 88058
rect 506480 87994 506532 88000
rect 505376 3392 505428 3398
rect 505376 3334 505428 3340
rect 504364 3052 504416 3058
rect 504364 2994 504416 3000
rect 504008 598 504220 626
rect 504008 490 504036 598
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 503732 462 504036 490
rect 504192 480 504220 598
rect 505388 480 505416 3334
rect 506492 480 506520 87994
rect 506572 79416 506624 79422
rect 506572 79358 506624 79364
rect 506584 16574 506612 79358
rect 507872 16574 507900 98738
rect 512000 98728 512052 98734
rect 512000 98670 512052 98676
rect 511264 87984 511316 87990
rect 511264 87926 511316 87932
rect 510620 78056 510672 78062
rect 510620 77998 510672 78004
rect 510632 16574 510660 77998
rect 506584 16546 507256 16574
rect 507872 16546 508912 16574
rect 510632 16546 511212 16574
rect 507228 490 507256 16546
rect 507504 598 507716 626
rect 507504 490 507532 598
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507228 462 507532 490
rect 507688 480 507716 598
rect 508884 480 508912 16546
rect 510068 3052 510120 3058
rect 510068 2994 510120 3000
rect 510080 480 510108 2994
rect 511184 2938 511212 16546
rect 511276 3058 511304 87926
rect 511264 3052 511316 3058
rect 511264 2994 511316 3000
rect 511184 2910 511304 2938
rect 511276 480 511304 2910
rect 512012 490 512040 98670
rect 529940 98660 529992 98666
rect 529940 98602 529992 98608
rect 518900 94580 518952 94586
rect 518900 94522 518952 94528
rect 515404 87848 515456 87854
rect 515404 87790 515456 87796
rect 514760 14476 514812 14482
rect 514760 14418 514812 14424
rect 513564 3052 513616 3058
rect 513564 2994 513616 3000
rect 512288 598 512500 626
rect 512288 490 512316 598
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512012 462 512316 490
rect 512472 480 512500 598
rect 513576 480 513604 2994
rect 514772 480 514800 14418
rect 515416 3602 515444 87790
rect 518164 87780 518216 87786
rect 518164 87722 518216 87728
rect 517520 76696 517572 76702
rect 517520 76638 517572 76644
rect 517532 16574 517560 76638
rect 517532 16546 517928 16574
rect 515036 3596 515088 3602
rect 515036 3538 515088 3544
rect 515404 3596 515456 3602
rect 515404 3538 515456 3544
rect 517152 3596 517204 3602
rect 517152 3538 517204 3544
rect 515048 2854 515076 3538
rect 515036 2848 515088 2854
rect 515036 2790 515088 2796
rect 515956 2848 516008 2854
rect 515956 2790 516008 2796
rect 515968 480 515996 2790
rect 517164 480 517192 3538
rect 517900 490 517928 16546
rect 518176 3874 518204 87722
rect 518912 16574 518940 94522
rect 520924 94512 520976 94518
rect 520924 94454 520976 94460
rect 518912 16546 519584 16574
rect 518164 3868 518216 3874
rect 518164 3810 518216 3816
rect 518176 598 518388 626
rect 518176 490 518204 598
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 517900 462 518204 490
rect 518360 480 518388 598
rect 519556 480 519584 16546
rect 520740 3868 520792 3874
rect 520740 3810 520792 3816
rect 520752 480 520780 3810
rect 520936 3398 520964 94454
rect 524420 93356 524472 93362
rect 524420 93298 524472 93304
rect 522304 89072 522356 89078
rect 522304 89014 522356 89020
rect 521844 6180 521896 6186
rect 521844 6122 521896 6128
rect 520924 3392 520976 3398
rect 520924 3334 520976 3340
rect 521856 480 521884 6122
rect 522316 3602 522344 89014
rect 524432 6914 524460 93298
rect 525064 93288 525116 93294
rect 525064 93230 525116 93236
rect 525076 16574 525104 93230
rect 529204 91792 529256 91798
rect 529204 91734 529256 91740
rect 525800 87916 525852 87922
rect 525800 87858 525852 87864
rect 525812 16574 525840 87858
rect 528560 85060 528612 85066
rect 528560 85002 528612 85008
rect 525076 16546 525196 16574
rect 525812 16546 526208 16574
rect 524432 6886 525104 6914
rect 522304 3596 522356 3602
rect 522304 3538 522356 3544
rect 524236 3596 524288 3602
rect 524236 3538 524288 3544
rect 523040 3392 523092 3398
rect 523040 3334 523092 3340
rect 523052 480 523080 3334
rect 524248 480 524276 3538
rect 525076 2802 525104 6886
rect 525168 2990 525196 16546
rect 525156 2984 525208 2990
rect 525156 2926 525208 2932
rect 525076 2774 525472 2802
rect 525444 480 525472 2774
rect 526180 490 526208 16546
rect 527824 2984 527876 2990
rect 527824 2926 527876 2932
rect 526456 598 526668 626
rect 526456 490 526484 598
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526180 462 526484 490
rect 526640 480 526668 598
rect 527836 480 527864 2926
rect 528572 490 528600 85002
rect 529216 3058 529244 91734
rect 529952 16574 529980 98602
rect 532700 95940 532752 95946
rect 532700 95882 532752 95888
rect 530584 79348 530636 79354
rect 530584 79290 530636 79296
rect 529952 16546 530164 16574
rect 529204 3052 529256 3058
rect 529204 2994 529256 3000
rect 528848 598 529060 626
rect 528848 490 528876 598
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528572 462 528876 490
rect 529032 480 529060 598
rect 530136 480 530164 16546
rect 530596 3534 530624 79290
rect 532712 16574 532740 95882
rect 536838 94752 536894 94761
rect 536838 94687 536894 94696
rect 536104 86556 536156 86562
rect 536104 86498 536156 86504
rect 535460 76628 535512 76634
rect 535460 76570 535512 76576
rect 535472 16574 535500 76570
rect 532712 16546 533752 16574
rect 535472 16546 536052 16574
rect 530584 3528 530636 3534
rect 530584 3470 530636 3476
rect 532516 3528 532568 3534
rect 532516 3470 532568 3476
rect 531320 3052 531372 3058
rect 531320 2994 531372 3000
rect 531332 480 531360 2994
rect 532528 480 532556 3470
rect 533724 480 533752 16546
rect 534908 3732 534960 3738
rect 534908 3674 534960 3680
rect 534920 480 534948 3674
rect 536024 3482 536052 16546
rect 536116 3874 536144 86498
rect 536852 16574 536880 94687
rect 538864 93220 538916 93226
rect 538864 93162 538916 93168
rect 536852 16546 537248 16574
rect 536104 3868 536156 3874
rect 536104 3810 536156 3816
rect 536024 3454 536144 3482
rect 536116 480 536144 3454
rect 537220 480 537248 16546
rect 538404 3868 538456 3874
rect 538404 3810 538456 3816
rect 538416 480 538444 3810
rect 538876 3670 538904 93162
rect 540244 90432 540296 90438
rect 540244 90374 540296 90380
rect 539600 10328 539652 10334
rect 539600 10270 539652 10276
rect 538864 3664 538916 3670
rect 538864 3606 538916 3612
rect 539612 480 539640 10270
rect 540256 3534 540284 90374
rect 543004 87712 543056 87718
rect 543004 87654 543056 87660
rect 542360 77988 542412 77994
rect 542360 77930 542412 77936
rect 542372 16574 542400 77930
rect 542372 16546 542768 16574
rect 540796 3596 540848 3602
rect 540796 3538 540848 3544
rect 540244 3528 540296 3534
rect 540244 3470 540296 3476
rect 540808 480 540836 3538
rect 541992 3528 542044 3534
rect 541992 3470 542044 3476
rect 542004 480 542032 3470
rect 542740 490 542768 16546
rect 543016 3126 543044 87654
rect 543752 16574 543780 98767
rect 550638 98696 550694 98705
rect 550638 98631 550694 98640
rect 547144 86488 547196 86494
rect 547144 86430 547196 86436
rect 543752 16546 544424 16574
rect 543004 3120 543056 3126
rect 543004 3062 543056 3068
rect 543016 598 543228 626
rect 543016 490 543044 598
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 542740 462 543044 490
rect 543200 480 543228 598
rect 544396 480 544424 16546
rect 546684 15904 546736 15910
rect 546684 15846 546736 15852
rect 545488 3120 545540 3126
rect 545488 3062 545540 3068
rect 545500 480 545528 3062
rect 546696 480 546724 15846
rect 547156 4146 547184 86430
rect 548524 76560 548576 76566
rect 548524 76502 548576 76508
rect 547144 4140 547196 4146
rect 547144 4082 547196 4088
rect 548536 3534 548564 76502
rect 550652 16574 550680 98631
rect 580262 97336 580318 97345
rect 580262 97271 580318 97280
rect 557538 95840 557594 95849
rect 557538 95775 557594 95784
rect 554780 93152 554832 93158
rect 554780 93094 554832 93100
rect 553400 89004 553452 89010
rect 553400 88946 553452 88952
rect 550652 16546 551048 16574
rect 549076 4140 549128 4146
rect 549076 4082 549128 4088
rect 548524 3528 548576 3534
rect 548524 3470 548576 3476
rect 547880 3460 547932 3466
rect 547880 3402 547932 3408
rect 547892 480 547920 3402
rect 549088 480 549116 4082
rect 550272 3528 550324 3534
rect 550272 3470 550324 3476
rect 550284 480 550312 3470
rect 551020 490 551048 16546
rect 553412 3534 553440 88946
rect 554792 16574 554820 93094
rect 556160 86420 556212 86426
rect 556160 86362 556212 86368
rect 554792 16546 555004 16574
rect 553768 4820 553820 4826
rect 553768 4762 553820 4768
rect 552664 3528 552716 3534
rect 552664 3470 552716 3476
rect 553400 3528 553452 3534
rect 553400 3470 553452 3476
rect 551296 598 551508 626
rect 551296 490 551324 598
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551020 462 551324 490
rect 551480 480 551508 598
rect 552676 480 552704 3470
rect 553780 480 553808 4762
rect 554976 480 555004 16546
rect 556172 480 556200 86362
rect 556252 25560 556304 25566
rect 556252 25502 556304 25508
rect 556264 16574 556292 25502
rect 557552 16574 557580 95775
rect 561678 94616 561734 94625
rect 561678 94551 561734 94560
rect 560392 86352 560444 86358
rect 560392 86294 560444 86300
rect 560300 75268 560352 75274
rect 560300 75210 560352 75216
rect 556264 16546 556936 16574
rect 557552 16546 558592 16574
rect 556908 490 556936 16546
rect 557184 598 557396 626
rect 557184 490 557212 598
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 556908 462 557212 490
rect 557368 480 557396 598
rect 558564 480 558592 16546
rect 560312 6914 560340 75210
rect 560404 16574 560432 86294
rect 561692 16574 561720 94551
rect 568578 94480 568634 94489
rect 568578 94415 568634 94424
rect 566464 90364 566516 90370
rect 566464 90306 566516 90312
rect 565820 84992 565872 84998
rect 565820 84934 565872 84940
rect 564532 84924 564584 84930
rect 564532 84866 564584 84872
rect 560404 16546 560524 16574
rect 561692 16546 562088 16574
rect 560312 6886 560432 6914
rect 559748 3528 559800 3534
rect 559748 3470 559800 3476
rect 559760 480 559788 3470
rect 560404 490 560432 6886
rect 560496 3534 560524 16546
rect 560484 3528 560536 3534
rect 560484 3470 560536 3476
rect 560680 598 560892 626
rect 560680 490 560708 598
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560404 462 560708 490
rect 560864 480 560892 598
rect 562060 480 562088 16546
rect 564544 3602 564572 84866
rect 564624 19984 564676 19990
rect 564624 19926 564676 19932
rect 563244 3596 563296 3602
rect 563244 3538 563296 3544
rect 564532 3596 564584 3602
rect 564532 3538 564584 3544
rect 563256 480 563284 3538
rect 564636 3482 564664 19926
rect 565832 6914 565860 84934
rect 566476 16574 566504 90306
rect 568592 16574 568620 94415
rect 575478 93120 575534 93129
rect 575478 93055 575534 93064
rect 569960 87644 570012 87650
rect 569960 87586 570012 87592
rect 569972 16574 570000 87586
rect 572812 84856 572864 84862
rect 572812 84798 572864 84804
rect 571340 82136 571392 82142
rect 571340 82078 571392 82084
rect 571352 16574 571380 82078
rect 572824 16574 572852 84798
rect 574100 80708 574152 80714
rect 574100 80650 574152 80656
rect 574112 16574 574140 80650
rect 575492 16574 575520 93055
rect 578240 75200 578292 75206
rect 578240 75142 578292 75148
rect 578252 16574 578280 75142
rect 579988 73160 580040 73166
rect 579988 73102 580040 73108
rect 580000 73001 580028 73102
rect 579986 72992 580042 73001
rect 579986 72927 580042 72936
rect 580172 60716 580224 60722
rect 580172 60658 580224 60664
rect 580184 59673 580212 60658
rect 580170 59664 580226 59673
rect 580170 59599 580226 59608
rect 580276 33998 580304 97271
rect 580264 33992 580316 33998
rect 580264 33934 580316 33940
rect 566476 16546 566596 16574
rect 568592 16546 568712 16574
rect 569972 16546 570368 16574
rect 571352 16546 571564 16574
rect 572824 16546 573496 16574
rect 574112 16546 575152 16574
rect 575492 16546 575888 16574
rect 578252 16546 578648 16574
rect 565832 6886 566504 6914
rect 564452 3454 564664 3482
rect 565636 3528 565688 3534
rect 565636 3470 565688 3476
rect 566476 3482 566504 6886
rect 566568 4146 566596 16546
rect 566556 4140 566608 4146
rect 566556 4082 566608 4088
rect 568028 4140 568080 4146
rect 568028 4082 568080 4088
rect 564452 480 564480 3454
rect 565648 480 565676 3470
rect 566476 3454 566872 3482
rect 566844 480 566872 3454
rect 568040 480 568068 4082
rect 568684 490 568712 16546
rect 568960 598 569172 626
rect 568960 490 568988 598
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 568684 462 568988 490
rect 569144 480 569172 598
rect 570340 480 570368 16546
rect 571536 480 571564 16546
rect 572720 3664 572772 3670
rect 572720 3606 572772 3612
rect 572732 480 572760 3606
rect 573468 490 573496 16546
rect 573744 598 573956 626
rect 573744 490 573772 598
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573468 462 573772 490
rect 573928 480 573956 598
rect 575124 480 575152 16546
rect 575860 490 575888 16546
rect 577412 3596 577464 3602
rect 577412 3538 577464 3544
rect 576136 598 576348 626
rect 576136 490 576164 598
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 575860 462 576164 490
rect 576320 480 576348 598
rect 577424 480 577452 3538
rect 578620 480 578648 16546
rect 582392 6633 582420 300902
rect 582484 19825 582512 303622
rect 582932 301096 582984 301102
rect 582932 301038 582984 301044
rect 582656 301028 582708 301034
rect 582656 300970 582708 300976
rect 582564 299532 582616 299538
rect 582564 299474 582616 299480
rect 582576 86193 582604 299474
rect 582562 86184 582618 86193
rect 582562 86119 582618 86128
rect 582668 46345 582696 300970
rect 582840 299600 582892 299606
rect 582840 299542 582892 299548
rect 582852 126041 582880 299542
rect 582944 165889 582972 301038
rect 583116 300892 583168 300898
rect 583116 300834 583168 300840
rect 583024 299668 583076 299674
rect 583024 299610 583076 299616
rect 583036 205737 583064 299610
rect 583022 205728 583078 205737
rect 583022 205663 583078 205672
rect 582930 165880 582986 165889
rect 582930 165815 582986 165824
rect 582838 126032 582894 126041
rect 582838 125967 582894 125976
rect 582838 97200 582894 97209
rect 582838 97135 582894 97144
rect 582748 86284 582800 86290
rect 582748 86226 582800 86232
rect 582654 46336 582710 46345
rect 582654 46271 582710 46280
rect 582564 33992 582616 33998
rect 582564 33934 582616 33940
rect 582470 19816 582526 19825
rect 582470 19751 582526 19760
rect 582576 16574 582604 33934
rect 582576 16546 582696 16574
rect 582378 6624 582434 6633
rect 582378 6559 582434 6568
rect 582196 3528 582248 3534
rect 582196 3470 582248 3476
rect 581000 3460 581052 3466
rect 581000 3402 581052 3408
rect 581012 480 581040 3402
rect 582208 480 582236 3470
rect 582668 3346 582696 16546
rect 582760 3602 582788 86226
rect 582748 3596 582800 3602
rect 582748 3538 582800 3544
rect 582852 3466 582880 97135
rect 582932 73840 582984 73846
rect 582932 73782 582984 73788
rect 582944 3534 582972 73782
rect 583128 33153 583156 300834
rect 583114 33144 583170 33153
rect 583114 33079 583170 33088
rect 582932 3528 582984 3534
rect 582932 3470 582984 3476
rect 582840 3460 582892 3466
rect 582840 3402 582892 3408
rect 582668 3318 583432 3346
rect 583404 480 583432 3318
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 3422 671200 3478 671256
rect 3330 579944 3386 580000
rect 3238 566888 3294 566944
rect 3330 553832 3386 553888
rect 2962 527856 3018 527912
rect 3054 501744 3110 501800
rect 3054 475632 3110 475688
rect 3146 449520 3202 449576
rect 2870 410488 2926 410544
rect 3146 358400 3202 358456
rect 3330 345344 3386 345400
rect 3330 319232 3386 319288
rect 3514 658144 3570 658200
rect 3514 632068 3516 632088
rect 3516 632068 3568 632088
rect 3568 632068 3570 632088
rect 3514 632032 3570 632068
rect 3514 619112 3570 619168
rect 3514 606056 3570 606112
rect 3514 514820 3570 514856
rect 3514 514800 3516 514820
rect 3516 514800 3568 514820
rect 3568 514800 3570 514820
rect 3514 462576 3570 462632
rect 3514 423544 3570 423600
rect 3514 397468 3516 397488
rect 3516 397468 3568 397488
rect 3568 397468 3570 397488
rect 3514 397432 3570 397468
rect 3514 371320 3570 371376
rect 3238 306176 3294 306232
rect 3054 293120 3110 293176
rect 3146 254088 3202 254144
rect 3330 214920 3386 214976
rect 3054 201864 3110 201920
rect 3238 162832 3294 162888
rect 3514 267144 3570 267200
rect 3514 241032 3570 241088
rect 3514 188808 3570 188864
rect 3514 149776 3570 149832
rect 3422 136720 3478 136776
rect 3422 110608 3478 110664
rect 3422 97552 3478 97608
rect 1306 94424 1362 94480
rect 4066 93064 4122 93120
rect 3146 84632 3202 84688
rect 3422 71576 3478 71632
rect 3054 58520 3110 58576
rect 3422 45500 3424 45520
rect 3424 45500 3476 45520
rect 3476 45500 3478 45520
rect 3422 45464 3478 45500
rect 2870 32408 2926 32464
rect 3422 19352 3478 19408
rect 3422 6432 3478 6488
rect 12346 95784 12402 95840
rect 17222 97144 17278 97200
rect 35254 97416 35310 97472
rect 29642 97280 29698 97336
rect 22742 95920 22798 95976
rect 28262 94560 28318 94616
rect 169666 186224 169722 186280
rect 171690 184184 171746 184240
rect 171782 170992 171838 171048
rect 172426 189896 172482 189952
rect 172058 188672 172114 188728
rect 172150 187620 172152 187640
rect 172152 187620 172204 187640
rect 172204 187620 172206 187640
rect 172150 187584 172206 187620
rect 171874 169224 171930 169280
rect 172426 184884 172482 184920
rect 172426 184864 172428 184884
rect 172428 184864 172480 184884
rect 172480 184864 172482 184884
rect 172426 182960 172482 183016
rect 172058 181736 172114 181792
rect 172426 180512 172482 180568
rect 172426 179152 172482 179208
rect 172426 177964 172428 177984
rect 172428 177964 172480 177984
rect 172480 177964 172482 177984
rect 172426 177928 172482 177964
rect 172334 177384 172390 177440
rect 172242 176024 172298 176080
rect 172426 174800 172482 174856
rect 172426 173612 172428 173632
rect 172428 173612 172480 173632
rect 172480 173612 172482 173632
rect 172426 173576 172482 173612
rect 172426 172388 172428 172408
rect 172428 172388 172480 172408
rect 172480 172388 172482 172408
rect 172426 172352 172482 172388
rect 172242 170448 172298 170504
rect 171966 166912 172022 166968
rect 171598 153720 171654 153776
rect 171690 153176 171746 153232
rect 171598 152632 171654 152688
rect 170494 152088 170550 152144
rect 171690 150456 171746 150512
rect 171506 149368 171562 149424
rect 171690 148316 171692 148336
rect 171692 148316 171744 148336
rect 171744 148316 171746 148336
rect 171690 148280 171746 148316
rect 171506 147736 171562 147792
rect 171690 147192 171746 147248
rect 171690 145016 171746 145072
rect 171690 144472 171746 144528
rect 172058 165144 172114 165200
rect 172426 167864 172482 167920
rect 172426 164056 172482 164112
rect 172242 163512 172298 163568
rect 172150 162288 172206 162344
rect 172426 160928 172482 160984
rect 171782 144064 171838 144120
rect 172426 151544 172482 151600
rect 172242 151000 172298 151056
rect 172426 149912 172482 149968
rect 172426 148860 172428 148880
rect 172428 148860 172480 148880
rect 172480 148860 172482 148880
rect 172426 148824 172482 148860
rect 172334 146648 172390 146704
rect 172426 146104 172482 146160
rect 172426 145560 172482 145616
rect 171966 143520 172022 143576
rect 171874 142976 171930 143032
rect 172426 142432 172482 142488
rect 171874 141344 171930 141400
rect 172426 141888 172482 141944
rect 172334 140800 172390 140856
rect 172150 140292 172152 140312
rect 172152 140292 172204 140312
rect 172204 140292 172206 140312
rect 172150 140256 172206 140292
rect 172426 139712 172482 139768
rect 172242 139204 172244 139224
rect 172244 139204 172296 139224
rect 172296 139204 172298 139224
rect 172242 139168 172298 139204
rect 172426 138624 172482 138680
rect 172334 138080 172390 138136
rect 172058 137536 172114 137592
rect 171690 136992 171746 137048
rect 171322 135360 171378 135416
rect 198554 298832 198610 298888
rect 197910 294480 197966 294536
rect 197542 292304 197598 292360
rect 198738 290128 198794 290184
rect 197542 288088 197598 288144
rect 198094 285912 198150 285968
rect 197358 283736 197414 283792
rect 197358 281580 197414 281616
rect 197358 281560 197360 281580
rect 197360 281560 197412 281580
rect 197412 281560 197414 281580
rect 197726 279384 197782 279440
rect 197358 277344 197414 277400
rect 172426 136484 172428 136504
rect 172428 136484 172480 136504
rect 172480 136484 172482 136504
rect 172426 136448 172482 136484
rect 172242 135904 172298 135960
rect 171874 134816 171930 134872
rect 171690 134272 171746 134328
rect 172426 133864 172482 133920
rect 172058 133320 172114 133376
rect 172426 132776 172482 132832
rect 171138 132232 171194 132288
rect 172426 131688 172482 131744
rect 171506 131144 171562 131200
rect 171874 130600 171930 130656
rect 172426 130076 172482 130112
rect 172426 130056 172428 130076
rect 172428 130056 172480 130076
rect 172480 130056 172482 130076
rect 171874 129512 171930 129568
rect 171506 128968 171562 129024
rect 171782 128424 171838 128480
rect 171690 127880 171746 127936
rect 171322 124636 171378 124672
rect 171322 124616 171324 124636
rect 171324 124616 171376 124636
rect 171376 124616 171378 124636
rect 172426 127336 172482 127392
rect 172058 126792 172114 126848
rect 172334 126248 172390 126304
rect 172426 125724 172482 125760
rect 172426 125704 172428 125724
rect 172428 125704 172480 125724
rect 172480 125704 172482 125724
rect 172426 125180 172482 125216
rect 172426 125160 172428 125180
rect 172428 125160 172480 125180
rect 172480 125160 172482 125180
rect 171966 124228 172022 124264
rect 171966 124208 171968 124228
rect 171968 124208 172020 124228
rect 172020 124208 172022 124228
rect 197542 272992 197598 273048
rect 197726 270816 197782 270872
rect 197818 268640 197874 268696
rect 197358 266484 197414 266520
rect 197358 266464 197360 266484
rect 197360 266464 197412 266484
rect 197412 266464 197414 266484
rect 197358 264424 197414 264480
rect 197358 262268 197414 262304
rect 197358 262248 197360 262268
rect 197360 262248 197412 262268
rect 197412 262248 197414 262268
rect 197726 260072 197782 260128
rect 197542 257896 197598 257952
rect 197910 255720 197966 255776
rect 197542 253680 197598 253736
rect 197358 251504 197414 251560
rect 197634 249328 197690 249384
rect 198002 247152 198058 247208
rect 197358 244976 197414 245032
rect 197910 242800 197966 242856
rect 197726 240760 197782 240816
rect 197542 238584 197598 238640
rect 197726 236408 197782 236464
rect 197726 234232 197782 234288
rect 197634 230016 197690 230072
rect 197358 227840 197414 227896
rect 197358 225664 197414 225720
rect 197358 223488 197414 223544
rect 197542 219136 197598 219192
rect 197358 217096 197414 217152
rect 197542 214920 197598 214976
rect 197358 212744 197414 212800
rect 197358 210568 197414 210624
rect 197358 206352 197414 206408
rect 197358 202000 197414 202056
rect 197358 197648 197414 197704
rect 197634 195472 197690 195528
rect 197358 193432 197414 193488
rect 197358 189100 197414 189136
rect 197358 189080 197360 189100
rect 197360 189080 197412 189100
rect 197412 189080 197414 189100
rect 197358 186904 197414 186960
rect 197358 184728 197414 184784
rect 197358 178336 197414 178392
rect 197634 176160 197690 176216
rect 197358 173984 197414 174040
rect 198646 275168 198702 275224
rect 198370 232056 198426 232112
rect 198186 208392 198242 208448
rect 198094 199824 198150 199880
rect 198278 204176 198334 204232
rect 198370 191256 198426 191312
rect 198094 182688 198150 182744
rect 198370 180512 198426 180568
rect 198186 171808 198242 171864
rect 197726 169768 197782 169824
rect 197542 167592 197598 167648
rect 198094 165416 198150 165472
rect 198002 163240 198058 163296
rect 197542 161064 197598 161120
rect 197358 159024 197414 159080
rect 197818 156848 197874 156904
rect 197358 154672 197414 154728
rect 197358 152496 197414 152552
rect 197358 150320 197414 150376
rect 197358 148144 197414 148200
rect 198830 221312 198886 221368
rect 198094 146104 198150 146160
rect 197358 143928 197414 143984
rect 197542 141752 197598 141808
rect 197726 139576 197782 139632
rect 197358 137400 197414 137456
rect 197358 135360 197414 135416
rect 197358 133184 197414 133240
rect 197358 131044 197360 131064
rect 197360 131044 197412 131064
rect 197412 131044 197414 131064
rect 197358 131008 197414 131044
rect 197358 128832 197414 128888
rect 197542 124480 197598 124536
rect 198462 126656 198518 126712
rect 217414 299376 217470 299432
rect 217966 299396 218022 299432
rect 217966 299376 217968 299396
rect 217968 299376 218020 299396
rect 218020 299376 218022 299396
rect 371882 369688 371938 369744
rect 371606 369144 371662 369200
rect 371698 368056 371754 368112
rect 371606 367512 371662 367568
rect 371238 366968 371294 367024
rect 371514 366424 371570 366480
rect 371606 365900 371662 365936
rect 371606 365880 371608 365900
rect 371608 365880 371660 365900
rect 371660 365880 371662 365900
rect 371238 365336 371294 365392
rect 371606 364792 371662 364848
rect 371698 364248 371754 364304
rect 371606 363704 371662 363760
rect 371698 362616 371754 362672
rect 371606 362072 371662 362128
rect 371606 361548 371662 361584
rect 371606 361528 371608 361548
rect 371608 361528 371660 361548
rect 371660 361528 371662 361548
rect 371422 360984 371478 361040
rect 371606 360460 371662 360496
rect 371606 360440 371608 360460
rect 371608 360440 371660 360460
rect 371660 360440 371662 360460
rect 372066 368600 372122 368656
rect 372526 363160 372582 363216
rect 372342 360032 372398 360088
rect 372158 359488 372214 359544
rect 371974 358944 372030 359000
rect 371698 358400 371754 358456
rect 371606 357856 371662 357912
rect 371606 357312 371662 357368
rect 371514 356768 371570 356824
rect 371238 356224 371294 356280
rect 371606 355680 371662 355736
rect 371514 355136 371570 355192
rect 371330 354592 371386 354648
rect 371698 354048 371754 354104
rect 371514 353504 371570 353560
rect 369306 350512 369362 350568
rect 370318 348744 370374 348800
rect 369398 347384 369454 347440
rect 217230 299240 217286 299296
rect 217690 299276 217692 299296
rect 217692 299276 217744 299296
rect 217744 299276 217746 299296
rect 217690 299240 217746 299276
rect 199842 296656 199898 296712
rect 302790 298424 302846 298480
rect 302790 295332 302792 295352
rect 302792 295332 302844 295352
rect 302844 295332 302846 295352
rect 302790 295296 302846 295332
rect 302238 292168 302294 292224
rect 302698 289040 302754 289096
rect 302790 285912 302846 285968
rect 302514 282784 302570 282840
rect 302790 279656 302846 279712
rect 302790 276528 302846 276584
rect 302974 273400 303030 273456
rect 302882 270272 302938 270328
rect 303250 267144 303306 267200
rect 302790 264016 302846 264072
rect 302790 260888 302846 260944
rect 302790 257760 302846 257816
rect 302330 254632 302386 254688
rect 302974 251504 303030 251560
rect 302790 248412 302792 248432
rect 302792 248412 302844 248432
rect 302844 248412 302846 248432
rect 302790 248376 302846 248412
rect 302882 245248 302938 245304
rect 302698 229608 302754 229664
rect 302698 226480 302754 226536
rect 303066 242120 303122 242176
rect 302974 235864 303030 235920
rect 303158 238992 303214 239048
rect 303250 232736 303306 232792
rect 302790 223352 302846 223408
rect 302790 220224 302846 220280
rect 302514 217096 302570 217152
rect 302790 213968 302846 214024
rect 302790 210840 302846 210896
rect 302330 207712 302386 207768
rect 302698 204584 302754 204640
rect 302790 201492 302792 201512
rect 302792 201492 302844 201512
rect 302844 201492 302846 201512
rect 302790 201456 302846 201492
rect 302790 198328 302846 198384
rect 302330 195200 302386 195256
rect 198002 122440 198058 122496
rect 197542 120264 197598 120320
rect 197910 118088 197966 118144
rect 198370 115912 198426 115968
rect 197358 113736 197414 113792
rect 197358 111732 197360 111752
rect 197360 111732 197412 111752
rect 197412 111732 197414 111752
rect 197358 111696 197414 111732
rect 197358 109520 197414 109576
rect 198554 107344 198610 107400
rect 197542 105168 197598 105224
rect 197910 102992 197966 103048
rect 302790 192072 302846 192128
rect 302790 188980 302792 189000
rect 302792 188980 302844 189000
rect 302844 188980 302846 189000
rect 302790 188944 302846 188980
rect 302698 185816 302754 185872
rect 302790 179560 302846 179616
rect 302790 176432 302846 176488
rect 302974 182688 303030 182744
rect 302882 173304 302938 173360
rect 302790 170176 302846 170232
rect 303066 167048 303122 167104
rect 302882 163920 302938 163976
rect 302514 160792 302570 160848
rect 302790 157664 302846 157720
rect 302606 154536 302662 154592
rect 302698 151408 302754 151464
rect 302330 148280 302386 148336
rect 302790 145152 302846 145208
rect 302790 142060 302792 142080
rect 302792 142060 302844 142080
rect 302844 142060 302846 142080
rect 302790 142024 302846 142060
rect 302698 138896 302754 138952
rect 302882 135768 302938 135824
rect 302606 129512 302662 129568
rect 302790 126384 302846 126440
rect 302974 132640 303030 132696
rect 302790 123256 302846 123312
rect 302514 120128 302570 120184
rect 302790 117000 302846 117056
rect 302790 110744 302846 110800
rect 302790 107616 302846 107672
rect 302974 113872 303030 113928
rect 302882 104488 302938 104544
rect 302790 101496 302846 101552
rect 197542 100952 197598 101008
rect 196622 97552 196678 97608
rect 199474 97824 199530 97880
rect 200118 94424 200174 94480
rect 199474 93064 199530 93120
rect 200670 97824 200726 97880
rect 202694 97144 202750 97200
rect 203338 97280 203394 97336
rect 203062 95920 203118 95976
rect 201866 95784 201922 95840
rect 204350 97416 204406 97472
rect 203890 94560 203946 94616
rect 204902 97552 204958 97608
rect 260286 3440 260342 3496
rect 260746 3304 260802 3360
rect 281906 97416 281962 97472
rect 284482 97144 284538 97200
rect 290002 97552 290058 97608
rect 289818 96872 289874 96928
rect 291658 94696 291714 94752
rect 291934 96872 291990 96928
rect 293038 98776 293094 98832
rect 294234 98640 294290 98696
rect 296074 94560 296130 94616
rect 296810 96872 296866 96928
rect 297454 97144 297510 97200
rect 297270 96736 297326 96792
rect 297822 98912 297878 98968
rect 299110 97280 299166 97336
rect 298374 95784 298430 95840
rect 299018 93064 299074 93120
rect 300306 97552 300362 97608
rect 299478 97280 299534 97336
rect 300122 96872 300178 96928
rect 300766 96736 300822 96792
rect 300766 94424 300822 94480
rect 353942 266192 353998 266248
rect 362866 337728 362922 337784
rect 364890 337728 364946 337784
rect 369858 345752 369914 345808
rect 369490 297336 369546 297392
rect 369398 296792 369454 296848
rect 369398 296248 369454 296304
rect 369398 295860 369454 295896
rect 369398 295840 369400 295860
rect 369400 295840 369452 295860
rect 369452 295840 369454 295860
rect 369490 278976 369546 279032
rect 369398 278604 369400 278624
rect 369400 278604 369452 278624
rect 369452 278604 369454 278624
rect 369398 278568 369454 278604
rect 369398 275340 369400 275360
rect 369400 275340 369452 275360
rect 369452 275340 369454 275360
rect 369398 275304 369454 275340
rect 356702 266056 356758 266112
rect 362866 266056 362922 266112
rect 364890 266056 364946 266112
rect 369398 222808 369454 222864
rect 370226 345480 370282 345536
rect 369858 274216 369914 274272
rect 370134 340604 370190 340640
rect 370134 340584 370136 340604
rect 370136 340584 370188 340604
rect 370188 340584 370190 340604
rect 370226 340176 370282 340232
rect 370134 295568 370190 295624
rect 370042 273264 370098 273320
rect 369950 268912 370006 268968
rect 369582 220632 369638 220688
rect 369858 220632 369914 220688
rect 369950 218456 370006 218512
rect 369674 208700 369676 208720
rect 369676 208700 369728 208720
rect 369728 208700 369730 208720
rect 369674 208664 369730 208700
rect 369582 206488 369638 206544
rect 369398 206116 369400 206136
rect 369400 206116 369452 206136
rect 369452 206116 369454 206136
rect 369398 206080 369454 206116
rect 369490 204040 369546 204096
rect 369766 207032 369822 207088
rect 364522 196016 364578 196072
rect 362866 194520 362922 194576
rect 364890 194520 364946 194576
rect 369306 152904 369362 152960
rect 370410 347112 370466 347168
rect 370318 276800 370374 276856
rect 371974 352960 372030 353016
rect 371606 349308 371662 349344
rect 371606 349288 371608 349308
rect 371608 349288 371660 349308
rect 371660 349288 371662 349308
rect 371606 348220 371662 348256
rect 371606 348200 371608 348220
rect 371608 348200 371660 348220
rect 371660 348200 371662 348220
rect 371422 344392 371478 344448
rect 371330 342216 371386 342272
rect 371238 293936 371294 293992
rect 371238 291760 371294 291816
rect 371238 290128 371294 290184
rect 371238 287000 371294 287056
rect 371238 281560 371294 281616
rect 370410 275168 370466 275224
rect 370594 274080 370650 274136
rect 370226 268232 370282 268288
rect 370134 221312 370190 221368
rect 370318 221856 370374 221912
rect 370502 222944 370558 223000
rect 370410 219136 370466 219192
rect 370226 217504 370282 217560
rect 370410 211656 370466 211712
rect 370318 209480 370374 209536
rect 370134 208936 370190 208992
rect 370042 201864 370098 201920
rect 370226 202000 370282 202056
rect 370502 203088 370558 203144
rect 369490 136584 369546 136640
rect 369398 132368 369454 132424
rect 369306 131960 369362 132016
rect 369950 134544 370006 134600
rect 369858 133592 369914 133648
rect 370686 268232 370742 268288
rect 370594 202000 370650 202056
rect 371514 342760 371570 342816
rect 371422 272448 371478 272504
rect 371882 344936 371938 344992
rect 371790 341672 371846 341728
rect 371698 295024 371754 295080
rect 371698 294480 371754 294536
rect 371698 292848 371754 292904
rect 371698 292340 371700 292360
rect 371700 292340 371752 292360
rect 371752 292340 371754 292360
rect 371698 292304 371754 292340
rect 371698 290672 371754 290728
rect 371698 289604 371754 289640
rect 371698 289584 371700 289604
rect 371700 289584 371752 289604
rect 371752 289584 371754 289604
rect 371698 289076 371700 289096
rect 371700 289076 371752 289096
rect 371752 289076 371754 289096
rect 371698 289040 371754 289076
rect 371698 288516 371754 288552
rect 371698 288496 371700 288516
rect 371700 288496 371752 288516
rect 371752 288496 371754 288516
rect 371698 288088 371754 288144
rect 371698 287544 371754 287600
rect 371698 286456 371754 286512
rect 371606 285912 371662 285968
rect 371606 285368 371662 285424
rect 371606 284824 371662 284880
rect 371698 284280 371754 284336
rect 371606 283736 371662 283792
rect 371698 283192 371754 283248
rect 371606 282684 371608 282704
rect 371608 282684 371660 282704
rect 371660 282684 371662 282704
rect 371606 282648 371662 282684
rect 371606 282140 371608 282160
rect 371608 282140 371660 282160
rect 371660 282140 371662 282160
rect 371606 282104 371662 282140
rect 371606 281016 371662 281072
rect 371514 270816 371570 270872
rect 371330 270272 371386 270328
rect 371422 270136 371478 270192
rect 371422 269184 371478 269240
rect 371330 224576 371386 224632
rect 371330 222944 371386 223000
rect 371238 222420 371294 222456
rect 371238 222400 371240 222420
rect 371240 222400 371292 222420
rect 371292 222400 371294 222420
rect 371238 221856 371294 221912
rect 371054 218084 371056 218104
rect 371056 218084 371108 218104
rect 371108 218084 371110 218104
rect 371054 218048 371110 218084
rect 371330 216416 371386 216472
rect 371330 213832 371386 213888
rect 371238 209480 371294 209536
rect 371330 208936 371386 208992
rect 371238 203632 371294 203688
rect 371238 198736 371294 198792
rect 371698 277364 371754 277400
rect 371698 277344 371700 277364
rect 371700 277344 371752 277364
rect 371752 277344 371754 277364
rect 371698 276256 371754 276312
rect 371698 272992 371754 273048
rect 371606 225120 371662 225176
rect 371606 224032 371662 224088
rect 371606 223488 371662 223544
rect 371606 216996 371608 217016
rect 371608 216996 371660 217016
rect 371660 216996 371662 217016
rect 371606 216960 371662 216996
rect 371606 216008 371662 216064
rect 371606 214920 371662 214976
rect 371606 214376 371662 214432
rect 371606 213288 371662 213344
rect 371606 211112 371662 211168
rect 371606 210604 371608 210624
rect 371608 210604 371660 210624
rect 371660 210604 371662 210624
rect 371606 210568 371662 210604
rect 371606 205828 371662 205864
rect 371606 205808 371608 205828
rect 371608 205808 371660 205828
rect 371660 205808 371662 205828
rect 371606 205300 371608 205320
rect 371608 205300 371660 205320
rect 371660 205300 371662 205320
rect 371606 205264 371662 205300
rect 371606 204756 371608 204776
rect 371608 204756 371660 204776
rect 371660 204756 371662 204776
rect 371606 204720 371662 204756
rect 371606 204212 371608 204232
rect 371608 204212 371660 204232
rect 371660 204212 371662 204232
rect 371606 204176 371662 204212
rect 372434 351872 372490 351928
rect 372066 343848 372122 343904
rect 371974 281560 372030 281616
rect 371974 279384 372030 279440
rect 371882 272992 371938 273048
rect 371974 272448 372030 272504
rect 371882 270816 371938 270872
rect 371790 269728 371846 269784
rect 371698 200912 371754 200968
rect 371606 198872 371662 198928
rect 371514 198192 371570 198248
rect 371330 197104 371386 197160
rect 370686 196152 370742 196208
rect 370318 137536 370374 137592
rect 370410 135904 370466 135960
rect 370226 135360 370282 135416
rect 370134 132776 370190 132832
rect 369582 131416 369638 131472
rect 369306 130872 369362 130928
rect 370502 130056 370558 130112
rect 369950 129784 370006 129840
rect 369858 129104 369914 129160
rect 369398 126384 369454 126440
rect 369306 124908 369362 124944
rect 369306 124888 369308 124908
rect 369308 124888 369360 124908
rect 369360 124888 369362 124908
rect 362774 123936 362830 123992
rect 365166 123936 365222 123992
rect 370226 129004 370228 129024
rect 370228 129004 370280 129024
rect 370280 129004 370282 129024
rect 370226 128968 370282 129004
rect 370042 128560 370098 128616
rect 370134 125704 370190 125760
rect 369858 124344 369914 124400
rect 370318 127336 370374 127392
rect 370226 124616 370282 124672
rect 370410 126248 370466 126304
rect 371238 196560 371294 196616
rect 370778 136992 370834 137048
rect 370870 134816 370926 134872
rect 371238 126384 371294 126440
rect 371422 153720 371478 153776
rect 371422 152632 371478 152688
rect 371422 151544 371478 151600
rect 371422 150456 371478 150512
rect 371422 149912 371478 149968
rect 371422 148824 371478 148880
rect 371422 147192 371478 147248
rect 371422 146140 371424 146160
rect 371424 146140 371476 146160
rect 371476 146140 371478 146160
rect 371422 146104 371478 146140
rect 371422 145016 371478 145072
rect 371422 144472 371478 144528
rect 371422 144064 371478 144120
rect 371422 143520 371478 143576
rect 371422 142432 371478 142488
rect 371422 141924 371424 141944
rect 371424 141924 371476 141944
rect 371476 141924 371478 141944
rect 371422 141888 371478 141924
rect 371422 139712 371478 139768
rect 371422 139168 371478 139224
rect 371422 138660 371424 138680
rect 371424 138660 371476 138680
rect 371476 138660 371478 138680
rect 371422 138624 371478 138660
rect 372250 341128 372306 341184
rect 372158 293428 372160 293448
rect 372160 293428 372212 293448
rect 372212 293428 372214 293448
rect 372158 293392 372214 293428
rect 372158 291216 372214 291272
rect 372158 281016 372214 281072
rect 372066 271904 372122 271960
rect 372526 346568 372582 346624
rect 372434 279928 372490 279984
rect 372802 349832 372858 349888
rect 372894 296656 372950 296712
rect 372802 277888 372858 277944
rect 372526 274624 372582 274680
rect 372250 270136 372306 270192
rect 372066 219680 372122 219736
rect 372066 212744 372122 212800
rect 372066 202544 372122 202600
rect 371974 200368 372030 200424
rect 371882 198736 371938 198792
rect 371790 197648 371846 197704
rect 371606 127880 371662 127936
rect 371514 126248 371570 126304
rect 371330 125160 371386 125216
rect 371238 124616 371294 124672
rect 370686 124208 370742 124264
rect 372250 225684 372306 225720
rect 372250 225664 372252 225684
rect 372252 225664 372304 225684
rect 372304 225664 372306 225684
rect 372526 225004 372582 225040
rect 372526 224984 372528 225004
rect 372528 224984 372580 225004
rect 372580 224984 372582 225004
rect 372618 218592 372674 218648
rect 372342 215484 372398 215520
rect 372342 215464 372344 215484
rect 372344 215464 372396 215484
rect 372396 215464 372398 215484
rect 372802 220224 372858 220280
rect 372250 212200 372306 212256
rect 372710 210060 372712 210080
rect 372712 210060 372764 210080
rect 372764 210060 372766 210080
rect 372710 210024 372766 210060
rect 372158 199824 372214 199880
rect 372066 199280 372122 199336
rect 372158 198872 372214 198928
rect 372066 159296 372122 159352
rect 371974 153176 372030 153232
rect 371882 152088 371938 152144
rect 371974 151000 372030 151056
rect 371974 149368 372030 149424
rect 372526 148280 372582 148336
rect 371974 147736 372030 147792
rect 371974 146648 372030 146704
rect 371974 145560 372030 145616
rect 371974 142976 372030 143032
rect 371974 141344 372030 141400
rect 372066 140800 372122 140856
rect 373262 153040 373318 153096
rect 371974 140292 371976 140312
rect 371976 140292 372028 140312
rect 372028 140292 372030 140312
rect 371974 140256 372030 140292
rect 371974 138080 372030 138136
rect 371882 128560 371938 128616
rect 371790 125704 371846 125760
rect 375746 208392 375802 208448
rect 445206 369416 445262 369472
rect 445666 368328 445722 368384
rect 445666 367124 445722 367160
rect 445666 367104 445668 367124
rect 445668 367104 445720 367124
rect 445720 367104 445722 367124
rect 445298 366016 445354 366072
rect 445666 364792 445722 364848
rect 444930 363704 444986 363760
rect 445206 362480 445262 362536
rect 445114 361392 445170 361448
rect 444562 360168 444618 360224
rect 444562 357856 444618 357912
rect 444378 356768 444434 356824
rect 444746 355544 444802 355600
rect 444746 353232 444802 353288
rect 444470 352144 444526 352200
rect 444378 350920 444434 350976
rect 441802 225020 441804 225040
rect 441804 225020 441856 225040
rect 441856 225020 441858 225040
rect 441802 224984 441858 225020
rect 441802 224204 441804 224224
rect 441804 224204 441856 224224
rect 441856 224204 441858 224224
rect 441802 224168 441858 224204
rect 444470 349832 444526 349888
rect 445666 348608 445722 348664
rect 444654 347520 444710 347576
rect 445298 346296 445354 346352
rect 445666 345208 445722 345264
rect 445666 343984 445722 344040
rect 445022 342896 445078 342952
rect 444562 341672 444618 341728
rect 444562 340584 444618 340640
rect 445666 297472 445722 297528
rect 445666 296384 445722 296440
rect 445850 359080 445906 359136
rect 445666 295160 445722 295216
rect 445666 294072 445722 294128
rect 445666 292848 445722 292904
rect 445666 291760 445722 291816
rect 445666 290536 445722 290592
rect 445666 289448 445722 289504
rect 445666 288224 445722 288280
rect 445482 287136 445538 287192
rect 445666 285948 445668 285968
rect 445668 285948 445720 285968
rect 445720 285948 445722 285968
rect 445666 285912 445722 285948
rect 445390 284844 445446 284880
rect 445390 284824 445392 284844
rect 445392 284824 445444 284844
rect 445444 284824 445446 284844
rect 445666 283620 445722 283656
rect 445666 283600 445668 283620
rect 445668 283600 445720 283620
rect 445720 283600 445722 283620
rect 445666 281324 445668 281344
rect 445668 281324 445720 281344
rect 445720 281324 445722 281344
rect 445666 281288 445722 281324
rect 445022 280236 445024 280256
rect 445024 280236 445076 280256
rect 445076 280236 445078 280256
rect 445022 280200 445078 280236
rect 444654 278976 444710 279032
rect 444470 277888 444526 277944
rect 444562 268676 444564 268696
rect 444564 268676 444616 268696
rect 444616 268676 444618 268696
rect 444562 268640 444618 268676
rect 444562 223080 444618 223136
rect 444562 210468 444564 210488
rect 444564 210468 444616 210488
rect 444616 210468 444618 210488
rect 444562 210432 444618 210468
rect 445666 276684 445722 276720
rect 445666 276664 445668 276684
rect 445668 276664 445720 276684
rect 445720 276664 445722 276684
rect 445666 275576 445722 275632
rect 445666 274352 445722 274408
rect 445022 273264 445078 273320
rect 445666 272040 445722 272096
rect 445666 270952 445722 271008
rect 445390 269764 445392 269784
rect 445392 269764 445444 269784
rect 445444 269764 445446 269784
rect 445390 269728 445446 269764
rect 445666 221992 445722 222048
rect 445114 220768 445170 220824
rect 445666 219680 445722 219736
rect 445666 218456 445722 218512
rect 445942 354456 445998 354512
rect 445850 282512 445906 282568
rect 445666 217368 445722 217424
rect 445666 216164 445722 216200
rect 445666 216144 445668 216164
rect 445668 216144 445720 216164
rect 445720 216144 445722 216164
rect 445666 215056 445722 215112
rect 445666 213868 445668 213888
rect 445668 213868 445720 213888
rect 445720 213868 445722 213888
rect 445666 213832 445722 213868
rect 445298 212780 445300 212800
rect 445300 212780 445352 212800
rect 445352 212780 445354 212800
rect 445298 212744 445354 212780
rect 445666 211556 445668 211576
rect 445668 211556 445720 211576
rect 445720 211556 445722 211576
rect 445666 211520 445722 211556
rect 445666 209228 445722 209264
rect 445666 209208 445668 209228
rect 445668 209208 445720 209228
rect 445720 209208 445722 209228
rect 445114 208156 445116 208176
rect 445116 208156 445168 208176
rect 445168 208156 445170 208176
rect 445114 208120 445170 208156
rect 444746 206896 444802 206952
rect 444470 205808 444526 205864
rect 372526 125160 372582 125216
rect 372434 124208 372490 124264
rect 441802 148960 441858 149016
rect 441802 129784 441858 129840
rect 442998 129240 443054 129296
rect 441894 126384 441950 126440
rect 441802 125468 441804 125488
rect 441804 125468 441856 125488
rect 441856 125468 441858 125488
rect 441802 125432 441858 125468
rect 441802 124908 441858 124944
rect 441802 124888 441804 124908
rect 441804 124888 441856 124908
rect 441856 124888 441858 124908
rect 444378 147736 444434 147792
rect 444378 146548 444380 146568
rect 444380 146548 444432 146568
rect 444432 146548 444434 146568
rect 444378 146512 444434 146548
rect 444378 136176 444434 136232
rect 444562 140800 444618 140856
rect 444470 133864 444526 133920
rect 444470 132640 444526 132696
rect 443642 128016 443698 128072
rect 443274 125704 443330 125760
rect 445298 204584 445354 204640
rect 445022 203496 445078 203552
rect 445666 202272 445722 202328
rect 445666 201184 445722 201240
rect 445666 199960 445722 200016
rect 445666 198872 445722 198928
rect 445390 197668 445446 197704
rect 445390 197648 445392 197668
rect 445392 197648 445444 197668
rect 445444 197648 445446 197668
rect 444930 153448 444986 153504
rect 444930 151136 444986 151192
rect 444930 150048 444986 150104
rect 445666 152360 445722 152416
rect 445666 145424 445722 145480
rect 445298 144200 445354 144256
rect 445206 143112 445262 143168
rect 445114 141924 445116 141944
rect 445116 141924 445168 141944
rect 445168 141924 445170 141944
rect 445114 141888 445170 141924
rect 445114 139576 445170 139632
rect 444838 137264 444894 137320
rect 444746 134952 444802 135008
rect 445666 131552 445722 131608
rect 444838 130328 444894 130384
rect 444838 129240 444894 129296
rect 445666 126928 445722 126984
rect 445850 196560 445906 196616
rect 445942 138488 445998 138544
rect 454222 159296 454278 159352
rect 580170 697176 580226 697232
rect 580170 683848 580226 683904
rect 580170 670692 580172 670712
rect 580172 670692 580224 670712
rect 580224 670692 580226 670712
rect 580170 670656 580226 670692
rect 580170 644000 580226 644056
rect 580170 630808 580226 630864
rect 580170 617480 580226 617536
rect 579802 590960 579858 591016
rect 580170 577632 580226 577688
rect 579802 564304 579858 564360
rect 580170 537784 580226 537840
rect 580170 524476 580226 524512
rect 580170 524456 580172 524476
rect 580172 524456 580224 524476
rect 580224 524456 580226 524476
rect 580170 511264 580226 511320
rect 580170 484608 580226 484664
rect 579986 471416 580042 471472
rect 580170 458088 580226 458144
rect 580170 431568 580226 431624
rect 580170 418240 580226 418296
rect 580170 404912 580226 404968
rect 582378 378392 582434 378448
rect 580170 325216 580226 325272
rect 580170 312024 580226 312080
rect 582470 365064 582526 365120
rect 582562 351872 582618 351928
rect 579894 298696 579950 298752
rect 579894 272176 579950 272232
rect 580262 258848 580318 258904
rect 580170 245556 580172 245576
rect 580172 245556 580224 245576
rect 580224 245556 580226 245576
rect 580170 245520 580226 245556
rect 579986 232328 580042 232384
rect 579894 219000 579950 219056
rect 580262 192480 580318 192536
rect 580170 179152 580226 179208
rect 579618 152632 579674 152688
rect 580170 139340 580172 139360
rect 580172 139340 580224 139360
rect 580224 139340 580226 139360
rect 580170 139304 580226 139340
rect 579802 112784 579858 112840
rect 350446 3440 350502 3496
rect 349250 3304 349306 3360
rect 580170 99456 580226 99512
rect 458822 98912 458878 98968
rect 461582 97416 461638 97472
rect 543738 98776 543794 98832
rect 536838 94696 536894 94752
rect 550638 98640 550694 98696
rect 580262 97280 580318 97336
rect 557538 95784 557594 95840
rect 561678 94560 561734 94616
rect 568578 94424 568634 94480
rect 575478 93064 575534 93120
rect 579986 72936 580042 72992
rect 580170 59608 580226 59664
rect 582562 86128 582618 86184
rect 583022 205672 583078 205728
rect 582930 165824 582986 165880
rect 582838 125976 582894 126032
rect 582838 97144 582894 97200
rect 582654 46280 582710 46336
rect 582470 19760 582526 19816
rect 582378 6568 582434 6624
rect 583114 33088 583170 33144
<< metal3 >>
rect -960 697220 480 697460
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 580165 683906 580231 683909
rect 583520 683906 584960 683996
rect 580165 683904 584960 683906
rect 580165 683848 580170 683904
rect 580226 683848 584960 683904
rect 580165 683846 584960 683848
rect 580165 683843 580231 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3417 671258 3483 671261
rect -960 671256 3483 671258
rect -960 671200 3422 671256
rect 3478 671200 3483 671256
rect -960 671198 3483 671200
rect -960 671108 480 671198
rect 3417 671195 3483 671198
rect 580165 670714 580231 670717
rect 583520 670714 584960 670804
rect 580165 670712 584960 670714
rect 580165 670656 580170 670712
rect 580226 670656 584960 670712
rect 580165 670654 584960 670656
rect 580165 670651 580231 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3509 658202 3575 658205
rect -960 658200 3575 658202
rect -960 658144 3514 658200
rect 3570 658144 3575 658200
rect -960 658142 3575 658144
rect -960 658052 480 658142
rect 3509 658139 3575 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 580165 644058 580231 644061
rect 583520 644058 584960 644148
rect 580165 644056 584960 644058
rect 580165 644000 580170 644056
rect 580226 644000 584960 644056
rect 580165 643998 584960 644000
rect 580165 643995 580231 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 3509 632090 3575 632093
rect -960 632088 3575 632090
rect -960 632032 3514 632088
rect 3570 632032 3575 632088
rect -960 632030 3575 632032
rect -960 631940 480 632030
rect 3509 632027 3575 632030
rect 580165 630866 580231 630869
rect 583520 630866 584960 630956
rect 580165 630864 584960 630866
rect 580165 630808 580170 630864
rect 580226 630808 584960 630864
rect 580165 630806 584960 630808
rect 580165 630803 580231 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3509 619170 3575 619173
rect -960 619168 3575 619170
rect -960 619112 3514 619168
rect 3570 619112 3575 619168
rect -960 619110 3575 619112
rect -960 619020 480 619110
rect 3509 619107 3575 619110
rect 580165 617538 580231 617541
rect 583520 617538 584960 617628
rect 580165 617536 584960 617538
rect 580165 617480 580170 617536
rect 580226 617480 584960 617536
rect 580165 617478 584960 617480
rect 580165 617475 580231 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3509 606114 3575 606117
rect -960 606112 3575 606114
rect -960 606056 3514 606112
rect 3570 606056 3575 606112
rect -960 606054 3575 606056
rect -960 605964 480 606054
rect 3509 606051 3575 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 579797 591018 579863 591021
rect 583520 591018 584960 591108
rect 579797 591016 584960 591018
rect 579797 590960 579802 591016
rect 579858 590960 584960 591016
rect 579797 590958 584960 590960
rect 579797 590955 579863 590958
rect 583520 590868 584960 590958
rect -960 580002 480 580092
rect 3325 580002 3391 580005
rect -960 580000 3391 580002
rect -960 579944 3330 580000
rect 3386 579944 3391 580000
rect -960 579942 3391 579944
rect -960 579852 480 579942
rect 3325 579939 3391 579942
rect 580165 577690 580231 577693
rect 583520 577690 584960 577780
rect 580165 577688 584960 577690
rect 580165 577632 580170 577688
rect 580226 577632 584960 577688
rect 580165 577630 584960 577632
rect 580165 577627 580231 577630
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 3233 566946 3299 566949
rect -960 566944 3299 566946
rect -960 566888 3238 566944
rect 3294 566888 3299 566944
rect -960 566886 3299 566888
rect -960 566796 480 566886
rect 3233 566883 3299 566886
rect 579797 564362 579863 564365
rect 583520 564362 584960 564452
rect 579797 564360 584960 564362
rect 579797 564304 579802 564360
rect 579858 564304 584960 564360
rect 579797 564302 584960 564304
rect 579797 564299 579863 564302
rect 583520 564212 584960 564302
rect -960 553890 480 553980
rect 3325 553890 3391 553893
rect -960 553888 3391 553890
rect -960 553832 3330 553888
rect 3386 553832 3391 553888
rect -960 553830 3391 553832
rect -960 553740 480 553830
rect 3325 553827 3391 553830
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 580165 537842 580231 537845
rect 583520 537842 584960 537932
rect 580165 537840 584960 537842
rect 580165 537784 580170 537840
rect 580226 537784 584960 537840
rect 580165 537782 584960 537784
rect 580165 537779 580231 537782
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect 2957 527914 3023 527917
rect -960 527912 3023 527914
rect -960 527856 2962 527912
rect 3018 527856 3023 527912
rect -960 527854 3023 527856
rect -960 527764 480 527854
rect 2957 527851 3023 527854
rect 580165 524514 580231 524517
rect 583520 524514 584960 524604
rect 580165 524512 584960 524514
rect 580165 524456 580170 524512
rect 580226 524456 584960 524512
rect 580165 524454 584960 524456
rect 580165 524451 580231 524454
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 3509 514858 3575 514861
rect -960 514856 3575 514858
rect -960 514800 3514 514856
rect 3570 514800 3575 514856
rect -960 514798 3575 514800
rect -960 514708 480 514798
rect 3509 514795 3575 514798
rect 580165 511322 580231 511325
rect 583520 511322 584960 511412
rect 580165 511320 584960 511322
rect 580165 511264 580170 511320
rect 580226 511264 584960 511320
rect 580165 511262 584960 511264
rect 580165 511259 580231 511262
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect 3049 501802 3115 501805
rect -960 501800 3115 501802
rect -960 501744 3054 501800
rect 3110 501744 3115 501800
rect -960 501742 3115 501744
rect -960 501652 480 501742
rect 3049 501739 3115 501742
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 580165 484666 580231 484669
rect 583520 484666 584960 484756
rect 580165 484664 584960 484666
rect 580165 484608 580170 484664
rect 580226 484608 584960 484664
rect 580165 484606 584960 484608
rect 580165 484603 580231 484606
rect 583520 484516 584960 484606
rect -960 475690 480 475780
rect 3049 475690 3115 475693
rect -960 475688 3115 475690
rect -960 475632 3054 475688
rect 3110 475632 3115 475688
rect -960 475630 3115 475632
rect -960 475540 480 475630
rect 3049 475627 3115 475630
rect 579981 471474 580047 471477
rect 583520 471474 584960 471564
rect 579981 471472 584960 471474
rect 579981 471416 579986 471472
rect 580042 471416 584960 471472
rect 579981 471414 584960 471416
rect 579981 471411 580047 471414
rect 583520 471324 584960 471414
rect -960 462634 480 462724
rect 3509 462634 3575 462637
rect -960 462632 3575 462634
rect -960 462576 3514 462632
rect 3570 462576 3575 462632
rect -960 462574 3575 462576
rect -960 462484 480 462574
rect 3509 462571 3575 462574
rect 580165 458146 580231 458149
rect 583520 458146 584960 458236
rect 580165 458144 584960 458146
rect 580165 458088 580170 458144
rect 580226 458088 584960 458144
rect 580165 458086 584960 458088
rect 580165 458083 580231 458086
rect 583520 457996 584960 458086
rect -960 449578 480 449668
rect 3141 449578 3207 449581
rect -960 449576 3207 449578
rect -960 449520 3146 449576
rect 3202 449520 3207 449576
rect -960 449518 3207 449520
rect -960 449428 480 449518
rect 3141 449515 3207 449518
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 580165 431626 580231 431629
rect 583520 431626 584960 431716
rect 580165 431624 584960 431626
rect 580165 431568 580170 431624
rect 580226 431568 584960 431624
rect 580165 431566 584960 431568
rect 580165 431563 580231 431566
rect 583520 431476 584960 431566
rect -960 423602 480 423692
rect 3509 423602 3575 423605
rect -960 423600 3575 423602
rect -960 423544 3514 423600
rect 3570 423544 3575 423600
rect -960 423542 3575 423544
rect -960 423452 480 423542
rect 3509 423539 3575 423542
rect 580165 418298 580231 418301
rect 583520 418298 584960 418388
rect 580165 418296 584960 418298
rect 580165 418240 580170 418296
rect 580226 418240 584960 418296
rect 580165 418238 584960 418240
rect 580165 418235 580231 418238
rect 583520 418148 584960 418238
rect -960 410546 480 410636
rect 2865 410546 2931 410549
rect -960 410544 2931 410546
rect -960 410488 2870 410544
rect 2926 410488 2931 410544
rect -960 410486 2931 410488
rect -960 410396 480 410486
rect 2865 410483 2931 410486
rect 580165 404970 580231 404973
rect 583520 404970 584960 405060
rect 580165 404968 584960 404970
rect 580165 404912 580170 404968
rect 580226 404912 584960 404968
rect 580165 404910 584960 404912
rect 580165 404907 580231 404910
rect 583520 404820 584960 404910
rect -960 397490 480 397580
rect 3509 397490 3575 397493
rect -960 397488 3575 397490
rect -960 397432 3514 397488
rect 3570 397432 3575 397488
rect -960 397430 3575 397432
rect -960 397340 480 397430
rect 3509 397427 3575 397430
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 582373 378450 582439 378453
rect 583520 378450 584960 378540
rect 582373 378448 584960 378450
rect 582373 378392 582378 378448
rect 582434 378392 584960 378448
rect 582373 378390 584960 378392
rect 582373 378387 582439 378390
rect 583520 378300 584960 378390
rect -960 371378 480 371468
rect 3509 371378 3575 371381
rect -960 371376 3575 371378
rect -960 371320 3514 371376
rect 3570 371320 3575 371376
rect -960 371318 3575 371320
rect -960 371228 480 371318
rect 3509 371315 3575 371318
rect 371877 369746 371943 369749
rect 369932 369744 371943 369746
rect 369932 369688 371882 369744
rect 371938 369688 371943 369744
rect 369932 369686 371943 369688
rect 371877 369683 371943 369686
rect 445201 369474 445267 369477
rect 441876 369472 445267 369474
rect 441876 369416 445206 369472
rect 445262 369416 445267 369472
rect 441876 369414 445267 369416
rect 445201 369411 445267 369414
rect 371601 369202 371667 369205
rect 369932 369200 371667 369202
rect 369932 369144 371606 369200
rect 371662 369144 371667 369200
rect 369932 369142 371667 369144
rect 371601 369139 371667 369142
rect 372061 368658 372127 368661
rect 369932 368656 372127 368658
rect 369932 368600 372066 368656
rect 372122 368600 372127 368656
rect 369932 368598 372127 368600
rect 372061 368595 372127 368598
rect 445661 368386 445727 368389
rect 441876 368384 445727 368386
rect 441876 368328 445666 368384
rect 445722 368328 445727 368384
rect 441876 368326 445727 368328
rect 445661 368323 445727 368326
rect 371693 368114 371759 368117
rect 369932 368112 371759 368114
rect 369932 368056 371698 368112
rect 371754 368056 371759 368112
rect 369932 368054 371759 368056
rect 371693 368051 371759 368054
rect 371601 367570 371667 367573
rect 369932 367568 371667 367570
rect 369932 367512 371606 367568
rect 371662 367512 371667 367568
rect 369932 367510 371667 367512
rect 371601 367507 371667 367510
rect 445661 367162 445727 367165
rect 441876 367160 445727 367162
rect 441876 367104 445666 367160
rect 445722 367104 445727 367160
rect 441876 367102 445727 367104
rect 445661 367099 445727 367102
rect 371233 367026 371299 367029
rect 369932 367024 371299 367026
rect 369932 366968 371238 367024
rect 371294 366968 371299 367024
rect 369932 366966 371299 366968
rect 371233 366963 371299 366966
rect 371509 366482 371575 366485
rect 369932 366480 371575 366482
rect 369932 366424 371514 366480
rect 371570 366424 371575 366480
rect 369932 366422 371575 366424
rect 371509 366419 371575 366422
rect 445293 366074 445359 366077
rect 441876 366072 445359 366074
rect 441876 366016 445298 366072
rect 445354 366016 445359 366072
rect 441876 366014 445359 366016
rect 445293 366011 445359 366014
rect 371601 365938 371667 365941
rect 369932 365936 371667 365938
rect 369932 365880 371606 365936
rect 371662 365880 371667 365936
rect 369932 365878 371667 365880
rect 371601 365875 371667 365878
rect 371233 365394 371299 365397
rect 369932 365392 371299 365394
rect 369932 365336 371238 365392
rect 371294 365336 371299 365392
rect 369932 365334 371299 365336
rect 371233 365331 371299 365334
rect 582465 365122 582531 365125
rect 583520 365122 584960 365212
rect 582465 365120 584960 365122
rect 582465 365064 582470 365120
rect 582526 365064 584960 365120
rect 582465 365062 584960 365064
rect 582465 365059 582531 365062
rect 583520 364972 584960 365062
rect 371601 364850 371667 364853
rect 445661 364850 445727 364853
rect 369932 364848 371667 364850
rect 369932 364792 371606 364848
rect 371662 364792 371667 364848
rect 369932 364790 371667 364792
rect 441876 364848 445727 364850
rect 441876 364792 445666 364848
rect 445722 364792 445727 364848
rect 441876 364790 445727 364792
rect 371601 364787 371667 364790
rect 445661 364787 445727 364790
rect 371693 364306 371759 364309
rect 369932 364304 371759 364306
rect 369932 364248 371698 364304
rect 371754 364248 371759 364304
rect 369932 364246 371759 364248
rect 371693 364243 371759 364246
rect 371601 363762 371667 363765
rect 444925 363762 444991 363765
rect 369932 363760 371667 363762
rect 369932 363704 371606 363760
rect 371662 363704 371667 363760
rect 369932 363702 371667 363704
rect 441876 363760 444991 363762
rect 441876 363704 444930 363760
rect 444986 363704 444991 363760
rect 441876 363702 444991 363704
rect 371601 363699 371667 363702
rect 444925 363699 444991 363702
rect 372521 363218 372587 363221
rect 369932 363216 372587 363218
rect 369932 363160 372526 363216
rect 372582 363160 372587 363216
rect 369932 363158 372587 363160
rect 372521 363155 372587 363158
rect 371693 362674 371759 362677
rect 369932 362672 371759 362674
rect 369932 362616 371698 362672
rect 371754 362616 371759 362672
rect 369932 362614 371759 362616
rect 371693 362611 371759 362614
rect 445201 362538 445267 362541
rect 441876 362536 445267 362538
rect 441876 362480 445206 362536
rect 445262 362480 445267 362536
rect 441876 362478 445267 362480
rect 445201 362475 445267 362478
rect 371601 362130 371667 362133
rect 369932 362128 371667 362130
rect 369932 362072 371606 362128
rect 371662 362072 371667 362128
rect 369932 362070 371667 362072
rect 371601 362067 371667 362070
rect 371601 361586 371667 361589
rect 369932 361584 371667 361586
rect 369932 361528 371606 361584
rect 371662 361528 371667 361584
rect 369932 361526 371667 361528
rect 371601 361523 371667 361526
rect 445109 361450 445175 361453
rect 441876 361448 445175 361450
rect 441876 361392 445114 361448
rect 445170 361392 445175 361448
rect 441876 361390 445175 361392
rect 445109 361387 445175 361390
rect 371417 361042 371483 361045
rect 369932 361040 371483 361042
rect 369932 360984 371422 361040
rect 371478 360984 371483 361040
rect 369932 360982 371483 360984
rect 371417 360979 371483 360982
rect 371601 360498 371667 360501
rect 369932 360496 371667 360498
rect 369932 360440 371606 360496
rect 371662 360440 371667 360496
rect 369932 360438 371667 360440
rect 371601 360435 371667 360438
rect 444557 360226 444623 360229
rect 441876 360224 444623 360226
rect 441876 360168 444562 360224
rect 444618 360168 444623 360224
rect 441876 360166 444623 360168
rect 444557 360163 444623 360166
rect 372337 360090 372403 360093
rect 369932 360088 372403 360090
rect 369932 360032 372342 360088
rect 372398 360032 372403 360088
rect 369932 360030 372403 360032
rect 372337 360027 372403 360030
rect 372153 359546 372219 359549
rect 369932 359544 372219 359546
rect 369932 359488 372158 359544
rect 372214 359488 372219 359544
rect 369932 359486 372219 359488
rect 372153 359483 372219 359486
rect 445845 359138 445911 359141
rect 441876 359136 445911 359138
rect 441876 359080 445850 359136
rect 445906 359080 445911 359136
rect 441876 359078 445911 359080
rect 445845 359075 445911 359078
rect 371969 359002 372035 359005
rect 369932 359000 372035 359002
rect 369932 358944 371974 359000
rect 372030 358944 372035 359000
rect 369932 358942 372035 358944
rect 371969 358939 372035 358942
rect -960 358458 480 358548
rect 3141 358458 3207 358461
rect 371693 358458 371759 358461
rect -960 358456 3207 358458
rect -960 358400 3146 358456
rect 3202 358400 3207 358456
rect -960 358398 3207 358400
rect 369932 358456 371759 358458
rect 369932 358400 371698 358456
rect 371754 358400 371759 358456
rect 369932 358398 371759 358400
rect -960 358308 480 358398
rect 3141 358395 3207 358398
rect 371693 358395 371759 358398
rect 371601 357914 371667 357917
rect 444557 357914 444623 357917
rect 369932 357912 371667 357914
rect 369932 357856 371606 357912
rect 371662 357856 371667 357912
rect 369932 357854 371667 357856
rect 441876 357912 444623 357914
rect 441876 357856 444562 357912
rect 444618 357856 444623 357912
rect 441876 357854 444623 357856
rect 371601 357851 371667 357854
rect 444557 357851 444623 357854
rect 371601 357370 371667 357373
rect 369932 357368 371667 357370
rect 369932 357312 371606 357368
rect 371662 357312 371667 357368
rect 369932 357310 371667 357312
rect 371601 357307 371667 357310
rect 371509 356826 371575 356829
rect 444373 356826 444439 356829
rect 369932 356824 371575 356826
rect 369932 356768 371514 356824
rect 371570 356768 371575 356824
rect 369932 356766 371575 356768
rect 441876 356824 444439 356826
rect 441876 356768 444378 356824
rect 444434 356768 444439 356824
rect 441876 356766 444439 356768
rect 371509 356763 371575 356766
rect 444373 356763 444439 356766
rect 371233 356282 371299 356285
rect 369932 356280 371299 356282
rect 369932 356224 371238 356280
rect 371294 356224 371299 356280
rect 369932 356222 371299 356224
rect 371233 356219 371299 356222
rect 371601 355738 371667 355741
rect 369932 355736 371667 355738
rect 369932 355680 371606 355736
rect 371662 355680 371667 355736
rect 369932 355678 371667 355680
rect 371601 355675 371667 355678
rect 444741 355602 444807 355605
rect 441876 355600 444807 355602
rect 441876 355544 444746 355600
rect 444802 355544 444807 355600
rect 441876 355542 444807 355544
rect 444741 355539 444807 355542
rect 371509 355194 371575 355197
rect 369932 355192 371575 355194
rect 369932 355136 371514 355192
rect 371570 355136 371575 355192
rect 369932 355134 371575 355136
rect 371509 355131 371575 355134
rect 371325 354650 371391 354653
rect 369932 354648 371391 354650
rect 369932 354592 371330 354648
rect 371386 354592 371391 354648
rect 369932 354590 371391 354592
rect 371325 354587 371391 354590
rect 445937 354514 446003 354517
rect 441876 354512 446003 354514
rect 441876 354456 445942 354512
rect 445998 354456 446003 354512
rect 441876 354454 446003 354456
rect 445937 354451 446003 354454
rect 371693 354106 371759 354109
rect 369932 354104 371759 354106
rect 369932 354048 371698 354104
rect 371754 354048 371759 354104
rect 369932 354046 371759 354048
rect 371693 354043 371759 354046
rect 371509 353562 371575 353565
rect 369932 353560 371575 353562
rect 369932 353504 371514 353560
rect 371570 353504 371575 353560
rect 369932 353502 371575 353504
rect 371509 353499 371575 353502
rect 444741 353290 444807 353293
rect 441876 353288 444807 353290
rect 441876 353232 444746 353288
rect 444802 353232 444807 353288
rect 441876 353230 444807 353232
rect 444741 353227 444807 353230
rect 371969 353018 372035 353021
rect 369932 353016 372035 353018
rect 369932 352960 371974 353016
rect 372030 352960 372035 353016
rect 369932 352958 372035 352960
rect 371969 352955 372035 352958
rect 372102 352474 372108 352476
rect 369932 352414 372108 352474
rect 372102 352412 372108 352414
rect 372172 352412 372178 352476
rect 444465 352202 444531 352205
rect 441876 352200 444531 352202
rect 441876 352144 444470 352200
rect 444526 352144 444531 352200
rect 441876 352142 444531 352144
rect 444465 352139 444531 352142
rect 372429 351930 372495 351933
rect 369932 351928 372495 351930
rect 369932 351872 372434 351928
rect 372490 351872 372495 351928
rect 369932 351870 372495 351872
rect 372429 351867 372495 351870
rect 582557 351930 582623 351933
rect 583520 351930 584960 352020
rect 582557 351928 584960 351930
rect 582557 351872 582562 351928
rect 582618 351872 584960 351928
rect 582557 351870 584960 351872
rect 582557 351867 582623 351870
rect 583520 351780 584960 351870
rect 371734 351386 371740 351388
rect 369932 351326 371740 351386
rect 371734 351324 371740 351326
rect 371804 351324 371810 351388
rect 444373 350978 444439 350981
rect 441876 350976 444439 350978
rect 441876 350920 444378 350976
rect 444434 350920 444439 350976
rect 441876 350918 444439 350920
rect 444373 350915 444439 350918
rect 371366 350842 371372 350844
rect 369932 350782 371372 350842
rect 371366 350780 371372 350782
rect 371436 350780 371442 350844
rect 369301 350570 369367 350573
rect 369301 350568 369410 350570
rect 369301 350512 369306 350568
rect 369362 350512 369410 350568
rect 369301 350507 369410 350512
rect 369350 350268 369410 350507
rect 372797 349890 372863 349893
rect 444465 349890 444531 349893
rect 369932 349888 372863 349890
rect 369932 349832 372802 349888
rect 372858 349832 372863 349888
rect 369932 349830 372863 349832
rect 441876 349888 444531 349890
rect 441876 349832 444470 349888
rect 444526 349832 444531 349888
rect 441876 349830 444531 349832
rect 372797 349827 372863 349830
rect 444465 349827 444531 349830
rect 371601 349346 371667 349349
rect 369932 349344 371667 349346
rect 369932 349288 371606 349344
rect 371662 349288 371667 349344
rect 369932 349286 371667 349288
rect 371601 349283 371667 349286
rect 370313 348802 370379 348805
rect 369932 348800 370379 348802
rect 369932 348744 370318 348800
rect 370374 348744 370379 348800
rect 369932 348742 370379 348744
rect 370313 348739 370379 348742
rect 445661 348666 445727 348669
rect 441876 348664 445727 348666
rect 441876 348608 445666 348664
rect 445722 348608 445727 348664
rect 441876 348606 445727 348608
rect 445661 348603 445727 348606
rect 371601 348258 371667 348261
rect 369932 348256 371667 348258
rect 369932 348200 371606 348256
rect 371662 348200 371667 348256
rect 369932 348198 371667 348200
rect 371601 348195 371667 348198
rect 369350 347445 369410 347684
rect 444649 347578 444715 347581
rect 441876 347576 444715 347578
rect 441876 347520 444654 347576
rect 444710 347520 444715 347576
rect 441876 347518 444715 347520
rect 444649 347515 444715 347518
rect 369350 347440 369459 347445
rect 369350 347384 369398 347440
rect 369454 347384 369459 347440
rect 369350 347382 369459 347384
rect 369393 347379 369459 347382
rect 370405 347170 370471 347173
rect 369932 347168 370471 347170
rect 369932 347112 370410 347168
rect 370466 347112 370471 347168
rect 369932 347110 370471 347112
rect 370405 347107 370471 347110
rect 372521 346626 372587 346629
rect 369932 346624 372587 346626
rect 369932 346568 372526 346624
rect 372582 346568 372587 346624
rect 369932 346566 372587 346568
rect 372521 346563 372587 346566
rect 445293 346354 445359 346357
rect 441876 346352 445359 346354
rect 441876 346296 445298 346352
rect 445354 346296 445359 346352
rect 441876 346294 445359 346296
rect 445293 346291 445359 346294
rect 369902 345813 369962 346052
rect 369853 345808 369962 345813
rect 369853 345752 369858 345808
rect 369914 345752 369962 345808
rect 369853 345750 369962 345752
rect 369853 345747 369919 345750
rect 370221 345538 370287 345541
rect 369932 345536 370287 345538
rect -960 345402 480 345492
rect 369932 345480 370226 345536
rect 370282 345480 370287 345536
rect 369932 345478 370287 345480
rect 370221 345475 370287 345478
rect 3325 345402 3391 345405
rect -960 345400 3391 345402
rect -960 345344 3330 345400
rect 3386 345344 3391 345400
rect -960 345342 3391 345344
rect -960 345252 480 345342
rect 3325 345339 3391 345342
rect 445661 345266 445727 345269
rect 441876 345264 445727 345266
rect 441876 345208 445666 345264
rect 445722 345208 445727 345264
rect 441876 345206 445727 345208
rect 445661 345203 445727 345206
rect 371877 344994 371943 344997
rect 369932 344992 371943 344994
rect 369932 344936 371882 344992
rect 371938 344936 371943 344992
rect 369932 344934 371943 344936
rect 371877 344931 371943 344934
rect 371417 344450 371483 344453
rect 369932 344448 371483 344450
rect 369932 344392 371422 344448
rect 371478 344392 371483 344448
rect 369932 344390 371483 344392
rect 371417 344387 371483 344390
rect 445661 344042 445727 344045
rect 441876 344040 445727 344042
rect 441876 343984 445666 344040
rect 445722 343984 445727 344040
rect 441876 343982 445727 343984
rect 445661 343979 445727 343982
rect 372061 343906 372127 343909
rect 369932 343904 372127 343906
rect 369932 343848 372066 343904
rect 372122 343848 372127 343904
rect 369932 343846 372127 343848
rect 372061 343843 372127 343846
rect 371182 343362 371188 343364
rect 369932 343302 371188 343362
rect 371182 343300 371188 343302
rect 371252 343300 371258 343364
rect 445017 342954 445083 342957
rect 441876 342952 445083 342954
rect 441876 342896 445022 342952
rect 445078 342896 445083 342952
rect 441876 342894 445083 342896
rect 445017 342891 445083 342894
rect 371509 342818 371575 342821
rect 369932 342816 371575 342818
rect 369932 342760 371514 342816
rect 371570 342760 371575 342816
rect 369932 342758 371575 342760
rect 371509 342755 371575 342758
rect 371325 342274 371391 342277
rect 369932 342272 371391 342274
rect 369932 342216 371330 342272
rect 371386 342216 371391 342272
rect 369932 342214 371391 342216
rect 371325 342211 371391 342214
rect 371785 341730 371851 341733
rect 444557 341730 444623 341733
rect 369932 341728 371851 341730
rect 369932 341672 371790 341728
rect 371846 341672 371851 341728
rect 369932 341670 371851 341672
rect 441876 341728 444623 341730
rect 441876 341672 444562 341728
rect 444618 341672 444623 341728
rect 441876 341670 444623 341672
rect 371785 341667 371851 341670
rect 444557 341667 444623 341670
rect 372245 341186 372311 341189
rect 369932 341184 372311 341186
rect 369932 341128 372250 341184
rect 372306 341128 372311 341184
rect 369932 341126 372311 341128
rect 372245 341123 372311 341126
rect 370129 340642 370195 340645
rect 444557 340642 444623 340645
rect 369932 340640 370195 340642
rect 369932 340584 370134 340640
rect 370190 340584 370195 340640
rect 369932 340582 370195 340584
rect 441876 340640 444623 340642
rect 441876 340584 444562 340640
rect 444618 340584 444623 340640
rect 441876 340582 444623 340584
rect 370129 340579 370195 340582
rect 444557 340579 444623 340582
rect 370221 340234 370287 340237
rect 369932 340232 370287 340234
rect 369932 340176 370226 340232
rect 370282 340176 370287 340232
rect 369932 340174 370287 340176
rect 370221 340171 370287 340174
rect 583520 338452 584960 338692
rect 361614 337724 361620 337788
rect 361684 337786 361690 337788
rect 362861 337786 362927 337789
rect 361684 337784 362927 337786
rect 361684 337728 362866 337784
rect 362922 337728 362927 337784
rect 361684 337726 362927 337728
rect 361684 337724 361690 337726
rect 362861 337723 362927 337726
rect 364374 337724 364380 337788
rect 364444 337786 364450 337788
rect 364885 337786 364951 337789
rect 364444 337784 364951 337786
rect 364444 337728 364890 337784
rect 364946 337728 364951 337784
rect 364444 337726 364951 337728
rect 364444 337724 364450 337726
rect 364885 337723 364951 337726
rect -960 332196 480 332436
rect 580165 325274 580231 325277
rect 583520 325274 584960 325364
rect 580165 325272 584960 325274
rect 580165 325216 580170 325272
rect 580226 325216 584960 325272
rect 580165 325214 584960 325216
rect 580165 325211 580231 325214
rect 583520 325124 584960 325214
rect -960 319290 480 319380
rect 3325 319290 3391 319293
rect -960 319288 3391 319290
rect -960 319232 3330 319288
rect 3386 319232 3391 319288
rect -960 319230 3391 319232
rect -960 319140 480 319230
rect 3325 319227 3391 319230
rect 580165 312082 580231 312085
rect 583520 312082 584960 312172
rect 580165 312080 584960 312082
rect 580165 312024 580170 312080
rect 580226 312024 584960 312080
rect 580165 312022 584960 312024
rect 580165 312019 580231 312022
rect 583520 311932 584960 312022
rect -960 306234 480 306324
rect 3233 306234 3299 306237
rect -960 306232 3299 306234
rect -960 306176 3238 306232
rect 3294 306176 3299 306232
rect -960 306174 3299 306176
rect -960 306084 480 306174
rect 3233 306171 3299 306174
rect 217409 299434 217475 299437
rect 217961 299434 218027 299437
rect 217409 299432 218027 299434
rect 217409 299376 217414 299432
rect 217470 299376 217966 299432
rect 218022 299376 218027 299432
rect 217409 299374 218027 299376
rect 217409 299371 217475 299374
rect 217961 299371 218027 299374
rect 217225 299298 217291 299301
rect 217685 299298 217751 299301
rect 217225 299296 217751 299298
rect 217225 299240 217230 299296
rect 217286 299240 217690 299296
rect 217746 299240 217751 299296
rect 217225 299238 217751 299240
rect 217225 299235 217291 299238
rect 217685 299235 217751 299238
rect 198549 298890 198615 298893
rect 198549 298888 200100 298890
rect 198549 298832 198554 298888
rect 198610 298832 200100 298888
rect 198549 298830 200100 298832
rect 198549 298827 198615 298830
rect 579889 298754 579955 298757
rect 583520 298754 584960 298844
rect 579889 298752 584960 298754
rect 579889 298696 579894 298752
rect 579950 298696 584960 298752
rect 579889 298694 584960 298696
rect 579889 298691 579955 298694
rect 583520 298604 584960 298694
rect 302785 298482 302851 298485
rect 299828 298480 302851 298482
rect 299828 298424 302790 298480
rect 302846 298424 302851 298480
rect 299828 298422 302851 298424
rect 302785 298419 302851 298422
rect 369534 297397 369594 297772
rect 445661 297530 445727 297533
rect 441876 297528 445727 297530
rect 441876 297472 445666 297528
rect 445722 297472 445727 297528
rect 441876 297470 445727 297472
rect 445661 297467 445727 297470
rect 369485 297392 369594 297397
rect 369485 297336 369490 297392
rect 369546 297336 369594 297392
rect 369485 297334 369594 297336
rect 369485 297331 369551 297334
rect 369350 296853 369410 297228
rect 369350 296848 369459 296853
rect 369350 296792 369398 296848
rect 369454 296792 369459 296848
rect 369350 296790 369459 296792
rect 369393 296787 369459 296790
rect 199837 296714 199903 296717
rect 372889 296714 372955 296717
rect 199837 296712 200100 296714
rect 199837 296656 199842 296712
rect 199898 296656 200100 296712
rect 369380 296712 372955 296714
rect 369380 296684 372894 296712
rect 199837 296654 200100 296656
rect 369350 296656 372894 296684
rect 372950 296656 372955 296712
rect 369350 296654 372955 296656
rect 199837 296651 199903 296654
rect 369350 296309 369410 296654
rect 372889 296651 372955 296654
rect 445661 296442 445727 296445
rect 441876 296440 445727 296442
rect 441876 296384 445666 296440
rect 445722 296384 445727 296440
rect 441876 296382 445727 296384
rect 445661 296379 445727 296382
rect 369350 296304 369459 296309
rect 369350 296248 369398 296304
rect 369454 296248 369459 296304
rect 369350 296246 369459 296248
rect 369393 296243 369459 296246
rect 369350 295901 369410 296140
rect 369350 295896 369459 295901
rect 369350 295840 369398 295896
rect 369454 295840 369459 295896
rect 369350 295838 369459 295840
rect 369393 295835 369459 295838
rect 370129 295626 370195 295629
rect 369932 295624 370195 295626
rect 369932 295568 370134 295624
rect 370190 295568 370195 295624
rect 369932 295566 370195 295568
rect 370129 295563 370195 295566
rect 302785 295354 302851 295357
rect 299828 295352 302851 295354
rect 299828 295296 302790 295352
rect 302846 295296 302851 295352
rect 299828 295294 302851 295296
rect 302785 295291 302851 295294
rect 445661 295218 445727 295221
rect 441876 295216 445727 295218
rect 441876 295160 445666 295216
rect 445722 295160 445727 295216
rect 441876 295158 445727 295160
rect 445661 295155 445727 295158
rect 371693 295082 371759 295085
rect 369932 295080 371759 295082
rect 369932 295024 371698 295080
rect 371754 295024 371759 295080
rect 369932 295022 371759 295024
rect 371693 295019 371759 295022
rect 197905 294538 197971 294541
rect 371693 294538 371759 294541
rect 197905 294536 200100 294538
rect 197905 294480 197910 294536
rect 197966 294480 200100 294536
rect 197905 294478 200100 294480
rect 369932 294536 371759 294538
rect 369932 294480 371698 294536
rect 371754 294480 371759 294536
rect 369932 294478 371759 294480
rect 197905 294475 197971 294478
rect 371693 294475 371759 294478
rect 445661 294130 445727 294133
rect 441876 294128 445727 294130
rect 441876 294072 445666 294128
rect 445722 294072 445727 294128
rect 441876 294070 445727 294072
rect 445661 294067 445727 294070
rect 371233 293994 371299 293997
rect 369932 293992 371299 293994
rect 369932 293936 371238 293992
rect 371294 293936 371299 293992
rect 369932 293934 371299 293936
rect 371233 293931 371299 293934
rect 372153 293450 372219 293453
rect 369932 293448 372219 293450
rect 369932 293392 372158 293448
rect 372214 293392 372219 293448
rect 369932 293390 372219 293392
rect 372153 293387 372219 293390
rect -960 293178 480 293268
rect 3049 293178 3115 293181
rect -960 293176 3115 293178
rect -960 293120 3054 293176
rect 3110 293120 3115 293176
rect -960 293118 3115 293120
rect -960 293028 480 293118
rect 3049 293115 3115 293118
rect 371693 292906 371759 292909
rect 445661 292906 445727 292909
rect 369932 292904 371759 292906
rect 369932 292848 371698 292904
rect 371754 292848 371759 292904
rect 369932 292846 371759 292848
rect 441876 292904 445727 292906
rect 441876 292848 445666 292904
rect 445722 292848 445727 292904
rect 441876 292846 445727 292848
rect 371693 292843 371759 292846
rect 445661 292843 445727 292846
rect 197537 292362 197603 292365
rect 371693 292362 371759 292365
rect 197537 292360 200100 292362
rect 197537 292304 197542 292360
rect 197598 292304 200100 292360
rect 197537 292302 200100 292304
rect 369932 292360 371759 292362
rect 369932 292304 371698 292360
rect 371754 292304 371759 292360
rect 369932 292302 371759 292304
rect 197537 292299 197603 292302
rect 371693 292299 371759 292302
rect 302233 292226 302299 292229
rect 299828 292224 302299 292226
rect 299828 292168 302238 292224
rect 302294 292168 302299 292224
rect 299828 292166 302299 292168
rect 302233 292163 302299 292166
rect 371233 291818 371299 291821
rect 445661 291818 445727 291821
rect 369932 291816 371299 291818
rect 369932 291760 371238 291816
rect 371294 291760 371299 291816
rect 369932 291758 371299 291760
rect 441876 291816 445727 291818
rect 441876 291760 445666 291816
rect 445722 291760 445727 291816
rect 441876 291758 445727 291760
rect 371233 291755 371299 291758
rect 445661 291755 445727 291758
rect 372153 291274 372219 291277
rect 369932 291272 372219 291274
rect 369932 291216 372158 291272
rect 372214 291216 372219 291272
rect 369932 291214 372219 291216
rect 372153 291211 372219 291214
rect 371693 290730 371759 290733
rect 369932 290728 371759 290730
rect 369932 290672 371698 290728
rect 371754 290672 371759 290728
rect 369932 290670 371759 290672
rect 371693 290667 371759 290670
rect 445661 290594 445727 290597
rect 441876 290592 445727 290594
rect 441876 290536 445666 290592
rect 445722 290536 445727 290592
rect 441876 290534 445727 290536
rect 445661 290531 445727 290534
rect 198733 290186 198799 290189
rect 371233 290186 371299 290189
rect 198733 290184 200100 290186
rect 198733 290128 198738 290184
rect 198794 290128 200100 290184
rect 198733 290126 200100 290128
rect 369932 290184 371299 290186
rect 369932 290128 371238 290184
rect 371294 290128 371299 290184
rect 369932 290126 371299 290128
rect 198733 290123 198799 290126
rect 371233 290123 371299 290126
rect 371693 289642 371759 289645
rect 369932 289640 371759 289642
rect 369932 289584 371698 289640
rect 371754 289584 371759 289640
rect 369932 289582 371759 289584
rect 371693 289579 371759 289582
rect 445661 289506 445727 289509
rect 441876 289504 445727 289506
rect 441876 289448 445666 289504
rect 445722 289448 445727 289504
rect 441876 289446 445727 289448
rect 445661 289443 445727 289446
rect 302693 289098 302759 289101
rect 371693 289098 371759 289101
rect 299828 289096 302759 289098
rect 299828 289040 302698 289096
rect 302754 289040 302759 289096
rect 299828 289038 302759 289040
rect 369932 289096 371759 289098
rect 369932 289040 371698 289096
rect 371754 289040 371759 289096
rect 369932 289038 371759 289040
rect 302693 289035 302759 289038
rect 371693 289035 371759 289038
rect 371693 288554 371759 288557
rect 369932 288552 371759 288554
rect 369932 288496 371698 288552
rect 371754 288496 371759 288552
rect 369932 288494 371759 288496
rect 371693 288491 371759 288494
rect 445661 288282 445727 288285
rect 441876 288280 445727 288282
rect 441876 288224 445666 288280
rect 445722 288224 445727 288280
rect 441876 288222 445727 288224
rect 445661 288219 445727 288222
rect 197537 288146 197603 288149
rect 371693 288146 371759 288149
rect 197537 288144 200100 288146
rect 197537 288088 197542 288144
rect 197598 288088 200100 288144
rect 197537 288086 200100 288088
rect 369932 288144 371759 288146
rect 369932 288088 371698 288144
rect 371754 288088 371759 288144
rect 369932 288086 371759 288088
rect 197537 288083 197603 288086
rect 371693 288083 371759 288086
rect 371693 287602 371759 287605
rect 369932 287600 371759 287602
rect 369932 287544 371698 287600
rect 371754 287544 371759 287600
rect 369932 287542 371759 287544
rect 371693 287539 371759 287542
rect 445477 287194 445543 287197
rect 441876 287192 445543 287194
rect 441876 287136 445482 287192
rect 445538 287136 445543 287192
rect 441876 287134 445543 287136
rect 445477 287131 445543 287134
rect 371233 287058 371299 287061
rect 369932 287056 371299 287058
rect 369932 287000 371238 287056
rect 371294 287000 371299 287056
rect 369932 286998 371299 287000
rect 371233 286995 371299 286998
rect 371693 286514 371759 286517
rect 369932 286512 371759 286514
rect 369932 286456 371698 286512
rect 371754 286456 371759 286512
rect 369932 286454 371759 286456
rect 371693 286451 371759 286454
rect 198089 285970 198155 285973
rect 302785 285970 302851 285973
rect 371601 285970 371667 285973
rect 445661 285970 445727 285973
rect 198089 285968 200100 285970
rect 198089 285912 198094 285968
rect 198150 285912 200100 285968
rect 198089 285910 200100 285912
rect 299828 285968 302851 285970
rect 299828 285912 302790 285968
rect 302846 285912 302851 285968
rect 299828 285910 302851 285912
rect 369932 285968 371667 285970
rect 369932 285912 371606 285968
rect 371662 285912 371667 285968
rect 369932 285910 371667 285912
rect 441876 285968 445727 285970
rect 441876 285912 445666 285968
rect 445722 285912 445727 285968
rect 441876 285910 445727 285912
rect 198089 285907 198155 285910
rect 302785 285907 302851 285910
rect 371601 285907 371667 285910
rect 445661 285907 445727 285910
rect 371601 285426 371667 285429
rect 369932 285424 371667 285426
rect 369932 285368 371606 285424
rect 371662 285368 371667 285424
rect 369932 285366 371667 285368
rect 371601 285363 371667 285366
rect 583520 285276 584960 285516
rect 371601 284882 371667 284885
rect 445385 284882 445451 284885
rect 369932 284880 371667 284882
rect 369932 284824 371606 284880
rect 371662 284824 371667 284880
rect 369932 284822 371667 284824
rect 441876 284880 445451 284882
rect 441876 284824 445390 284880
rect 445446 284824 445451 284880
rect 441876 284822 445451 284824
rect 371601 284819 371667 284822
rect 445385 284819 445451 284822
rect 371693 284338 371759 284341
rect 369932 284336 371759 284338
rect 369932 284280 371698 284336
rect 371754 284280 371759 284336
rect 369932 284278 371759 284280
rect 371693 284275 371759 284278
rect 197353 283794 197419 283797
rect 371601 283794 371667 283797
rect 197353 283792 200100 283794
rect 197353 283736 197358 283792
rect 197414 283736 200100 283792
rect 197353 283734 200100 283736
rect 369932 283792 371667 283794
rect 369932 283736 371606 283792
rect 371662 283736 371667 283792
rect 369932 283734 371667 283736
rect 197353 283731 197419 283734
rect 371601 283731 371667 283734
rect 445661 283658 445727 283661
rect 441876 283656 445727 283658
rect 441876 283600 445666 283656
rect 445722 283600 445727 283656
rect 441876 283598 445727 283600
rect 445661 283595 445727 283598
rect 371693 283250 371759 283253
rect 369932 283248 371759 283250
rect 369932 283192 371698 283248
rect 371754 283192 371759 283248
rect 369932 283190 371759 283192
rect 371693 283187 371759 283190
rect 302509 282842 302575 282845
rect 299828 282840 302575 282842
rect 299828 282784 302514 282840
rect 302570 282784 302575 282840
rect 299828 282782 302575 282784
rect 302509 282779 302575 282782
rect 371601 282706 371667 282709
rect 369932 282704 371667 282706
rect 369932 282648 371606 282704
rect 371662 282648 371667 282704
rect 369932 282646 371667 282648
rect 371601 282643 371667 282646
rect 445845 282570 445911 282573
rect 441876 282568 445911 282570
rect 441876 282512 445850 282568
rect 445906 282512 445911 282568
rect 441876 282510 445911 282512
rect 445845 282507 445911 282510
rect 371601 282162 371667 282165
rect 369932 282160 371667 282162
rect 369932 282104 371606 282160
rect 371662 282104 371667 282160
rect 369932 282102 371667 282104
rect 371601 282099 371667 282102
rect 197353 281618 197419 281621
rect 371233 281618 371299 281621
rect 371969 281618 372035 281621
rect 197353 281616 200100 281618
rect 197353 281560 197358 281616
rect 197414 281560 200100 281616
rect 197353 281558 200100 281560
rect 369932 281616 372035 281618
rect 369932 281560 371238 281616
rect 371294 281560 371974 281616
rect 372030 281560 372035 281616
rect 369932 281558 372035 281560
rect 197353 281555 197419 281558
rect 371233 281555 371299 281558
rect 371969 281555 372035 281558
rect 445661 281346 445727 281349
rect 441876 281344 445727 281346
rect 441876 281288 445666 281344
rect 445722 281288 445727 281344
rect 441876 281286 445727 281288
rect 445661 281283 445727 281286
rect 371601 281074 371667 281077
rect 372153 281074 372219 281077
rect 369932 281072 372219 281074
rect 369932 281016 371606 281072
rect 371662 281016 372158 281072
rect 372214 281016 372219 281072
rect 369932 281014 372219 281016
rect 371601 281011 371667 281014
rect 372153 281011 372219 281014
rect 372102 280530 372108 280532
rect 369932 280470 372108 280530
rect 372102 280468 372108 280470
rect 372172 280468 372178 280532
rect 445017 280258 445083 280261
rect 441876 280256 445083 280258
rect -960 279972 480 280212
rect 441876 280200 445022 280256
rect 445078 280200 445083 280256
rect 441876 280198 445083 280200
rect 445017 280195 445083 280198
rect 371918 279986 371924 279988
rect 369932 279926 371924 279986
rect 371918 279924 371924 279926
rect 371988 279986 371994 279988
rect 372429 279986 372495 279989
rect 371988 279984 372495 279986
rect 371988 279928 372434 279984
rect 372490 279928 372495 279984
rect 371988 279926 372495 279928
rect 371988 279924 371994 279926
rect 372429 279923 372495 279926
rect 302785 279714 302851 279717
rect 299828 279712 302851 279714
rect 299828 279656 302790 279712
rect 302846 279656 302851 279712
rect 299828 279654 302851 279656
rect 302785 279651 302851 279654
rect 197721 279442 197787 279445
rect 371734 279442 371740 279444
rect 197721 279440 200100 279442
rect 197721 279384 197726 279440
rect 197782 279384 200100 279440
rect 197721 279382 200100 279384
rect 369932 279382 371740 279442
rect 197721 279379 197787 279382
rect 371734 279380 371740 279382
rect 371804 279442 371810 279444
rect 371969 279442 372035 279445
rect 371804 279440 372035 279442
rect 371804 279384 371974 279440
rect 372030 279384 372035 279440
rect 371804 279382 372035 279384
rect 371804 279380 371810 279382
rect 371969 279379 372035 279382
rect 369485 279034 369551 279037
rect 444649 279034 444715 279037
rect 369485 279032 369962 279034
rect 369485 278976 369490 279032
rect 369546 278976 369962 279032
rect 369485 278974 369962 278976
rect 441876 279032 444715 279034
rect 441876 278976 444654 279032
rect 444710 278976 444715 279032
rect 441876 278974 444715 278976
rect 369485 278971 369551 278974
rect 369902 278898 369962 278974
rect 444649 278971 444715 278974
rect 371366 278898 371372 278900
rect 369902 278868 371372 278898
rect 369932 278838 371372 278868
rect 371366 278836 371372 278838
rect 371436 278836 371442 278900
rect 369393 278626 369459 278629
rect 369350 278624 369459 278626
rect 369350 278568 369398 278624
rect 369454 278568 369459 278624
rect 369350 278563 369459 278568
rect 369350 278324 369410 278563
rect 372797 277946 372863 277949
rect 444465 277946 444531 277949
rect 369932 277944 372863 277946
rect 369932 277888 372802 277944
rect 372858 277888 372863 277944
rect 369932 277886 372863 277888
rect 441876 277944 444531 277946
rect 441876 277888 444470 277944
rect 444526 277888 444531 277944
rect 441876 277886 444531 277888
rect 372797 277883 372863 277886
rect 444465 277883 444531 277886
rect 197353 277402 197419 277405
rect 371693 277402 371759 277405
rect 197353 277400 200100 277402
rect 197353 277344 197358 277400
rect 197414 277344 200100 277400
rect 197353 277342 200100 277344
rect 369932 277400 371759 277402
rect 369932 277344 371698 277400
rect 371754 277344 371759 277400
rect 369932 277342 371759 277344
rect 197353 277339 197419 277342
rect 371693 277339 371759 277342
rect 370313 276858 370379 276861
rect 369932 276856 370379 276858
rect 369932 276800 370318 276856
rect 370374 276800 370379 276856
rect 369932 276798 370379 276800
rect 370313 276795 370379 276798
rect 445661 276722 445727 276725
rect 441876 276720 445727 276722
rect 441876 276664 445666 276720
rect 445722 276664 445727 276720
rect 441876 276662 445727 276664
rect 445661 276659 445727 276662
rect 302785 276586 302851 276589
rect 299828 276584 302851 276586
rect 299828 276528 302790 276584
rect 302846 276528 302851 276584
rect 299828 276526 302851 276528
rect 302785 276523 302851 276526
rect 371693 276314 371759 276317
rect 369932 276312 371759 276314
rect 369932 276256 371698 276312
rect 371754 276256 371759 276312
rect 369932 276254 371759 276256
rect 371693 276251 371759 276254
rect 369350 275365 369410 275740
rect 445661 275634 445727 275637
rect 441876 275632 445727 275634
rect 441876 275576 445666 275632
rect 445722 275576 445727 275632
rect 441876 275574 445727 275576
rect 445661 275571 445727 275574
rect 369350 275360 369459 275365
rect 369350 275304 369398 275360
rect 369454 275304 369459 275360
rect 369350 275302 369459 275304
rect 369393 275299 369459 275302
rect 198641 275226 198707 275229
rect 370405 275226 370471 275229
rect 198641 275224 200100 275226
rect 198641 275168 198646 275224
rect 198702 275168 200100 275224
rect 369932 275224 370471 275226
rect 369932 275196 370410 275224
rect 198641 275166 200100 275168
rect 369902 275168 370410 275196
rect 370466 275168 370471 275224
rect 369902 275166 370471 275168
rect 198641 275163 198707 275166
rect 369902 274818 369962 275166
rect 370405 275163 370471 275166
rect 370262 274818 370268 274820
rect 369902 274758 370268 274818
rect 370262 274756 370268 274758
rect 370332 274756 370338 274820
rect 372521 274682 372587 274685
rect 369932 274680 372587 274682
rect 369932 274624 372526 274680
rect 372582 274624 372587 274680
rect 369932 274622 372587 274624
rect 372521 274619 372587 274622
rect 445661 274410 445727 274413
rect 441876 274408 445727 274410
rect 441876 274352 445666 274408
rect 445722 274352 445727 274408
rect 441876 274350 445727 274352
rect 445661 274347 445727 274350
rect 369853 274274 369919 274277
rect 369853 274272 369962 274274
rect 369853 274216 369858 274272
rect 369914 274216 369962 274272
rect 369853 274211 369962 274216
rect 369902 274138 369962 274211
rect 370589 274138 370655 274141
rect 369902 274136 370655 274138
rect 369902 274108 370594 274136
rect 369932 274080 370594 274108
rect 370650 274080 370655 274136
rect 369932 274078 370655 274080
rect 370589 274075 370655 274078
rect 302969 273458 303035 273461
rect 299828 273456 303035 273458
rect 299828 273400 302974 273456
rect 303030 273400 303035 273456
rect 299828 273398 303035 273400
rect 302969 273395 303035 273398
rect 369902 273322 369962 273564
rect 370037 273322 370103 273325
rect 445017 273322 445083 273325
rect 369902 273320 370103 273322
rect 369902 273264 370042 273320
rect 370098 273264 370103 273320
rect 369902 273262 370103 273264
rect 441876 273320 445083 273322
rect 441876 273264 445022 273320
rect 445078 273264 445083 273320
rect 441876 273262 445083 273264
rect 370037 273259 370103 273262
rect 445017 273259 445083 273262
rect 197537 273050 197603 273053
rect 371693 273050 371759 273053
rect 371877 273050 371943 273053
rect 197537 273048 200100 273050
rect 197537 272992 197542 273048
rect 197598 272992 200100 273048
rect 197537 272990 200100 272992
rect 369932 273048 371943 273050
rect 369932 272992 371698 273048
rect 371754 272992 371882 273048
rect 371938 272992 371943 273048
rect 369932 272990 371943 272992
rect 197537 272987 197603 272990
rect 371693 272987 371759 272990
rect 371877 272987 371943 272990
rect 371417 272506 371483 272509
rect 371969 272506 372035 272509
rect 369932 272504 372035 272506
rect 369932 272448 371422 272504
rect 371478 272448 371974 272504
rect 372030 272448 372035 272504
rect 369932 272446 372035 272448
rect 371417 272443 371483 272446
rect 371969 272443 372035 272446
rect 579889 272234 579955 272237
rect 583520 272234 584960 272324
rect 579889 272232 584960 272234
rect 579889 272176 579894 272232
rect 579950 272176 584960 272232
rect 579889 272174 584960 272176
rect 579889 272171 579955 272174
rect 445661 272098 445727 272101
rect 441876 272096 445727 272098
rect 441876 272040 445666 272096
rect 445722 272040 445727 272096
rect 583520 272084 584960 272174
rect 441876 272038 445727 272040
rect 445661 272035 445727 272038
rect 372061 271962 372127 271965
rect 369932 271960 372127 271962
rect 369932 271904 372066 271960
rect 372122 271904 372127 271960
rect 369932 271902 372127 271904
rect 372061 271899 372127 271902
rect 371182 271418 371188 271420
rect 369932 271358 371188 271418
rect 371182 271356 371188 271358
rect 371252 271356 371258 271420
rect 445661 271010 445727 271013
rect 441876 271008 445727 271010
rect 441876 270952 445666 271008
rect 445722 270952 445727 271008
rect 441876 270950 445727 270952
rect 445661 270947 445727 270950
rect 197721 270874 197787 270877
rect 371509 270874 371575 270877
rect 371877 270874 371943 270877
rect 197721 270872 200100 270874
rect 197721 270816 197726 270872
rect 197782 270816 200100 270872
rect 197721 270814 200100 270816
rect 369932 270872 371943 270874
rect 369932 270816 371514 270872
rect 371570 270816 371882 270872
rect 371938 270816 371943 270872
rect 369932 270814 371943 270816
rect 197721 270811 197787 270814
rect 371509 270811 371575 270814
rect 371877 270811 371943 270814
rect 302877 270330 302943 270333
rect 371325 270330 371391 270333
rect 299828 270328 302943 270330
rect 299828 270272 302882 270328
rect 302938 270272 302943 270328
rect 299828 270270 302943 270272
rect 369932 270328 371391 270330
rect 369932 270272 371330 270328
rect 371386 270272 371391 270328
rect 369932 270270 371391 270272
rect 302877 270267 302943 270270
rect 371325 270267 371391 270270
rect 371417 270194 371483 270197
rect 372245 270194 372311 270197
rect 371417 270192 372311 270194
rect 371417 270136 371422 270192
rect 371478 270136 372250 270192
rect 372306 270136 372311 270192
rect 371417 270134 372311 270136
rect 371417 270131 371483 270134
rect 372245 270131 372311 270134
rect 371785 269786 371851 269789
rect 445385 269786 445451 269789
rect 369932 269784 371851 269786
rect 369932 269728 371790 269784
rect 371846 269728 371851 269784
rect 369932 269726 371851 269728
rect 441876 269784 445451 269786
rect 441876 269728 445390 269784
rect 445446 269728 445451 269784
rect 441876 269726 445451 269728
rect 371785 269723 371851 269726
rect 445385 269723 445451 269726
rect 371417 269242 371483 269245
rect 369932 269240 371483 269242
rect 369932 269184 371422 269240
rect 371478 269184 371483 269240
rect 369932 269182 371483 269184
rect 371417 269179 371483 269182
rect 369945 268970 370011 268973
rect 369902 268968 370011 268970
rect 369902 268912 369950 268968
rect 370006 268912 370011 268968
rect 369902 268907 370011 268912
rect 197813 268698 197879 268701
rect 197813 268696 200100 268698
rect 197813 268640 197818 268696
rect 197874 268640 200100 268696
rect 197813 268638 200100 268640
rect 197813 268635 197879 268638
rect 369902 268426 369962 268907
rect 444557 268698 444623 268701
rect 441876 268696 444623 268698
rect 441876 268640 444562 268696
rect 444618 268640 444623 268696
rect 441876 268638 444623 268640
rect 444557 268635 444623 268638
rect 370078 268426 370084 268428
rect 369902 268366 370084 268426
rect 370078 268364 370084 268366
rect 370148 268364 370154 268428
rect 370221 268290 370287 268293
rect 370681 268290 370747 268293
rect 369932 268288 370747 268290
rect 369932 268232 370226 268288
rect 370282 268232 370686 268288
rect 370742 268232 370747 268288
rect 369932 268230 370747 268232
rect 370221 268227 370287 268230
rect 370681 268227 370747 268230
rect -960 267202 480 267292
rect 3509 267202 3575 267205
rect 303245 267202 303311 267205
rect -960 267200 3575 267202
rect -960 267144 3514 267200
rect 3570 267144 3575 267200
rect -960 267142 3575 267144
rect 299828 267200 303311 267202
rect 299828 267144 303250 267200
rect 303306 267144 303311 267200
rect 299828 267142 303311 267144
rect -960 267052 480 267142
rect 3509 267139 3575 267142
rect 303245 267139 303311 267142
rect 197353 266522 197419 266525
rect 197353 266520 200100 266522
rect 197353 266464 197358 266520
rect 197414 266464 200100 266520
rect 197353 266462 200100 266464
rect 197353 266459 197419 266462
rect 353937 266250 354003 266253
rect 353937 266248 364442 266250
rect 353937 266192 353942 266248
rect 353998 266192 364442 266248
rect 353937 266190 364442 266192
rect 353937 266187 354003 266190
rect 356697 266114 356763 266117
rect 361614 266114 361620 266116
rect 356697 266112 361620 266114
rect 356697 266056 356702 266112
rect 356758 266056 361620 266112
rect 356697 266054 361620 266056
rect 356697 266051 356763 266054
rect 361614 266052 361620 266054
rect 361684 266114 361690 266116
rect 362861 266114 362927 266117
rect 364382 266116 364442 266190
rect 361684 266112 362927 266114
rect 361684 266056 362866 266112
rect 362922 266056 362927 266112
rect 361684 266054 362927 266056
rect 361684 266052 361690 266054
rect 362861 266051 362927 266054
rect 364374 266052 364380 266116
rect 364444 266114 364450 266116
rect 364885 266114 364951 266117
rect 364444 266112 364951 266114
rect 364444 266056 364890 266112
rect 364946 266056 364951 266112
rect 364444 266054 364951 266056
rect 364444 266052 364450 266054
rect 364885 266051 364951 266054
rect 197353 264482 197419 264485
rect 197353 264480 200100 264482
rect 197353 264424 197358 264480
rect 197414 264424 200100 264480
rect 197353 264422 200100 264424
rect 197353 264419 197419 264422
rect 302785 264074 302851 264077
rect 299828 264072 302851 264074
rect 299828 264016 302790 264072
rect 302846 264016 302851 264072
rect 299828 264014 302851 264016
rect 302785 264011 302851 264014
rect 197353 262306 197419 262309
rect 197353 262304 200100 262306
rect 197353 262248 197358 262304
rect 197414 262248 200100 262304
rect 197353 262246 200100 262248
rect 197353 262243 197419 262246
rect 302785 260946 302851 260949
rect 299828 260944 302851 260946
rect 299828 260888 302790 260944
rect 302846 260888 302851 260944
rect 299828 260886 302851 260888
rect 302785 260883 302851 260886
rect 197721 260130 197787 260133
rect 197721 260128 200100 260130
rect 197721 260072 197726 260128
rect 197782 260072 200100 260128
rect 197721 260070 200100 260072
rect 197721 260067 197787 260070
rect 580257 258906 580323 258909
rect 583520 258906 584960 258996
rect 580257 258904 584960 258906
rect 580257 258848 580262 258904
rect 580318 258848 584960 258904
rect 580257 258846 584960 258848
rect 580257 258843 580323 258846
rect 583520 258756 584960 258846
rect 197537 257954 197603 257957
rect 197537 257952 200100 257954
rect 197537 257896 197542 257952
rect 197598 257896 200100 257952
rect 197537 257894 200100 257896
rect 197537 257891 197603 257894
rect 302785 257818 302851 257821
rect 299828 257816 302851 257818
rect 299828 257760 302790 257816
rect 302846 257760 302851 257816
rect 299828 257758 302851 257760
rect 302785 257755 302851 257758
rect 197905 255778 197971 255781
rect 197905 255776 200100 255778
rect 197905 255720 197910 255776
rect 197966 255720 200100 255776
rect 197905 255718 200100 255720
rect 197905 255715 197971 255718
rect 302325 254690 302391 254693
rect 299828 254688 302391 254690
rect 299828 254632 302330 254688
rect 302386 254632 302391 254688
rect 299828 254630 302391 254632
rect 302325 254627 302391 254630
rect -960 254146 480 254236
rect 3141 254146 3207 254149
rect -960 254144 3207 254146
rect -960 254088 3146 254144
rect 3202 254088 3207 254144
rect -960 254086 3207 254088
rect -960 253996 480 254086
rect 3141 254083 3207 254086
rect 197537 253738 197603 253741
rect 197537 253736 200100 253738
rect 197537 253680 197542 253736
rect 197598 253680 200100 253736
rect 197537 253678 200100 253680
rect 197537 253675 197603 253678
rect 197353 251562 197419 251565
rect 302969 251562 303035 251565
rect 197353 251560 200100 251562
rect 197353 251504 197358 251560
rect 197414 251504 200100 251560
rect 197353 251502 200100 251504
rect 299828 251560 303035 251562
rect 299828 251504 302974 251560
rect 303030 251504 303035 251560
rect 299828 251502 303035 251504
rect 197353 251499 197419 251502
rect 302969 251499 303035 251502
rect 197629 249386 197695 249389
rect 197629 249384 200100 249386
rect 197629 249328 197634 249384
rect 197690 249328 200100 249384
rect 197629 249326 200100 249328
rect 197629 249323 197695 249326
rect 302785 248434 302851 248437
rect 299828 248432 302851 248434
rect 299828 248376 302790 248432
rect 302846 248376 302851 248432
rect 299828 248374 302851 248376
rect 302785 248371 302851 248374
rect 197997 247210 198063 247213
rect 197997 247208 200100 247210
rect 197997 247152 198002 247208
rect 198058 247152 200100 247208
rect 197997 247150 200100 247152
rect 197997 247147 198063 247150
rect 580165 245578 580231 245581
rect 583520 245578 584960 245668
rect 580165 245576 584960 245578
rect 580165 245520 580170 245576
rect 580226 245520 584960 245576
rect 580165 245518 584960 245520
rect 580165 245515 580231 245518
rect 583520 245428 584960 245518
rect 302877 245306 302943 245309
rect 299828 245304 302943 245306
rect 299828 245248 302882 245304
rect 302938 245248 302943 245304
rect 299828 245246 302943 245248
rect 302877 245243 302943 245246
rect 197353 245034 197419 245037
rect 197353 245032 200100 245034
rect 197353 244976 197358 245032
rect 197414 244976 200100 245032
rect 197353 244974 200100 244976
rect 197353 244971 197419 244974
rect 197905 242858 197971 242861
rect 197905 242856 200100 242858
rect 197905 242800 197910 242856
rect 197966 242800 200100 242856
rect 197905 242798 200100 242800
rect 197905 242795 197971 242798
rect 303061 242178 303127 242181
rect 299828 242176 303127 242178
rect 299828 242120 303066 242176
rect 303122 242120 303127 242176
rect 299828 242118 303127 242120
rect 303061 242115 303127 242118
rect -960 241090 480 241180
rect 3509 241090 3575 241093
rect -960 241088 3575 241090
rect -960 241032 3514 241088
rect 3570 241032 3575 241088
rect -960 241030 3575 241032
rect -960 240940 480 241030
rect 3509 241027 3575 241030
rect 197721 240818 197787 240821
rect 197721 240816 200100 240818
rect 197721 240760 197726 240816
rect 197782 240760 200100 240816
rect 197721 240758 200100 240760
rect 197721 240755 197787 240758
rect 303153 239050 303219 239053
rect 299828 239048 303219 239050
rect 299828 238992 303158 239048
rect 303214 238992 303219 239048
rect 299828 238990 303219 238992
rect 303153 238987 303219 238990
rect 197537 238642 197603 238645
rect 197537 238640 200100 238642
rect 197537 238584 197542 238640
rect 197598 238584 200100 238640
rect 197537 238582 200100 238584
rect 197537 238579 197603 238582
rect 197721 236466 197787 236469
rect 197721 236464 200100 236466
rect 197721 236408 197726 236464
rect 197782 236408 200100 236464
rect 197721 236406 200100 236408
rect 197721 236403 197787 236406
rect 302969 235922 303035 235925
rect 299828 235920 303035 235922
rect 299828 235864 302974 235920
rect 303030 235864 303035 235920
rect 299828 235862 303035 235864
rect 302969 235859 303035 235862
rect 197721 234290 197787 234293
rect 197721 234288 200100 234290
rect 197721 234232 197726 234288
rect 197782 234232 200100 234288
rect 197721 234230 200100 234232
rect 197721 234227 197787 234230
rect 303245 232794 303311 232797
rect 299828 232792 303311 232794
rect 299828 232736 303250 232792
rect 303306 232736 303311 232792
rect 299828 232734 303311 232736
rect 303245 232731 303311 232734
rect 579981 232386 580047 232389
rect 583520 232386 584960 232476
rect 579981 232384 584960 232386
rect 579981 232328 579986 232384
rect 580042 232328 584960 232384
rect 579981 232326 584960 232328
rect 579981 232323 580047 232326
rect 583520 232236 584960 232326
rect 198365 232114 198431 232117
rect 198365 232112 200100 232114
rect 198365 232056 198370 232112
rect 198426 232056 200100 232112
rect 198365 232054 200100 232056
rect 198365 232051 198431 232054
rect 197629 230074 197695 230077
rect 197629 230072 200100 230074
rect 197629 230016 197634 230072
rect 197690 230016 200100 230072
rect 197629 230014 200100 230016
rect 197629 230011 197695 230014
rect 302693 229666 302759 229669
rect 299828 229664 302759 229666
rect 299828 229608 302698 229664
rect 302754 229608 302759 229664
rect 299828 229606 302759 229608
rect 302693 229603 302759 229606
rect -960 227884 480 228124
rect 197353 227898 197419 227901
rect 197353 227896 200100 227898
rect 197353 227840 197358 227896
rect 197414 227840 200100 227896
rect 197353 227838 200100 227840
rect 197353 227835 197419 227838
rect 302693 226538 302759 226541
rect 299828 226536 302759 226538
rect 299828 226480 302698 226536
rect 302754 226480 302759 226536
rect 299828 226478 302759 226480
rect 302693 226475 302759 226478
rect 197353 225722 197419 225725
rect 372245 225722 372311 225725
rect 197353 225720 200100 225722
rect 197353 225664 197358 225720
rect 197414 225664 200100 225720
rect 197353 225662 200100 225664
rect 369932 225720 372311 225722
rect 369932 225664 372250 225720
rect 372306 225664 372311 225720
rect 369932 225662 372311 225664
rect 197353 225659 197419 225662
rect 372245 225659 372311 225662
rect 371601 225178 371667 225181
rect 369932 225176 371667 225178
rect 369932 225120 371606 225176
rect 371662 225120 371667 225176
rect 369932 225118 371667 225120
rect 371601 225115 371667 225118
rect 441846 225045 441906 225420
rect 372102 224980 372108 225044
rect 372172 225042 372178 225044
rect 372521 225042 372587 225045
rect 372172 225040 372587 225042
rect 372172 224984 372526 225040
rect 372582 224984 372587 225040
rect 372172 224982 372587 224984
rect 372172 224980 372178 224982
rect 372521 224979 372587 224982
rect 441797 225040 441906 225045
rect 441797 224984 441802 225040
rect 441858 224984 441906 225040
rect 441797 224982 441906 224984
rect 441797 224979 441863 224982
rect 371325 224634 371391 224637
rect 369932 224632 371391 224634
rect 369932 224576 371330 224632
rect 371386 224576 371391 224632
rect 369932 224574 371391 224576
rect 371325 224571 371391 224574
rect 441846 224229 441906 224332
rect 441797 224224 441906 224229
rect 441797 224168 441802 224224
rect 441858 224168 441906 224224
rect 441797 224166 441906 224168
rect 441797 224163 441863 224166
rect 371601 224090 371667 224093
rect 369932 224088 371667 224090
rect 369932 224032 371606 224088
rect 371662 224032 371667 224088
rect 369932 224030 371667 224032
rect 371601 224027 371667 224030
rect 197353 223546 197419 223549
rect 371601 223546 371667 223549
rect 197353 223544 200100 223546
rect 197353 223488 197358 223544
rect 197414 223488 200100 223544
rect 197353 223486 200100 223488
rect 369932 223544 371667 223546
rect 369932 223488 371606 223544
rect 371662 223488 371667 223544
rect 369932 223486 371667 223488
rect 197353 223483 197419 223486
rect 371601 223483 371667 223486
rect 302785 223410 302851 223413
rect 299828 223408 302851 223410
rect 299828 223352 302790 223408
rect 302846 223352 302851 223408
rect 299828 223350 302851 223352
rect 302785 223347 302851 223350
rect 444557 223138 444623 223141
rect 441876 223136 444623 223138
rect 441876 223080 444562 223136
rect 444618 223080 444623 223136
rect 441876 223078 444623 223080
rect 444557 223075 444623 223078
rect 370497 223002 370563 223005
rect 371325 223002 371391 223005
rect 369932 223000 371391 223002
rect 369932 222944 370502 223000
rect 370558 222944 371330 223000
rect 371386 222944 371391 223000
rect 369932 222942 371391 222944
rect 370497 222939 370563 222942
rect 371325 222939 371391 222942
rect 369393 222866 369459 222869
rect 369350 222864 369459 222866
rect 369350 222808 369398 222864
rect 369454 222808 369459 222864
rect 369350 222803 369459 222808
rect 369350 222458 369410 222803
rect 371233 222458 371299 222461
rect 369350 222456 371299 222458
rect 369350 222428 371238 222456
rect 369380 222400 371238 222428
rect 371294 222400 371299 222456
rect 369380 222398 371299 222400
rect 371233 222395 371299 222398
rect 445661 222050 445727 222053
rect 441876 222048 445727 222050
rect 441876 221992 445666 222048
rect 445722 221992 445727 222048
rect 441876 221990 445727 221992
rect 445661 221987 445727 221990
rect 370313 221914 370379 221917
rect 371233 221914 371299 221917
rect 369932 221912 371299 221914
rect 369932 221856 370318 221912
rect 370374 221856 371238 221912
rect 371294 221856 371299 221912
rect 369932 221854 371299 221856
rect 370313 221851 370379 221854
rect 371233 221851 371299 221854
rect 198825 221370 198891 221373
rect 370129 221370 370195 221373
rect 198825 221368 200100 221370
rect 198825 221312 198830 221368
rect 198886 221312 200100 221368
rect 198825 221310 200100 221312
rect 369932 221368 370195 221370
rect 369932 221312 370134 221368
rect 370190 221312 370195 221368
rect 369932 221310 370195 221312
rect 198825 221307 198891 221310
rect 370129 221307 370195 221310
rect 445109 220826 445175 220829
rect 441876 220824 445175 220826
rect 369902 220693 369962 220796
rect 441876 220768 445114 220824
rect 445170 220768 445175 220824
rect 441876 220766 445175 220768
rect 445109 220763 445175 220766
rect 369577 220690 369643 220693
rect 369534 220688 369643 220690
rect 369534 220632 369582 220688
rect 369638 220632 369643 220688
rect 369534 220627 369643 220632
rect 369853 220688 369962 220693
rect 369853 220632 369858 220688
rect 369914 220632 369962 220688
rect 369853 220630 369962 220632
rect 369853 220627 369919 220630
rect 302785 220282 302851 220285
rect 299828 220280 302851 220282
rect 299828 220224 302790 220280
rect 302846 220224 302851 220280
rect 369534 220282 369594 220627
rect 372797 220282 372863 220285
rect 369534 220280 372863 220282
rect 369534 220252 372802 220280
rect 299828 220222 302851 220224
rect 369564 220224 372802 220252
rect 372858 220224 372863 220280
rect 369564 220222 372863 220224
rect 302785 220219 302851 220222
rect 372797 220219 372863 220222
rect 372061 219738 372127 219741
rect 445661 219738 445727 219741
rect 369932 219736 372127 219738
rect 369932 219680 372066 219736
rect 372122 219680 372127 219736
rect 369932 219678 372127 219680
rect 441876 219736 445727 219738
rect 441876 219680 445666 219736
rect 445722 219680 445727 219736
rect 441876 219678 445727 219680
rect 372061 219675 372127 219678
rect 445661 219675 445727 219678
rect 197537 219194 197603 219197
rect 370405 219194 370471 219197
rect 197537 219192 200100 219194
rect 197537 219136 197542 219192
rect 197598 219136 200100 219192
rect 197537 219134 200100 219136
rect 369932 219192 370471 219194
rect 369932 219136 370410 219192
rect 370466 219136 370471 219192
rect 369932 219134 370471 219136
rect 197537 219131 197603 219134
rect 370405 219131 370471 219134
rect 579889 219058 579955 219061
rect 583520 219058 584960 219148
rect 579889 219056 584960 219058
rect 579889 219000 579894 219056
rect 579950 219000 584960 219056
rect 579889 218998 584960 219000
rect 579889 218995 579955 218998
rect 583520 218908 584960 218998
rect 372613 218650 372679 218653
rect 369932 218648 372679 218650
rect 369932 218592 372618 218648
rect 372674 218592 372679 218648
rect 369932 218590 372679 218592
rect 372613 218587 372679 218590
rect 369945 218514 370011 218517
rect 445661 218514 445727 218517
rect 369902 218512 370011 218514
rect 369902 218456 369950 218512
rect 370006 218456 370011 218512
rect 369902 218451 370011 218456
rect 441876 218512 445727 218514
rect 441876 218456 445666 218512
rect 445722 218456 445727 218512
rect 441876 218454 445727 218456
rect 445661 218451 445727 218454
rect 369902 218106 369962 218451
rect 371049 218106 371115 218109
rect 369902 218104 371115 218106
rect 369902 218076 371054 218104
rect 369932 218048 371054 218076
rect 371110 218048 371115 218104
rect 369932 218046 371115 218048
rect 371049 218043 371115 218046
rect 370221 217562 370287 217565
rect 369932 217560 370287 217562
rect 369932 217504 370226 217560
rect 370282 217504 370287 217560
rect 369932 217502 370287 217504
rect 370221 217499 370287 217502
rect 445661 217426 445727 217429
rect 441876 217424 445727 217426
rect 441876 217368 445666 217424
rect 445722 217368 445727 217424
rect 441876 217366 445727 217368
rect 445661 217363 445727 217366
rect 197353 217154 197419 217157
rect 302509 217154 302575 217157
rect 197353 217152 200100 217154
rect 197353 217096 197358 217152
rect 197414 217096 200100 217152
rect 197353 217094 200100 217096
rect 299828 217152 302575 217154
rect 299828 217096 302514 217152
rect 302570 217096 302575 217152
rect 299828 217094 302575 217096
rect 197353 217091 197419 217094
rect 302509 217091 302575 217094
rect 371601 217018 371667 217021
rect 369932 217016 371667 217018
rect 369932 216960 371606 217016
rect 371662 216960 371667 217016
rect 369932 216958 371667 216960
rect 371601 216955 371667 216958
rect 371325 216474 371391 216477
rect 369932 216472 371391 216474
rect 369932 216416 371330 216472
rect 371386 216416 371391 216472
rect 369932 216414 371391 216416
rect 371325 216411 371391 216414
rect 445661 216202 445727 216205
rect 441876 216200 445727 216202
rect 441876 216144 445666 216200
rect 445722 216144 445727 216200
rect 441876 216142 445727 216144
rect 445661 216139 445727 216142
rect 371601 216066 371667 216069
rect 369932 216064 371667 216066
rect 369932 216008 371606 216064
rect 371662 216008 371667 216064
rect 369932 216006 371667 216008
rect 371601 216003 371667 216006
rect 372337 215522 372403 215525
rect 369932 215520 372403 215522
rect 369932 215464 372342 215520
rect 372398 215464 372403 215520
rect 369932 215462 372403 215464
rect 372337 215459 372403 215462
rect 445661 215114 445727 215117
rect 441876 215112 445727 215114
rect -960 214978 480 215068
rect 441876 215056 445666 215112
rect 445722 215056 445727 215112
rect 441876 215054 445727 215056
rect 445661 215051 445727 215054
rect 3325 214978 3391 214981
rect -960 214976 3391 214978
rect -960 214920 3330 214976
rect 3386 214920 3391 214976
rect -960 214918 3391 214920
rect -960 214828 480 214918
rect 3325 214915 3391 214918
rect 197537 214978 197603 214981
rect 371601 214978 371667 214981
rect 197537 214976 200100 214978
rect 197537 214920 197542 214976
rect 197598 214920 200100 214976
rect 197537 214918 200100 214920
rect 369932 214976 371667 214978
rect 369932 214920 371606 214976
rect 371662 214920 371667 214976
rect 369932 214918 371667 214920
rect 197537 214915 197603 214918
rect 371601 214915 371667 214918
rect 371601 214434 371667 214437
rect 369932 214432 371667 214434
rect 369932 214376 371606 214432
rect 371662 214376 371667 214432
rect 369932 214374 371667 214376
rect 371601 214371 371667 214374
rect 302785 214026 302851 214029
rect 299828 214024 302851 214026
rect 299828 213968 302790 214024
rect 302846 213968 302851 214024
rect 299828 213966 302851 213968
rect 302785 213963 302851 213966
rect 371325 213890 371391 213893
rect 445661 213890 445727 213893
rect 369932 213888 371391 213890
rect 369932 213832 371330 213888
rect 371386 213832 371391 213888
rect 369932 213830 371391 213832
rect 441876 213888 445727 213890
rect 441876 213832 445666 213888
rect 445722 213832 445727 213888
rect 441876 213830 445727 213832
rect 371325 213827 371391 213830
rect 445661 213827 445727 213830
rect 371601 213346 371667 213349
rect 369932 213344 371667 213346
rect 369932 213288 371606 213344
rect 371662 213288 371667 213344
rect 369932 213286 371667 213288
rect 371601 213283 371667 213286
rect 197353 212802 197419 212805
rect 372061 212802 372127 212805
rect 445293 212802 445359 212805
rect 197353 212800 200100 212802
rect 197353 212744 197358 212800
rect 197414 212744 200100 212800
rect 197353 212742 200100 212744
rect 369932 212800 372127 212802
rect 369932 212744 372066 212800
rect 372122 212744 372127 212800
rect 369932 212742 372127 212744
rect 441876 212800 445359 212802
rect 441876 212744 445298 212800
rect 445354 212744 445359 212800
rect 441876 212742 445359 212744
rect 197353 212739 197419 212742
rect 372061 212739 372127 212742
rect 445293 212739 445359 212742
rect 372245 212258 372311 212261
rect 369932 212256 372311 212258
rect 369932 212200 372250 212256
rect 372306 212200 372311 212256
rect 369932 212198 372311 212200
rect 372245 212195 372311 212198
rect 370405 211714 370471 211717
rect 369932 211712 370471 211714
rect 369932 211656 370410 211712
rect 370466 211656 370471 211712
rect 369932 211654 370471 211656
rect 370405 211651 370471 211654
rect 445661 211578 445727 211581
rect 441876 211576 445727 211578
rect 441876 211520 445666 211576
rect 445722 211520 445727 211576
rect 441876 211518 445727 211520
rect 445661 211515 445727 211518
rect 371601 211170 371667 211173
rect 369932 211168 371667 211170
rect 369932 211112 371606 211168
rect 371662 211112 371667 211168
rect 369932 211110 371667 211112
rect 371601 211107 371667 211110
rect 302785 210898 302851 210901
rect 299828 210896 302851 210898
rect 299828 210840 302790 210896
rect 302846 210840 302851 210896
rect 299828 210838 302851 210840
rect 302785 210835 302851 210838
rect 197353 210626 197419 210629
rect 371601 210626 371667 210629
rect 197353 210624 200100 210626
rect 197353 210568 197358 210624
rect 197414 210568 200100 210624
rect 197353 210566 200100 210568
rect 369932 210624 371667 210626
rect 369932 210568 371606 210624
rect 371662 210568 371667 210624
rect 369932 210566 371667 210568
rect 197353 210563 197419 210566
rect 371601 210563 371667 210566
rect 444557 210490 444623 210493
rect 441876 210488 444623 210490
rect 441876 210432 444562 210488
rect 444618 210432 444623 210488
rect 441876 210430 444623 210432
rect 444557 210427 444623 210430
rect 372705 210082 372771 210085
rect 369932 210080 372771 210082
rect 369932 210024 372710 210080
rect 372766 210024 372771 210080
rect 369932 210022 372771 210024
rect 372705 210019 372771 210022
rect 370313 209538 370379 209541
rect 371233 209538 371299 209541
rect 369932 209536 371299 209538
rect 369932 209480 370318 209536
rect 370374 209480 371238 209536
rect 371294 209480 371299 209536
rect 369932 209478 371299 209480
rect 370313 209475 370379 209478
rect 371233 209475 371299 209478
rect 445661 209266 445727 209269
rect 441876 209264 445727 209266
rect 441876 209208 445666 209264
rect 445722 209208 445727 209264
rect 441876 209206 445727 209208
rect 445661 209203 445727 209206
rect 370129 208994 370195 208997
rect 371325 208994 371391 208997
rect 369932 208992 371391 208994
rect 369932 208936 370134 208992
rect 370190 208936 371330 208992
rect 371386 208936 371391 208992
rect 369932 208934 371391 208936
rect 370129 208931 370195 208934
rect 371325 208931 371391 208934
rect 369669 208722 369735 208725
rect 369669 208720 369778 208722
rect 369669 208664 369674 208720
rect 369730 208664 369778 208720
rect 369669 208659 369778 208664
rect 198181 208450 198247 208453
rect 198181 208448 200100 208450
rect 198181 208392 198186 208448
rect 198242 208392 200100 208448
rect 369718 208420 369778 208659
rect 371918 208450 371924 208452
rect 198181 208390 200100 208392
rect 371742 208390 371924 208450
rect 198181 208387 198247 208390
rect 371742 208314 371802 208390
rect 371918 208388 371924 208390
rect 371988 208450 371994 208452
rect 375741 208450 375807 208453
rect 371988 208448 375807 208450
rect 371988 208392 375746 208448
rect 375802 208392 375807 208448
rect 371988 208390 375807 208392
rect 371988 208388 371994 208390
rect 375741 208387 375807 208390
rect 369902 208254 371802 208314
rect 369902 207876 369962 208254
rect 445109 208178 445175 208181
rect 441876 208176 445175 208178
rect 441876 208120 445114 208176
rect 445170 208120 445175 208176
rect 441876 208118 445175 208120
rect 445109 208115 445175 208118
rect 302325 207770 302391 207773
rect 299828 207768 302391 207770
rect 299828 207712 302330 207768
rect 302386 207712 302391 207768
rect 299828 207710 302391 207712
rect 302325 207707 302391 207710
rect 369718 207093 369778 207332
rect 369718 207088 369827 207093
rect 369718 207032 369766 207088
rect 369822 207032 369827 207088
rect 369718 207030 369827 207032
rect 369761 207027 369827 207030
rect 444741 206954 444807 206957
rect 441876 206952 444807 206954
rect 441876 206896 444746 206952
rect 444802 206896 444807 206952
rect 441876 206894 444807 206896
rect 444741 206891 444807 206894
rect 369534 206549 369594 206788
rect 369534 206544 369643 206549
rect 369534 206488 369582 206544
rect 369638 206488 369643 206544
rect 369534 206486 369643 206488
rect 369577 206483 369643 206486
rect 197353 206410 197419 206413
rect 197353 206408 200100 206410
rect 197353 206352 197358 206408
rect 197414 206352 200100 206408
rect 197353 206350 200100 206352
rect 197353 206347 197419 206350
rect 369350 206141 369410 206244
rect 369350 206136 369459 206141
rect 369350 206080 369398 206136
rect 369454 206080 369459 206136
rect 369350 206078 369459 206080
rect 369393 206075 369459 206078
rect 371601 205866 371667 205869
rect 444465 205866 444531 205869
rect 369932 205864 371667 205866
rect 369932 205808 371606 205864
rect 371662 205808 371667 205864
rect 369932 205806 371667 205808
rect 441876 205864 444531 205866
rect 441876 205808 444470 205864
rect 444526 205808 444531 205864
rect 441876 205806 444531 205808
rect 371601 205803 371667 205806
rect 444465 205803 444531 205806
rect 583017 205730 583083 205733
rect 583520 205730 584960 205820
rect 583017 205728 584960 205730
rect 583017 205672 583022 205728
rect 583078 205672 584960 205728
rect 583017 205670 584960 205672
rect 583017 205667 583083 205670
rect 583520 205580 584960 205670
rect 371601 205322 371667 205325
rect 369932 205320 371667 205322
rect 369932 205264 371606 205320
rect 371662 205264 371667 205320
rect 369932 205262 371667 205264
rect 371601 205259 371667 205262
rect 371601 204778 371667 204781
rect 369932 204776 371667 204778
rect 369932 204720 371606 204776
rect 371662 204720 371667 204776
rect 369932 204718 371667 204720
rect 371601 204715 371667 204718
rect 302693 204642 302759 204645
rect 445293 204642 445359 204645
rect 299828 204640 302759 204642
rect 299828 204584 302698 204640
rect 302754 204584 302759 204640
rect 299828 204582 302759 204584
rect 441876 204640 445359 204642
rect 441876 204584 445298 204640
rect 445354 204584 445359 204640
rect 441876 204582 445359 204584
rect 302693 204579 302759 204582
rect 445293 204579 445359 204582
rect 198273 204234 198339 204237
rect 371601 204234 371667 204237
rect 198273 204232 200100 204234
rect 198273 204176 198278 204232
rect 198334 204176 200100 204232
rect 198273 204174 200100 204176
rect 369932 204232 371667 204234
rect 369932 204176 371606 204232
rect 371662 204176 371667 204232
rect 369932 204174 371667 204176
rect 198273 204171 198339 204174
rect 371601 204171 371667 204174
rect 369485 204098 369551 204101
rect 369485 204096 369962 204098
rect 369485 204040 369490 204096
rect 369546 204040 369962 204096
rect 369485 204038 369962 204040
rect 369485 204035 369551 204038
rect 369902 203690 369962 204038
rect 371233 203690 371299 203693
rect 369902 203688 371299 203690
rect 369902 203660 371238 203688
rect 369932 203632 371238 203660
rect 371294 203632 371299 203688
rect 369932 203630 371299 203632
rect 371233 203627 371299 203630
rect 445017 203554 445083 203557
rect 441876 203552 445083 203554
rect 441876 203496 445022 203552
rect 445078 203496 445083 203552
rect 441876 203494 445083 203496
rect 445017 203491 445083 203494
rect 370262 203146 370268 203148
rect 369932 203086 370268 203146
rect 370262 203084 370268 203086
rect 370332 203146 370338 203148
rect 370497 203146 370563 203149
rect 370332 203144 370563 203146
rect 370332 203088 370502 203144
rect 370558 203088 370563 203144
rect 370332 203086 370563 203088
rect 370332 203084 370338 203086
rect 370497 203083 370563 203086
rect 372061 202602 372127 202605
rect 369932 202600 372127 202602
rect 369932 202544 372066 202600
rect 372122 202544 372127 202600
rect 369932 202542 372127 202544
rect 372061 202539 372127 202542
rect 445661 202330 445727 202333
rect 441876 202328 445727 202330
rect 441876 202272 445666 202328
rect 445722 202272 445727 202328
rect 441876 202270 445727 202272
rect 445661 202267 445727 202270
rect 197353 202058 197419 202061
rect 370221 202058 370287 202061
rect 370589 202058 370655 202061
rect 197353 202056 200100 202058
rect -960 201922 480 202012
rect 197353 202000 197358 202056
rect 197414 202000 200100 202056
rect 197353 201998 200100 202000
rect 369932 202056 370655 202058
rect 369932 202000 370226 202056
rect 370282 202000 370594 202056
rect 370650 202000 370655 202056
rect 369932 201998 370655 202000
rect 197353 201995 197419 201998
rect 370221 201995 370287 201998
rect 370589 201995 370655 201998
rect 3049 201922 3115 201925
rect 370037 201922 370103 201925
rect -960 201920 3115 201922
rect -960 201864 3054 201920
rect 3110 201864 3115 201920
rect -960 201862 3115 201864
rect -960 201772 480 201862
rect 3049 201859 3115 201862
rect 369902 201920 370103 201922
rect 369902 201864 370042 201920
rect 370098 201864 370103 201920
rect 369902 201862 370103 201864
rect 302785 201514 302851 201517
rect 299828 201512 302851 201514
rect 299828 201456 302790 201512
rect 302846 201456 302851 201512
rect 369902 201484 369962 201862
rect 370037 201859 370103 201862
rect 299828 201454 302851 201456
rect 302785 201451 302851 201454
rect 445661 201242 445727 201245
rect 441876 201240 445727 201242
rect 441876 201184 445666 201240
rect 445722 201184 445727 201240
rect 441876 201182 445727 201184
rect 445661 201179 445727 201182
rect 371693 200970 371759 200973
rect 369932 200968 371759 200970
rect 369932 200912 371698 200968
rect 371754 200912 371759 200968
rect 369932 200910 371759 200912
rect 371693 200907 371759 200910
rect 371969 200426 372035 200429
rect 369932 200424 372035 200426
rect 369932 200368 371974 200424
rect 372030 200368 372035 200424
rect 369932 200366 372035 200368
rect 371969 200363 372035 200366
rect 445661 200018 445727 200021
rect 441876 200016 445727 200018
rect 441876 199960 445666 200016
rect 445722 199960 445727 200016
rect 441876 199958 445727 199960
rect 445661 199955 445727 199958
rect 198089 199882 198155 199885
rect 372153 199882 372219 199885
rect 198089 199880 200100 199882
rect 198089 199824 198094 199880
rect 198150 199824 200100 199880
rect 198089 199822 200100 199824
rect 369932 199880 372219 199882
rect 369932 199824 372158 199880
rect 372214 199824 372219 199880
rect 369932 199822 372219 199824
rect 198089 199819 198155 199822
rect 372153 199819 372219 199822
rect 371366 199338 371372 199340
rect 369932 199278 371372 199338
rect 371366 199276 371372 199278
rect 371436 199338 371442 199340
rect 372061 199338 372127 199341
rect 371436 199336 372127 199338
rect 371436 199280 372066 199336
rect 372122 199280 372127 199336
rect 371436 199278 372127 199280
rect 371436 199276 371442 199278
rect 372061 199275 372127 199278
rect 371601 198930 371667 198933
rect 372153 198930 372219 198933
rect 445661 198930 445727 198933
rect 371601 198928 372219 198930
rect 371601 198872 371606 198928
rect 371662 198872 372158 198928
rect 372214 198872 372219 198928
rect 371601 198870 372219 198872
rect 441876 198928 445727 198930
rect 441876 198872 445666 198928
rect 445722 198872 445727 198928
rect 441876 198870 445727 198872
rect 371601 198867 371667 198870
rect 372153 198867 372219 198870
rect 445661 198867 445727 198870
rect 371233 198794 371299 198797
rect 371877 198794 371943 198797
rect 369932 198792 371943 198794
rect 369932 198736 371238 198792
rect 371294 198736 371882 198792
rect 371938 198736 371943 198792
rect 369932 198734 371943 198736
rect 371233 198731 371299 198734
rect 371877 198731 371943 198734
rect 302785 198386 302851 198389
rect 299828 198384 302851 198386
rect 299828 198328 302790 198384
rect 302846 198328 302851 198384
rect 299828 198326 302851 198328
rect 302785 198323 302851 198326
rect 371509 198250 371575 198253
rect 369932 198248 371575 198250
rect 369932 198192 371514 198248
rect 371570 198192 371575 198248
rect 369932 198190 371575 198192
rect 371509 198187 371575 198190
rect 197353 197706 197419 197709
rect 371785 197706 371851 197709
rect 445385 197706 445451 197709
rect 197353 197704 200100 197706
rect 197353 197648 197358 197704
rect 197414 197648 200100 197704
rect 197353 197646 200100 197648
rect 369932 197704 371851 197706
rect 369932 197648 371790 197704
rect 371846 197648 371851 197704
rect 369932 197646 371851 197648
rect 441876 197704 445451 197706
rect 441876 197648 445390 197704
rect 445446 197648 445451 197704
rect 441876 197646 445451 197648
rect 197353 197643 197419 197646
rect 371785 197643 371851 197646
rect 445385 197643 445451 197646
rect 371325 197162 371391 197165
rect 369932 197160 371391 197162
rect 369932 197104 371330 197160
rect 371386 197104 371391 197160
rect 369932 197102 371391 197104
rect 371325 197099 371391 197102
rect 370078 196618 370084 196620
rect 369932 196558 370084 196618
rect 370078 196556 370084 196558
rect 370148 196618 370154 196620
rect 371233 196618 371299 196621
rect 445845 196618 445911 196621
rect 370148 196616 371299 196618
rect 370148 196560 371238 196616
rect 371294 196560 371299 196616
rect 370148 196558 371299 196560
rect 441876 196616 445911 196618
rect 441876 196560 445850 196616
rect 445906 196560 445911 196616
rect 441876 196558 445911 196560
rect 370148 196556 370154 196558
rect 371233 196555 371299 196558
rect 445845 196555 445911 196558
rect 370681 196210 370747 196213
rect 369932 196208 370747 196210
rect 369932 196152 370686 196208
rect 370742 196152 370747 196208
rect 369932 196150 370747 196152
rect 370681 196147 370747 196150
rect 364374 196012 364380 196076
rect 364444 196074 364450 196076
rect 364517 196074 364583 196077
rect 364444 196072 364583 196074
rect 364444 196016 364522 196072
rect 364578 196016 364583 196072
rect 364444 196014 364583 196016
rect 364444 196012 364450 196014
rect 364517 196011 364583 196014
rect 197629 195530 197695 195533
rect 197629 195528 200100 195530
rect 197629 195472 197634 195528
rect 197690 195472 200100 195528
rect 197629 195470 200100 195472
rect 197629 195467 197695 195470
rect 302325 195258 302391 195261
rect 299828 195256 302391 195258
rect 299828 195200 302330 195256
rect 302386 195200 302391 195256
rect 299828 195198 302391 195200
rect 302325 195195 302391 195198
rect 361614 194516 361620 194580
rect 361684 194578 361690 194580
rect 362718 194578 362724 194580
rect 361684 194518 362724 194578
rect 361684 194516 361690 194518
rect 362718 194516 362724 194518
rect 362788 194578 362794 194580
rect 362861 194578 362927 194581
rect 362788 194576 362927 194578
rect 362788 194520 362866 194576
rect 362922 194520 362927 194576
rect 362788 194518 362927 194520
rect 362788 194516 362794 194518
rect 362861 194515 362927 194518
rect 364885 194578 364951 194581
rect 365294 194578 365300 194580
rect 364885 194576 365300 194578
rect 364885 194520 364890 194576
rect 364946 194520 365300 194576
rect 364885 194518 365300 194520
rect 364885 194515 364951 194518
rect 365294 194516 365300 194518
rect 365364 194516 365370 194580
rect 197353 193490 197419 193493
rect 197353 193488 200100 193490
rect 197353 193432 197358 193488
rect 197414 193432 200100 193488
rect 197353 193430 200100 193432
rect 197353 193427 197419 193430
rect 580257 192538 580323 192541
rect 583520 192538 584960 192628
rect 580257 192536 584960 192538
rect 580257 192480 580262 192536
rect 580318 192480 584960 192536
rect 580257 192478 584960 192480
rect 580257 192475 580323 192478
rect 583520 192388 584960 192478
rect 302785 192130 302851 192133
rect 299828 192128 302851 192130
rect 299828 192072 302790 192128
rect 302846 192072 302851 192128
rect 299828 192070 302851 192072
rect 302785 192067 302851 192070
rect 198365 191314 198431 191317
rect 198365 191312 200100 191314
rect 198365 191256 198370 191312
rect 198426 191256 200100 191312
rect 198365 191254 200100 191256
rect 198365 191251 198431 191254
rect 172421 189954 172487 189957
rect 169894 189952 172487 189954
rect 169894 189896 172426 189952
rect 172482 189896 172487 189952
rect 169894 189894 172487 189896
rect 169894 189448 169954 189894
rect 172421 189891 172487 189894
rect 197353 189138 197419 189141
rect 197353 189136 200100 189138
rect 197353 189080 197358 189136
rect 197414 189080 200100 189136
rect 197353 189078 200100 189080
rect 197353 189075 197419 189078
rect 302785 189002 302851 189005
rect 299828 189000 302851 189002
rect -960 188866 480 188956
rect 299828 188944 302790 189000
rect 302846 188944 302851 189000
rect 299828 188942 302851 188944
rect 302785 188939 302851 188942
rect 3509 188866 3575 188869
rect -960 188864 3575 188866
rect -960 188808 3514 188864
rect 3570 188808 3575 188864
rect -960 188806 3575 188808
rect -960 188716 480 188806
rect 3509 188803 3575 188806
rect 172053 188730 172119 188733
rect 169894 188728 172119 188730
rect 169894 188672 172058 188728
rect 172114 188672 172119 188728
rect 169894 188670 172119 188672
rect 169894 188360 169954 188670
rect 172053 188667 172119 188670
rect 172145 187642 172211 187645
rect 169894 187640 172211 187642
rect 169894 187584 172150 187640
rect 172206 187584 172211 187640
rect 169894 187582 172211 187584
rect 169894 187136 169954 187582
rect 172145 187579 172211 187582
rect 197353 186962 197419 186965
rect 197353 186960 200100 186962
rect 197353 186904 197358 186960
rect 197414 186904 200100 186960
rect 197353 186902 200100 186904
rect 197353 186899 197419 186902
rect 169661 186282 169727 186285
rect 169661 186280 169770 186282
rect 169661 186224 169666 186280
rect 169722 186224 169770 186280
rect 169661 186219 169770 186224
rect 169710 186048 169770 186219
rect 302693 185874 302759 185877
rect 299828 185872 302759 185874
rect 299828 185816 302698 185872
rect 302754 185816 302759 185872
rect 299828 185814 302759 185816
rect 302693 185811 302759 185814
rect 172421 184922 172487 184925
rect 169894 184920 172487 184922
rect 169894 184864 172426 184920
rect 172482 184864 172487 184920
rect 169894 184862 172487 184864
rect 169894 184824 169954 184862
rect 172421 184859 172487 184862
rect 197353 184786 197419 184789
rect 197353 184784 200100 184786
rect 197353 184728 197358 184784
rect 197414 184728 200100 184784
rect 197353 184726 200100 184728
rect 197353 184723 197419 184726
rect 171685 184242 171751 184245
rect 169894 184240 171751 184242
rect 169894 184184 171690 184240
rect 171746 184184 171751 184240
rect 169894 184182 171751 184184
rect 169894 183736 169954 184182
rect 171685 184179 171751 184182
rect 172421 183018 172487 183021
rect 169894 183016 172487 183018
rect 169894 182960 172426 183016
rect 172482 182960 172487 183016
rect 169894 182958 172487 182960
rect 169894 182512 169954 182958
rect 172421 182955 172487 182958
rect 198089 182746 198155 182749
rect 302969 182746 303035 182749
rect 198089 182744 200100 182746
rect 198089 182688 198094 182744
rect 198150 182688 200100 182744
rect 198089 182686 200100 182688
rect 299828 182744 303035 182746
rect 299828 182688 302974 182744
rect 303030 182688 303035 182744
rect 299828 182686 303035 182688
rect 198089 182683 198155 182686
rect 302969 182683 303035 182686
rect 172053 181794 172119 181797
rect 169894 181792 172119 181794
rect 169894 181736 172058 181792
rect 172114 181736 172119 181792
rect 169894 181734 172119 181736
rect 169894 181424 169954 181734
rect 172053 181731 172119 181734
rect 172421 180570 172487 180573
rect 169894 180568 172487 180570
rect 169894 180512 172426 180568
rect 172482 180512 172487 180568
rect 169894 180510 172487 180512
rect 169894 180200 169954 180510
rect 172421 180507 172487 180510
rect 198365 180570 198431 180573
rect 198365 180568 200100 180570
rect 198365 180512 198370 180568
rect 198426 180512 200100 180568
rect 198365 180510 200100 180512
rect 198365 180507 198431 180510
rect 302785 179618 302851 179621
rect 299828 179616 302851 179618
rect 299828 179560 302790 179616
rect 302846 179560 302851 179616
rect 299828 179558 302851 179560
rect 302785 179555 302851 179558
rect 172421 179210 172487 179213
rect 169894 179208 172487 179210
rect 169894 179152 172426 179208
rect 172482 179152 172487 179208
rect 169894 179150 172487 179152
rect 169894 179112 169954 179150
rect 172421 179147 172487 179150
rect 580165 179210 580231 179213
rect 583520 179210 584960 179300
rect 580165 179208 584960 179210
rect 580165 179152 580170 179208
rect 580226 179152 584960 179208
rect 580165 179150 584960 179152
rect 580165 179147 580231 179150
rect 583520 179060 584960 179150
rect 197353 178394 197419 178397
rect 197353 178392 200100 178394
rect 197353 178336 197358 178392
rect 197414 178336 200100 178392
rect 197353 178334 200100 178336
rect 197353 178331 197419 178334
rect 172421 177986 172487 177989
rect 169894 177984 172487 177986
rect 169894 177928 172426 177984
rect 172482 177928 172487 177984
rect 169894 177926 172487 177928
rect 169894 177888 169954 177926
rect 172421 177923 172487 177926
rect 172329 177442 172395 177445
rect 169894 177440 172395 177442
rect 169894 177384 172334 177440
rect 172390 177384 172395 177440
rect 169894 177382 172395 177384
rect 169894 176800 169954 177382
rect 172329 177379 172395 177382
rect 302785 176490 302851 176493
rect 299828 176488 302851 176490
rect 299828 176432 302790 176488
rect 302846 176432 302851 176488
rect 299828 176430 302851 176432
rect 302785 176427 302851 176430
rect 197629 176218 197695 176221
rect 197629 176216 200100 176218
rect 197629 176160 197634 176216
rect 197690 176160 200100 176216
rect 197629 176158 200100 176160
rect 197629 176155 197695 176158
rect 172237 176082 172303 176085
rect 169894 176080 172303 176082
rect -960 175796 480 176036
rect 169894 176024 172242 176080
rect 172298 176024 172303 176080
rect 169894 176022 172303 176024
rect 169894 175576 169954 176022
rect 172237 176019 172303 176022
rect 172421 174858 172487 174861
rect 169894 174856 172487 174858
rect 169894 174800 172426 174856
rect 172482 174800 172487 174856
rect 169894 174798 172487 174800
rect 169894 174488 169954 174798
rect 172421 174795 172487 174798
rect 197353 174042 197419 174045
rect 197353 174040 200100 174042
rect 197353 173984 197358 174040
rect 197414 173984 200100 174040
rect 197353 173982 200100 173984
rect 197353 173979 197419 173982
rect 172421 173634 172487 173637
rect 169894 173632 172487 173634
rect 169894 173576 172426 173632
rect 172482 173576 172487 173632
rect 169894 173574 172487 173576
rect 169894 173264 169954 173574
rect 172421 173571 172487 173574
rect 302877 173362 302943 173365
rect 299828 173360 302943 173362
rect 299828 173304 302882 173360
rect 302938 173304 302943 173360
rect 299828 173302 302943 173304
rect 302877 173299 302943 173302
rect 172421 172410 172487 172413
rect 169894 172408 172487 172410
rect 169894 172352 172426 172408
rect 172482 172352 172487 172408
rect 169894 172350 172487 172352
rect 169894 172176 169954 172350
rect 172421 172347 172487 172350
rect 198181 171866 198247 171869
rect 198181 171864 200100 171866
rect 198181 171808 198186 171864
rect 198242 171808 200100 171864
rect 198181 171806 200100 171808
rect 198181 171803 198247 171806
rect 171777 171050 171843 171053
rect 169894 171048 171843 171050
rect 169894 170992 171782 171048
rect 171838 170992 171843 171048
rect 169894 170990 171843 170992
rect 169894 170952 169954 170990
rect 171777 170987 171843 170990
rect 172237 170506 172303 170509
rect 169894 170504 172303 170506
rect 169894 170448 172242 170504
rect 172298 170448 172303 170504
rect 169894 170446 172303 170448
rect 169894 169864 169954 170446
rect 172237 170443 172303 170446
rect 302785 170234 302851 170237
rect 299828 170232 302851 170234
rect 299828 170176 302790 170232
rect 302846 170176 302851 170232
rect 299828 170174 302851 170176
rect 302785 170171 302851 170174
rect 197721 169826 197787 169829
rect 197721 169824 200100 169826
rect 197721 169768 197726 169824
rect 197782 169768 200100 169824
rect 197721 169766 200100 169768
rect 197721 169763 197787 169766
rect 171869 169282 171935 169285
rect 169894 169280 171935 169282
rect 169894 169224 171874 169280
rect 171930 169224 171935 169280
rect 169894 169222 171935 169224
rect 169894 168640 169954 169222
rect 171869 169219 171935 169222
rect 172421 167922 172487 167925
rect 169894 167920 172487 167922
rect 169894 167864 172426 167920
rect 172482 167864 172487 167920
rect 169894 167862 172487 167864
rect 169894 167552 169954 167862
rect 172421 167859 172487 167862
rect 197537 167650 197603 167653
rect 197537 167648 200100 167650
rect 197537 167592 197542 167648
rect 197598 167592 200100 167648
rect 197537 167590 200100 167592
rect 197537 167587 197603 167590
rect 303061 167106 303127 167109
rect 299828 167104 303127 167106
rect 299828 167048 303066 167104
rect 303122 167048 303127 167104
rect 299828 167046 303127 167048
rect 303061 167043 303127 167046
rect 171961 166970 172027 166973
rect 169894 166968 172027 166970
rect 169894 166912 171966 166968
rect 172022 166912 172027 166968
rect 169894 166910 172027 166912
rect 169894 166328 169954 166910
rect 171961 166907 172027 166910
rect 582925 165882 582991 165885
rect 583520 165882 584960 165972
rect 582925 165880 584960 165882
rect 582925 165824 582930 165880
rect 582986 165824 584960 165880
rect 582925 165822 584960 165824
rect 582925 165819 582991 165822
rect 583520 165732 584960 165822
rect 198089 165474 198155 165477
rect 198089 165472 200100 165474
rect 198089 165416 198094 165472
rect 198150 165416 200100 165472
rect 198089 165414 200100 165416
rect 198089 165411 198155 165414
rect 169894 165202 169954 165240
rect 172053 165202 172119 165205
rect 169894 165200 172119 165202
rect 169894 165144 172058 165200
rect 172114 165144 172119 165200
rect 169894 165142 172119 165144
rect 172053 165139 172119 165142
rect 172421 164114 172487 164117
rect 169894 164112 172487 164114
rect 169894 164056 172426 164112
rect 172482 164056 172487 164112
rect 169894 164054 172487 164056
rect 169894 164016 169954 164054
rect 172421 164051 172487 164054
rect 302877 163978 302943 163981
rect 299828 163976 302943 163978
rect 299828 163920 302882 163976
rect 302938 163920 302943 163976
rect 299828 163918 302943 163920
rect 302877 163915 302943 163918
rect 172237 163570 172303 163573
rect 169894 163568 172303 163570
rect 169894 163512 172242 163568
rect 172298 163512 172303 163568
rect 169894 163510 172303 163512
rect -960 162890 480 162980
rect 169894 162928 169954 163510
rect 172237 163507 172303 163510
rect 197997 163298 198063 163301
rect 197997 163296 200100 163298
rect 197997 163240 198002 163296
rect 198058 163240 200100 163296
rect 197997 163238 200100 163240
rect 197997 163235 198063 163238
rect 3233 162890 3299 162893
rect -960 162888 3299 162890
rect -960 162832 3238 162888
rect 3294 162832 3299 162888
rect -960 162830 3299 162832
rect -960 162740 480 162830
rect 3233 162827 3299 162830
rect 172145 162346 172211 162349
rect 169894 162344 172211 162346
rect 169894 162288 172150 162344
rect 172206 162288 172211 162344
rect 169894 162286 172211 162288
rect 169894 161704 169954 162286
rect 172145 162283 172211 162286
rect 197537 161122 197603 161125
rect 197537 161120 200100 161122
rect 197537 161064 197542 161120
rect 197598 161064 200100 161120
rect 197537 161062 200100 161064
rect 197537 161059 197603 161062
rect 172421 160986 172487 160989
rect 169894 160984 172487 160986
rect 169894 160928 172426 160984
rect 172482 160928 172487 160984
rect 169894 160926 172487 160928
rect 169894 160616 169954 160926
rect 172421 160923 172487 160926
rect 302509 160850 302575 160853
rect 299828 160848 302575 160850
rect 299828 160792 302514 160848
rect 302570 160792 302575 160848
rect 299828 160790 302575 160792
rect 302509 160787 302575 160790
rect 371734 159292 371740 159356
rect 371804 159354 371810 159356
rect 372061 159354 372127 159357
rect 454217 159354 454283 159357
rect 371804 159352 454283 159354
rect 371804 159296 372066 159352
rect 372122 159296 454222 159352
rect 454278 159296 454283 159352
rect 371804 159294 454283 159296
rect 371804 159292 371810 159294
rect 372061 159291 372127 159294
rect 454217 159291 454283 159294
rect 197353 159082 197419 159085
rect 197353 159080 200100 159082
rect 197353 159024 197358 159080
rect 197414 159024 200100 159080
rect 197353 159022 200100 159024
rect 197353 159019 197419 159022
rect 302785 157722 302851 157725
rect 299828 157720 302851 157722
rect 299828 157664 302790 157720
rect 302846 157664 302851 157720
rect 299828 157662 302851 157664
rect 302785 157659 302851 157662
rect 197813 156906 197879 156909
rect 197813 156904 200100 156906
rect 197813 156848 197818 156904
rect 197874 156848 200100 156904
rect 197813 156846 200100 156848
rect 197813 156843 197879 156846
rect 197353 154730 197419 154733
rect 197353 154728 200100 154730
rect 197353 154672 197358 154728
rect 197414 154672 200100 154728
rect 197353 154670 200100 154672
rect 197353 154667 197419 154670
rect 302601 154594 302667 154597
rect 299828 154592 302667 154594
rect 299828 154536 302606 154592
rect 302662 154536 302667 154592
rect 299828 154534 302667 154536
rect 302601 154531 302667 154534
rect 171593 153778 171659 153781
rect 371417 153778 371483 153781
rect 169924 153776 171659 153778
rect 169924 153720 171598 153776
rect 171654 153720 171659 153776
rect 169924 153718 171659 153720
rect 369932 153776 371483 153778
rect 369932 153720 371422 153776
rect 371478 153720 371483 153776
rect 369932 153718 371483 153720
rect 171593 153715 171659 153718
rect 371417 153715 371483 153718
rect 444925 153506 444991 153509
rect 441876 153504 444991 153506
rect 441876 153448 444930 153504
rect 444986 153448 444991 153504
rect 441876 153446 444991 153448
rect 444925 153443 444991 153446
rect 171685 153234 171751 153237
rect 371969 153234 372035 153237
rect 169924 153232 171751 153234
rect 169924 153176 171690 153232
rect 171746 153176 171751 153232
rect 169924 153174 171751 153176
rect 369932 153232 372035 153234
rect 369932 153176 371974 153232
rect 372030 153176 372035 153232
rect 369932 153174 372035 153176
rect 171685 153171 171751 153174
rect 371969 153171 372035 153174
rect 370078 153036 370084 153100
rect 370148 153098 370154 153100
rect 373257 153098 373323 153101
rect 370148 153096 373323 153098
rect 370148 153040 373262 153096
rect 373318 153040 373323 153096
rect 370148 153038 373323 153040
rect 370148 153036 370154 153038
rect 369301 152962 369367 152965
rect 370086 152962 370146 153036
rect 373257 153035 373323 153038
rect 369301 152960 370146 152962
rect 369301 152904 369306 152960
rect 369362 152904 370146 152960
rect 369301 152902 370146 152904
rect 369301 152899 369367 152902
rect 171593 152690 171659 152693
rect 371417 152690 371483 152693
rect 169924 152688 171659 152690
rect 169924 152632 171598 152688
rect 171654 152632 171659 152688
rect 169924 152630 171659 152632
rect 369932 152688 371483 152690
rect 369932 152632 371422 152688
rect 371478 152632 371483 152688
rect 369932 152630 371483 152632
rect 171593 152627 171659 152630
rect 371417 152627 371483 152630
rect 579613 152690 579679 152693
rect 583520 152690 584960 152780
rect 579613 152688 584960 152690
rect 579613 152632 579618 152688
rect 579674 152632 584960 152688
rect 579613 152630 584960 152632
rect 579613 152627 579679 152630
rect 197353 152554 197419 152557
rect 197353 152552 200100 152554
rect 197353 152496 197358 152552
rect 197414 152496 200100 152552
rect 583520 152540 584960 152630
rect 197353 152494 200100 152496
rect 197353 152491 197419 152494
rect 445661 152418 445727 152421
rect 441876 152416 445727 152418
rect 441876 152360 445666 152416
rect 445722 152360 445727 152416
rect 441876 152358 445727 152360
rect 445661 152355 445727 152358
rect 170489 152146 170555 152149
rect 371877 152146 371943 152149
rect 169924 152144 170555 152146
rect 169924 152088 170494 152144
rect 170550 152088 170555 152144
rect 169924 152086 170555 152088
rect 369932 152144 371943 152146
rect 369932 152088 371882 152144
rect 371938 152088 371943 152144
rect 369932 152086 371943 152088
rect 170489 152083 170555 152086
rect 371877 152083 371943 152086
rect 172421 151602 172487 151605
rect 371417 151602 371483 151605
rect 169924 151600 172487 151602
rect 169924 151544 172426 151600
rect 172482 151544 172487 151600
rect 169924 151542 172487 151544
rect 369932 151600 371483 151602
rect 369932 151544 371422 151600
rect 371478 151544 371483 151600
rect 369932 151542 371483 151544
rect 172421 151539 172487 151542
rect 371417 151539 371483 151542
rect 302693 151466 302759 151469
rect 299828 151464 302759 151466
rect 299828 151408 302698 151464
rect 302754 151408 302759 151464
rect 299828 151406 302759 151408
rect 302693 151403 302759 151406
rect 444925 151194 444991 151197
rect 441876 151192 444991 151194
rect 441876 151136 444930 151192
rect 444986 151136 444991 151192
rect 441876 151134 444991 151136
rect 444925 151131 444991 151134
rect 172237 151058 172303 151061
rect 371969 151058 372035 151061
rect 169924 151056 172303 151058
rect 169924 151000 172242 151056
rect 172298 151000 172303 151056
rect 169924 150998 172303 151000
rect 369932 151056 372035 151058
rect 369932 151000 371974 151056
rect 372030 151000 372035 151056
rect 369932 150998 372035 151000
rect 172237 150995 172303 150998
rect 371969 150995 372035 150998
rect 171685 150514 171751 150517
rect 371417 150514 371483 150517
rect 169924 150512 171751 150514
rect 169924 150456 171690 150512
rect 171746 150456 171751 150512
rect 169924 150454 171751 150456
rect 369932 150512 371483 150514
rect 369932 150456 371422 150512
rect 371478 150456 371483 150512
rect 369932 150454 371483 150456
rect 171685 150451 171751 150454
rect 371417 150451 371483 150454
rect 197353 150378 197419 150381
rect 197353 150376 200100 150378
rect 197353 150320 197358 150376
rect 197414 150320 200100 150376
rect 197353 150318 200100 150320
rect 197353 150315 197419 150318
rect 444925 150106 444991 150109
rect 441876 150104 444991 150106
rect 441876 150048 444930 150104
rect 444986 150048 444991 150104
rect 441876 150046 444991 150048
rect 444925 150043 444991 150046
rect 172421 149970 172487 149973
rect 371417 149970 371483 149973
rect 169924 149968 172487 149970
rect -960 149834 480 149924
rect 169924 149912 172426 149968
rect 172482 149912 172487 149968
rect 169924 149910 172487 149912
rect 369932 149968 371483 149970
rect 369932 149912 371422 149968
rect 371478 149912 371483 149968
rect 369932 149910 371483 149912
rect 172421 149907 172487 149910
rect 371417 149907 371483 149910
rect 3509 149834 3575 149837
rect -960 149832 3575 149834
rect -960 149776 3514 149832
rect 3570 149776 3575 149832
rect -960 149774 3575 149776
rect -960 149684 480 149774
rect 3509 149771 3575 149774
rect 171501 149426 171567 149429
rect 371969 149426 372035 149429
rect 169924 149424 171567 149426
rect 169924 149368 171506 149424
rect 171562 149368 171567 149424
rect 169924 149366 171567 149368
rect 369932 149424 372035 149426
rect 369932 149368 371974 149424
rect 372030 149368 372035 149424
rect 369932 149366 372035 149368
rect 171501 149363 171567 149366
rect 371969 149363 372035 149366
rect 441797 149018 441863 149021
rect 441797 149016 441906 149018
rect 441797 148960 441802 149016
rect 441858 148960 441906 149016
rect 441797 148955 441906 148960
rect 172421 148882 172487 148885
rect 371417 148882 371483 148885
rect 169924 148880 172487 148882
rect 169924 148824 172426 148880
rect 172482 148824 172487 148880
rect 169924 148822 172487 148824
rect 369932 148880 371483 148882
rect 369932 148824 371422 148880
rect 371478 148824 371483 148880
rect 441846 148852 441906 148955
rect 369932 148822 371483 148824
rect 172421 148819 172487 148822
rect 371417 148819 371483 148822
rect 171685 148338 171751 148341
rect 302325 148338 302391 148341
rect 372521 148338 372587 148341
rect 169924 148336 171751 148338
rect 169924 148280 171690 148336
rect 171746 148280 171751 148336
rect 169924 148278 171751 148280
rect 299828 148336 302391 148338
rect 299828 148280 302330 148336
rect 302386 148280 302391 148336
rect 299828 148278 302391 148280
rect 369932 148336 372587 148338
rect 369932 148280 372526 148336
rect 372582 148280 372587 148336
rect 369932 148278 372587 148280
rect 171685 148275 171751 148278
rect 302325 148275 302391 148278
rect 372521 148275 372587 148278
rect 197353 148202 197419 148205
rect 197353 148200 200100 148202
rect 197353 148144 197358 148200
rect 197414 148144 200100 148200
rect 197353 148142 200100 148144
rect 197353 148139 197419 148142
rect 171501 147794 171567 147797
rect 371969 147794 372035 147797
rect 444373 147794 444439 147797
rect 169924 147792 171567 147794
rect 169924 147736 171506 147792
rect 171562 147736 171567 147792
rect 169924 147734 171567 147736
rect 369932 147792 372035 147794
rect 369932 147736 371974 147792
rect 372030 147736 372035 147792
rect 369932 147734 372035 147736
rect 441876 147792 444439 147794
rect 441876 147736 444378 147792
rect 444434 147736 444439 147792
rect 441876 147734 444439 147736
rect 171501 147731 171567 147734
rect 371969 147731 372035 147734
rect 444373 147731 444439 147734
rect 171685 147250 171751 147253
rect 371417 147250 371483 147253
rect 169924 147248 171751 147250
rect 169924 147192 171690 147248
rect 171746 147192 171751 147248
rect 169924 147190 171751 147192
rect 369932 147248 371483 147250
rect 369932 147192 371422 147248
rect 371478 147192 371483 147248
rect 369932 147190 371483 147192
rect 171685 147187 171751 147190
rect 371417 147187 371483 147190
rect 172329 146706 172395 146709
rect 371969 146706 372035 146709
rect 169924 146704 172395 146706
rect 169924 146648 172334 146704
rect 172390 146648 172395 146704
rect 169924 146646 172395 146648
rect 369932 146704 372035 146706
rect 369932 146648 371974 146704
rect 372030 146648 372035 146704
rect 369932 146646 372035 146648
rect 172329 146643 172395 146646
rect 371969 146643 372035 146646
rect 444373 146570 444439 146573
rect 441876 146568 444439 146570
rect 441876 146512 444378 146568
rect 444434 146512 444439 146568
rect 441876 146510 444439 146512
rect 444373 146507 444439 146510
rect 172421 146162 172487 146165
rect 169924 146160 172487 146162
rect 169924 146104 172426 146160
rect 172482 146104 172487 146160
rect 169924 146102 172487 146104
rect 172421 146099 172487 146102
rect 198089 146162 198155 146165
rect 371417 146162 371483 146165
rect 198089 146160 200100 146162
rect 198089 146104 198094 146160
rect 198150 146104 200100 146160
rect 198089 146102 200100 146104
rect 369932 146160 371483 146162
rect 369932 146104 371422 146160
rect 371478 146104 371483 146160
rect 369932 146102 371483 146104
rect 198089 146099 198155 146102
rect 371417 146099 371483 146102
rect 172421 145618 172487 145621
rect 371969 145618 372035 145621
rect 169924 145616 172487 145618
rect 169924 145560 172426 145616
rect 172482 145560 172487 145616
rect 169924 145558 172487 145560
rect 369932 145616 372035 145618
rect 369932 145560 371974 145616
rect 372030 145560 372035 145616
rect 369932 145558 372035 145560
rect 172421 145555 172487 145558
rect 371969 145555 372035 145558
rect 445661 145482 445727 145485
rect 441876 145480 445727 145482
rect 441876 145424 445666 145480
rect 445722 145424 445727 145480
rect 441876 145422 445727 145424
rect 445661 145419 445727 145422
rect 302785 145210 302851 145213
rect 299828 145208 302851 145210
rect 299828 145152 302790 145208
rect 302846 145152 302851 145208
rect 299828 145150 302851 145152
rect 302785 145147 302851 145150
rect 171685 145074 171751 145077
rect 371417 145074 371483 145077
rect 169924 145072 171751 145074
rect 169924 145016 171690 145072
rect 171746 145016 171751 145072
rect 169924 145014 171751 145016
rect 369932 145072 371483 145074
rect 369932 145016 371422 145072
rect 371478 145016 371483 145072
rect 369932 145014 371483 145016
rect 171685 145011 171751 145014
rect 371417 145011 371483 145014
rect 171685 144530 171751 144533
rect 371417 144530 371483 144533
rect 169924 144528 171751 144530
rect 169924 144472 171690 144528
rect 171746 144472 171751 144528
rect 169924 144470 171751 144472
rect 369932 144528 371483 144530
rect 369932 144472 371422 144528
rect 371478 144472 371483 144528
rect 369932 144470 371483 144472
rect 171685 144467 171751 144470
rect 371417 144467 371483 144470
rect 445293 144258 445359 144261
rect 441876 144256 445359 144258
rect 441876 144200 445298 144256
rect 445354 144200 445359 144256
rect 441876 144198 445359 144200
rect 445293 144195 445359 144198
rect 171777 144122 171843 144125
rect 371417 144122 371483 144125
rect 169924 144120 171843 144122
rect 169924 144064 171782 144120
rect 171838 144064 171843 144120
rect 169924 144062 171843 144064
rect 369932 144120 371483 144122
rect 369932 144064 371422 144120
rect 371478 144064 371483 144120
rect 369932 144062 371483 144064
rect 171777 144059 171843 144062
rect 371417 144059 371483 144062
rect 197353 143986 197419 143989
rect 197353 143984 200100 143986
rect 197353 143928 197358 143984
rect 197414 143928 200100 143984
rect 197353 143926 200100 143928
rect 197353 143923 197419 143926
rect 171961 143578 172027 143581
rect 371417 143578 371483 143581
rect 169924 143576 172027 143578
rect 169924 143520 171966 143576
rect 172022 143520 172027 143576
rect 169924 143518 172027 143520
rect 369932 143576 371483 143578
rect 369932 143520 371422 143576
rect 371478 143520 371483 143576
rect 369932 143518 371483 143520
rect 171961 143515 172027 143518
rect 371417 143515 371483 143518
rect 445201 143170 445267 143173
rect 441876 143168 445267 143170
rect 441876 143112 445206 143168
rect 445262 143112 445267 143168
rect 441876 143110 445267 143112
rect 445201 143107 445267 143110
rect 171869 143034 171935 143037
rect 371969 143034 372035 143037
rect 169924 143032 171935 143034
rect 169924 142976 171874 143032
rect 171930 142976 171935 143032
rect 169924 142974 171935 142976
rect 369932 143032 372035 143034
rect 369932 142976 371974 143032
rect 372030 142976 372035 143032
rect 369932 142974 372035 142976
rect 171869 142971 171935 142974
rect 371969 142971 372035 142974
rect 172421 142490 172487 142493
rect 371417 142490 371483 142493
rect 169924 142488 172487 142490
rect 169924 142432 172426 142488
rect 172482 142432 172487 142488
rect 169924 142430 172487 142432
rect 369932 142488 371483 142490
rect 369932 142432 371422 142488
rect 371478 142432 371483 142488
rect 369932 142430 371483 142432
rect 172421 142427 172487 142430
rect 371417 142427 371483 142430
rect 302785 142082 302851 142085
rect 299828 142080 302851 142082
rect 299828 142024 302790 142080
rect 302846 142024 302851 142080
rect 299828 142022 302851 142024
rect 302785 142019 302851 142022
rect 172421 141946 172487 141949
rect 371417 141946 371483 141949
rect 445109 141946 445175 141949
rect 169924 141944 172487 141946
rect 169924 141888 172426 141944
rect 172482 141888 172487 141944
rect 169924 141886 172487 141888
rect 369932 141944 371483 141946
rect 369932 141888 371422 141944
rect 371478 141888 371483 141944
rect 369932 141886 371483 141888
rect 441876 141944 445175 141946
rect 441876 141888 445114 141944
rect 445170 141888 445175 141944
rect 441876 141886 445175 141888
rect 172421 141883 172487 141886
rect 371417 141883 371483 141886
rect 445109 141883 445175 141886
rect 197537 141810 197603 141813
rect 197537 141808 200100 141810
rect 197537 141752 197542 141808
rect 197598 141752 200100 141808
rect 197537 141750 200100 141752
rect 197537 141747 197603 141750
rect 171869 141402 171935 141405
rect 371969 141402 372035 141405
rect 169924 141400 171935 141402
rect 169924 141344 171874 141400
rect 171930 141344 171935 141400
rect 169924 141342 171935 141344
rect 369932 141400 372035 141402
rect 369932 141344 371974 141400
rect 372030 141344 372035 141400
rect 369932 141342 372035 141344
rect 171869 141339 171935 141342
rect 371969 141339 372035 141342
rect 172329 140858 172395 140861
rect 372061 140858 372127 140861
rect 444557 140858 444623 140861
rect 169924 140856 172395 140858
rect 169924 140800 172334 140856
rect 172390 140800 172395 140856
rect 169924 140798 172395 140800
rect 369932 140856 372127 140858
rect 369932 140800 372066 140856
rect 372122 140800 372127 140856
rect 369932 140798 372127 140800
rect 441876 140856 444623 140858
rect 441876 140800 444562 140856
rect 444618 140800 444623 140856
rect 441876 140798 444623 140800
rect 172329 140795 172395 140798
rect 372061 140795 372127 140798
rect 444557 140795 444623 140798
rect 172145 140314 172211 140317
rect 371969 140314 372035 140317
rect 169924 140312 172211 140314
rect 169924 140256 172150 140312
rect 172206 140256 172211 140312
rect 169924 140254 172211 140256
rect 369932 140312 372035 140314
rect 369932 140256 371974 140312
rect 372030 140256 372035 140312
rect 369932 140254 372035 140256
rect 172145 140251 172211 140254
rect 371969 140251 372035 140254
rect 172421 139770 172487 139773
rect 371417 139770 371483 139773
rect 169924 139768 172487 139770
rect 169924 139712 172426 139768
rect 172482 139712 172487 139768
rect 169924 139710 172487 139712
rect 369932 139768 371483 139770
rect 369932 139712 371422 139768
rect 371478 139712 371483 139768
rect 369932 139710 371483 139712
rect 172421 139707 172487 139710
rect 371417 139707 371483 139710
rect 197721 139634 197787 139637
rect 445109 139634 445175 139637
rect 197721 139632 200100 139634
rect 197721 139576 197726 139632
rect 197782 139576 200100 139632
rect 197721 139574 200100 139576
rect 441876 139632 445175 139634
rect 441876 139576 445114 139632
rect 445170 139576 445175 139632
rect 441876 139574 445175 139576
rect 197721 139571 197787 139574
rect 445109 139571 445175 139574
rect 580165 139362 580231 139365
rect 583520 139362 584960 139452
rect 580165 139360 584960 139362
rect 580165 139304 580170 139360
rect 580226 139304 584960 139360
rect 580165 139302 584960 139304
rect 580165 139299 580231 139302
rect 172237 139226 172303 139229
rect 371417 139226 371483 139229
rect 169924 139224 172303 139226
rect 169924 139168 172242 139224
rect 172298 139168 172303 139224
rect 169924 139166 172303 139168
rect 369932 139224 371483 139226
rect 369932 139168 371422 139224
rect 371478 139168 371483 139224
rect 583520 139212 584960 139302
rect 369932 139166 371483 139168
rect 172237 139163 172303 139166
rect 371417 139163 371483 139166
rect 302693 138954 302759 138957
rect 299828 138952 302759 138954
rect 299828 138896 302698 138952
rect 302754 138896 302759 138952
rect 299828 138894 302759 138896
rect 302693 138891 302759 138894
rect 172421 138682 172487 138685
rect 371417 138682 371483 138685
rect 169924 138680 172487 138682
rect 169924 138624 172426 138680
rect 172482 138624 172487 138680
rect 169924 138622 172487 138624
rect 369932 138680 371483 138682
rect 369932 138624 371422 138680
rect 371478 138624 371483 138680
rect 369932 138622 371483 138624
rect 172421 138619 172487 138622
rect 371417 138619 371483 138622
rect 445937 138546 446003 138549
rect 441876 138544 446003 138546
rect 441876 138488 445942 138544
rect 445998 138488 446003 138544
rect 441876 138486 446003 138488
rect 445937 138483 446003 138486
rect 172329 138138 172395 138141
rect 371969 138138 372035 138141
rect 169924 138136 172395 138138
rect 169924 138080 172334 138136
rect 172390 138080 172395 138136
rect 169924 138078 172395 138080
rect 369932 138136 372035 138138
rect 369932 138080 371974 138136
rect 372030 138080 372035 138136
rect 369932 138078 372035 138080
rect 172329 138075 172395 138078
rect 371969 138075 372035 138078
rect 172053 137594 172119 137597
rect 370313 137594 370379 137597
rect 169924 137592 172119 137594
rect 169924 137536 172058 137592
rect 172114 137536 172119 137592
rect 169924 137534 172119 137536
rect 369932 137592 370379 137594
rect 369932 137536 370318 137592
rect 370374 137536 370379 137592
rect 369932 137534 370379 137536
rect 172053 137531 172119 137534
rect 370313 137531 370379 137534
rect 197353 137458 197419 137461
rect 197353 137456 200100 137458
rect 197353 137400 197358 137456
rect 197414 137400 200100 137456
rect 197353 137398 200100 137400
rect 197353 137395 197419 137398
rect 444833 137322 444899 137325
rect 441876 137320 444899 137322
rect 441876 137264 444838 137320
rect 444894 137264 444899 137320
rect 441876 137262 444899 137264
rect 444833 137259 444899 137262
rect 171685 137050 171751 137053
rect 370773 137050 370839 137053
rect 169924 137048 171751 137050
rect 169924 136992 171690 137048
rect 171746 136992 171751 137048
rect 169924 136990 171751 136992
rect 369932 137048 370839 137050
rect 369932 136992 370778 137048
rect 370834 136992 370839 137048
rect 369932 136990 370839 136992
rect 171685 136987 171751 136990
rect 370773 136987 370839 136990
rect -960 136778 480 136868
rect 3417 136778 3483 136781
rect -960 136776 3483 136778
rect -960 136720 3422 136776
rect 3478 136720 3483 136776
rect -960 136718 3483 136720
rect -960 136628 480 136718
rect 3417 136715 3483 136718
rect 369485 136642 369551 136645
rect 369485 136640 369594 136642
rect 369485 136584 369490 136640
rect 369546 136584 369594 136640
rect 369485 136579 369594 136584
rect 172421 136506 172487 136509
rect 169924 136504 172487 136506
rect 169924 136448 172426 136504
rect 172482 136448 172487 136504
rect 369534 136476 369594 136579
rect 169924 136446 172487 136448
rect 172421 136443 172487 136446
rect 444373 136234 444439 136237
rect 441876 136232 444439 136234
rect 441876 136176 444378 136232
rect 444434 136176 444439 136232
rect 441876 136174 444439 136176
rect 444373 136171 444439 136174
rect 172237 135962 172303 135965
rect 370405 135962 370471 135965
rect 169924 135960 172303 135962
rect 169924 135904 172242 135960
rect 172298 135904 172303 135960
rect 169924 135902 172303 135904
rect 369932 135960 370471 135962
rect 369932 135904 370410 135960
rect 370466 135904 370471 135960
rect 369932 135902 370471 135904
rect 172237 135899 172303 135902
rect 370405 135899 370471 135902
rect 302877 135826 302943 135829
rect 299828 135824 302943 135826
rect 299828 135768 302882 135824
rect 302938 135768 302943 135824
rect 299828 135766 302943 135768
rect 302877 135763 302943 135766
rect 171317 135418 171383 135421
rect 169924 135416 171383 135418
rect 169924 135360 171322 135416
rect 171378 135360 171383 135416
rect 169924 135358 171383 135360
rect 171317 135355 171383 135358
rect 197353 135418 197419 135421
rect 370221 135418 370287 135421
rect 197353 135416 200100 135418
rect 197353 135360 197358 135416
rect 197414 135360 200100 135416
rect 197353 135358 200100 135360
rect 369932 135416 370287 135418
rect 369932 135360 370226 135416
rect 370282 135360 370287 135416
rect 369932 135358 370287 135360
rect 197353 135355 197419 135358
rect 370221 135355 370287 135358
rect 444741 135010 444807 135013
rect 441876 135008 444807 135010
rect 441876 134952 444746 135008
rect 444802 134952 444807 135008
rect 441876 134950 444807 134952
rect 444741 134947 444807 134950
rect 171869 134874 171935 134877
rect 370865 134874 370931 134877
rect 169924 134872 171935 134874
rect 169924 134816 171874 134872
rect 171930 134816 171935 134872
rect 169924 134814 171935 134816
rect 369932 134872 370931 134874
rect 369932 134816 370870 134872
rect 370926 134816 370931 134872
rect 369932 134814 370931 134816
rect 171869 134811 171935 134814
rect 370865 134811 370931 134814
rect 369945 134602 370011 134605
rect 369902 134600 370011 134602
rect 369902 134544 369950 134600
rect 370006 134544 370011 134600
rect 369902 134539 370011 134544
rect 171685 134330 171751 134333
rect 169924 134328 171751 134330
rect 169924 134272 171690 134328
rect 171746 134272 171751 134328
rect 369902 134300 369962 134539
rect 169924 134270 171751 134272
rect 171685 134267 171751 134270
rect 369894 133996 369900 134060
rect 369964 133996 369970 134060
rect 172421 133922 172487 133925
rect 169924 133920 172487 133922
rect 169924 133864 172426 133920
rect 172482 133864 172487 133920
rect 369902 133892 369962 133996
rect 444465 133922 444531 133925
rect 441876 133920 444531 133922
rect 169924 133862 172487 133864
rect 441876 133864 444470 133920
rect 444526 133864 444531 133920
rect 441876 133862 444531 133864
rect 172421 133859 172487 133862
rect 444465 133859 444531 133862
rect 369853 133650 369919 133653
rect 369853 133648 369962 133650
rect 369853 133592 369858 133648
rect 369914 133592 369962 133648
rect 369853 133587 369962 133592
rect 172053 133378 172119 133381
rect 169924 133376 172119 133378
rect 169924 133320 172058 133376
rect 172114 133320 172119 133376
rect 369902 133348 369962 133587
rect 169924 133318 172119 133320
rect 172053 133315 172119 133318
rect 197353 133242 197419 133245
rect 197353 133240 200100 133242
rect 197353 133184 197358 133240
rect 197414 133184 200100 133240
rect 197353 133182 200100 133184
rect 197353 133179 197419 133182
rect 172421 132834 172487 132837
rect 370129 132834 370195 132837
rect 169924 132832 172487 132834
rect 169924 132776 172426 132832
rect 172482 132776 172487 132832
rect 169924 132774 172487 132776
rect 369932 132832 370195 132834
rect 369932 132776 370134 132832
rect 370190 132776 370195 132832
rect 369932 132774 370195 132776
rect 172421 132771 172487 132774
rect 370129 132771 370195 132774
rect 302969 132698 303035 132701
rect 444465 132698 444531 132701
rect 299828 132696 303035 132698
rect 299828 132640 302974 132696
rect 303030 132640 303035 132696
rect 299828 132638 303035 132640
rect 441876 132696 444531 132698
rect 441876 132640 444470 132696
rect 444526 132640 444531 132696
rect 441876 132638 444531 132640
rect 302969 132635 303035 132638
rect 444465 132635 444531 132638
rect 369393 132426 369459 132429
rect 369350 132424 369459 132426
rect 369350 132368 369398 132424
rect 369454 132368 369459 132424
rect 369350 132363 369459 132368
rect 171133 132290 171199 132293
rect 169924 132288 171199 132290
rect 169924 132232 171138 132288
rect 171194 132232 171199 132288
rect 369350 132260 369410 132363
rect 169924 132230 171199 132232
rect 171133 132227 171199 132230
rect 369301 132018 369367 132021
rect 369301 132016 369410 132018
rect 369301 131960 369306 132016
rect 369362 131960 369410 132016
rect 369301 131955 369410 131960
rect 172421 131746 172487 131749
rect 169924 131744 172487 131746
rect 169924 131688 172426 131744
rect 172482 131688 172487 131744
rect 369350 131716 369410 131955
rect 169924 131686 172487 131688
rect 172421 131683 172487 131686
rect 445661 131610 445727 131613
rect 441876 131608 445727 131610
rect 441876 131552 445666 131608
rect 445722 131552 445727 131608
rect 441876 131550 445727 131552
rect 445661 131547 445727 131550
rect 369577 131474 369643 131477
rect 369534 131472 369643 131474
rect 369534 131416 369582 131472
rect 369638 131416 369643 131472
rect 369534 131411 369643 131416
rect 171501 131202 171567 131205
rect 169924 131200 171567 131202
rect 169924 131144 171506 131200
rect 171562 131144 171567 131200
rect 369534 131172 369594 131411
rect 169924 131142 171567 131144
rect 171501 131139 171567 131142
rect 197353 131066 197419 131069
rect 197353 131064 200100 131066
rect 197353 131008 197358 131064
rect 197414 131008 200100 131064
rect 197353 131006 200100 131008
rect 197353 131003 197419 131006
rect 369301 130930 369367 130933
rect 369301 130928 369410 130930
rect 369301 130872 369306 130928
rect 369362 130872 369410 130928
rect 369301 130867 369410 130872
rect 171869 130658 171935 130661
rect 169924 130656 171935 130658
rect 169924 130600 171874 130656
rect 171930 130600 171935 130656
rect 369350 130628 369410 130867
rect 169924 130598 171935 130600
rect 171869 130595 171935 130598
rect 444833 130386 444899 130389
rect 441876 130384 444899 130386
rect 441876 130356 444838 130384
rect 441846 130328 444838 130356
rect 444894 130328 444899 130384
rect 441846 130326 444899 130328
rect 172421 130114 172487 130117
rect 370497 130114 370563 130117
rect 169924 130112 172487 130114
rect 169924 130056 172426 130112
rect 172482 130056 172487 130112
rect 369932 130112 370563 130114
rect 369932 130084 370502 130112
rect 169924 130054 172487 130056
rect 172421 130051 172487 130054
rect 369902 130056 370502 130084
rect 370558 130056 370563 130112
rect 369902 130054 370563 130056
rect 369902 129845 369962 130054
rect 370497 130051 370563 130054
rect 441846 129845 441906 130326
rect 444833 130323 444899 130326
rect 369902 129840 370011 129845
rect 369902 129784 369950 129840
rect 370006 129784 370011 129840
rect 369902 129782 370011 129784
rect 369945 129779 370011 129782
rect 441797 129840 441906 129845
rect 441797 129784 441802 129840
rect 441858 129784 441906 129840
rect 441797 129782 441906 129784
rect 441797 129779 441863 129782
rect 171869 129570 171935 129573
rect 302601 129570 302667 129573
rect 169924 129568 171935 129570
rect 169924 129512 171874 129568
rect 171930 129512 171935 129568
rect 169924 129510 171935 129512
rect 299828 129568 302667 129570
rect 299828 129512 302606 129568
rect 302662 129512 302667 129568
rect 299828 129510 302667 129512
rect 171869 129507 171935 129510
rect 302601 129507 302667 129510
rect 369902 129165 369962 129540
rect 442993 129298 443059 129301
rect 444833 129298 444899 129301
rect 441876 129296 444899 129298
rect 441876 129240 442998 129296
rect 443054 129240 444838 129296
rect 444894 129240 444899 129296
rect 441876 129238 444899 129240
rect 442993 129235 443059 129238
rect 444833 129235 444899 129238
rect 369853 129160 369962 129165
rect 369853 129104 369858 129160
rect 369914 129104 369962 129160
rect 369853 129102 369962 129104
rect 369853 129099 369919 129102
rect 171501 129026 171567 129029
rect 370221 129026 370287 129029
rect 169924 129024 171567 129026
rect 169924 128968 171506 129024
rect 171562 128968 171567 129024
rect 169924 128966 171567 128968
rect 369932 129024 370287 129026
rect 369932 128968 370226 129024
rect 370282 128968 370287 129024
rect 369932 128966 370287 128968
rect 171501 128963 171567 128966
rect 370221 128963 370287 128966
rect 197353 128890 197419 128893
rect 197353 128888 200100 128890
rect 197353 128832 197358 128888
rect 197414 128832 200100 128888
rect 197353 128830 200100 128832
rect 197353 128827 197419 128830
rect 370037 128618 370103 128621
rect 371877 128618 371943 128621
rect 369902 128616 371943 128618
rect 369902 128560 370042 128616
rect 370098 128560 371882 128616
rect 371938 128560 371943 128616
rect 369902 128558 371943 128560
rect 171777 128482 171843 128485
rect 169924 128480 171843 128482
rect 169924 128424 171782 128480
rect 171838 128424 171843 128480
rect 369902 128452 369962 128558
rect 370037 128555 370103 128558
rect 371877 128555 371943 128558
rect 169924 128422 171843 128424
rect 171777 128419 171843 128422
rect 443637 128074 443703 128077
rect 441876 128072 443703 128074
rect 441876 128016 443642 128072
rect 443698 128016 443703 128072
rect 441876 128014 443703 128016
rect 443637 128011 443703 128014
rect 171685 127938 171751 127941
rect 371601 127938 371667 127941
rect 169924 127936 171751 127938
rect 169924 127880 171690 127936
rect 171746 127880 171751 127936
rect 169924 127878 171751 127880
rect 369932 127936 371667 127938
rect 369932 127880 371606 127936
rect 371662 127880 371667 127936
rect 369932 127878 371667 127880
rect 171685 127875 171751 127878
rect 371601 127875 371667 127878
rect 172421 127394 172487 127397
rect 370313 127394 370379 127397
rect 371734 127394 371740 127396
rect 169924 127392 172487 127394
rect 169924 127336 172426 127392
rect 172482 127336 172487 127392
rect 169924 127334 172487 127336
rect 369932 127392 371740 127394
rect 369932 127336 370318 127392
rect 370374 127336 371740 127392
rect 369932 127334 371740 127336
rect 172421 127331 172487 127334
rect 370313 127331 370379 127334
rect 371734 127332 371740 127334
rect 371804 127332 371810 127396
rect 445661 126986 445727 126989
rect 441876 126984 445727 126986
rect 441876 126956 445666 126984
rect 441846 126928 445666 126956
rect 445722 126928 445727 126984
rect 441846 126926 445727 126928
rect 172053 126850 172119 126853
rect 169924 126848 172119 126850
rect 169924 126792 172058 126848
rect 172114 126792 172119 126848
rect 169924 126790 172119 126792
rect 172053 126787 172119 126790
rect 198457 126714 198523 126717
rect 198457 126712 200100 126714
rect 198457 126656 198462 126712
rect 198518 126656 200100 126712
rect 198457 126654 200100 126656
rect 198457 126651 198523 126654
rect 369350 126445 369410 126820
rect 441846 126445 441906 126926
rect 445661 126923 445727 126926
rect 302785 126442 302851 126445
rect 299828 126440 302851 126442
rect 299828 126384 302790 126440
rect 302846 126384 302851 126440
rect 299828 126382 302851 126384
rect 369350 126442 369459 126445
rect 371233 126442 371299 126445
rect 369350 126440 371299 126442
rect 369350 126384 369398 126440
rect 369454 126384 371238 126440
rect 371294 126384 371299 126440
rect 369350 126382 371299 126384
rect 441846 126440 441955 126445
rect 441846 126384 441894 126440
rect 441950 126384 441955 126440
rect 441846 126382 441955 126384
rect 302785 126379 302851 126382
rect 369393 126379 369459 126382
rect 371233 126379 371299 126382
rect 441889 126379 441955 126382
rect 172329 126306 172395 126309
rect 370405 126306 370471 126309
rect 371509 126306 371575 126309
rect 169924 126304 172395 126306
rect 169924 126248 172334 126304
rect 172390 126248 172395 126304
rect 169924 126246 172395 126248
rect 369932 126304 371575 126306
rect 369932 126248 370410 126304
rect 370466 126248 371514 126304
rect 371570 126248 371575 126304
rect 369932 126246 371575 126248
rect 172329 126243 172395 126246
rect 370405 126243 370471 126246
rect 371509 126243 371575 126246
rect 582833 126034 582899 126037
rect 583520 126034 584960 126124
rect 582833 126032 584960 126034
rect 582833 125976 582838 126032
rect 582894 125976 584960 126032
rect 582833 125974 584960 125976
rect 582833 125971 582899 125974
rect 583520 125884 584960 125974
rect 172421 125762 172487 125765
rect 370129 125762 370195 125765
rect 371785 125762 371851 125765
rect 443269 125762 443335 125765
rect 169924 125760 172487 125762
rect 169924 125704 172426 125760
rect 172482 125704 172487 125760
rect 169924 125702 172487 125704
rect 369932 125760 371851 125762
rect 369932 125704 370134 125760
rect 370190 125704 371790 125760
rect 371846 125704 371851 125760
rect 441876 125760 443335 125762
rect 441876 125732 443274 125760
rect 369932 125702 371851 125704
rect 172421 125699 172487 125702
rect 370129 125699 370195 125702
rect 371785 125699 371851 125702
rect 441846 125704 443274 125732
rect 443330 125704 443335 125760
rect 441846 125702 443335 125704
rect 441846 125493 441906 125702
rect 443269 125699 443335 125702
rect 441797 125488 441906 125493
rect 441797 125432 441802 125488
rect 441858 125432 441906 125488
rect 441797 125430 441906 125432
rect 441797 125427 441863 125430
rect 172421 125218 172487 125221
rect 371325 125218 371391 125221
rect 372521 125218 372587 125221
rect 169924 125216 172487 125218
rect 169924 125160 172426 125216
rect 172482 125160 172487 125216
rect 369380 125216 372587 125218
rect 369380 125188 371330 125216
rect 169924 125158 172487 125160
rect 172421 125155 172487 125158
rect 369350 125160 371330 125188
rect 371386 125160 372526 125216
rect 372582 125160 372587 125216
rect 369350 125158 372587 125160
rect 369350 124949 369410 125158
rect 371325 125155 371391 125158
rect 372521 125155 372587 125158
rect 369301 124944 369410 124949
rect 369301 124888 369306 124944
rect 369362 124888 369410 124944
rect 369301 124886 369410 124888
rect 441797 124946 441863 124949
rect 441797 124944 441906 124946
rect 441797 124888 441802 124944
rect 441858 124888 441906 124944
rect 369301 124883 369367 124886
rect 441797 124883 441906 124888
rect 171317 124674 171383 124677
rect 370221 124674 370287 124677
rect 371233 124674 371299 124677
rect 169924 124672 171383 124674
rect 169924 124616 171322 124672
rect 171378 124616 171383 124672
rect 169924 124614 171383 124616
rect 369932 124672 371299 124674
rect 369932 124616 370226 124672
rect 370282 124616 371238 124672
rect 371294 124616 371299 124672
rect 441846 124644 441906 124883
rect 369932 124614 371299 124616
rect 171317 124611 171383 124614
rect 370221 124611 370287 124614
rect 371233 124611 371299 124614
rect 197537 124538 197603 124541
rect 197537 124536 200100 124538
rect 197537 124480 197542 124536
rect 197598 124480 200100 124536
rect 197537 124478 200100 124480
rect 197537 124475 197603 124478
rect 369853 124402 369919 124405
rect 369853 124400 369962 124402
rect 369853 124344 369858 124400
rect 369914 124344 369962 124400
rect 369853 124339 369962 124344
rect 171961 124266 172027 124269
rect 169924 124264 172027 124266
rect 169924 124208 171966 124264
rect 172022 124208 172027 124264
rect 369902 124266 369962 124339
rect 370681 124266 370747 124269
rect 372429 124266 372495 124269
rect 369902 124264 372495 124266
rect 369902 124236 370686 124264
rect 169924 124206 172027 124208
rect 369932 124208 370686 124236
rect 370742 124208 372434 124264
rect 372490 124208 372495 124264
rect 369932 124206 372495 124208
rect 171961 124203 172027 124206
rect 370681 124203 370747 124206
rect 372429 124203 372495 124206
rect 362769 123996 362835 123997
rect 362718 123932 362724 123996
rect 362788 123994 362835 123996
rect 365161 123994 365227 123997
rect 365294 123994 365300 123996
rect 362788 123992 362880 123994
rect 362830 123936 362880 123992
rect 362788 123934 362880 123936
rect 365161 123992 365300 123994
rect 365161 123936 365166 123992
rect 365222 123936 365300 123992
rect 365161 123934 365300 123936
rect 362788 123932 362835 123934
rect 362769 123931 362835 123932
rect 365161 123931 365227 123934
rect 365294 123932 365300 123934
rect 365364 123932 365370 123996
rect -960 123572 480 123812
rect 302785 123314 302851 123317
rect 299828 123312 302851 123314
rect 299828 123256 302790 123312
rect 302846 123256 302851 123312
rect 299828 123254 302851 123256
rect 302785 123251 302851 123254
rect 197997 122498 198063 122501
rect 197997 122496 200100 122498
rect 197997 122440 198002 122496
rect 198058 122440 200100 122496
rect 197997 122438 200100 122440
rect 197997 122435 198063 122438
rect 197537 120322 197603 120325
rect 197537 120320 200100 120322
rect 197537 120264 197542 120320
rect 197598 120264 200100 120320
rect 197537 120262 200100 120264
rect 197537 120259 197603 120262
rect 302509 120186 302575 120189
rect 299828 120184 302575 120186
rect 299828 120128 302514 120184
rect 302570 120128 302575 120184
rect 299828 120126 302575 120128
rect 302509 120123 302575 120126
rect 197905 118146 197971 118149
rect 197905 118144 200100 118146
rect 197905 118088 197910 118144
rect 197966 118088 200100 118144
rect 197905 118086 200100 118088
rect 197905 118083 197971 118086
rect 302785 117058 302851 117061
rect 299828 117056 302851 117058
rect 299828 117000 302790 117056
rect 302846 117000 302851 117056
rect 299828 116998 302851 117000
rect 302785 116995 302851 116998
rect 198365 115970 198431 115973
rect 198365 115968 200100 115970
rect 198365 115912 198370 115968
rect 198426 115912 200100 115968
rect 198365 115910 200100 115912
rect 198365 115907 198431 115910
rect 302969 113930 303035 113933
rect 299828 113928 303035 113930
rect 299828 113872 302974 113928
rect 303030 113872 303035 113928
rect 299828 113870 303035 113872
rect 302969 113867 303035 113870
rect 197353 113794 197419 113797
rect 197353 113792 200100 113794
rect 197353 113736 197358 113792
rect 197414 113736 200100 113792
rect 197353 113734 200100 113736
rect 197353 113731 197419 113734
rect 579797 112842 579863 112845
rect 583520 112842 584960 112932
rect 579797 112840 584960 112842
rect 579797 112784 579802 112840
rect 579858 112784 584960 112840
rect 579797 112782 584960 112784
rect 579797 112779 579863 112782
rect 583520 112692 584960 112782
rect 197353 111754 197419 111757
rect 197353 111752 200100 111754
rect 197353 111696 197358 111752
rect 197414 111696 200100 111752
rect 197353 111694 200100 111696
rect 197353 111691 197419 111694
rect 302785 110802 302851 110805
rect 299828 110800 302851 110802
rect -960 110666 480 110756
rect 299828 110744 302790 110800
rect 302846 110744 302851 110800
rect 299828 110742 302851 110744
rect 302785 110739 302851 110742
rect 3417 110666 3483 110669
rect -960 110664 3483 110666
rect -960 110608 3422 110664
rect 3478 110608 3483 110664
rect -960 110606 3483 110608
rect -960 110516 480 110606
rect 3417 110603 3483 110606
rect 197353 109578 197419 109581
rect 197353 109576 200100 109578
rect 197353 109520 197358 109576
rect 197414 109520 200100 109576
rect 197353 109518 200100 109520
rect 197353 109515 197419 109518
rect 302785 107674 302851 107677
rect 299828 107672 302851 107674
rect 299828 107616 302790 107672
rect 302846 107616 302851 107672
rect 299828 107614 302851 107616
rect 302785 107611 302851 107614
rect 198549 107402 198615 107405
rect 198549 107400 200100 107402
rect 198549 107344 198554 107400
rect 198610 107344 200100 107400
rect 198549 107342 200100 107344
rect 198549 107339 198615 107342
rect 197537 105226 197603 105229
rect 197537 105224 200100 105226
rect 197537 105168 197542 105224
rect 197598 105168 200100 105224
rect 197537 105166 200100 105168
rect 197537 105163 197603 105166
rect 302877 104546 302943 104549
rect 299828 104544 302943 104546
rect 299828 104488 302882 104544
rect 302938 104488 302943 104544
rect 299828 104486 302943 104488
rect 302877 104483 302943 104486
rect 197905 103050 197971 103053
rect 197905 103048 200100 103050
rect 197905 102992 197910 103048
rect 197966 102992 200100 103048
rect 197905 102990 200100 102992
rect 197905 102987 197971 102990
rect 302785 101554 302851 101557
rect 299828 101552 302851 101554
rect 299828 101496 302790 101552
rect 302846 101496 302851 101552
rect 299828 101494 302851 101496
rect 302785 101491 302851 101494
rect 197537 101010 197603 101013
rect 197537 101008 200100 101010
rect 197537 100952 197542 101008
rect 197598 100952 200100 101008
rect 197537 100950 200100 100952
rect 197537 100947 197603 100950
rect 580165 99514 580231 99517
rect 583520 99514 584960 99604
rect 580165 99512 584960 99514
rect 580165 99456 580170 99512
rect 580226 99456 584960 99512
rect 580165 99454 584960 99456
rect 580165 99451 580231 99454
rect 583520 99364 584960 99454
rect 297817 98970 297883 98973
rect 458817 98970 458883 98973
rect 297817 98968 458883 98970
rect 297817 98912 297822 98968
rect 297878 98912 458822 98968
rect 458878 98912 458883 98968
rect 297817 98910 458883 98912
rect 297817 98907 297883 98910
rect 458817 98907 458883 98910
rect 293033 98834 293099 98837
rect 543733 98834 543799 98837
rect 293033 98832 543799 98834
rect 293033 98776 293038 98832
rect 293094 98776 543738 98832
rect 543794 98776 543799 98832
rect 293033 98774 543799 98776
rect 293033 98771 293099 98774
rect 543733 98771 543799 98774
rect 294229 98698 294295 98701
rect 550633 98698 550699 98701
rect 294229 98696 550699 98698
rect 294229 98640 294234 98696
rect 294290 98640 550638 98696
rect 550694 98640 550699 98696
rect 294229 98638 550699 98640
rect 294229 98635 294295 98638
rect 550633 98635 550699 98638
rect 199469 97882 199535 97885
rect 200665 97882 200731 97885
rect 199469 97880 200731 97882
rect 199469 97824 199474 97880
rect 199530 97824 200670 97880
rect 200726 97824 200731 97880
rect 199469 97822 200731 97824
rect 199469 97819 199535 97822
rect 200665 97819 200731 97822
rect -960 97610 480 97700
rect 3417 97610 3483 97613
rect -960 97608 3483 97610
rect -960 97552 3422 97608
rect 3478 97552 3483 97608
rect -960 97550 3483 97552
rect -960 97460 480 97550
rect 3417 97547 3483 97550
rect 196617 97610 196683 97613
rect 204897 97610 204963 97613
rect 196617 97608 204963 97610
rect 196617 97552 196622 97608
rect 196678 97552 204902 97608
rect 204958 97552 204963 97608
rect 196617 97550 204963 97552
rect 196617 97547 196683 97550
rect 204897 97547 204963 97550
rect 289997 97610 290063 97613
rect 300301 97610 300367 97613
rect 289997 97608 300367 97610
rect 289997 97552 290002 97608
rect 290058 97552 300306 97608
rect 300362 97552 300367 97608
rect 289997 97550 300367 97552
rect 289997 97547 290063 97550
rect 300301 97547 300367 97550
rect 35249 97474 35315 97477
rect 204345 97474 204411 97477
rect 35249 97472 204411 97474
rect 35249 97416 35254 97472
rect 35310 97416 204350 97472
rect 204406 97416 204411 97472
rect 35249 97414 204411 97416
rect 35249 97411 35315 97414
rect 204345 97411 204411 97414
rect 281901 97474 281967 97477
rect 461577 97474 461643 97477
rect 281901 97472 461643 97474
rect 281901 97416 281906 97472
rect 281962 97416 461582 97472
rect 461638 97416 461643 97472
rect 281901 97414 461643 97416
rect 281901 97411 281967 97414
rect 461577 97411 461643 97414
rect 29637 97338 29703 97341
rect 203333 97338 203399 97341
rect 29637 97336 203399 97338
rect 29637 97280 29642 97336
rect 29698 97280 203338 97336
rect 203394 97280 203399 97336
rect 29637 97278 203399 97280
rect 29637 97275 29703 97278
rect 203333 97275 203399 97278
rect 299105 97338 299171 97341
rect 299473 97338 299539 97341
rect 580257 97338 580323 97341
rect 299105 97336 299306 97338
rect 299105 97280 299110 97336
rect 299166 97280 299306 97336
rect 299105 97278 299306 97280
rect 299105 97275 299171 97278
rect 17217 97202 17283 97205
rect 202689 97202 202755 97205
rect 17217 97200 202755 97202
rect 17217 97144 17222 97200
rect 17278 97144 202694 97200
rect 202750 97144 202755 97200
rect 17217 97142 202755 97144
rect 17217 97139 17283 97142
rect 202689 97139 202755 97142
rect 284477 97202 284543 97205
rect 297449 97202 297515 97205
rect 284477 97200 297515 97202
rect 284477 97144 284482 97200
rect 284538 97144 297454 97200
rect 297510 97144 297515 97200
rect 284477 97142 297515 97144
rect 299246 97202 299306 97278
rect 299473 97336 580323 97338
rect 299473 97280 299478 97336
rect 299534 97280 580262 97336
rect 580318 97280 580323 97336
rect 299473 97278 580323 97280
rect 299473 97275 299539 97278
rect 580257 97275 580323 97278
rect 582833 97202 582899 97205
rect 299246 97200 582899 97202
rect 299246 97144 582838 97200
rect 582894 97144 582899 97200
rect 299246 97142 582899 97144
rect 284477 97139 284543 97142
rect 297449 97139 297515 97142
rect 582833 97139 582899 97142
rect 289813 96930 289879 96933
rect 291929 96930 291995 96933
rect 289813 96928 291995 96930
rect 289813 96872 289818 96928
rect 289874 96872 291934 96928
rect 291990 96872 291995 96928
rect 289813 96870 291995 96872
rect 289813 96867 289879 96870
rect 291929 96867 291995 96870
rect 296805 96930 296871 96933
rect 300117 96930 300183 96933
rect 296805 96928 300183 96930
rect 296805 96872 296810 96928
rect 296866 96872 300122 96928
rect 300178 96872 300183 96928
rect 296805 96870 300183 96872
rect 296805 96867 296871 96870
rect 300117 96867 300183 96870
rect 297265 96794 297331 96797
rect 300761 96794 300827 96797
rect 297265 96792 300827 96794
rect 297265 96736 297270 96792
rect 297326 96736 300766 96792
rect 300822 96736 300827 96792
rect 297265 96734 300827 96736
rect 297265 96731 297331 96734
rect 300761 96731 300827 96734
rect 22737 95978 22803 95981
rect 203057 95978 203123 95981
rect 22737 95976 203123 95978
rect 22737 95920 22742 95976
rect 22798 95920 203062 95976
rect 203118 95920 203123 95976
rect 22737 95918 203123 95920
rect 22737 95915 22803 95918
rect 203057 95915 203123 95918
rect 12341 95842 12407 95845
rect 201861 95842 201927 95845
rect 12341 95840 201927 95842
rect 12341 95784 12346 95840
rect 12402 95784 201866 95840
rect 201922 95784 201927 95840
rect 12341 95782 201927 95784
rect 12341 95779 12407 95782
rect 201861 95779 201927 95782
rect 298369 95842 298435 95845
rect 557533 95842 557599 95845
rect 298369 95840 557599 95842
rect 298369 95784 298374 95840
rect 298430 95784 557538 95840
rect 557594 95784 557599 95840
rect 298369 95782 557599 95784
rect 298369 95779 298435 95782
rect 557533 95779 557599 95782
rect 291653 94754 291719 94757
rect 536833 94754 536899 94757
rect 291653 94752 536899 94754
rect 291653 94696 291658 94752
rect 291714 94696 536838 94752
rect 536894 94696 536899 94752
rect 291653 94694 536899 94696
rect 291653 94691 291719 94694
rect 536833 94691 536899 94694
rect 28257 94618 28323 94621
rect 203885 94618 203951 94621
rect 28257 94616 203951 94618
rect 28257 94560 28262 94616
rect 28318 94560 203890 94616
rect 203946 94560 203951 94616
rect 28257 94558 203951 94560
rect 28257 94555 28323 94558
rect 203885 94555 203951 94558
rect 296069 94618 296135 94621
rect 561673 94618 561739 94621
rect 296069 94616 561739 94618
rect 296069 94560 296074 94616
rect 296130 94560 561678 94616
rect 561734 94560 561739 94616
rect 296069 94558 561739 94560
rect 296069 94555 296135 94558
rect 561673 94555 561739 94558
rect 1301 94482 1367 94485
rect 200113 94482 200179 94485
rect 1301 94480 200179 94482
rect 1301 94424 1306 94480
rect 1362 94424 200118 94480
rect 200174 94424 200179 94480
rect 1301 94422 200179 94424
rect 1301 94419 1367 94422
rect 200113 94419 200179 94422
rect 300761 94482 300827 94485
rect 568573 94482 568639 94485
rect 300761 94480 568639 94482
rect 300761 94424 300766 94480
rect 300822 94424 568578 94480
rect 568634 94424 568639 94480
rect 300761 94422 568639 94424
rect 300761 94419 300827 94422
rect 568573 94419 568639 94422
rect 4061 93122 4127 93125
rect 199469 93122 199535 93125
rect 4061 93120 199535 93122
rect 4061 93064 4066 93120
rect 4122 93064 199474 93120
rect 199530 93064 199535 93120
rect 4061 93062 199535 93064
rect 4061 93059 4127 93062
rect 199469 93059 199535 93062
rect 299013 93122 299079 93125
rect 575473 93122 575539 93125
rect 299013 93120 575539 93122
rect 299013 93064 299018 93120
rect 299074 93064 575478 93120
rect 575534 93064 575539 93120
rect 299013 93062 575539 93064
rect 299013 93059 299079 93062
rect 575473 93059 575539 93062
rect 582557 86186 582623 86189
rect 583520 86186 584960 86276
rect 582557 86184 584960 86186
rect 582557 86128 582562 86184
rect 582618 86128 584960 86184
rect 582557 86126 584960 86128
rect 582557 86123 582623 86126
rect 583520 86036 584960 86126
rect -960 84690 480 84780
rect 3141 84690 3207 84693
rect -960 84688 3207 84690
rect -960 84632 3146 84688
rect 3202 84632 3207 84688
rect -960 84630 3207 84632
rect -960 84540 480 84630
rect 3141 84627 3207 84630
rect 579981 72994 580047 72997
rect 583520 72994 584960 73084
rect 579981 72992 584960 72994
rect 579981 72936 579986 72992
rect 580042 72936 584960 72992
rect 579981 72934 584960 72936
rect 579981 72931 580047 72934
rect 583520 72844 584960 72934
rect -960 71634 480 71724
rect 3417 71634 3483 71637
rect -960 71632 3483 71634
rect -960 71576 3422 71632
rect 3478 71576 3483 71632
rect -960 71574 3483 71576
rect -960 71484 480 71574
rect 3417 71571 3483 71574
rect 580165 59666 580231 59669
rect 583520 59666 584960 59756
rect 580165 59664 584960 59666
rect 580165 59608 580170 59664
rect 580226 59608 584960 59664
rect 580165 59606 584960 59608
rect 580165 59603 580231 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 3049 58578 3115 58581
rect -960 58576 3115 58578
rect -960 58520 3054 58576
rect 3110 58520 3115 58576
rect -960 58518 3115 58520
rect -960 58428 480 58518
rect 3049 58515 3115 58518
rect 582649 46338 582715 46341
rect 583520 46338 584960 46428
rect 582649 46336 584960 46338
rect 582649 46280 582654 46336
rect 582710 46280 584960 46336
rect 582649 46278 584960 46280
rect 582649 46275 582715 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 3417 45522 3483 45525
rect -960 45520 3483 45522
rect -960 45464 3422 45520
rect 3478 45464 3483 45520
rect -960 45462 3483 45464
rect -960 45372 480 45462
rect 3417 45459 3483 45462
rect 583109 33146 583175 33149
rect 583520 33146 584960 33236
rect 583109 33144 584960 33146
rect 583109 33088 583114 33144
rect 583170 33088 584960 33144
rect 583109 33086 584960 33088
rect 583109 33083 583175 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 2865 32466 2931 32469
rect -960 32464 2931 32466
rect -960 32408 2870 32464
rect 2926 32408 2931 32464
rect -960 32406 2931 32408
rect -960 32316 480 32406
rect 2865 32403 2931 32406
rect 582465 19818 582531 19821
rect 583520 19818 584960 19908
rect 582465 19816 584960 19818
rect 582465 19760 582470 19816
rect 582526 19760 584960 19816
rect 582465 19758 584960 19760
rect 582465 19755 582531 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3417 19410 3483 19413
rect -960 19408 3483 19410
rect -960 19352 3422 19408
rect 3478 19352 3483 19408
rect -960 19350 3483 19352
rect -960 19260 480 19350
rect 3417 19347 3483 19350
rect 582373 6626 582439 6629
rect 583520 6626 584960 6716
rect 582373 6624 584960 6626
rect -960 6490 480 6580
rect 582373 6568 582378 6624
rect 582434 6568 584960 6624
rect 582373 6566 584960 6568
rect 582373 6563 582439 6566
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect 583520 6476 584960 6566
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
rect 260281 3498 260347 3501
rect 350441 3498 350507 3501
rect 260281 3496 350507 3498
rect 260281 3440 260286 3496
rect 260342 3440 350446 3496
rect 350502 3440 350507 3496
rect 260281 3438 350507 3440
rect 260281 3435 260347 3438
rect 350441 3435 350507 3438
rect 260741 3362 260807 3365
rect 349245 3362 349311 3365
rect 260741 3360 349311 3362
rect 260741 3304 260746 3360
rect 260802 3304 349250 3360
rect 349306 3304 349311 3360
rect 260741 3302 349311 3304
rect 260741 3299 260807 3302
rect 349245 3299 349311 3302
<< via3 >>
rect 372108 352412 372172 352476
rect 371740 351324 371804 351388
rect 371372 350780 371436 350844
rect 371188 343300 371252 343364
rect 361620 337724 361684 337788
rect 364380 337724 364444 337788
rect 372108 280468 372172 280532
rect 371924 279924 371988 279988
rect 371740 279380 371804 279444
rect 371372 278836 371436 278900
rect 370268 274756 370332 274820
rect 371188 271356 371252 271420
rect 370084 268364 370148 268428
rect 361620 266052 361684 266116
rect 364380 266052 364444 266116
rect 372108 224980 372172 225044
rect 371924 208388 371988 208452
rect 370268 203084 370332 203148
rect 371372 199276 371436 199340
rect 370084 196556 370148 196620
rect 364380 196012 364444 196076
rect 361620 194516 361684 194580
rect 362724 194516 362788 194580
rect 365300 194516 365364 194580
rect 371740 159292 371804 159356
rect 370084 153036 370148 153100
rect 369900 133996 369964 134060
rect 371740 127332 371804 127396
rect 362724 123992 362788 123996
rect 362724 123936 362774 123992
rect 362774 123936 362788 123992
rect 362724 123932 362788 123936
rect 365300 123932 365364 123996
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 680614 -8106 711002
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 -8106 680614
rect -8726 680294 -8106 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 -8106 680294
rect -8726 644614 -8106 680058
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 -8106 644614
rect -8726 644294 -8106 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 -8106 644294
rect -8726 608614 -8106 644058
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 -8106 608614
rect -8726 608294 -8106 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 -8106 608294
rect -8726 572614 -8106 608058
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 -8106 572614
rect -8726 572294 -8106 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 -8106 572294
rect -8726 536614 -8106 572058
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 -8106 536614
rect -8726 536294 -8106 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 -8106 536294
rect -8726 500614 -8106 536058
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 -8106 500614
rect -8726 500294 -8106 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 -8106 500294
rect -8726 464614 -8106 500058
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 -8106 464614
rect -8726 464294 -8106 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 -8106 464294
rect -8726 428614 -8106 464058
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 -8106 428614
rect -8726 428294 -8106 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 -8106 428294
rect -8726 392614 -8106 428058
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 -8106 392614
rect -8726 392294 -8106 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 -8106 392294
rect -8726 356614 -8106 392058
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 -8106 356614
rect -8726 356294 -8106 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 -8106 356294
rect -8726 320614 -8106 356058
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 -8106 320614
rect -8726 320294 -8106 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 -8106 320294
rect -8726 284614 -8106 320058
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 -8106 284614
rect -8726 284294 -8106 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 -8106 284294
rect -8726 248614 -8106 284058
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 -8106 248614
rect -8726 248294 -8106 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 -8106 248294
rect -8726 212614 -8106 248058
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 -8106 212614
rect -8726 212294 -8106 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 -8106 212294
rect -8726 176614 -8106 212058
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 -8106 176614
rect -8726 176294 -8106 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 -8106 176294
rect -8726 140614 -8106 176058
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 -8106 140614
rect -8726 140294 -8106 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 -8106 140294
rect -8726 104614 -8106 140058
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 -8106 104614
rect -8726 104294 -8106 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 -8106 104294
rect -8726 68614 -8106 104058
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 -8106 68614
rect -8726 68294 -8106 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 -8106 68294
rect -8726 32614 -8106 68058
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 -8106 32614
rect -8726 32294 -8106 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 -8106 32294
rect -8726 -7066 -8106 32058
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 698614 -7146 710042
rect 12954 710598 13574 711590
rect 12954 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 13574 710598
rect 12954 710278 13574 710362
rect 12954 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 13574 710278
rect -7766 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 -7146 698614
rect -7766 698294 -7146 698378
rect -7766 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 -7146 698294
rect -7766 662614 -7146 698058
rect -7766 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 -7146 662614
rect -7766 662294 -7146 662378
rect -7766 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 -7146 662294
rect -7766 626614 -7146 662058
rect -7766 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 -7146 626614
rect -7766 626294 -7146 626378
rect -7766 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 -7146 626294
rect -7766 590614 -7146 626058
rect -7766 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 -7146 590614
rect -7766 590294 -7146 590378
rect -7766 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 -7146 590294
rect -7766 554614 -7146 590058
rect -7766 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 -7146 554614
rect -7766 554294 -7146 554378
rect -7766 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 -7146 554294
rect -7766 518614 -7146 554058
rect -7766 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 -7146 518614
rect -7766 518294 -7146 518378
rect -7766 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 -7146 518294
rect -7766 482614 -7146 518058
rect -7766 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 -7146 482614
rect -7766 482294 -7146 482378
rect -7766 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 -7146 482294
rect -7766 446614 -7146 482058
rect -7766 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 -7146 446614
rect -7766 446294 -7146 446378
rect -7766 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 -7146 446294
rect -7766 410614 -7146 446058
rect -7766 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 -7146 410614
rect -7766 410294 -7146 410378
rect -7766 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 -7146 410294
rect -7766 374614 -7146 410058
rect -7766 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 -7146 374614
rect -7766 374294 -7146 374378
rect -7766 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 -7146 374294
rect -7766 338614 -7146 374058
rect -7766 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 -7146 338614
rect -7766 338294 -7146 338378
rect -7766 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 -7146 338294
rect -7766 302614 -7146 338058
rect -7766 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 -7146 302614
rect -7766 302294 -7146 302378
rect -7766 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 -7146 302294
rect -7766 266614 -7146 302058
rect -7766 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 -7146 266614
rect -7766 266294 -7146 266378
rect -7766 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 -7146 266294
rect -7766 230614 -7146 266058
rect -7766 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 -7146 230614
rect -7766 230294 -7146 230378
rect -7766 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 -7146 230294
rect -7766 194614 -7146 230058
rect -7766 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 -7146 194614
rect -7766 194294 -7146 194378
rect -7766 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 -7146 194294
rect -7766 158614 -7146 194058
rect -7766 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 -7146 158614
rect -7766 158294 -7146 158378
rect -7766 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 -7146 158294
rect -7766 122614 -7146 158058
rect -7766 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 -7146 122614
rect -7766 122294 -7146 122378
rect -7766 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 -7146 122294
rect -7766 86614 -7146 122058
rect -7766 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 -7146 86614
rect -7766 86294 -7146 86378
rect -7766 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 -7146 86294
rect -7766 50614 -7146 86058
rect -7766 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 -7146 50614
rect -7766 50294 -7146 50378
rect -7766 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 -7146 50294
rect -7766 14614 -7146 50058
rect -7766 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 -7146 14614
rect -7766 14294 -7146 14378
rect -7766 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 -7146 14294
rect -7766 -6106 -7146 14058
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 676894 -6186 709082
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 -6186 676894
rect -6806 676574 -6186 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 -6186 676574
rect -6806 640894 -6186 676338
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 -6186 640894
rect -6806 640574 -6186 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 -6186 640574
rect -6806 604894 -6186 640338
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 -6186 604894
rect -6806 604574 -6186 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 -6186 604574
rect -6806 568894 -6186 604338
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 -6186 568894
rect -6806 568574 -6186 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 -6186 568574
rect -6806 532894 -6186 568338
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 -6186 532894
rect -6806 532574 -6186 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 -6186 532574
rect -6806 496894 -6186 532338
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 -6186 496894
rect -6806 496574 -6186 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 -6186 496574
rect -6806 460894 -6186 496338
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 -6186 460894
rect -6806 460574 -6186 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 -6186 460574
rect -6806 424894 -6186 460338
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 -6186 424894
rect -6806 424574 -6186 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 -6186 424574
rect -6806 388894 -6186 424338
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 -6186 388894
rect -6806 388574 -6186 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 -6186 388574
rect -6806 352894 -6186 388338
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 -6186 352894
rect -6806 352574 -6186 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 -6186 352574
rect -6806 316894 -6186 352338
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 -6186 316894
rect -6806 316574 -6186 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 -6186 316574
rect -6806 280894 -6186 316338
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 -6186 280894
rect -6806 280574 -6186 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 -6186 280574
rect -6806 244894 -6186 280338
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 -6186 244894
rect -6806 244574 -6186 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 -6186 244574
rect -6806 208894 -6186 244338
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 -6186 208894
rect -6806 208574 -6186 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 -6186 208574
rect -6806 172894 -6186 208338
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 -6186 172894
rect -6806 172574 -6186 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 -6186 172574
rect -6806 136894 -6186 172338
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 -6186 136894
rect -6806 136574 -6186 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 -6186 136574
rect -6806 100894 -6186 136338
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 -6186 100894
rect -6806 100574 -6186 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 -6186 100574
rect -6806 64894 -6186 100338
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 -6186 64894
rect -6806 64574 -6186 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 -6186 64574
rect -6806 28894 -6186 64338
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 -6186 28894
rect -6806 28574 -6186 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 -6186 28574
rect -6806 -5146 -6186 28338
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 694894 -5226 708122
rect 9234 708678 9854 709670
rect 9234 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 9854 708678
rect 9234 708358 9854 708442
rect 9234 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 9854 708358
rect -5846 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 -5226 694894
rect -5846 694574 -5226 694658
rect -5846 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 -5226 694574
rect -5846 658894 -5226 694338
rect -5846 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 -5226 658894
rect -5846 658574 -5226 658658
rect -5846 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 -5226 658574
rect -5846 622894 -5226 658338
rect -5846 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 -5226 622894
rect -5846 622574 -5226 622658
rect -5846 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 -5226 622574
rect -5846 586894 -5226 622338
rect -5846 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 -5226 586894
rect -5846 586574 -5226 586658
rect -5846 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 -5226 586574
rect -5846 550894 -5226 586338
rect -5846 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 -5226 550894
rect -5846 550574 -5226 550658
rect -5846 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 -5226 550574
rect -5846 514894 -5226 550338
rect -5846 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 -5226 514894
rect -5846 514574 -5226 514658
rect -5846 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 -5226 514574
rect -5846 478894 -5226 514338
rect -5846 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 -5226 478894
rect -5846 478574 -5226 478658
rect -5846 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 -5226 478574
rect -5846 442894 -5226 478338
rect -5846 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 -5226 442894
rect -5846 442574 -5226 442658
rect -5846 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 -5226 442574
rect -5846 406894 -5226 442338
rect -5846 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 -5226 406894
rect -5846 406574 -5226 406658
rect -5846 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 -5226 406574
rect -5846 370894 -5226 406338
rect -5846 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 -5226 370894
rect -5846 370574 -5226 370658
rect -5846 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 -5226 370574
rect -5846 334894 -5226 370338
rect -5846 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 -5226 334894
rect -5846 334574 -5226 334658
rect -5846 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 -5226 334574
rect -5846 298894 -5226 334338
rect -5846 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 -5226 298894
rect -5846 298574 -5226 298658
rect -5846 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 -5226 298574
rect -5846 262894 -5226 298338
rect -5846 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 -5226 262894
rect -5846 262574 -5226 262658
rect -5846 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 -5226 262574
rect -5846 226894 -5226 262338
rect -5846 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 -5226 226894
rect -5846 226574 -5226 226658
rect -5846 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 -5226 226574
rect -5846 190894 -5226 226338
rect -5846 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 -5226 190894
rect -5846 190574 -5226 190658
rect -5846 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 -5226 190574
rect -5846 154894 -5226 190338
rect -5846 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 -5226 154894
rect -5846 154574 -5226 154658
rect -5846 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 -5226 154574
rect -5846 118894 -5226 154338
rect -5846 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 -5226 118894
rect -5846 118574 -5226 118658
rect -5846 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 -5226 118574
rect -5846 82894 -5226 118338
rect -5846 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 -5226 82894
rect -5846 82574 -5226 82658
rect -5846 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 -5226 82574
rect -5846 46894 -5226 82338
rect -5846 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 -5226 46894
rect -5846 46574 -5226 46658
rect -5846 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 -5226 46574
rect -5846 10894 -5226 46338
rect -5846 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 -5226 10894
rect -5846 10574 -5226 10658
rect -5846 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 -5226 10574
rect -5846 -4186 -5226 10338
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 673174 -4266 707162
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 -4266 673174
rect -4886 672854 -4266 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 -4266 672854
rect -4886 637174 -4266 672618
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 -4266 637174
rect -4886 636854 -4266 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 -4266 636854
rect -4886 601174 -4266 636618
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 -4266 601174
rect -4886 600854 -4266 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 -4266 600854
rect -4886 565174 -4266 600618
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 -4266 565174
rect -4886 564854 -4266 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 -4266 564854
rect -4886 529174 -4266 564618
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 -4266 529174
rect -4886 528854 -4266 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 -4266 528854
rect -4886 493174 -4266 528618
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 -4266 493174
rect -4886 492854 -4266 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 -4266 492854
rect -4886 457174 -4266 492618
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 -4266 457174
rect -4886 456854 -4266 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 -4266 456854
rect -4886 421174 -4266 456618
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 -4266 421174
rect -4886 420854 -4266 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 -4266 420854
rect -4886 385174 -4266 420618
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 -4266 385174
rect -4886 384854 -4266 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 -4266 384854
rect -4886 349174 -4266 384618
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 -4266 349174
rect -4886 348854 -4266 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 -4266 348854
rect -4886 313174 -4266 348618
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 -4266 313174
rect -4886 312854 -4266 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 -4266 312854
rect -4886 277174 -4266 312618
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 -4266 277174
rect -4886 276854 -4266 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 -4266 276854
rect -4886 241174 -4266 276618
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 -4266 241174
rect -4886 240854 -4266 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 -4266 240854
rect -4886 205174 -4266 240618
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 -4266 205174
rect -4886 204854 -4266 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 -4266 204854
rect -4886 169174 -4266 204618
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 -4266 169174
rect -4886 168854 -4266 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 -4266 168854
rect -4886 133174 -4266 168618
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 -4266 133174
rect -4886 132854 -4266 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 -4266 132854
rect -4886 97174 -4266 132618
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 -4266 97174
rect -4886 96854 -4266 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 -4266 96854
rect -4886 61174 -4266 96618
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 -4266 61174
rect -4886 60854 -4266 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 -4266 60854
rect -4886 25174 -4266 60618
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 -4266 25174
rect -4886 24854 -4266 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 -4266 24854
rect -4886 -3226 -4266 24618
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 691174 -3306 706202
rect 5514 706758 6134 707750
rect 5514 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 6134 706758
rect 5514 706438 6134 706522
rect 5514 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 6134 706438
rect -3926 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 -3306 691174
rect -3926 690854 -3306 690938
rect -3926 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 -3306 690854
rect -3926 655174 -3306 690618
rect -3926 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 -3306 655174
rect -3926 654854 -3306 654938
rect -3926 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 -3306 654854
rect -3926 619174 -3306 654618
rect -3926 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 -3306 619174
rect -3926 618854 -3306 618938
rect -3926 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 -3306 618854
rect -3926 583174 -3306 618618
rect -3926 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 -3306 583174
rect -3926 582854 -3306 582938
rect -3926 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 -3306 582854
rect -3926 547174 -3306 582618
rect -3926 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 -3306 547174
rect -3926 546854 -3306 546938
rect -3926 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 -3306 546854
rect -3926 511174 -3306 546618
rect -3926 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 -3306 511174
rect -3926 510854 -3306 510938
rect -3926 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 -3306 510854
rect -3926 475174 -3306 510618
rect -3926 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 -3306 475174
rect -3926 474854 -3306 474938
rect -3926 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 -3306 474854
rect -3926 439174 -3306 474618
rect -3926 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 -3306 439174
rect -3926 438854 -3306 438938
rect -3926 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 -3306 438854
rect -3926 403174 -3306 438618
rect -3926 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 -3306 403174
rect -3926 402854 -3306 402938
rect -3926 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 -3306 402854
rect -3926 367174 -3306 402618
rect -3926 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 -3306 367174
rect -3926 366854 -3306 366938
rect -3926 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 -3306 366854
rect -3926 331174 -3306 366618
rect -3926 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 -3306 331174
rect -3926 330854 -3306 330938
rect -3926 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 -3306 330854
rect -3926 295174 -3306 330618
rect -3926 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 -3306 295174
rect -3926 294854 -3306 294938
rect -3926 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 -3306 294854
rect -3926 259174 -3306 294618
rect -3926 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 -3306 259174
rect -3926 258854 -3306 258938
rect -3926 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 -3306 258854
rect -3926 223174 -3306 258618
rect -3926 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 -3306 223174
rect -3926 222854 -3306 222938
rect -3926 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 -3306 222854
rect -3926 187174 -3306 222618
rect -3926 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 -3306 187174
rect -3926 186854 -3306 186938
rect -3926 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 -3306 186854
rect -3926 151174 -3306 186618
rect -3926 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 -3306 151174
rect -3926 150854 -3306 150938
rect -3926 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 -3306 150854
rect -3926 115174 -3306 150618
rect -3926 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 -3306 115174
rect -3926 114854 -3306 114938
rect -3926 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 -3306 114854
rect -3926 79174 -3306 114618
rect -3926 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 -3306 79174
rect -3926 78854 -3306 78938
rect -3926 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 -3306 78854
rect -3926 43174 -3306 78618
rect -3926 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 -3306 43174
rect -3926 42854 -3306 42938
rect -3926 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 -3306 42854
rect -3926 7174 -3306 42618
rect -3926 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 -3306 7174
rect -3926 6854 -3306 6938
rect -3926 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 -3306 6854
rect -3926 -2266 -3306 6618
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 669454 -2346 705242
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 -2346 669454
rect -2966 669134 -2346 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 -2346 669134
rect -2966 633454 -2346 668898
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 -2346 633454
rect -2966 633134 -2346 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 -2346 633134
rect -2966 597454 -2346 632898
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 -2346 597454
rect -2966 597134 -2346 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 -2346 597134
rect -2966 561454 -2346 596898
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 -2346 561454
rect -2966 561134 -2346 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 -2346 561134
rect -2966 525454 -2346 560898
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 -2346 525454
rect -2966 525134 -2346 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 -2346 525134
rect -2966 489454 -2346 524898
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 -2346 489454
rect -2966 489134 -2346 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 -2346 489134
rect -2966 453454 -2346 488898
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 -2346 453454
rect -2966 453134 -2346 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 -2346 453134
rect -2966 417454 -2346 452898
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 -2346 417454
rect -2966 417134 -2346 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 -2346 417134
rect -2966 381454 -2346 416898
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 -2346 381454
rect -2966 381134 -2346 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 -2346 381134
rect -2966 345454 -2346 380898
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 -2346 345454
rect -2966 345134 -2346 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 -2346 345134
rect -2966 309454 -2346 344898
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 -2346 309454
rect -2966 309134 -2346 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 -2346 309134
rect -2966 273454 -2346 308898
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 -2346 273454
rect -2966 273134 -2346 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 -2346 273134
rect -2966 237454 -2346 272898
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 -2346 237454
rect -2966 237134 -2346 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 -2346 237134
rect -2966 201454 -2346 236898
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 -2346 201454
rect -2966 201134 -2346 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 -2346 201134
rect -2966 165454 -2346 200898
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 -2346 165454
rect -2966 165134 -2346 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 -2346 165134
rect -2966 129454 -2346 164898
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 -2346 129454
rect -2966 129134 -2346 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 -2346 129134
rect -2966 93454 -2346 128898
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 -2346 93454
rect -2966 93134 -2346 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 -2346 93134
rect -2966 57454 -2346 92898
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 -2346 57454
rect -2966 57134 -2346 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 -2346 57134
rect -2966 21454 -2346 56898
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 -2346 21454
rect -2966 21134 -2346 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 -2346 21134
rect -2966 -1306 -2346 20898
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 705830
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 1794 -1894 2414 -902
rect 5514 691174 6134 706202
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 5514 619174 6134 654618
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 5514 259174 6134 294618
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 5514 223174 6134 258618
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 5514 187174 6134 222618
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 5514 151174 6134 186618
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 5514 115174 6134 150618
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 5514 79174 6134 114618
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 5514 43174 6134 78618
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 5514 7174 6134 42618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect 5514 -2266 6134 6618
rect 5514 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 6134 -2266
rect 5514 -2586 6134 -2502
rect 5514 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 6134 -2586
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect 5514 -3814 6134 -2822
rect 9234 694894 9854 708122
rect 9234 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 9854 694894
rect 9234 694574 9854 694658
rect 9234 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 9854 694574
rect 9234 658894 9854 694338
rect 9234 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 9854 658894
rect 9234 658574 9854 658658
rect 9234 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 9854 658574
rect 9234 622894 9854 658338
rect 9234 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 9854 622894
rect 9234 622574 9854 622658
rect 9234 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 9854 622574
rect 9234 586894 9854 622338
rect 9234 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 9854 586894
rect 9234 586574 9854 586658
rect 9234 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 9854 586574
rect 9234 550894 9854 586338
rect 9234 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 9854 550894
rect 9234 550574 9854 550658
rect 9234 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 9854 550574
rect 9234 514894 9854 550338
rect 9234 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 9854 514894
rect 9234 514574 9854 514658
rect 9234 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 9854 514574
rect 9234 478894 9854 514338
rect 9234 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 9854 478894
rect 9234 478574 9854 478658
rect 9234 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 9854 478574
rect 9234 442894 9854 478338
rect 9234 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 9854 442894
rect 9234 442574 9854 442658
rect 9234 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 9854 442574
rect 9234 406894 9854 442338
rect 9234 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 9854 406894
rect 9234 406574 9854 406658
rect 9234 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 9854 406574
rect 9234 370894 9854 406338
rect 9234 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 9854 370894
rect 9234 370574 9854 370658
rect 9234 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 9854 370574
rect 9234 334894 9854 370338
rect 9234 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 9854 334894
rect 9234 334574 9854 334658
rect 9234 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 9854 334574
rect 9234 298894 9854 334338
rect 9234 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 9854 298894
rect 9234 298574 9854 298658
rect 9234 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 9854 298574
rect 9234 262894 9854 298338
rect 9234 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 9854 262894
rect 9234 262574 9854 262658
rect 9234 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 9854 262574
rect 9234 226894 9854 262338
rect 9234 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 9854 226894
rect 9234 226574 9854 226658
rect 9234 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 9854 226574
rect 9234 190894 9854 226338
rect 9234 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 9854 190894
rect 9234 190574 9854 190658
rect 9234 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 9854 190574
rect 9234 154894 9854 190338
rect 9234 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 9854 154894
rect 9234 154574 9854 154658
rect 9234 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 9854 154574
rect 9234 118894 9854 154338
rect 9234 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 9854 118894
rect 9234 118574 9854 118658
rect 9234 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 9854 118574
rect 9234 82894 9854 118338
rect 9234 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 9854 82894
rect 9234 82574 9854 82658
rect 9234 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 9854 82574
rect 9234 46894 9854 82338
rect 9234 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 9854 46894
rect 9234 46574 9854 46658
rect 9234 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 9854 46574
rect 9234 10894 9854 46338
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect 9234 -4186 9854 10338
rect 9234 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 9854 -4186
rect 9234 -4506 9854 -4422
rect 9234 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 9854 -4506
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect 9234 -5734 9854 -4742
rect 12954 698614 13574 710042
rect 30954 711558 31574 711590
rect 30954 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 31574 711558
rect 30954 711238 31574 711322
rect 30954 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 31574 711238
rect 27234 709638 27854 709670
rect 27234 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 27854 709638
rect 27234 709318 27854 709402
rect 27234 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 27854 709318
rect 23514 707718 24134 707750
rect 23514 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 24134 707718
rect 23514 707398 24134 707482
rect 23514 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 24134 707398
rect 12954 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 13574 698614
rect 12954 698294 13574 698378
rect 12954 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 13574 698294
rect 12954 662614 13574 698058
rect 12954 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 13574 662614
rect 12954 662294 13574 662378
rect 12954 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 13574 662294
rect 12954 626614 13574 662058
rect 12954 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 13574 626614
rect 12954 626294 13574 626378
rect 12954 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 13574 626294
rect 12954 590614 13574 626058
rect 12954 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 13574 590614
rect 12954 590294 13574 590378
rect 12954 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 13574 590294
rect 12954 554614 13574 590058
rect 12954 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 13574 554614
rect 12954 554294 13574 554378
rect 12954 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 13574 554294
rect 12954 518614 13574 554058
rect 12954 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 13574 518614
rect 12954 518294 13574 518378
rect 12954 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 13574 518294
rect 12954 482614 13574 518058
rect 12954 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 13574 482614
rect 12954 482294 13574 482378
rect 12954 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 13574 482294
rect 12954 446614 13574 482058
rect 12954 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 13574 446614
rect 12954 446294 13574 446378
rect 12954 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 13574 446294
rect 12954 410614 13574 446058
rect 12954 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 13574 410614
rect 12954 410294 13574 410378
rect 12954 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 13574 410294
rect 12954 374614 13574 410058
rect 12954 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 13574 374614
rect 12954 374294 13574 374378
rect 12954 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 13574 374294
rect 12954 338614 13574 374058
rect 12954 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 13574 338614
rect 12954 338294 13574 338378
rect 12954 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 13574 338294
rect 12954 302614 13574 338058
rect 12954 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 13574 302614
rect 12954 302294 13574 302378
rect 12954 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 13574 302294
rect 12954 266614 13574 302058
rect 12954 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 13574 266614
rect 12954 266294 13574 266378
rect 12954 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 13574 266294
rect 12954 230614 13574 266058
rect 12954 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 13574 230614
rect 12954 230294 13574 230378
rect 12954 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 13574 230294
rect 12954 194614 13574 230058
rect 12954 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 13574 194614
rect 12954 194294 13574 194378
rect 12954 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 13574 194294
rect 12954 158614 13574 194058
rect 12954 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 13574 158614
rect 12954 158294 13574 158378
rect 12954 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 13574 158294
rect 12954 122614 13574 158058
rect 12954 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 13574 122614
rect 12954 122294 13574 122378
rect 12954 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 13574 122294
rect 12954 86614 13574 122058
rect 12954 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 13574 86614
rect 12954 86294 13574 86378
rect 12954 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 13574 86294
rect 12954 50614 13574 86058
rect 12954 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 13574 50614
rect 12954 50294 13574 50378
rect 12954 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 13574 50294
rect 12954 14614 13574 50058
rect 12954 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 13574 14614
rect 12954 14294 13574 14378
rect 12954 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 13574 14294
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect 12954 -6106 13574 14058
rect 19794 705798 20414 705830
rect 19794 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 20414 705798
rect 19794 705478 20414 705562
rect 19794 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 20414 705478
rect 19794 669454 20414 705242
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -1306 20414 20898
rect 19794 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 20414 -1306
rect 19794 -1626 20414 -1542
rect 19794 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 20414 -1626
rect 19794 -1894 20414 -1862
rect 23514 673174 24134 707162
rect 23514 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 24134 673174
rect 23514 672854 24134 672938
rect 23514 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 24134 672854
rect 23514 637174 24134 672618
rect 23514 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 24134 637174
rect 23514 636854 24134 636938
rect 23514 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 24134 636854
rect 23514 601174 24134 636618
rect 23514 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 24134 601174
rect 23514 600854 24134 600938
rect 23514 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 24134 600854
rect 23514 565174 24134 600618
rect 23514 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 24134 565174
rect 23514 564854 24134 564938
rect 23514 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 24134 564854
rect 23514 529174 24134 564618
rect 23514 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 24134 529174
rect 23514 528854 24134 528938
rect 23514 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 24134 528854
rect 23514 493174 24134 528618
rect 23514 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 24134 493174
rect 23514 492854 24134 492938
rect 23514 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 24134 492854
rect 23514 457174 24134 492618
rect 23514 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 24134 457174
rect 23514 456854 24134 456938
rect 23514 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 24134 456854
rect 23514 421174 24134 456618
rect 23514 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 24134 421174
rect 23514 420854 24134 420938
rect 23514 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 24134 420854
rect 23514 385174 24134 420618
rect 23514 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 24134 385174
rect 23514 384854 24134 384938
rect 23514 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 24134 384854
rect 23514 349174 24134 384618
rect 23514 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 24134 349174
rect 23514 348854 24134 348938
rect 23514 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 24134 348854
rect 23514 313174 24134 348618
rect 23514 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 24134 313174
rect 23514 312854 24134 312938
rect 23514 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 24134 312854
rect 23514 277174 24134 312618
rect 23514 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 24134 277174
rect 23514 276854 24134 276938
rect 23514 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 24134 276854
rect 23514 241174 24134 276618
rect 23514 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 24134 241174
rect 23514 240854 24134 240938
rect 23514 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 24134 240854
rect 23514 205174 24134 240618
rect 23514 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 24134 205174
rect 23514 204854 24134 204938
rect 23514 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 24134 204854
rect 23514 169174 24134 204618
rect 23514 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 24134 169174
rect 23514 168854 24134 168938
rect 23514 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 24134 168854
rect 23514 133174 24134 168618
rect 23514 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 24134 133174
rect 23514 132854 24134 132938
rect 23514 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 24134 132854
rect 23514 97174 24134 132618
rect 23514 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 24134 97174
rect 23514 96854 24134 96938
rect 23514 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 24134 96854
rect 23514 61174 24134 96618
rect 23514 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 24134 61174
rect 23514 60854 24134 60938
rect 23514 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 24134 60854
rect 23514 25174 24134 60618
rect 23514 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 24134 25174
rect 23514 24854 24134 24938
rect 23514 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 24134 24854
rect 23514 -3226 24134 24618
rect 23514 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 24134 -3226
rect 23514 -3546 24134 -3462
rect 23514 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 24134 -3546
rect 23514 -3814 24134 -3782
rect 27234 676894 27854 709082
rect 27234 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 27854 676894
rect 27234 676574 27854 676658
rect 27234 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 27854 676574
rect 27234 640894 27854 676338
rect 27234 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 27854 640894
rect 27234 640574 27854 640658
rect 27234 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 27854 640574
rect 27234 604894 27854 640338
rect 27234 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 27854 604894
rect 27234 604574 27854 604658
rect 27234 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 27854 604574
rect 27234 568894 27854 604338
rect 27234 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 27854 568894
rect 27234 568574 27854 568658
rect 27234 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 27854 568574
rect 27234 532894 27854 568338
rect 27234 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 27854 532894
rect 27234 532574 27854 532658
rect 27234 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 27854 532574
rect 27234 496894 27854 532338
rect 27234 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 27854 496894
rect 27234 496574 27854 496658
rect 27234 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 27854 496574
rect 27234 460894 27854 496338
rect 27234 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 27854 460894
rect 27234 460574 27854 460658
rect 27234 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 27854 460574
rect 27234 424894 27854 460338
rect 27234 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 27854 424894
rect 27234 424574 27854 424658
rect 27234 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 27854 424574
rect 27234 388894 27854 424338
rect 27234 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 27854 388894
rect 27234 388574 27854 388658
rect 27234 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 27854 388574
rect 27234 352894 27854 388338
rect 27234 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 27854 352894
rect 27234 352574 27854 352658
rect 27234 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 27854 352574
rect 27234 316894 27854 352338
rect 27234 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 27854 316894
rect 27234 316574 27854 316658
rect 27234 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 27854 316574
rect 27234 280894 27854 316338
rect 27234 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 27854 280894
rect 27234 280574 27854 280658
rect 27234 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 27854 280574
rect 27234 244894 27854 280338
rect 27234 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 27854 244894
rect 27234 244574 27854 244658
rect 27234 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 27854 244574
rect 27234 208894 27854 244338
rect 27234 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 27854 208894
rect 27234 208574 27854 208658
rect 27234 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 27854 208574
rect 27234 172894 27854 208338
rect 27234 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 27854 172894
rect 27234 172574 27854 172658
rect 27234 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 27854 172574
rect 27234 136894 27854 172338
rect 27234 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 27854 136894
rect 27234 136574 27854 136658
rect 27234 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 27854 136574
rect 27234 100894 27854 136338
rect 27234 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 27854 100894
rect 27234 100574 27854 100658
rect 27234 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 27854 100574
rect 27234 64894 27854 100338
rect 27234 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 27854 64894
rect 27234 64574 27854 64658
rect 27234 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 27854 64574
rect 27234 28894 27854 64338
rect 27234 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 27854 28894
rect 27234 28574 27854 28658
rect 27234 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 27854 28574
rect 27234 -5146 27854 28338
rect 27234 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 27854 -5146
rect 27234 -5466 27854 -5382
rect 27234 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 27854 -5466
rect 27234 -5734 27854 -5702
rect 30954 680614 31574 711002
rect 48954 710598 49574 711590
rect 48954 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 49574 710598
rect 48954 710278 49574 710362
rect 48954 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 49574 710278
rect 45234 708678 45854 709670
rect 45234 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 45854 708678
rect 45234 708358 45854 708442
rect 45234 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 45854 708358
rect 41514 706758 42134 707750
rect 41514 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 42134 706758
rect 41514 706438 42134 706522
rect 41514 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 42134 706438
rect 30954 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 31574 680614
rect 30954 680294 31574 680378
rect 30954 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 31574 680294
rect 30954 644614 31574 680058
rect 30954 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 31574 644614
rect 30954 644294 31574 644378
rect 30954 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 31574 644294
rect 30954 608614 31574 644058
rect 30954 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 31574 608614
rect 30954 608294 31574 608378
rect 30954 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 31574 608294
rect 30954 572614 31574 608058
rect 30954 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 31574 572614
rect 30954 572294 31574 572378
rect 30954 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 31574 572294
rect 30954 536614 31574 572058
rect 30954 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 31574 536614
rect 30954 536294 31574 536378
rect 30954 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 31574 536294
rect 30954 500614 31574 536058
rect 30954 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 31574 500614
rect 30954 500294 31574 500378
rect 30954 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 31574 500294
rect 30954 464614 31574 500058
rect 30954 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 31574 464614
rect 30954 464294 31574 464378
rect 30954 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 31574 464294
rect 30954 428614 31574 464058
rect 30954 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 31574 428614
rect 30954 428294 31574 428378
rect 30954 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 31574 428294
rect 30954 392614 31574 428058
rect 30954 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 31574 392614
rect 30954 392294 31574 392378
rect 30954 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 31574 392294
rect 30954 356614 31574 392058
rect 30954 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 31574 356614
rect 30954 356294 31574 356378
rect 30954 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 31574 356294
rect 30954 320614 31574 356058
rect 30954 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 31574 320614
rect 30954 320294 31574 320378
rect 30954 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 31574 320294
rect 30954 284614 31574 320058
rect 30954 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 31574 284614
rect 30954 284294 31574 284378
rect 30954 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 31574 284294
rect 30954 248614 31574 284058
rect 30954 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 31574 248614
rect 30954 248294 31574 248378
rect 30954 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 31574 248294
rect 30954 212614 31574 248058
rect 30954 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 31574 212614
rect 30954 212294 31574 212378
rect 30954 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 31574 212294
rect 30954 176614 31574 212058
rect 30954 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 31574 176614
rect 30954 176294 31574 176378
rect 30954 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 31574 176294
rect 30954 140614 31574 176058
rect 30954 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 31574 140614
rect 30954 140294 31574 140378
rect 30954 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 31574 140294
rect 30954 104614 31574 140058
rect 30954 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 31574 104614
rect 30954 104294 31574 104378
rect 30954 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 31574 104294
rect 30954 68614 31574 104058
rect 30954 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 31574 68614
rect 30954 68294 31574 68378
rect 30954 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 31574 68294
rect 30954 32614 31574 68058
rect 30954 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 31574 32614
rect 30954 32294 31574 32378
rect 30954 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 31574 32294
rect 12954 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 13574 -6106
rect 12954 -6426 13574 -6342
rect 12954 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 13574 -6426
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 12954 -7654 13574 -6662
rect 30954 -7066 31574 32058
rect 37794 704838 38414 705830
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -1894 38414 -902
rect 41514 691174 42134 706202
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 41514 655174 42134 690618
rect 41514 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 42134 655174
rect 41514 654854 42134 654938
rect 41514 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 42134 654854
rect 41514 619174 42134 654618
rect 41514 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 42134 619174
rect 41514 618854 42134 618938
rect 41514 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 42134 618854
rect 41514 583174 42134 618618
rect 41514 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 42134 583174
rect 41514 582854 42134 582938
rect 41514 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 42134 582854
rect 41514 547174 42134 582618
rect 41514 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 42134 547174
rect 41514 546854 42134 546938
rect 41514 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 42134 546854
rect 41514 511174 42134 546618
rect 41514 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 42134 511174
rect 41514 510854 42134 510938
rect 41514 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 42134 510854
rect 41514 475174 42134 510618
rect 41514 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 42134 475174
rect 41514 474854 42134 474938
rect 41514 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 42134 474854
rect 41514 439174 42134 474618
rect 41514 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 42134 439174
rect 41514 438854 42134 438938
rect 41514 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 42134 438854
rect 41514 403174 42134 438618
rect 41514 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 42134 403174
rect 41514 402854 42134 402938
rect 41514 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 42134 402854
rect 41514 367174 42134 402618
rect 41514 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 42134 367174
rect 41514 366854 42134 366938
rect 41514 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 42134 366854
rect 41514 331174 42134 366618
rect 41514 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 42134 331174
rect 41514 330854 42134 330938
rect 41514 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 42134 330854
rect 41514 295174 42134 330618
rect 41514 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 42134 295174
rect 41514 294854 42134 294938
rect 41514 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 42134 294854
rect 41514 259174 42134 294618
rect 41514 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 42134 259174
rect 41514 258854 42134 258938
rect 41514 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 42134 258854
rect 41514 223174 42134 258618
rect 41514 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 42134 223174
rect 41514 222854 42134 222938
rect 41514 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 42134 222854
rect 41514 187174 42134 222618
rect 41514 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 42134 187174
rect 41514 186854 42134 186938
rect 41514 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 42134 186854
rect 41514 151174 42134 186618
rect 41514 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 42134 151174
rect 41514 150854 42134 150938
rect 41514 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 42134 150854
rect 41514 115174 42134 150618
rect 41514 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 42134 115174
rect 41514 114854 42134 114938
rect 41514 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 42134 114854
rect 41514 79174 42134 114618
rect 41514 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 42134 79174
rect 41514 78854 42134 78938
rect 41514 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 42134 78854
rect 41514 43174 42134 78618
rect 41514 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 42134 43174
rect 41514 42854 42134 42938
rect 41514 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 42134 42854
rect 41514 7174 42134 42618
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -2266 42134 6618
rect 41514 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 42134 -2266
rect 41514 -2586 42134 -2502
rect 41514 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 42134 -2586
rect 41514 -3814 42134 -2822
rect 45234 694894 45854 708122
rect 45234 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 45854 694894
rect 45234 694574 45854 694658
rect 45234 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 45854 694574
rect 45234 658894 45854 694338
rect 45234 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 45854 658894
rect 45234 658574 45854 658658
rect 45234 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 45854 658574
rect 45234 622894 45854 658338
rect 45234 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 45854 622894
rect 45234 622574 45854 622658
rect 45234 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 45854 622574
rect 45234 586894 45854 622338
rect 45234 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 45854 586894
rect 45234 586574 45854 586658
rect 45234 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 45854 586574
rect 45234 550894 45854 586338
rect 45234 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 45854 550894
rect 45234 550574 45854 550658
rect 45234 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 45854 550574
rect 45234 514894 45854 550338
rect 45234 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 45854 514894
rect 45234 514574 45854 514658
rect 45234 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 45854 514574
rect 45234 478894 45854 514338
rect 45234 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 45854 478894
rect 45234 478574 45854 478658
rect 45234 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 45854 478574
rect 45234 442894 45854 478338
rect 45234 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 45854 442894
rect 45234 442574 45854 442658
rect 45234 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 45854 442574
rect 45234 406894 45854 442338
rect 45234 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 45854 406894
rect 45234 406574 45854 406658
rect 45234 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 45854 406574
rect 45234 370894 45854 406338
rect 45234 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 45854 370894
rect 45234 370574 45854 370658
rect 45234 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 45854 370574
rect 45234 334894 45854 370338
rect 45234 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 45854 334894
rect 45234 334574 45854 334658
rect 45234 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 45854 334574
rect 45234 298894 45854 334338
rect 45234 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 45854 298894
rect 45234 298574 45854 298658
rect 45234 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 45854 298574
rect 45234 262894 45854 298338
rect 45234 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 45854 262894
rect 45234 262574 45854 262658
rect 45234 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 45854 262574
rect 45234 226894 45854 262338
rect 45234 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 45854 226894
rect 45234 226574 45854 226658
rect 45234 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 45854 226574
rect 45234 190894 45854 226338
rect 45234 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 45854 190894
rect 45234 190574 45854 190658
rect 45234 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 45854 190574
rect 45234 154894 45854 190338
rect 45234 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 45854 154894
rect 45234 154574 45854 154658
rect 45234 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 45854 154574
rect 45234 118894 45854 154338
rect 45234 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 45854 118894
rect 45234 118574 45854 118658
rect 45234 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 45854 118574
rect 45234 82894 45854 118338
rect 45234 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 45854 82894
rect 45234 82574 45854 82658
rect 45234 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 45854 82574
rect 45234 46894 45854 82338
rect 45234 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 45854 46894
rect 45234 46574 45854 46658
rect 45234 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 45854 46574
rect 45234 10894 45854 46338
rect 45234 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 45854 10894
rect 45234 10574 45854 10658
rect 45234 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 45854 10574
rect 45234 -4186 45854 10338
rect 45234 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 45854 -4186
rect 45234 -4506 45854 -4422
rect 45234 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 45854 -4506
rect 45234 -5734 45854 -4742
rect 48954 698614 49574 710042
rect 66954 711558 67574 711590
rect 66954 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 67574 711558
rect 66954 711238 67574 711322
rect 66954 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 67574 711238
rect 63234 709638 63854 709670
rect 63234 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 63854 709638
rect 63234 709318 63854 709402
rect 63234 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 63854 709318
rect 59514 707718 60134 707750
rect 59514 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 60134 707718
rect 59514 707398 60134 707482
rect 59514 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 60134 707398
rect 48954 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 49574 698614
rect 48954 698294 49574 698378
rect 48954 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 49574 698294
rect 48954 662614 49574 698058
rect 48954 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 49574 662614
rect 48954 662294 49574 662378
rect 48954 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 49574 662294
rect 48954 626614 49574 662058
rect 48954 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 49574 626614
rect 48954 626294 49574 626378
rect 48954 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 49574 626294
rect 48954 590614 49574 626058
rect 48954 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 49574 590614
rect 48954 590294 49574 590378
rect 48954 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 49574 590294
rect 48954 554614 49574 590058
rect 48954 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 49574 554614
rect 48954 554294 49574 554378
rect 48954 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 49574 554294
rect 48954 518614 49574 554058
rect 48954 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 49574 518614
rect 48954 518294 49574 518378
rect 48954 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 49574 518294
rect 48954 482614 49574 518058
rect 48954 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 49574 482614
rect 48954 482294 49574 482378
rect 48954 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 49574 482294
rect 48954 446614 49574 482058
rect 48954 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 49574 446614
rect 48954 446294 49574 446378
rect 48954 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 49574 446294
rect 48954 410614 49574 446058
rect 48954 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 49574 410614
rect 48954 410294 49574 410378
rect 48954 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 49574 410294
rect 48954 374614 49574 410058
rect 48954 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 49574 374614
rect 48954 374294 49574 374378
rect 48954 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 49574 374294
rect 48954 338614 49574 374058
rect 48954 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 49574 338614
rect 48954 338294 49574 338378
rect 48954 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 49574 338294
rect 48954 302614 49574 338058
rect 48954 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 49574 302614
rect 48954 302294 49574 302378
rect 48954 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 49574 302294
rect 48954 266614 49574 302058
rect 48954 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 49574 266614
rect 48954 266294 49574 266378
rect 48954 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 49574 266294
rect 48954 230614 49574 266058
rect 48954 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 49574 230614
rect 48954 230294 49574 230378
rect 48954 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 49574 230294
rect 48954 194614 49574 230058
rect 48954 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 49574 194614
rect 48954 194294 49574 194378
rect 48954 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 49574 194294
rect 48954 158614 49574 194058
rect 48954 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 49574 158614
rect 48954 158294 49574 158378
rect 48954 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 49574 158294
rect 48954 122614 49574 158058
rect 48954 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 49574 122614
rect 48954 122294 49574 122378
rect 48954 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 49574 122294
rect 48954 86614 49574 122058
rect 48954 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 49574 86614
rect 48954 86294 49574 86378
rect 48954 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 49574 86294
rect 48954 50614 49574 86058
rect 48954 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 49574 50614
rect 48954 50294 49574 50378
rect 48954 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 49574 50294
rect 48954 14614 49574 50058
rect 48954 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 49574 14614
rect 48954 14294 49574 14378
rect 48954 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 49574 14294
rect 30954 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 31574 -7066
rect 30954 -7386 31574 -7302
rect 30954 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 31574 -7386
rect 30954 -7654 31574 -7622
rect 48954 -6106 49574 14058
rect 55794 705798 56414 705830
rect 55794 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 56414 705798
rect 55794 705478 56414 705562
rect 55794 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 56414 705478
rect 55794 669454 56414 705242
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 273454 56414 308898
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 237454 56414 272898
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55794 201454 56414 236898
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -1306 56414 20898
rect 55794 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 56414 -1306
rect 55794 -1626 56414 -1542
rect 55794 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 56414 -1626
rect 55794 -1894 56414 -1862
rect 59514 673174 60134 707162
rect 59514 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 60134 673174
rect 59514 672854 60134 672938
rect 59514 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 60134 672854
rect 59514 637174 60134 672618
rect 59514 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 60134 637174
rect 59514 636854 60134 636938
rect 59514 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 60134 636854
rect 59514 601174 60134 636618
rect 59514 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 60134 601174
rect 59514 600854 60134 600938
rect 59514 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 60134 600854
rect 59514 565174 60134 600618
rect 59514 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 60134 565174
rect 59514 564854 60134 564938
rect 59514 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 60134 564854
rect 59514 529174 60134 564618
rect 59514 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 60134 529174
rect 59514 528854 60134 528938
rect 59514 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 60134 528854
rect 59514 493174 60134 528618
rect 59514 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 60134 493174
rect 59514 492854 60134 492938
rect 59514 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 60134 492854
rect 59514 457174 60134 492618
rect 59514 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 60134 457174
rect 59514 456854 60134 456938
rect 59514 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 60134 456854
rect 59514 421174 60134 456618
rect 59514 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 60134 421174
rect 59514 420854 60134 420938
rect 59514 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 60134 420854
rect 59514 385174 60134 420618
rect 59514 384938 59546 385174
rect 59782 384938 59866 385174
rect 60102 384938 60134 385174
rect 59514 384854 60134 384938
rect 59514 384618 59546 384854
rect 59782 384618 59866 384854
rect 60102 384618 60134 384854
rect 59514 349174 60134 384618
rect 59514 348938 59546 349174
rect 59782 348938 59866 349174
rect 60102 348938 60134 349174
rect 59514 348854 60134 348938
rect 59514 348618 59546 348854
rect 59782 348618 59866 348854
rect 60102 348618 60134 348854
rect 59514 313174 60134 348618
rect 59514 312938 59546 313174
rect 59782 312938 59866 313174
rect 60102 312938 60134 313174
rect 59514 312854 60134 312938
rect 59514 312618 59546 312854
rect 59782 312618 59866 312854
rect 60102 312618 60134 312854
rect 59514 277174 60134 312618
rect 59514 276938 59546 277174
rect 59782 276938 59866 277174
rect 60102 276938 60134 277174
rect 59514 276854 60134 276938
rect 59514 276618 59546 276854
rect 59782 276618 59866 276854
rect 60102 276618 60134 276854
rect 59514 241174 60134 276618
rect 59514 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 60134 241174
rect 59514 240854 60134 240938
rect 59514 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 60134 240854
rect 59514 205174 60134 240618
rect 59514 204938 59546 205174
rect 59782 204938 59866 205174
rect 60102 204938 60134 205174
rect 59514 204854 60134 204938
rect 59514 204618 59546 204854
rect 59782 204618 59866 204854
rect 60102 204618 60134 204854
rect 59514 169174 60134 204618
rect 59514 168938 59546 169174
rect 59782 168938 59866 169174
rect 60102 168938 60134 169174
rect 59514 168854 60134 168938
rect 59514 168618 59546 168854
rect 59782 168618 59866 168854
rect 60102 168618 60134 168854
rect 59514 133174 60134 168618
rect 59514 132938 59546 133174
rect 59782 132938 59866 133174
rect 60102 132938 60134 133174
rect 59514 132854 60134 132938
rect 59514 132618 59546 132854
rect 59782 132618 59866 132854
rect 60102 132618 60134 132854
rect 59514 97174 60134 132618
rect 59514 96938 59546 97174
rect 59782 96938 59866 97174
rect 60102 96938 60134 97174
rect 59514 96854 60134 96938
rect 59514 96618 59546 96854
rect 59782 96618 59866 96854
rect 60102 96618 60134 96854
rect 59514 61174 60134 96618
rect 59514 60938 59546 61174
rect 59782 60938 59866 61174
rect 60102 60938 60134 61174
rect 59514 60854 60134 60938
rect 59514 60618 59546 60854
rect 59782 60618 59866 60854
rect 60102 60618 60134 60854
rect 59514 25174 60134 60618
rect 59514 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 60134 25174
rect 59514 24854 60134 24938
rect 59514 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 60134 24854
rect 59514 -3226 60134 24618
rect 59514 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 60134 -3226
rect 59514 -3546 60134 -3462
rect 59514 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 60134 -3546
rect 59514 -3814 60134 -3782
rect 63234 676894 63854 709082
rect 63234 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 63854 676894
rect 63234 676574 63854 676658
rect 63234 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 63854 676574
rect 63234 640894 63854 676338
rect 63234 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 63854 640894
rect 63234 640574 63854 640658
rect 63234 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 63854 640574
rect 63234 604894 63854 640338
rect 63234 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 63854 604894
rect 63234 604574 63854 604658
rect 63234 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 63854 604574
rect 63234 568894 63854 604338
rect 63234 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 63854 568894
rect 63234 568574 63854 568658
rect 63234 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 63854 568574
rect 63234 532894 63854 568338
rect 63234 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 63854 532894
rect 63234 532574 63854 532658
rect 63234 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 63854 532574
rect 63234 496894 63854 532338
rect 63234 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 63854 496894
rect 63234 496574 63854 496658
rect 63234 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 63854 496574
rect 63234 460894 63854 496338
rect 63234 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 63854 460894
rect 63234 460574 63854 460658
rect 63234 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 63854 460574
rect 63234 424894 63854 460338
rect 63234 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 63854 424894
rect 63234 424574 63854 424658
rect 63234 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 63854 424574
rect 63234 388894 63854 424338
rect 63234 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 63854 388894
rect 63234 388574 63854 388658
rect 63234 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 63854 388574
rect 63234 352894 63854 388338
rect 63234 352658 63266 352894
rect 63502 352658 63586 352894
rect 63822 352658 63854 352894
rect 63234 352574 63854 352658
rect 63234 352338 63266 352574
rect 63502 352338 63586 352574
rect 63822 352338 63854 352574
rect 63234 316894 63854 352338
rect 63234 316658 63266 316894
rect 63502 316658 63586 316894
rect 63822 316658 63854 316894
rect 63234 316574 63854 316658
rect 63234 316338 63266 316574
rect 63502 316338 63586 316574
rect 63822 316338 63854 316574
rect 63234 280894 63854 316338
rect 63234 280658 63266 280894
rect 63502 280658 63586 280894
rect 63822 280658 63854 280894
rect 63234 280574 63854 280658
rect 63234 280338 63266 280574
rect 63502 280338 63586 280574
rect 63822 280338 63854 280574
rect 63234 244894 63854 280338
rect 63234 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 63854 244894
rect 63234 244574 63854 244658
rect 63234 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 63854 244574
rect 63234 208894 63854 244338
rect 63234 208658 63266 208894
rect 63502 208658 63586 208894
rect 63822 208658 63854 208894
rect 63234 208574 63854 208658
rect 63234 208338 63266 208574
rect 63502 208338 63586 208574
rect 63822 208338 63854 208574
rect 63234 172894 63854 208338
rect 63234 172658 63266 172894
rect 63502 172658 63586 172894
rect 63822 172658 63854 172894
rect 63234 172574 63854 172658
rect 63234 172338 63266 172574
rect 63502 172338 63586 172574
rect 63822 172338 63854 172574
rect 63234 136894 63854 172338
rect 63234 136658 63266 136894
rect 63502 136658 63586 136894
rect 63822 136658 63854 136894
rect 63234 136574 63854 136658
rect 63234 136338 63266 136574
rect 63502 136338 63586 136574
rect 63822 136338 63854 136574
rect 63234 100894 63854 136338
rect 63234 100658 63266 100894
rect 63502 100658 63586 100894
rect 63822 100658 63854 100894
rect 63234 100574 63854 100658
rect 63234 100338 63266 100574
rect 63502 100338 63586 100574
rect 63822 100338 63854 100574
rect 63234 64894 63854 100338
rect 63234 64658 63266 64894
rect 63502 64658 63586 64894
rect 63822 64658 63854 64894
rect 63234 64574 63854 64658
rect 63234 64338 63266 64574
rect 63502 64338 63586 64574
rect 63822 64338 63854 64574
rect 63234 28894 63854 64338
rect 63234 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 63854 28894
rect 63234 28574 63854 28658
rect 63234 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 63854 28574
rect 63234 -5146 63854 28338
rect 63234 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 63854 -5146
rect 63234 -5466 63854 -5382
rect 63234 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 63854 -5466
rect 63234 -5734 63854 -5702
rect 66954 680614 67574 711002
rect 84954 710598 85574 711590
rect 84954 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 85574 710598
rect 84954 710278 85574 710362
rect 84954 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 85574 710278
rect 81234 708678 81854 709670
rect 81234 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 81854 708678
rect 81234 708358 81854 708442
rect 81234 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 81854 708358
rect 77514 706758 78134 707750
rect 77514 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 78134 706758
rect 77514 706438 78134 706522
rect 77514 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 78134 706438
rect 66954 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 67574 680614
rect 66954 680294 67574 680378
rect 66954 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 67574 680294
rect 66954 644614 67574 680058
rect 66954 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 67574 644614
rect 66954 644294 67574 644378
rect 66954 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 67574 644294
rect 66954 608614 67574 644058
rect 66954 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 67574 608614
rect 66954 608294 67574 608378
rect 66954 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 67574 608294
rect 66954 572614 67574 608058
rect 66954 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 67574 572614
rect 66954 572294 67574 572378
rect 66954 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 67574 572294
rect 66954 536614 67574 572058
rect 66954 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 67574 536614
rect 66954 536294 67574 536378
rect 66954 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 67574 536294
rect 66954 500614 67574 536058
rect 66954 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 67574 500614
rect 66954 500294 67574 500378
rect 66954 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 67574 500294
rect 66954 464614 67574 500058
rect 66954 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 67574 464614
rect 66954 464294 67574 464378
rect 66954 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 67574 464294
rect 66954 428614 67574 464058
rect 66954 428378 66986 428614
rect 67222 428378 67306 428614
rect 67542 428378 67574 428614
rect 66954 428294 67574 428378
rect 66954 428058 66986 428294
rect 67222 428058 67306 428294
rect 67542 428058 67574 428294
rect 66954 392614 67574 428058
rect 66954 392378 66986 392614
rect 67222 392378 67306 392614
rect 67542 392378 67574 392614
rect 66954 392294 67574 392378
rect 66954 392058 66986 392294
rect 67222 392058 67306 392294
rect 67542 392058 67574 392294
rect 66954 356614 67574 392058
rect 66954 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 67574 356614
rect 66954 356294 67574 356378
rect 66954 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 67574 356294
rect 66954 320614 67574 356058
rect 66954 320378 66986 320614
rect 67222 320378 67306 320614
rect 67542 320378 67574 320614
rect 66954 320294 67574 320378
rect 66954 320058 66986 320294
rect 67222 320058 67306 320294
rect 67542 320058 67574 320294
rect 66954 284614 67574 320058
rect 66954 284378 66986 284614
rect 67222 284378 67306 284614
rect 67542 284378 67574 284614
rect 66954 284294 67574 284378
rect 66954 284058 66986 284294
rect 67222 284058 67306 284294
rect 67542 284058 67574 284294
rect 66954 248614 67574 284058
rect 66954 248378 66986 248614
rect 67222 248378 67306 248614
rect 67542 248378 67574 248614
rect 66954 248294 67574 248378
rect 66954 248058 66986 248294
rect 67222 248058 67306 248294
rect 67542 248058 67574 248294
rect 66954 212614 67574 248058
rect 66954 212378 66986 212614
rect 67222 212378 67306 212614
rect 67542 212378 67574 212614
rect 66954 212294 67574 212378
rect 66954 212058 66986 212294
rect 67222 212058 67306 212294
rect 67542 212058 67574 212294
rect 66954 176614 67574 212058
rect 66954 176378 66986 176614
rect 67222 176378 67306 176614
rect 67542 176378 67574 176614
rect 66954 176294 67574 176378
rect 66954 176058 66986 176294
rect 67222 176058 67306 176294
rect 67542 176058 67574 176294
rect 66954 140614 67574 176058
rect 66954 140378 66986 140614
rect 67222 140378 67306 140614
rect 67542 140378 67574 140614
rect 66954 140294 67574 140378
rect 66954 140058 66986 140294
rect 67222 140058 67306 140294
rect 67542 140058 67574 140294
rect 66954 104614 67574 140058
rect 66954 104378 66986 104614
rect 67222 104378 67306 104614
rect 67542 104378 67574 104614
rect 66954 104294 67574 104378
rect 66954 104058 66986 104294
rect 67222 104058 67306 104294
rect 67542 104058 67574 104294
rect 66954 68614 67574 104058
rect 66954 68378 66986 68614
rect 67222 68378 67306 68614
rect 67542 68378 67574 68614
rect 66954 68294 67574 68378
rect 66954 68058 66986 68294
rect 67222 68058 67306 68294
rect 67542 68058 67574 68294
rect 66954 32614 67574 68058
rect 66954 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 67574 32614
rect 66954 32294 67574 32378
rect 66954 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 67574 32294
rect 48954 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 49574 -6106
rect 48954 -6426 49574 -6342
rect 48954 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 49574 -6426
rect 48954 -7654 49574 -6662
rect 66954 -7066 67574 32058
rect 73794 704838 74414 705830
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 579454 74414 614898
rect 73794 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 74414 579454
rect 73794 579134 74414 579218
rect 73794 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 74414 579134
rect 73794 543454 74414 578898
rect 73794 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 74414 543454
rect 73794 543134 74414 543218
rect 73794 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 74414 543134
rect 73794 507454 74414 542898
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 471454 74414 506898
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73794 435454 74414 470898
rect 73794 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 74414 435454
rect 73794 435134 74414 435218
rect 73794 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 74414 435134
rect 73794 399454 74414 434898
rect 73794 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 74414 399454
rect 73794 399134 74414 399218
rect 73794 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 74414 399134
rect 73794 363454 74414 398898
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 73794 327454 74414 362898
rect 73794 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 74414 327454
rect 73794 327134 74414 327218
rect 73794 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 74414 327134
rect 73794 291454 74414 326898
rect 73794 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 74414 291454
rect 73794 291134 74414 291218
rect 73794 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 74414 291134
rect 73794 255454 74414 290898
rect 73794 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 74414 255454
rect 73794 255134 74414 255218
rect 73794 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 74414 255134
rect 73794 219454 74414 254898
rect 73794 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 74414 219454
rect 73794 219134 74414 219218
rect 73794 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 74414 219134
rect 73794 183454 74414 218898
rect 73794 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 74414 183454
rect 73794 183134 74414 183218
rect 73794 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 74414 183134
rect 73794 147454 74414 182898
rect 73794 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 74414 147454
rect 73794 147134 74414 147218
rect 73794 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 74414 147134
rect 73794 111454 74414 146898
rect 73794 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 74414 111454
rect 73794 111134 74414 111218
rect 73794 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 74414 111134
rect 73794 75454 74414 110898
rect 73794 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 74414 75454
rect 73794 75134 74414 75218
rect 73794 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 74414 75134
rect 73794 39454 74414 74898
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -1894 74414 -902
rect 77514 691174 78134 706202
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 655174 78134 690618
rect 77514 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 78134 655174
rect 77514 654854 78134 654938
rect 77514 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 78134 654854
rect 77514 619174 78134 654618
rect 77514 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 78134 619174
rect 77514 618854 78134 618938
rect 77514 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 78134 618854
rect 77514 583174 78134 618618
rect 77514 582938 77546 583174
rect 77782 582938 77866 583174
rect 78102 582938 78134 583174
rect 77514 582854 78134 582938
rect 77514 582618 77546 582854
rect 77782 582618 77866 582854
rect 78102 582618 78134 582854
rect 77514 547174 78134 582618
rect 77514 546938 77546 547174
rect 77782 546938 77866 547174
rect 78102 546938 78134 547174
rect 77514 546854 78134 546938
rect 77514 546618 77546 546854
rect 77782 546618 77866 546854
rect 78102 546618 78134 546854
rect 77514 511174 78134 546618
rect 77514 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 78134 511174
rect 77514 510854 78134 510938
rect 77514 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 78134 510854
rect 77514 475174 78134 510618
rect 77514 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 78134 475174
rect 77514 474854 78134 474938
rect 77514 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 78134 474854
rect 77514 439174 78134 474618
rect 77514 438938 77546 439174
rect 77782 438938 77866 439174
rect 78102 438938 78134 439174
rect 77514 438854 78134 438938
rect 77514 438618 77546 438854
rect 77782 438618 77866 438854
rect 78102 438618 78134 438854
rect 77514 403174 78134 438618
rect 77514 402938 77546 403174
rect 77782 402938 77866 403174
rect 78102 402938 78134 403174
rect 77514 402854 78134 402938
rect 77514 402618 77546 402854
rect 77782 402618 77866 402854
rect 78102 402618 78134 402854
rect 77514 367174 78134 402618
rect 77514 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 78134 367174
rect 77514 366854 78134 366938
rect 77514 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 78134 366854
rect 77514 331174 78134 366618
rect 77514 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 78134 331174
rect 77514 330854 78134 330938
rect 77514 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 78134 330854
rect 77514 295174 78134 330618
rect 77514 294938 77546 295174
rect 77782 294938 77866 295174
rect 78102 294938 78134 295174
rect 77514 294854 78134 294938
rect 77514 294618 77546 294854
rect 77782 294618 77866 294854
rect 78102 294618 78134 294854
rect 77514 259174 78134 294618
rect 77514 258938 77546 259174
rect 77782 258938 77866 259174
rect 78102 258938 78134 259174
rect 77514 258854 78134 258938
rect 77514 258618 77546 258854
rect 77782 258618 77866 258854
rect 78102 258618 78134 258854
rect 77514 223174 78134 258618
rect 77514 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 78134 223174
rect 77514 222854 78134 222938
rect 77514 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 78134 222854
rect 77514 187174 78134 222618
rect 77514 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 78134 187174
rect 77514 186854 78134 186938
rect 77514 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 78134 186854
rect 77514 151174 78134 186618
rect 77514 150938 77546 151174
rect 77782 150938 77866 151174
rect 78102 150938 78134 151174
rect 77514 150854 78134 150938
rect 77514 150618 77546 150854
rect 77782 150618 77866 150854
rect 78102 150618 78134 150854
rect 77514 115174 78134 150618
rect 77514 114938 77546 115174
rect 77782 114938 77866 115174
rect 78102 114938 78134 115174
rect 77514 114854 78134 114938
rect 77514 114618 77546 114854
rect 77782 114618 77866 114854
rect 78102 114618 78134 114854
rect 77514 79174 78134 114618
rect 77514 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 78134 79174
rect 77514 78854 78134 78938
rect 77514 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 78134 78854
rect 77514 43174 78134 78618
rect 77514 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 78134 43174
rect 77514 42854 78134 42938
rect 77514 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 78134 42854
rect 77514 7174 78134 42618
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 77514 -2266 78134 6618
rect 77514 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 78134 -2266
rect 77514 -2586 78134 -2502
rect 77514 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 78134 -2586
rect 77514 -3814 78134 -2822
rect 81234 694894 81854 708122
rect 81234 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 81854 694894
rect 81234 694574 81854 694658
rect 81234 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 81854 694574
rect 81234 658894 81854 694338
rect 81234 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 81854 658894
rect 81234 658574 81854 658658
rect 81234 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 81854 658574
rect 81234 622894 81854 658338
rect 81234 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 81854 622894
rect 81234 622574 81854 622658
rect 81234 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 81854 622574
rect 81234 586894 81854 622338
rect 81234 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 81854 586894
rect 81234 586574 81854 586658
rect 81234 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 81854 586574
rect 81234 550894 81854 586338
rect 81234 550658 81266 550894
rect 81502 550658 81586 550894
rect 81822 550658 81854 550894
rect 81234 550574 81854 550658
rect 81234 550338 81266 550574
rect 81502 550338 81586 550574
rect 81822 550338 81854 550574
rect 81234 514894 81854 550338
rect 81234 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 81854 514894
rect 81234 514574 81854 514658
rect 81234 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 81854 514574
rect 81234 478894 81854 514338
rect 81234 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 81854 478894
rect 81234 478574 81854 478658
rect 81234 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 81854 478574
rect 81234 442894 81854 478338
rect 81234 442658 81266 442894
rect 81502 442658 81586 442894
rect 81822 442658 81854 442894
rect 81234 442574 81854 442658
rect 81234 442338 81266 442574
rect 81502 442338 81586 442574
rect 81822 442338 81854 442574
rect 81234 406894 81854 442338
rect 81234 406658 81266 406894
rect 81502 406658 81586 406894
rect 81822 406658 81854 406894
rect 81234 406574 81854 406658
rect 81234 406338 81266 406574
rect 81502 406338 81586 406574
rect 81822 406338 81854 406574
rect 81234 370894 81854 406338
rect 81234 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 81854 370894
rect 81234 370574 81854 370658
rect 81234 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 81854 370574
rect 81234 334894 81854 370338
rect 81234 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 81854 334894
rect 81234 334574 81854 334658
rect 81234 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 81854 334574
rect 81234 298894 81854 334338
rect 81234 298658 81266 298894
rect 81502 298658 81586 298894
rect 81822 298658 81854 298894
rect 81234 298574 81854 298658
rect 81234 298338 81266 298574
rect 81502 298338 81586 298574
rect 81822 298338 81854 298574
rect 81234 262894 81854 298338
rect 81234 262658 81266 262894
rect 81502 262658 81586 262894
rect 81822 262658 81854 262894
rect 81234 262574 81854 262658
rect 81234 262338 81266 262574
rect 81502 262338 81586 262574
rect 81822 262338 81854 262574
rect 81234 226894 81854 262338
rect 81234 226658 81266 226894
rect 81502 226658 81586 226894
rect 81822 226658 81854 226894
rect 81234 226574 81854 226658
rect 81234 226338 81266 226574
rect 81502 226338 81586 226574
rect 81822 226338 81854 226574
rect 81234 190894 81854 226338
rect 81234 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 81854 190894
rect 81234 190574 81854 190658
rect 81234 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 81854 190574
rect 81234 154894 81854 190338
rect 81234 154658 81266 154894
rect 81502 154658 81586 154894
rect 81822 154658 81854 154894
rect 81234 154574 81854 154658
rect 81234 154338 81266 154574
rect 81502 154338 81586 154574
rect 81822 154338 81854 154574
rect 81234 118894 81854 154338
rect 81234 118658 81266 118894
rect 81502 118658 81586 118894
rect 81822 118658 81854 118894
rect 81234 118574 81854 118658
rect 81234 118338 81266 118574
rect 81502 118338 81586 118574
rect 81822 118338 81854 118574
rect 81234 82894 81854 118338
rect 81234 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 81854 82894
rect 81234 82574 81854 82658
rect 81234 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 81854 82574
rect 81234 46894 81854 82338
rect 81234 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 81854 46894
rect 81234 46574 81854 46658
rect 81234 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 81854 46574
rect 81234 10894 81854 46338
rect 81234 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 81854 10894
rect 81234 10574 81854 10658
rect 81234 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 81854 10574
rect 81234 -4186 81854 10338
rect 81234 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 81854 -4186
rect 81234 -4506 81854 -4422
rect 81234 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 81854 -4506
rect 81234 -5734 81854 -4742
rect 84954 698614 85574 710042
rect 102954 711558 103574 711590
rect 102954 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 103574 711558
rect 102954 711238 103574 711322
rect 102954 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 103574 711238
rect 99234 709638 99854 709670
rect 99234 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 99854 709638
rect 99234 709318 99854 709402
rect 99234 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 99854 709318
rect 95514 707718 96134 707750
rect 95514 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 96134 707718
rect 95514 707398 96134 707482
rect 95514 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 96134 707398
rect 84954 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 85574 698614
rect 84954 698294 85574 698378
rect 84954 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 85574 698294
rect 84954 662614 85574 698058
rect 84954 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 85574 662614
rect 84954 662294 85574 662378
rect 84954 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 85574 662294
rect 84954 626614 85574 662058
rect 84954 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 85574 626614
rect 84954 626294 85574 626378
rect 84954 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 85574 626294
rect 84954 590614 85574 626058
rect 84954 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 85574 590614
rect 84954 590294 85574 590378
rect 84954 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 85574 590294
rect 84954 554614 85574 590058
rect 84954 554378 84986 554614
rect 85222 554378 85306 554614
rect 85542 554378 85574 554614
rect 84954 554294 85574 554378
rect 84954 554058 84986 554294
rect 85222 554058 85306 554294
rect 85542 554058 85574 554294
rect 84954 518614 85574 554058
rect 84954 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 85574 518614
rect 84954 518294 85574 518378
rect 84954 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 85574 518294
rect 84954 482614 85574 518058
rect 84954 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 85574 482614
rect 84954 482294 85574 482378
rect 84954 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 85574 482294
rect 84954 446614 85574 482058
rect 84954 446378 84986 446614
rect 85222 446378 85306 446614
rect 85542 446378 85574 446614
rect 84954 446294 85574 446378
rect 84954 446058 84986 446294
rect 85222 446058 85306 446294
rect 85542 446058 85574 446294
rect 84954 410614 85574 446058
rect 84954 410378 84986 410614
rect 85222 410378 85306 410614
rect 85542 410378 85574 410614
rect 84954 410294 85574 410378
rect 84954 410058 84986 410294
rect 85222 410058 85306 410294
rect 85542 410058 85574 410294
rect 84954 374614 85574 410058
rect 84954 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 85574 374614
rect 84954 374294 85574 374378
rect 84954 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 85574 374294
rect 84954 338614 85574 374058
rect 84954 338378 84986 338614
rect 85222 338378 85306 338614
rect 85542 338378 85574 338614
rect 84954 338294 85574 338378
rect 84954 338058 84986 338294
rect 85222 338058 85306 338294
rect 85542 338058 85574 338294
rect 84954 302614 85574 338058
rect 84954 302378 84986 302614
rect 85222 302378 85306 302614
rect 85542 302378 85574 302614
rect 84954 302294 85574 302378
rect 84954 302058 84986 302294
rect 85222 302058 85306 302294
rect 85542 302058 85574 302294
rect 84954 266614 85574 302058
rect 84954 266378 84986 266614
rect 85222 266378 85306 266614
rect 85542 266378 85574 266614
rect 84954 266294 85574 266378
rect 84954 266058 84986 266294
rect 85222 266058 85306 266294
rect 85542 266058 85574 266294
rect 84954 230614 85574 266058
rect 84954 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 85574 230614
rect 84954 230294 85574 230378
rect 84954 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 85574 230294
rect 84954 194614 85574 230058
rect 84954 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 85574 194614
rect 84954 194294 85574 194378
rect 84954 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 85574 194294
rect 84954 158614 85574 194058
rect 84954 158378 84986 158614
rect 85222 158378 85306 158614
rect 85542 158378 85574 158614
rect 84954 158294 85574 158378
rect 84954 158058 84986 158294
rect 85222 158058 85306 158294
rect 85542 158058 85574 158294
rect 84954 122614 85574 158058
rect 84954 122378 84986 122614
rect 85222 122378 85306 122614
rect 85542 122378 85574 122614
rect 84954 122294 85574 122378
rect 84954 122058 84986 122294
rect 85222 122058 85306 122294
rect 85542 122058 85574 122294
rect 84954 86614 85574 122058
rect 84954 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 85574 86614
rect 84954 86294 85574 86378
rect 84954 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 85574 86294
rect 84954 50614 85574 86058
rect 84954 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 85574 50614
rect 84954 50294 85574 50378
rect 84954 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 85574 50294
rect 84954 14614 85574 50058
rect 84954 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 85574 14614
rect 84954 14294 85574 14378
rect 84954 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 85574 14294
rect 66954 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 67574 -7066
rect 66954 -7386 67574 -7302
rect 66954 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 67574 -7386
rect 66954 -7654 67574 -7622
rect 84954 -6106 85574 14058
rect 91794 705798 92414 705830
rect 91794 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 92414 705798
rect 91794 705478 92414 705562
rect 91794 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 92414 705478
rect 91794 669454 92414 705242
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 91794 561454 92414 596898
rect 91794 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 92414 561454
rect 91794 561134 92414 561218
rect 91794 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 92414 561134
rect 91794 525454 92414 560898
rect 91794 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 92414 525454
rect 91794 525134 92414 525218
rect 91794 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 92414 525134
rect 91794 489454 92414 524898
rect 91794 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 92414 489454
rect 91794 489134 92414 489218
rect 91794 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 92414 489134
rect 91794 453454 92414 488898
rect 91794 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 92414 453454
rect 91794 453134 92414 453218
rect 91794 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 92414 453134
rect 91794 417454 92414 452898
rect 91794 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 92414 417454
rect 91794 417134 92414 417218
rect 91794 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 92414 417134
rect 91794 381454 92414 416898
rect 91794 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 92414 381454
rect 91794 381134 92414 381218
rect 91794 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 92414 381134
rect 91794 345454 92414 380898
rect 91794 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 92414 345454
rect 91794 345134 92414 345218
rect 91794 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 92414 345134
rect 91794 309454 92414 344898
rect 91794 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 92414 309454
rect 91794 309134 92414 309218
rect 91794 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 92414 309134
rect 91794 273454 92414 308898
rect 91794 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 92414 273454
rect 91794 273134 92414 273218
rect 91794 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 92414 273134
rect 91794 237454 92414 272898
rect 91794 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 92414 237454
rect 91794 237134 92414 237218
rect 91794 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 92414 237134
rect 91794 201454 92414 236898
rect 91794 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 92414 201454
rect 91794 201134 92414 201218
rect 91794 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 92414 201134
rect 91794 165454 92414 200898
rect 91794 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 92414 165454
rect 91794 165134 92414 165218
rect 91794 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 92414 165134
rect 91794 129454 92414 164898
rect 91794 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 92414 129454
rect 91794 129134 92414 129218
rect 91794 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 92414 129134
rect 91794 93454 92414 128898
rect 91794 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 92414 93454
rect 91794 93134 92414 93218
rect 91794 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 92414 93134
rect 91794 57454 92414 92898
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -1306 92414 20898
rect 91794 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 92414 -1306
rect 91794 -1626 92414 -1542
rect 91794 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 92414 -1626
rect 91794 -1894 92414 -1862
rect 95514 673174 96134 707162
rect 95514 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 96134 673174
rect 95514 672854 96134 672938
rect 95514 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 96134 672854
rect 95514 637174 96134 672618
rect 95514 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 96134 637174
rect 95514 636854 96134 636938
rect 95514 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 96134 636854
rect 95514 601174 96134 636618
rect 95514 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 96134 601174
rect 95514 600854 96134 600938
rect 95514 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 96134 600854
rect 95514 565174 96134 600618
rect 95514 564938 95546 565174
rect 95782 564938 95866 565174
rect 96102 564938 96134 565174
rect 95514 564854 96134 564938
rect 95514 564618 95546 564854
rect 95782 564618 95866 564854
rect 96102 564618 96134 564854
rect 95514 529174 96134 564618
rect 95514 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 96134 529174
rect 95514 528854 96134 528938
rect 95514 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 96134 528854
rect 95514 493174 96134 528618
rect 95514 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 96134 493174
rect 95514 492854 96134 492938
rect 95514 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 96134 492854
rect 95514 457174 96134 492618
rect 95514 456938 95546 457174
rect 95782 456938 95866 457174
rect 96102 456938 96134 457174
rect 95514 456854 96134 456938
rect 95514 456618 95546 456854
rect 95782 456618 95866 456854
rect 96102 456618 96134 456854
rect 95514 421174 96134 456618
rect 95514 420938 95546 421174
rect 95782 420938 95866 421174
rect 96102 420938 96134 421174
rect 95514 420854 96134 420938
rect 95514 420618 95546 420854
rect 95782 420618 95866 420854
rect 96102 420618 96134 420854
rect 95514 385174 96134 420618
rect 95514 384938 95546 385174
rect 95782 384938 95866 385174
rect 96102 384938 96134 385174
rect 95514 384854 96134 384938
rect 95514 384618 95546 384854
rect 95782 384618 95866 384854
rect 96102 384618 96134 384854
rect 95514 349174 96134 384618
rect 95514 348938 95546 349174
rect 95782 348938 95866 349174
rect 96102 348938 96134 349174
rect 95514 348854 96134 348938
rect 95514 348618 95546 348854
rect 95782 348618 95866 348854
rect 96102 348618 96134 348854
rect 95514 313174 96134 348618
rect 95514 312938 95546 313174
rect 95782 312938 95866 313174
rect 96102 312938 96134 313174
rect 95514 312854 96134 312938
rect 95514 312618 95546 312854
rect 95782 312618 95866 312854
rect 96102 312618 96134 312854
rect 95514 277174 96134 312618
rect 95514 276938 95546 277174
rect 95782 276938 95866 277174
rect 96102 276938 96134 277174
rect 95514 276854 96134 276938
rect 95514 276618 95546 276854
rect 95782 276618 95866 276854
rect 96102 276618 96134 276854
rect 95514 241174 96134 276618
rect 95514 240938 95546 241174
rect 95782 240938 95866 241174
rect 96102 240938 96134 241174
rect 95514 240854 96134 240938
rect 95514 240618 95546 240854
rect 95782 240618 95866 240854
rect 96102 240618 96134 240854
rect 95514 205174 96134 240618
rect 95514 204938 95546 205174
rect 95782 204938 95866 205174
rect 96102 204938 96134 205174
rect 95514 204854 96134 204938
rect 95514 204618 95546 204854
rect 95782 204618 95866 204854
rect 96102 204618 96134 204854
rect 95514 169174 96134 204618
rect 95514 168938 95546 169174
rect 95782 168938 95866 169174
rect 96102 168938 96134 169174
rect 95514 168854 96134 168938
rect 95514 168618 95546 168854
rect 95782 168618 95866 168854
rect 96102 168618 96134 168854
rect 95514 133174 96134 168618
rect 95514 132938 95546 133174
rect 95782 132938 95866 133174
rect 96102 132938 96134 133174
rect 95514 132854 96134 132938
rect 95514 132618 95546 132854
rect 95782 132618 95866 132854
rect 96102 132618 96134 132854
rect 95514 97174 96134 132618
rect 95514 96938 95546 97174
rect 95782 96938 95866 97174
rect 96102 96938 96134 97174
rect 95514 96854 96134 96938
rect 95514 96618 95546 96854
rect 95782 96618 95866 96854
rect 96102 96618 96134 96854
rect 95514 61174 96134 96618
rect 95514 60938 95546 61174
rect 95782 60938 95866 61174
rect 96102 60938 96134 61174
rect 95514 60854 96134 60938
rect 95514 60618 95546 60854
rect 95782 60618 95866 60854
rect 96102 60618 96134 60854
rect 95514 25174 96134 60618
rect 95514 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 96134 25174
rect 95514 24854 96134 24938
rect 95514 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 96134 24854
rect 95514 -3226 96134 24618
rect 95514 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 96134 -3226
rect 95514 -3546 96134 -3462
rect 95514 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 96134 -3546
rect 95514 -3814 96134 -3782
rect 99234 676894 99854 709082
rect 99234 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 99854 676894
rect 99234 676574 99854 676658
rect 99234 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 99854 676574
rect 99234 640894 99854 676338
rect 99234 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 99854 640894
rect 99234 640574 99854 640658
rect 99234 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 99854 640574
rect 99234 604894 99854 640338
rect 99234 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 99854 604894
rect 99234 604574 99854 604658
rect 99234 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 99854 604574
rect 99234 568894 99854 604338
rect 99234 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 99854 568894
rect 99234 568574 99854 568658
rect 99234 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 99854 568574
rect 99234 532894 99854 568338
rect 99234 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 99854 532894
rect 99234 532574 99854 532658
rect 99234 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 99854 532574
rect 99234 496894 99854 532338
rect 99234 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 99854 496894
rect 99234 496574 99854 496658
rect 99234 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 99854 496574
rect 99234 460894 99854 496338
rect 99234 460658 99266 460894
rect 99502 460658 99586 460894
rect 99822 460658 99854 460894
rect 99234 460574 99854 460658
rect 99234 460338 99266 460574
rect 99502 460338 99586 460574
rect 99822 460338 99854 460574
rect 99234 424894 99854 460338
rect 99234 424658 99266 424894
rect 99502 424658 99586 424894
rect 99822 424658 99854 424894
rect 99234 424574 99854 424658
rect 99234 424338 99266 424574
rect 99502 424338 99586 424574
rect 99822 424338 99854 424574
rect 99234 388894 99854 424338
rect 99234 388658 99266 388894
rect 99502 388658 99586 388894
rect 99822 388658 99854 388894
rect 99234 388574 99854 388658
rect 99234 388338 99266 388574
rect 99502 388338 99586 388574
rect 99822 388338 99854 388574
rect 99234 352894 99854 388338
rect 99234 352658 99266 352894
rect 99502 352658 99586 352894
rect 99822 352658 99854 352894
rect 99234 352574 99854 352658
rect 99234 352338 99266 352574
rect 99502 352338 99586 352574
rect 99822 352338 99854 352574
rect 99234 316894 99854 352338
rect 99234 316658 99266 316894
rect 99502 316658 99586 316894
rect 99822 316658 99854 316894
rect 99234 316574 99854 316658
rect 99234 316338 99266 316574
rect 99502 316338 99586 316574
rect 99822 316338 99854 316574
rect 99234 280894 99854 316338
rect 99234 280658 99266 280894
rect 99502 280658 99586 280894
rect 99822 280658 99854 280894
rect 99234 280574 99854 280658
rect 99234 280338 99266 280574
rect 99502 280338 99586 280574
rect 99822 280338 99854 280574
rect 99234 244894 99854 280338
rect 99234 244658 99266 244894
rect 99502 244658 99586 244894
rect 99822 244658 99854 244894
rect 99234 244574 99854 244658
rect 99234 244338 99266 244574
rect 99502 244338 99586 244574
rect 99822 244338 99854 244574
rect 99234 208894 99854 244338
rect 99234 208658 99266 208894
rect 99502 208658 99586 208894
rect 99822 208658 99854 208894
rect 99234 208574 99854 208658
rect 99234 208338 99266 208574
rect 99502 208338 99586 208574
rect 99822 208338 99854 208574
rect 99234 172894 99854 208338
rect 99234 172658 99266 172894
rect 99502 172658 99586 172894
rect 99822 172658 99854 172894
rect 99234 172574 99854 172658
rect 99234 172338 99266 172574
rect 99502 172338 99586 172574
rect 99822 172338 99854 172574
rect 99234 136894 99854 172338
rect 99234 136658 99266 136894
rect 99502 136658 99586 136894
rect 99822 136658 99854 136894
rect 99234 136574 99854 136658
rect 99234 136338 99266 136574
rect 99502 136338 99586 136574
rect 99822 136338 99854 136574
rect 99234 100894 99854 136338
rect 99234 100658 99266 100894
rect 99502 100658 99586 100894
rect 99822 100658 99854 100894
rect 99234 100574 99854 100658
rect 99234 100338 99266 100574
rect 99502 100338 99586 100574
rect 99822 100338 99854 100574
rect 99234 64894 99854 100338
rect 99234 64658 99266 64894
rect 99502 64658 99586 64894
rect 99822 64658 99854 64894
rect 99234 64574 99854 64658
rect 99234 64338 99266 64574
rect 99502 64338 99586 64574
rect 99822 64338 99854 64574
rect 99234 28894 99854 64338
rect 99234 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 99854 28894
rect 99234 28574 99854 28658
rect 99234 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 99854 28574
rect 99234 -5146 99854 28338
rect 99234 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 99854 -5146
rect 99234 -5466 99854 -5382
rect 99234 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 99854 -5466
rect 99234 -5734 99854 -5702
rect 102954 680614 103574 711002
rect 120954 710598 121574 711590
rect 120954 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 121574 710598
rect 120954 710278 121574 710362
rect 120954 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 121574 710278
rect 117234 708678 117854 709670
rect 117234 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 117854 708678
rect 117234 708358 117854 708442
rect 117234 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 117854 708358
rect 113514 706758 114134 707750
rect 113514 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 114134 706758
rect 113514 706438 114134 706522
rect 113514 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 114134 706438
rect 102954 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 103574 680614
rect 102954 680294 103574 680378
rect 102954 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 103574 680294
rect 102954 644614 103574 680058
rect 102954 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 103574 644614
rect 102954 644294 103574 644378
rect 102954 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 103574 644294
rect 102954 608614 103574 644058
rect 102954 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 103574 608614
rect 102954 608294 103574 608378
rect 102954 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 103574 608294
rect 102954 572614 103574 608058
rect 102954 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 103574 572614
rect 102954 572294 103574 572378
rect 102954 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 103574 572294
rect 102954 536614 103574 572058
rect 102954 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 103574 536614
rect 102954 536294 103574 536378
rect 102954 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 103574 536294
rect 102954 500614 103574 536058
rect 102954 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 103574 500614
rect 102954 500294 103574 500378
rect 102954 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 103574 500294
rect 102954 464614 103574 500058
rect 102954 464378 102986 464614
rect 103222 464378 103306 464614
rect 103542 464378 103574 464614
rect 102954 464294 103574 464378
rect 102954 464058 102986 464294
rect 103222 464058 103306 464294
rect 103542 464058 103574 464294
rect 102954 428614 103574 464058
rect 102954 428378 102986 428614
rect 103222 428378 103306 428614
rect 103542 428378 103574 428614
rect 102954 428294 103574 428378
rect 102954 428058 102986 428294
rect 103222 428058 103306 428294
rect 103542 428058 103574 428294
rect 102954 392614 103574 428058
rect 102954 392378 102986 392614
rect 103222 392378 103306 392614
rect 103542 392378 103574 392614
rect 102954 392294 103574 392378
rect 102954 392058 102986 392294
rect 103222 392058 103306 392294
rect 103542 392058 103574 392294
rect 102954 356614 103574 392058
rect 102954 356378 102986 356614
rect 103222 356378 103306 356614
rect 103542 356378 103574 356614
rect 102954 356294 103574 356378
rect 102954 356058 102986 356294
rect 103222 356058 103306 356294
rect 103542 356058 103574 356294
rect 102954 320614 103574 356058
rect 102954 320378 102986 320614
rect 103222 320378 103306 320614
rect 103542 320378 103574 320614
rect 102954 320294 103574 320378
rect 102954 320058 102986 320294
rect 103222 320058 103306 320294
rect 103542 320058 103574 320294
rect 102954 284614 103574 320058
rect 102954 284378 102986 284614
rect 103222 284378 103306 284614
rect 103542 284378 103574 284614
rect 102954 284294 103574 284378
rect 102954 284058 102986 284294
rect 103222 284058 103306 284294
rect 103542 284058 103574 284294
rect 102954 248614 103574 284058
rect 102954 248378 102986 248614
rect 103222 248378 103306 248614
rect 103542 248378 103574 248614
rect 102954 248294 103574 248378
rect 102954 248058 102986 248294
rect 103222 248058 103306 248294
rect 103542 248058 103574 248294
rect 102954 212614 103574 248058
rect 102954 212378 102986 212614
rect 103222 212378 103306 212614
rect 103542 212378 103574 212614
rect 102954 212294 103574 212378
rect 102954 212058 102986 212294
rect 103222 212058 103306 212294
rect 103542 212058 103574 212294
rect 102954 176614 103574 212058
rect 102954 176378 102986 176614
rect 103222 176378 103306 176614
rect 103542 176378 103574 176614
rect 102954 176294 103574 176378
rect 102954 176058 102986 176294
rect 103222 176058 103306 176294
rect 103542 176058 103574 176294
rect 102954 140614 103574 176058
rect 102954 140378 102986 140614
rect 103222 140378 103306 140614
rect 103542 140378 103574 140614
rect 102954 140294 103574 140378
rect 102954 140058 102986 140294
rect 103222 140058 103306 140294
rect 103542 140058 103574 140294
rect 102954 104614 103574 140058
rect 102954 104378 102986 104614
rect 103222 104378 103306 104614
rect 103542 104378 103574 104614
rect 102954 104294 103574 104378
rect 102954 104058 102986 104294
rect 103222 104058 103306 104294
rect 103542 104058 103574 104294
rect 102954 68614 103574 104058
rect 102954 68378 102986 68614
rect 103222 68378 103306 68614
rect 103542 68378 103574 68614
rect 102954 68294 103574 68378
rect 102954 68058 102986 68294
rect 103222 68058 103306 68294
rect 103542 68058 103574 68294
rect 102954 32614 103574 68058
rect 102954 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 103574 32614
rect 102954 32294 103574 32378
rect 102954 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 103574 32294
rect 84954 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 85574 -6106
rect 84954 -6426 85574 -6342
rect 84954 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 85574 -6426
rect 84954 -7654 85574 -6662
rect 102954 -7066 103574 32058
rect 109794 704838 110414 705830
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 109794 543454 110414 578898
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 109794 507454 110414 542898
rect 109794 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 110414 507454
rect 109794 507134 110414 507218
rect 109794 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 110414 507134
rect 109794 471454 110414 506898
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 109794 435454 110414 470898
rect 109794 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 110414 435454
rect 109794 435134 110414 435218
rect 109794 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 110414 435134
rect 109794 399454 110414 434898
rect 109794 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 110414 399454
rect 109794 399134 110414 399218
rect 109794 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 110414 399134
rect 109794 363454 110414 398898
rect 109794 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 110414 363454
rect 109794 363134 110414 363218
rect 109794 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 110414 363134
rect 109794 327454 110414 362898
rect 109794 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 110414 327454
rect 109794 327134 110414 327218
rect 109794 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 110414 327134
rect 109794 291454 110414 326898
rect 109794 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 110414 291454
rect 109794 291134 110414 291218
rect 109794 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 110414 291134
rect 109794 255454 110414 290898
rect 109794 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 110414 255454
rect 109794 255134 110414 255218
rect 109794 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 110414 255134
rect 109794 219454 110414 254898
rect 109794 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 110414 219454
rect 109794 219134 110414 219218
rect 109794 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 110414 219134
rect 109794 183454 110414 218898
rect 109794 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 110414 183454
rect 109794 183134 110414 183218
rect 109794 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 110414 183134
rect 109794 147454 110414 182898
rect 109794 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 110414 147454
rect 109794 147134 110414 147218
rect 109794 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 110414 147134
rect 109794 111454 110414 146898
rect 109794 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 110414 111454
rect 109794 111134 110414 111218
rect 109794 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 110414 111134
rect 109794 75454 110414 110898
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 109794 75134 110414 75218
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 109794 39454 110414 74898
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -1894 110414 -902
rect 113514 691174 114134 706202
rect 113514 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 114134 691174
rect 113514 690854 114134 690938
rect 113514 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 114134 690854
rect 113514 655174 114134 690618
rect 113514 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 114134 655174
rect 113514 654854 114134 654938
rect 113514 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 114134 654854
rect 113514 619174 114134 654618
rect 113514 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 114134 619174
rect 113514 618854 114134 618938
rect 113514 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 114134 618854
rect 113514 583174 114134 618618
rect 113514 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 114134 583174
rect 113514 582854 114134 582938
rect 113514 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 114134 582854
rect 113514 547174 114134 582618
rect 113514 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 114134 547174
rect 113514 546854 114134 546938
rect 113514 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 114134 546854
rect 113514 511174 114134 546618
rect 113514 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 114134 511174
rect 113514 510854 114134 510938
rect 113514 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 114134 510854
rect 113514 475174 114134 510618
rect 113514 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 114134 475174
rect 113514 474854 114134 474938
rect 113514 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 114134 474854
rect 113514 439174 114134 474618
rect 113514 438938 113546 439174
rect 113782 438938 113866 439174
rect 114102 438938 114134 439174
rect 113514 438854 114134 438938
rect 113514 438618 113546 438854
rect 113782 438618 113866 438854
rect 114102 438618 114134 438854
rect 113514 403174 114134 438618
rect 113514 402938 113546 403174
rect 113782 402938 113866 403174
rect 114102 402938 114134 403174
rect 113514 402854 114134 402938
rect 113514 402618 113546 402854
rect 113782 402618 113866 402854
rect 114102 402618 114134 402854
rect 113514 367174 114134 402618
rect 113514 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 114134 367174
rect 113514 366854 114134 366938
rect 113514 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 114134 366854
rect 113514 331174 114134 366618
rect 113514 330938 113546 331174
rect 113782 330938 113866 331174
rect 114102 330938 114134 331174
rect 113514 330854 114134 330938
rect 113514 330618 113546 330854
rect 113782 330618 113866 330854
rect 114102 330618 114134 330854
rect 113514 295174 114134 330618
rect 113514 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 114134 295174
rect 113514 294854 114134 294938
rect 113514 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 114134 294854
rect 113514 259174 114134 294618
rect 113514 258938 113546 259174
rect 113782 258938 113866 259174
rect 114102 258938 114134 259174
rect 113514 258854 114134 258938
rect 113514 258618 113546 258854
rect 113782 258618 113866 258854
rect 114102 258618 114134 258854
rect 113514 223174 114134 258618
rect 113514 222938 113546 223174
rect 113782 222938 113866 223174
rect 114102 222938 114134 223174
rect 113514 222854 114134 222938
rect 113514 222618 113546 222854
rect 113782 222618 113866 222854
rect 114102 222618 114134 222854
rect 113514 187174 114134 222618
rect 113514 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 114134 187174
rect 113514 186854 114134 186938
rect 113514 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 114134 186854
rect 113514 151174 114134 186618
rect 113514 150938 113546 151174
rect 113782 150938 113866 151174
rect 114102 150938 114134 151174
rect 113514 150854 114134 150938
rect 113514 150618 113546 150854
rect 113782 150618 113866 150854
rect 114102 150618 114134 150854
rect 113514 115174 114134 150618
rect 113514 114938 113546 115174
rect 113782 114938 113866 115174
rect 114102 114938 114134 115174
rect 113514 114854 114134 114938
rect 113514 114618 113546 114854
rect 113782 114618 113866 114854
rect 114102 114618 114134 114854
rect 113514 79174 114134 114618
rect 113514 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 114134 79174
rect 113514 78854 114134 78938
rect 113514 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 114134 78854
rect 113514 43174 114134 78618
rect 113514 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 114134 43174
rect 113514 42854 114134 42938
rect 113514 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 114134 42854
rect 113514 7174 114134 42618
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 113514 -2266 114134 6618
rect 113514 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 114134 -2266
rect 113514 -2586 114134 -2502
rect 113514 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 114134 -2586
rect 113514 -3814 114134 -2822
rect 117234 694894 117854 708122
rect 117234 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 117854 694894
rect 117234 694574 117854 694658
rect 117234 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 117854 694574
rect 117234 658894 117854 694338
rect 117234 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 117854 658894
rect 117234 658574 117854 658658
rect 117234 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 117854 658574
rect 117234 622894 117854 658338
rect 117234 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 117854 622894
rect 117234 622574 117854 622658
rect 117234 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 117854 622574
rect 117234 586894 117854 622338
rect 117234 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 117854 586894
rect 117234 586574 117854 586658
rect 117234 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 117854 586574
rect 117234 550894 117854 586338
rect 117234 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 117854 550894
rect 117234 550574 117854 550658
rect 117234 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 117854 550574
rect 117234 514894 117854 550338
rect 117234 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 117854 514894
rect 117234 514574 117854 514658
rect 117234 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 117854 514574
rect 117234 478894 117854 514338
rect 117234 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 117854 478894
rect 117234 478574 117854 478658
rect 117234 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 117854 478574
rect 117234 442894 117854 478338
rect 117234 442658 117266 442894
rect 117502 442658 117586 442894
rect 117822 442658 117854 442894
rect 117234 442574 117854 442658
rect 117234 442338 117266 442574
rect 117502 442338 117586 442574
rect 117822 442338 117854 442574
rect 117234 406894 117854 442338
rect 117234 406658 117266 406894
rect 117502 406658 117586 406894
rect 117822 406658 117854 406894
rect 117234 406574 117854 406658
rect 117234 406338 117266 406574
rect 117502 406338 117586 406574
rect 117822 406338 117854 406574
rect 117234 370894 117854 406338
rect 117234 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 117854 370894
rect 117234 370574 117854 370658
rect 117234 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 117854 370574
rect 117234 334894 117854 370338
rect 117234 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 117854 334894
rect 117234 334574 117854 334658
rect 117234 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 117854 334574
rect 117234 298894 117854 334338
rect 117234 298658 117266 298894
rect 117502 298658 117586 298894
rect 117822 298658 117854 298894
rect 117234 298574 117854 298658
rect 117234 298338 117266 298574
rect 117502 298338 117586 298574
rect 117822 298338 117854 298574
rect 117234 262894 117854 298338
rect 117234 262658 117266 262894
rect 117502 262658 117586 262894
rect 117822 262658 117854 262894
rect 117234 262574 117854 262658
rect 117234 262338 117266 262574
rect 117502 262338 117586 262574
rect 117822 262338 117854 262574
rect 117234 226894 117854 262338
rect 117234 226658 117266 226894
rect 117502 226658 117586 226894
rect 117822 226658 117854 226894
rect 117234 226574 117854 226658
rect 117234 226338 117266 226574
rect 117502 226338 117586 226574
rect 117822 226338 117854 226574
rect 117234 190894 117854 226338
rect 117234 190658 117266 190894
rect 117502 190658 117586 190894
rect 117822 190658 117854 190894
rect 117234 190574 117854 190658
rect 117234 190338 117266 190574
rect 117502 190338 117586 190574
rect 117822 190338 117854 190574
rect 117234 154894 117854 190338
rect 117234 154658 117266 154894
rect 117502 154658 117586 154894
rect 117822 154658 117854 154894
rect 117234 154574 117854 154658
rect 117234 154338 117266 154574
rect 117502 154338 117586 154574
rect 117822 154338 117854 154574
rect 117234 118894 117854 154338
rect 117234 118658 117266 118894
rect 117502 118658 117586 118894
rect 117822 118658 117854 118894
rect 117234 118574 117854 118658
rect 117234 118338 117266 118574
rect 117502 118338 117586 118574
rect 117822 118338 117854 118574
rect 117234 82894 117854 118338
rect 117234 82658 117266 82894
rect 117502 82658 117586 82894
rect 117822 82658 117854 82894
rect 117234 82574 117854 82658
rect 117234 82338 117266 82574
rect 117502 82338 117586 82574
rect 117822 82338 117854 82574
rect 117234 46894 117854 82338
rect 117234 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 117854 46894
rect 117234 46574 117854 46658
rect 117234 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 117854 46574
rect 117234 10894 117854 46338
rect 117234 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 117854 10894
rect 117234 10574 117854 10658
rect 117234 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 117854 10574
rect 117234 -4186 117854 10338
rect 117234 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 117854 -4186
rect 117234 -4506 117854 -4422
rect 117234 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 117854 -4506
rect 117234 -5734 117854 -4742
rect 120954 698614 121574 710042
rect 138954 711558 139574 711590
rect 138954 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 139574 711558
rect 138954 711238 139574 711322
rect 138954 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 139574 711238
rect 135234 709638 135854 709670
rect 135234 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 135854 709638
rect 135234 709318 135854 709402
rect 135234 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 135854 709318
rect 131514 707718 132134 707750
rect 131514 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 132134 707718
rect 131514 707398 132134 707482
rect 131514 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 132134 707398
rect 120954 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 121574 698614
rect 120954 698294 121574 698378
rect 120954 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 121574 698294
rect 120954 662614 121574 698058
rect 120954 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 121574 662614
rect 120954 662294 121574 662378
rect 120954 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 121574 662294
rect 120954 626614 121574 662058
rect 120954 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 121574 626614
rect 120954 626294 121574 626378
rect 120954 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 121574 626294
rect 120954 590614 121574 626058
rect 120954 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 121574 590614
rect 120954 590294 121574 590378
rect 120954 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 121574 590294
rect 120954 554614 121574 590058
rect 120954 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 121574 554614
rect 120954 554294 121574 554378
rect 120954 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 121574 554294
rect 120954 518614 121574 554058
rect 120954 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 121574 518614
rect 120954 518294 121574 518378
rect 120954 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 121574 518294
rect 120954 482614 121574 518058
rect 120954 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 121574 482614
rect 120954 482294 121574 482378
rect 120954 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 121574 482294
rect 120954 446614 121574 482058
rect 120954 446378 120986 446614
rect 121222 446378 121306 446614
rect 121542 446378 121574 446614
rect 120954 446294 121574 446378
rect 120954 446058 120986 446294
rect 121222 446058 121306 446294
rect 121542 446058 121574 446294
rect 120954 410614 121574 446058
rect 120954 410378 120986 410614
rect 121222 410378 121306 410614
rect 121542 410378 121574 410614
rect 120954 410294 121574 410378
rect 120954 410058 120986 410294
rect 121222 410058 121306 410294
rect 121542 410058 121574 410294
rect 120954 374614 121574 410058
rect 120954 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 121574 374614
rect 120954 374294 121574 374378
rect 120954 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 121574 374294
rect 120954 338614 121574 374058
rect 120954 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 121574 338614
rect 120954 338294 121574 338378
rect 120954 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 121574 338294
rect 120954 302614 121574 338058
rect 120954 302378 120986 302614
rect 121222 302378 121306 302614
rect 121542 302378 121574 302614
rect 120954 302294 121574 302378
rect 120954 302058 120986 302294
rect 121222 302058 121306 302294
rect 121542 302058 121574 302294
rect 120954 266614 121574 302058
rect 120954 266378 120986 266614
rect 121222 266378 121306 266614
rect 121542 266378 121574 266614
rect 120954 266294 121574 266378
rect 120954 266058 120986 266294
rect 121222 266058 121306 266294
rect 121542 266058 121574 266294
rect 120954 230614 121574 266058
rect 120954 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 121574 230614
rect 120954 230294 121574 230378
rect 120954 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 121574 230294
rect 120954 194614 121574 230058
rect 120954 194378 120986 194614
rect 121222 194378 121306 194614
rect 121542 194378 121574 194614
rect 120954 194294 121574 194378
rect 120954 194058 120986 194294
rect 121222 194058 121306 194294
rect 121542 194058 121574 194294
rect 120954 158614 121574 194058
rect 120954 158378 120986 158614
rect 121222 158378 121306 158614
rect 121542 158378 121574 158614
rect 120954 158294 121574 158378
rect 120954 158058 120986 158294
rect 121222 158058 121306 158294
rect 121542 158058 121574 158294
rect 120954 122614 121574 158058
rect 120954 122378 120986 122614
rect 121222 122378 121306 122614
rect 121542 122378 121574 122614
rect 120954 122294 121574 122378
rect 120954 122058 120986 122294
rect 121222 122058 121306 122294
rect 121542 122058 121574 122294
rect 120954 86614 121574 122058
rect 120954 86378 120986 86614
rect 121222 86378 121306 86614
rect 121542 86378 121574 86614
rect 120954 86294 121574 86378
rect 120954 86058 120986 86294
rect 121222 86058 121306 86294
rect 121542 86058 121574 86294
rect 120954 50614 121574 86058
rect 120954 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 121574 50614
rect 120954 50294 121574 50378
rect 120954 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 121574 50294
rect 120954 14614 121574 50058
rect 120954 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 121574 14614
rect 120954 14294 121574 14378
rect 120954 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 121574 14294
rect 102954 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 103574 -7066
rect 102954 -7386 103574 -7302
rect 102954 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 103574 -7386
rect 102954 -7654 103574 -7622
rect 120954 -6106 121574 14058
rect 127794 705798 128414 705830
rect 127794 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 128414 705798
rect 127794 705478 128414 705562
rect 127794 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 128414 705478
rect 127794 669454 128414 705242
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 127794 561454 128414 596898
rect 127794 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 128414 561454
rect 127794 561134 128414 561218
rect 127794 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 128414 561134
rect 127794 525454 128414 560898
rect 127794 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 128414 525454
rect 127794 525134 128414 525218
rect 127794 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 128414 525134
rect 127794 489454 128414 524898
rect 127794 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 128414 489454
rect 127794 489134 128414 489218
rect 127794 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 128414 489134
rect 127794 453454 128414 488898
rect 127794 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 128414 453454
rect 127794 453134 128414 453218
rect 127794 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 128414 453134
rect 127794 417454 128414 452898
rect 127794 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 128414 417454
rect 127794 417134 128414 417218
rect 127794 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 128414 417134
rect 127794 381454 128414 416898
rect 127794 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 128414 381454
rect 127794 381134 128414 381218
rect 127794 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 128414 381134
rect 127794 345454 128414 380898
rect 127794 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 128414 345454
rect 127794 345134 128414 345218
rect 127794 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 128414 345134
rect 127794 309454 128414 344898
rect 127794 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 128414 309454
rect 127794 309134 128414 309218
rect 127794 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 128414 309134
rect 127794 273454 128414 308898
rect 127794 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 128414 273454
rect 127794 273134 128414 273218
rect 127794 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 128414 273134
rect 127794 237454 128414 272898
rect 127794 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 128414 237454
rect 127794 237134 128414 237218
rect 127794 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 128414 237134
rect 127794 201454 128414 236898
rect 127794 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 128414 201454
rect 127794 201134 128414 201218
rect 127794 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 128414 201134
rect 127794 165454 128414 200898
rect 127794 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 128414 165454
rect 127794 165134 128414 165218
rect 127794 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 128414 165134
rect 127794 129454 128414 164898
rect 127794 129218 127826 129454
rect 128062 129218 128146 129454
rect 128382 129218 128414 129454
rect 127794 129134 128414 129218
rect 127794 128898 127826 129134
rect 128062 128898 128146 129134
rect 128382 128898 128414 129134
rect 127794 93454 128414 128898
rect 127794 93218 127826 93454
rect 128062 93218 128146 93454
rect 128382 93218 128414 93454
rect 127794 93134 128414 93218
rect 127794 92898 127826 93134
rect 128062 92898 128146 93134
rect 128382 92898 128414 93134
rect 127794 57454 128414 92898
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -1306 128414 20898
rect 127794 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 128414 -1306
rect 127794 -1626 128414 -1542
rect 127794 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 128414 -1626
rect 127794 -1894 128414 -1862
rect 131514 673174 132134 707162
rect 131514 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 132134 673174
rect 131514 672854 132134 672938
rect 131514 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 132134 672854
rect 131514 637174 132134 672618
rect 131514 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 132134 637174
rect 131514 636854 132134 636938
rect 131514 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 132134 636854
rect 131514 601174 132134 636618
rect 131514 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 132134 601174
rect 131514 600854 132134 600938
rect 131514 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 132134 600854
rect 131514 565174 132134 600618
rect 131514 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 132134 565174
rect 131514 564854 132134 564938
rect 131514 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 132134 564854
rect 131514 529174 132134 564618
rect 131514 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 132134 529174
rect 131514 528854 132134 528938
rect 131514 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 132134 528854
rect 131514 493174 132134 528618
rect 131514 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 132134 493174
rect 131514 492854 132134 492938
rect 131514 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 132134 492854
rect 131514 457174 132134 492618
rect 131514 456938 131546 457174
rect 131782 456938 131866 457174
rect 132102 456938 132134 457174
rect 131514 456854 132134 456938
rect 131514 456618 131546 456854
rect 131782 456618 131866 456854
rect 132102 456618 132134 456854
rect 131514 421174 132134 456618
rect 131514 420938 131546 421174
rect 131782 420938 131866 421174
rect 132102 420938 132134 421174
rect 131514 420854 132134 420938
rect 131514 420618 131546 420854
rect 131782 420618 131866 420854
rect 132102 420618 132134 420854
rect 131514 385174 132134 420618
rect 131514 384938 131546 385174
rect 131782 384938 131866 385174
rect 132102 384938 132134 385174
rect 131514 384854 132134 384938
rect 131514 384618 131546 384854
rect 131782 384618 131866 384854
rect 132102 384618 132134 384854
rect 131514 349174 132134 384618
rect 131514 348938 131546 349174
rect 131782 348938 131866 349174
rect 132102 348938 132134 349174
rect 131514 348854 132134 348938
rect 131514 348618 131546 348854
rect 131782 348618 131866 348854
rect 132102 348618 132134 348854
rect 131514 313174 132134 348618
rect 131514 312938 131546 313174
rect 131782 312938 131866 313174
rect 132102 312938 132134 313174
rect 131514 312854 132134 312938
rect 131514 312618 131546 312854
rect 131782 312618 131866 312854
rect 132102 312618 132134 312854
rect 131514 277174 132134 312618
rect 131514 276938 131546 277174
rect 131782 276938 131866 277174
rect 132102 276938 132134 277174
rect 131514 276854 132134 276938
rect 131514 276618 131546 276854
rect 131782 276618 131866 276854
rect 132102 276618 132134 276854
rect 131514 241174 132134 276618
rect 131514 240938 131546 241174
rect 131782 240938 131866 241174
rect 132102 240938 132134 241174
rect 131514 240854 132134 240938
rect 131514 240618 131546 240854
rect 131782 240618 131866 240854
rect 132102 240618 132134 240854
rect 131514 205174 132134 240618
rect 131514 204938 131546 205174
rect 131782 204938 131866 205174
rect 132102 204938 132134 205174
rect 131514 204854 132134 204938
rect 131514 204618 131546 204854
rect 131782 204618 131866 204854
rect 132102 204618 132134 204854
rect 131514 169174 132134 204618
rect 131514 168938 131546 169174
rect 131782 168938 131866 169174
rect 132102 168938 132134 169174
rect 131514 168854 132134 168938
rect 131514 168618 131546 168854
rect 131782 168618 131866 168854
rect 132102 168618 132134 168854
rect 131514 133174 132134 168618
rect 131514 132938 131546 133174
rect 131782 132938 131866 133174
rect 132102 132938 132134 133174
rect 131514 132854 132134 132938
rect 131514 132618 131546 132854
rect 131782 132618 131866 132854
rect 132102 132618 132134 132854
rect 131514 97174 132134 132618
rect 131514 96938 131546 97174
rect 131782 96938 131866 97174
rect 132102 96938 132134 97174
rect 131514 96854 132134 96938
rect 131514 96618 131546 96854
rect 131782 96618 131866 96854
rect 132102 96618 132134 96854
rect 131514 61174 132134 96618
rect 131514 60938 131546 61174
rect 131782 60938 131866 61174
rect 132102 60938 132134 61174
rect 131514 60854 132134 60938
rect 131514 60618 131546 60854
rect 131782 60618 131866 60854
rect 132102 60618 132134 60854
rect 131514 25174 132134 60618
rect 131514 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 132134 25174
rect 131514 24854 132134 24938
rect 131514 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 132134 24854
rect 131514 -3226 132134 24618
rect 131514 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 132134 -3226
rect 131514 -3546 132134 -3462
rect 131514 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 132134 -3546
rect 131514 -3814 132134 -3782
rect 135234 676894 135854 709082
rect 135234 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 135854 676894
rect 135234 676574 135854 676658
rect 135234 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 135854 676574
rect 135234 640894 135854 676338
rect 135234 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 135854 640894
rect 135234 640574 135854 640658
rect 135234 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 135854 640574
rect 135234 604894 135854 640338
rect 135234 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 135854 604894
rect 135234 604574 135854 604658
rect 135234 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 135854 604574
rect 135234 568894 135854 604338
rect 135234 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 135854 568894
rect 135234 568574 135854 568658
rect 135234 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 135854 568574
rect 135234 532894 135854 568338
rect 135234 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 135854 532894
rect 135234 532574 135854 532658
rect 135234 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 135854 532574
rect 135234 496894 135854 532338
rect 135234 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 135854 496894
rect 135234 496574 135854 496658
rect 135234 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 135854 496574
rect 135234 460894 135854 496338
rect 135234 460658 135266 460894
rect 135502 460658 135586 460894
rect 135822 460658 135854 460894
rect 135234 460574 135854 460658
rect 135234 460338 135266 460574
rect 135502 460338 135586 460574
rect 135822 460338 135854 460574
rect 135234 424894 135854 460338
rect 135234 424658 135266 424894
rect 135502 424658 135586 424894
rect 135822 424658 135854 424894
rect 135234 424574 135854 424658
rect 135234 424338 135266 424574
rect 135502 424338 135586 424574
rect 135822 424338 135854 424574
rect 135234 388894 135854 424338
rect 135234 388658 135266 388894
rect 135502 388658 135586 388894
rect 135822 388658 135854 388894
rect 135234 388574 135854 388658
rect 135234 388338 135266 388574
rect 135502 388338 135586 388574
rect 135822 388338 135854 388574
rect 135234 352894 135854 388338
rect 135234 352658 135266 352894
rect 135502 352658 135586 352894
rect 135822 352658 135854 352894
rect 135234 352574 135854 352658
rect 135234 352338 135266 352574
rect 135502 352338 135586 352574
rect 135822 352338 135854 352574
rect 135234 316894 135854 352338
rect 135234 316658 135266 316894
rect 135502 316658 135586 316894
rect 135822 316658 135854 316894
rect 135234 316574 135854 316658
rect 135234 316338 135266 316574
rect 135502 316338 135586 316574
rect 135822 316338 135854 316574
rect 135234 280894 135854 316338
rect 135234 280658 135266 280894
rect 135502 280658 135586 280894
rect 135822 280658 135854 280894
rect 135234 280574 135854 280658
rect 135234 280338 135266 280574
rect 135502 280338 135586 280574
rect 135822 280338 135854 280574
rect 135234 244894 135854 280338
rect 135234 244658 135266 244894
rect 135502 244658 135586 244894
rect 135822 244658 135854 244894
rect 135234 244574 135854 244658
rect 135234 244338 135266 244574
rect 135502 244338 135586 244574
rect 135822 244338 135854 244574
rect 135234 208894 135854 244338
rect 135234 208658 135266 208894
rect 135502 208658 135586 208894
rect 135822 208658 135854 208894
rect 135234 208574 135854 208658
rect 135234 208338 135266 208574
rect 135502 208338 135586 208574
rect 135822 208338 135854 208574
rect 135234 172894 135854 208338
rect 135234 172658 135266 172894
rect 135502 172658 135586 172894
rect 135822 172658 135854 172894
rect 135234 172574 135854 172658
rect 135234 172338 135266 172574
rect 135502 172338 135586 172574
rect 135822 172338 135854 172574
rect 135234 136894 135854 172338
rect 135234 136658 135266 136894
rect 135502 136658 135586 136894
rect 135822 136658 135854 136894
rect 135234 136574 135854 136658
rect 135234 136338 135266 136574
rect 135502 136338 135586 136574
rect 135822 136338 135854 136574
rect 135234 100894 135854 136338
rect 135234 100658 135266 100894
rect 135502 100658 135586 100894
rect 135822 100658 135854 100894
rect 135234 100574 135854 100658
rect 135234 100338 135266 100574
rect 135502 100338 135586 100574
rect 135822 100338 135854 100574
rect 135234 64894 135854 100338
rect 135234 64658 135266 64894
rect 135502 64658 135586 64894
rect 135822 64658 135854 64894
rect 135234 64574 135854 64658
rect 135234 64338 135266 64574
rect 135502 64338 135586 64574
rect 135822 64338 135854 64574
rect 135234 28894 135854 64338
rect 135234 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 135854 28894
rect 135234 28574 135854 28658
rect 135234 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 135854 28574
rect 135234 -5146 135854 28338
rect 135234 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 135854 -5146
rect 135234 -5466 135854 -5382
rect 135234 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 135854 -5466
rect 135234 -5734 135854 -5702
rect 138954 680614 139574 711002
rect 156954 710598 157574 711590
rect 156954 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 157574 710598
rect 156954 710278 157574 710362
rect 156954 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 157574 710278
rect 153234 708678 153854 709670
rect 153234 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 153854 708678
rect 153234 708358 153854 708442
rect 153234 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 153854 708358
rect 149514 706758 150134 707750
rect 149514 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 150134 706758
rect 149514 706438 150134 706522
rect 149514 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 150134 706438
rect 138954 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 139574 680614
rect 138954 680294 139574 680378
rect 138954 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 139574 680294
rect 138954 644614 139574 680058
rect 138954 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 139574 644614
rect 138954 644294 139574 644378
rect 138954 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 139574 644294
rect 138954 608614 139574 644058
rect 138954 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 139574 608614
rect 138954 608294 139574 608378
rect 138954 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 139574 608294
rect 138954 572614 139574 608058
rect 138954 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 139574 572614
rect 138954 572294 139574 572378
rect 138954 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 139574 572294
rect 138954 536614 139574 572058
rect 138954 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 139574 536614
rect 138954 536294 139574 536378
rect 138954 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 139574 536294
rect 138954 500614 139574 536058
rect 138954 500378 138986 500614
rect 139222 500378 139306 500614
rect 139542 500378 139574 500614
rect 138954 500294 139574 500378
rect 138954 500058 138986 500294
rect 139222 500058 139306 500294
rect 139542 500058 139574 500294
rect 138954 464614 139574 500058
rect 138954 464378 138986 464614
rect 139222 464378 139306 464614
rect 139542 464378 139574 464614
rect 138954 464294 139574 464378
rect 138954 464058 138986 464294
rect 139222 464058 139306 464294
rect 139542 464058 139574 464294
rect 138954 428614 139574 464058
rect 138954 428378 138986 428614
rect 139222 428378 139306 428614
rect 139542 428378 139574 428614
rect 138954 428294 139574 428378
rect 138954 428058 138986 428294
rect 139222 428058 139306 428294
rect 139542 428058 139574 428294
rect 138954 392614 139574 428058
rect 138954 392378 138986 392614
rect 139222 392378 139306 392614
rect 139542 392378 139574 392614
rect 138954 392294 139574 392378
rect 138954 392058 138986 392294
rect 139222 392058 139306 392294
rect 139542 392058 139574 392294
rect 138954 356614 139574 392058
rect 138954 356378 138986 356614
rect 139222 356378 139306 356614
rect 139542 356378 139574 356614
rect 138954 356294 139574 356378
rect 138954 356058 138986 356294
rect 139222 356058 139306 356294
rect 139542 356058 139574 356294
rect 138954 320614 139574 356058
rect 138954 320378 138986 320614
rect 139222 320378 139306 320614
rect 139542 320378 139574 320614
rect 138954 320294 139574 320378
rect 138954 320058 138986 320294
rect 139222 320058 139306 320294
rect 139542 320058 139574 320294
rect 138954 284614 139574 320058
rect 138954 284378 138986 284614
rect 139222 284378 139306 284614
rect 139542 284378 139574 284614
rect 138954 284294 139574 284378
rect 138954 284058 138986 284294
rect 139222 284058 139306 284294
rect 139542 284058 139574 284294
rect 138954 248614 139574 284058
rect 138954 248378 138986 248614
rect 139222 248378 139306 248614
rect 139542 248378 139574 248614
rect 138954 248294 139574 248378
rect 138954 248058 138986 248294
rect 139222 248058 139306 248294
rect 139542 248058 139574 248294
rect 138954 212614 139574 248058
rect 138954 212378 138986 212614
rect 139222 212378 139306 212614
rect 139542 212378 139574 212614
rect 138954 212294 139574 212378
rect 138954 212058 138986 212294
rect 139222 212058 139306 212294
rect 139542 212058 139574 212294
rect 138954 176614 139574 212058
rect 138954 176378 138986 176614
rect 139222 176378 139306 176614
rect 139542 176378 139574 176614
rect 138954 176294 139574 176378
rect 138954 176058 138986 176294
rect 139222 176058 139306 176294
rect 139542 176058 139574 176294
rect 138954 140614 139574 176058
rect 138954 140378 138986 140614
rect 139222 140378 139306 140614
rect 139542 140378 139574 140614
rect 138954 140294 139574 140378
rect 138954 140058 138986 140294
rect 139222 140058 139306 140294
rect 139542 140058 139574 140294
rect 138954 104614 139574 140058
rect 138954 104378 138986 104614
rect 139222 104378 139306 104614
rect 139542 104378 139574 104614
rect 138954 104294 139574 104378
rect 138954 104058 138986 104294
rect 139222 104058 139306 104294
rect 139542 104058 139574 104294
rect 138954 68614 139574 104058
rect 138954 68378 138986 68614
rect 139222 68378 139306 68614
rect 139542 68378 139574 68614
rect 138954 68294 139574 68378
rect 138954 68058 138986 68294
rect 139222 68058 139306 68294
rect 139542 68058 139574 68294
rect 138954 32614 139574 68058
rect 138954 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 139574 32614
rect 138954 32294 139574 32378
rect 138954 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 139574 32294
rect 120954 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 121574 -6106
rect 120954 -6426 121574 -6342
rect 120954 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 121574 -6426
rect 120954 -7654 121574 -6662
rect 138954 -7066 139574 32058
rect 145794 704838 146414 705830
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 543454 146414 578898
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 507454 146414 542898
rect 145794 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 146414 507454
rect 145794 507134 146414 507218
rect 145794 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 146414 507134
rect 145794 471454 146414 506898
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 435454 146414 470898
rect 145794 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 146414 435454
rect 145794 435134 146414 435218
rect 145794 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 146414 435134
rect 145794 399454 146414 434898
rect 145794 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 146414 399454
rect 145794 399134 146414 399218
rect 145794 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 146414 399134
rect 145794 363454 146414 398898
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 145794 327454 146414 362898
rect 145794 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 146414 327454
rect 145794 327134 146414 327218
rect 145794 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 146414 327134
rect 145794 291454 146414 326898
rect 145794 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 146414 291454
rect 145794 291134 146414 291218
rect 145794 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 146414 291134
rect 145794 255454 146414 290898
rect 145794 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 146414 255454
rect 145794 255134 146414 255218
rect 145794 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 146414 255134
rect 145794 219454 146414 254898
rect 145794 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 146414 219454
rect 145794 219134 146414 219218
rect 145794 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 146414 219134
rect 145794 183454 146414 218898
rect 145794 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 146414 183454
rect 145794 183134 146414 183218
rect 145794 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 146414 183134
rect 145794 147454 146414 182898
rect 145794 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 146414 147454
rect 145794 147134 146414 147218
rect 145794 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 146414 147134
rect 145794 111454 146414 146898
rect 145794 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 146414 111454
rect 145794 111134 146414 111218
rect 145794 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 146414 111134
rect 145794 75454 146414 110898
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145794 75134 146414 75218
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 145794 39454 146414 74898
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -1894 146414 -902
rect 149514 691174 150134 706202
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 655174 150134 690618
rect 149514 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 150134 655174
rect 149514 654854 150134 654938
rect 149514 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 150134 654854
rect 149514 619174 150134 654618
rect 149514 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 150134 619174
rect 149514 618854 150134 618938
rect 149514 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 150134 618854
rect 149514 583174 150134 618618
rect 149514 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 150134 583174
rect 149514 582854 150134 582938
rect 149514 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 150134 582854
rect 149514 547174 150134 582618
rect 149514 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 150134 547174
rect 149514 546854 150134 546938
rect 149514 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 150134 546854
rect 149514 511174 150134 546618
rect 149514 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 150134 511174
rect 149514 510854 150134 510938
rect 149514 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 150134 510854
rect 149514 475174 150134 510618
rect 149514 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 150134 475174
rect 149514 474854 150134 474938
rect 149514 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 150134 474854
rect 149514 439174 150134 474618
rect 149514 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 150134 439174
rect 149514 438854 150134 438938
rect 149514 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 150134 438854
rect 149514 403174 150134 438618
rect 149514 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 150134 403174
rect 149514 402854 150134 402938
rect 149514 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 150134 402854
rect 149514 367174 150134 402618
rect 149514 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 150134 367174
rect 149514 366854 150134 366938
rect 149514 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 150134 366854
rect 149514 331174 150134 366618
rect 149514 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 150134 331174
rect 149514 330854 150134 330938
rect 149514 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 150134 330854
rect 149514 295174 150134 330618
rect 149514 294938 149546 295174
rect 149782 294938 149866 295174
rect 150102 294938 150134 295174
rect 149514 294854 150134 294938
rect 149514 294618 149546 294854
rect 149782 294618 149866 294854
rect 150102 294618 150134 294854
rect 149514 259174 150134 294618
rect 149514 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 150134 259174
rect 149514 258854 150134 258938
rect 149514 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 150134 258854
rect 149514 223174 150134 258618
rect 149514 222938 149546 223174
rect 149782 222938 149866 223174
rect 150102 222938 150134 223174
rect 149514 222854 150134 222938
rect 149514 222618 149546 222854
rect 149782 222618 149866 222854
rect 150102 222618 150134 222854
rect 149514 187174 150134 222618
rect 149514 186938 149546 187174
rect 149782 186938 149866 187174
rect 150102 186938 150134 187174
rect 149514 186854 150134 186938
rect 149514 186618 149546 186854
rect 149782 186618 149866 186854
rect 150102 186618 150134 186854
rect 149514 151174 150134 186618
rect 149514 150938 149546 151174
rect 149782 150938 149866 151174
rect 150102 150938 150134 151174
rect 149514 150854 150134 150938
rect 149514 150618 149546 150854
rect 149782 150618 149866 150854
rect 150102 150618 150134 150854
rect 149514 115174 150134 150618
rect 149514 114938 149546 115174
rect 149782 114938 149866 115174
rect 150102 114938 150134 115174
rect 149514 114854 150134 114938
rect 149514 114618 149546 114854
rect 149782 114618 149866 114854
rect 150102 114618 150134 114854
rect 149514 79174 150134 114618
rect 149514 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 150134 79174
rect 149514 78854 150134 78938
rect 149514 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 150134 78854
rect 149514 43174 150134 78618
rect 149514 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 150134 43174
rect 149514 42854 150134 42938
rect 149514 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 150134 42854
rect 149514 7174 150134 42618
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 149514 -2266 150134 6618
rect 149514 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 150134 -2266
rect 149514 -2586 150134 -2502
rect 149514 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 150134 -2586
rect 149514 -3814 150134 -2822
rect 153234 694894 153854 708122
rect 153234 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 153854 694894
rect 153234 694574 153854 694658
rect 153234 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 153854 694574
rect 153234 658894 153854 694338
rect 153234 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 153854 658894
rect 153234 658574 153854 658658
rect 153234 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 153854 658574
rect 153234 622894 153854 658338
rect 153234 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 153854 622894
rect 153234 622574 153854 622658
rect 153234 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 153854 622574
rect 153234 586894 153854 622338
rect 153234 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 153854 586894
rect 153234 586574 153854 586658
rect 153234 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 153854 586574
rect 153234 550894 153854 586338
rect 153234 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 153854 550894
rect 153234 550574 153854 550658
rect 153234 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 153854 550574
rect 153234 514894 153854 550338
rect 153234 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 153854 514894
rect 153234 514574 153854 514658
rect 153234 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 153854 514574
rect 153234 478894 153854 514338
rect 153234 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 153854 478894
rect 153234 478574 153854 478658
rect 153234 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 153854 478574
rect 153234 442894 153854 478338
rect 153234 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 153854 442894
rect 153234 442574 153854 442658
rect 153234 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 153854 442574
rect 153234 406894 153854 442338
rect 153234 406658 153266 406894
rect 153502 406658 153586 406894
rect 153822 406658 153854 406894
rect 153234 406574 153854 406658
rect 153234 406338 153266 406574
rect 153502 406338 153586 406574
rect 153822 406338 153854 406574
rect 153234 370894 153854 406338
rect 153234 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 153854 370894
rect 153234 370574 153854 370658
rect 153234 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 153854 370574
rect 153234 334894 153854 370338
rect 153234 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 153854 334894
rect 153234 334574 153854 334658
rect 153234 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 153854 334574
rect 153234 298894 153854 334338
rect 153234 298658 153266 298894
rect 153502 298658 153586 298894
rect 153822 298658 153854 298894
rect 153234 298574 153854 298658
rect 153234 298338 153266 298574
rect 153502 298338 153586 298574
rect 153822 298338 153854 298574
rect 153234 262894 153854 298338
rect 153234 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 153854 262894
rect 153234 262574 153854 262658
rect 153234 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 153854 262574
rect 153234 226894 153854 262338
rect 153234 226658 153266 226894
rect 153502 226658 153586 226894
rect 153822 226658 153854 226894
rect 153234 226574 153854 226658
rect 153234 226338 153266 226574
rect 153502 226338 153586 226574
rect 153822 226338 153854 226574
rect 153234 190894 153854 226338
rect 153234 190658 153266 190894
rect 153502 190658 153586 190894
rect 153822 190658 153854 190894
rect 153234 190574 153854 190658
rect 153234 190338 153266 190574
rect 153502 190338 153586 190574
rect 153822 190338 153854 190574
rect 153234 154894 153854 190338
rect 153234 154658 153266 154894
rect 153502 154658 153586 154894
rect 153822 154658 153854 154894
rect 153234 154574 153854 154658
rect 153234 154338 153266 154574
rect 153502 154338 153586 154574
rect 153822 154338 153854 154574
rect 153234 118894 153854 154338
rect 153234 118658 153266 118894
rect 153502 118658 153586 118894
rect 153822 118658 153854 118894
rect 153234 118574 153854 118658
rect 153234 118338 153266 118574
rect 153502 118338 153586 118574
rect 153822 118338 153854 118574
rect 153234 82894 153854 118338
rect 153234 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 153854 82894
rect 153234 82574 153854 82658
rect 153234 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 153854 82574
rect 153234 46894 153854 82338
rect 153234 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 153854 46894
rect 153234 46574 153854 46658
rect 153234 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 153854 46574
rect 153234 10894 153854 46338
rect 153234 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 153854 10894
rect 153234 10574 153854 10658
rect 153234 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 153854 10574
rect 153234 -4186 153854 10338
rect 153234 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 153854 -4186
rect 153234 -4506 153854 -4422
rect 153234 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 153854 -4506
rect 153234 -5734 153854 -4742
rect 156954 698614 157574 710042
rect 174954 711558 175574 711590
rect 174954 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 175574 711558
rect 174954 711238 175574 711322
rect 174954 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 175574 711238
rect 171234 709638 171854 709670
rect 171234 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 171854 709638
rect 171234 709318 171854 709402
rect 171234 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 171854 709318
rect 167514 707718 168134 707750
rect 167514 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 168134 707718
rect 167514 707398 168134 707482
rect 167514 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 168134 707398
rect 156954 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 157574 698614
rect 156954 698294 157574 698378
rect 156954 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 157574 698294
rect 156954 662614 157574 698058
rect 156954 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 157574 662614
rect 156954 662294 157574 662378
rect 156954 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 157574 662294
rect 156954 626614 157574 662058
rect 156954 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 157574 626614
rect 156954 626294 157574 626378
rect 156954 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 157574 626294
rect 156954 590614 157574 626058
rect 156954 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 157574 590614
rect 156954 590294 157574 590378
rect 156954 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 157574 590294
rect 156954 554614 157574 590058
rect 156954 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 157574 554614
rect 156954 554294 157574 554378
rect 156954 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 157574 554294
rect 156954 518614 157574 554058
rect 156954 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 157574 518614
rect 156954 518294 157574 518378
rect 156954 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 157574 518294
rect 156954 482614 157574 518058
rect 156954 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 157574 482614
rect 156954 482294 157574 482378
rect 156954 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 157574 482294
rect 156954 446614 157574 482058
rect 156954 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 157574 446614
rect 156954 446294 157574 446378
rect 156954 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 157574 446294
rect 156954 410614 157574 446058
rect 156954 410378 156986 410614
rect 157222 410378 157306 410614
rect 157542 410378 157574 410614
rect 156954 410294 157574 410378
rect 156954 410058 156986 410294
rect 157222 410058 157306 410294
rect 157542 410058 157574 410294
rect 156954 374614 157574 410058
rect 156954 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 157574 374614
rect 156954 374294 157574 374378
rect 156954 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 157574 374294
rect 156954 338614 157574 374058
rect 156954 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 157574 338614
rect 156954 338294 157574 338378
rect 156954 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 157574 338294
rect 156954 302614 157574 338058
rect 156954 302378 156986 302614
rect 157222 302378 157306 302614
rect 157542 302378 157574 302614
rect 156954 302294 157574 302378
rect 156954 302058 156986 302294
rect 157222 302058 157306 302294
rect 157542 302058 157574 302294
rect 156954 266614 157574 302058
rect 156954 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 157574 266614
rect 156954 266294 157574 266378
rect 156954 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 157574 266294
rect 156954 230614 157574 266058
rect 156954 230378 156986 230614
rect 157222 230378 157306 230614
rect 157542 230378 157574 230614
rect 156954 230294 157574 230378
rect 156954 230058 156986 230294
rect 157222 230058 157306 230294
rect 157542 230058 157574 230294
rect 156954 194614 157574 230058
rect 156954 194378 156986 194614
rect 157222 194378 157306 194614
rect 157542 194378 157574 194614
rect 156954 194294 157574 194378
rect 156954 194058 156986 194294
rect 157222 194058 157306 194294
rect 157542 194058 157574 194294
rect 156954 158614 157574 194058
rect 163794 705798 164414 705830
rect 163794 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 164414 705798
rect 163794 705478 164414 705562
rect 163794 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 164414 705478
rect 163794 669454 164414 705242
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 163794 561454 164414 596898
rect 163794 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 164414 561454
rect 163794 561134 164414 561218
rect 163794 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 164414 561134
rect 163794 525454 164414 560898
rect 163794 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 164414 525454
rect 163794 525134 164414 525218
rect 163794 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 164414 525134
rect 163794 489454 164414 524898
rect 163794 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 164414 489454
rect 163794 489134 164414 489218
rect 163794 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 164414 489134
rect 163794 453454 164414 488898
rect 163794 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 164414 453454
rect 163794 453134 164414 453218
rect 163794 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 164414 453134
rect 163794 417454 164414 452898
rect 163794 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 164414 417454
rect 163794 417134 164414 417218
rect 163794 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 164414 417134
rect 163794 381454 164414 416898
rect 163794 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 164414 381454
rect 163794 381134 164414 381218
rect 163794 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 164414 381134
rect 163794 345454 164414 380898
rect 163794 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 164414 345454
rect 163794 345134 164414 345218
rect 163794 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 164414 345134
rect 163794 309454 164414 344898
rect 163794 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 164414 309454
rect 163794 309134 164414 309218
rect 163794 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 164414 309134
rect 163794 273454 164414 308898
rect 163794 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 164414 273454
rect 163794 273134 164414 273218
rect 163794 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 164414 273134
rect 163794 237454 164414 272898
rect 163794 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 164414 237454
rect 163794 237134 164414 237218
rect 163794 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 164414 237134
rect 163794 201454 164414 236898
rect 163794 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 164414 201454
rect 163794 201134 164414 201218
rect 163794 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 164414 201134
rect 163794 192000 164414 200898
rect 167514 673174 168134 707162
rect 167514 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 168134 673174
rect 167514 672854 168134 672938
rect 167514 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 168134 672854
rect 167514 637174 168134 672618
rect 167514 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 168134 637174
rect 167514 636854 168134 636938
rect 167514 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 168134 636854
rect 167514 601174 168134 636618
rect 167514 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 168134 601174
rect 167514 600854 168134 600938
rect 167514 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 168134 600854
rect 167514 565174 168134 600618
rect 167514 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 168134 565174
rect 167514 564854 168134 564938
rect 167514 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 168134 564854
rect 167514 529174 168134 564618
rect 167514 528938 167546 529174
rect 167782 528938 167866 529174
rect 168102 528938 168134 529174
rect 167514 528854 168134 528938
rect 167514 528618 167546 528854
rect 167782 528618 167866 528854
rect 168102 528618 168134 528854
rect 167514 493174 168134 528618
rect 167514 492938 167546 493174
rect 167782 492938 167866 493174
rect 168102 492938 168134 493174
rect 167514 492854 168134 492938
rect 167514 492618 167546 492854
rect 167782 492618 167866 492854
rect 168102 492618 168134 492854
rect 167514 457174 168134 492618
rect 167514 456938 167546 457174
rect 167782 456938 167866 457174
rect 168102 456938 168134 457174
rect 167514 456854 168134 456938
rect 167514 456618 167546 456854
rect 167782 456618 167866 456854
rect 168102 456618 168134 456854
rect 167514 421174 168134 456618
rect 167514 420938 167546 421174
rect 167782 420938 167866 421174
rect 168102 420938 168134 421174
rect 167514 420854 168134 420938
rect 167514 420618 167546 420854
rect 167782 420618 167866 420854
rect 168102 420618 168134 420854
rect 167514 385174 168134 420618
rect 167514 384938 167546 385174
rect 167782 384938 167866 385174
rect 168102 384938 168134 385174
rect 167514 384854 168134 384938
rect 167514 384618 167546 384854
rect 167782 384618 167866 384854
rect 168102 384618 168134 384854
rect 167514 349174 168134 384618
rect 167514 348938 167546 349174
rect 167782 348938 167866 349174
rect 168102 348938 168134 349174
rect 167514 348854 168134 348938
rect 167514 348618 167546 348854
rect 167782 348618 167866 348854
rect 168102 348618 168134 348854
rect 167514 313174 168134 348618
rect 167514 312938 167546 313174
rect 167782 312938 167866 313174
rect 168102 312938 168134 313174
rect 167514 312854 168134 312938
rect 167514 312618 167546 312854
rect 167782 312618 167866 312854
rect 168102 312618 168134 312854
rect 167514 277174 168134 312618
rect 167514 276938 167546 277174
rect 167782 276938 167866 277174
rect 168102 276938 168134 277174
rect 167514 276854 168134 276938
rect 167514 276618 167546 276854
rect 167782 276618 167866 276854
rect 168102 276618 168134 276854
rect 167514 241174 168134 276618
rect 167514 240938 167546 241174
rect 167782 240938 167866 241174
rect 168102 240938 168134 241174
rect 167514 240854 168134 240938
rect 167514 240618 167546 240854
rect 167782 240618 167866 240854
rect 168102 240618 168134 240854
rect 167514 205174 168134 240618
rect 167514 204938 167546 205174
rect 167782 204938 167866 205174
rect 168102 204938 168134 205174
rect 167514 204854 168134 204938
rect 167514 204618 167546 204854
rect 167782 204618 167866 204854
rect 168102 204618 168134 204854
rect 167514 192000 168134 204618
rect 171234 676894 171854 709082
rect 171234 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 171854 676894
rect 171234 676574 171854 676658
rect 171234 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 171854 676574
rect 171234 640894 171854 676338
rect 171234 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 171854 640894
rect 171234 640574 171854 640658
rect 171234 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 171854 640574
rect 171234 604894 171854 640338
rect 171234 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 171854 604894
rect 171234 604574 171854 604658
rect 171234 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 171854 604574
rect 171234 568894 171854 604338
rect 171234 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 171854 568894
rect 171234 568574 171854 568658
rect 171234 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 171854 568574
rect 171234 532894 171854 568338
rect 171234 532658 171266 532894
rect 171502 532658 171586 532894
rect 171822 532658 171854 532894
rect 171234 532574 171854 532658
rect 171234 532338 171266 532574
rect 171502 532338 171586 532574
rect 171822 532338 171854 532574
rect 171234 496894 171854 532338
rect 171234 496658 171266 496894
rect 171502 496658 171586 496894
rect 171822 496658 171854 496894
rect 171234 496574 171854 496658
rect 171234 496338 171266 496574
rect 171502 496338 171586 496574
rect 171822 496338 171854 496574
rect 171234 460894 171854 496338
rect 171234 460658 171266 460894
rect 171502 460658 171586 460894
rect 171822 460658 171854 460894
rect 171234 460574 171854 460658
rect 171234 460338 171266 460574
rect 171502 460338 171586 460574
rect 171822 460338 171854 460574
rect 171234 424894 171854 460338
rect 171234 424658 171266 424894
rect 171502 424658 171586 424894
rect 171822 424658 171854 424894
rect 171234 424574 171854 424658
rect 171234 424338 171266 424574
rect 171502 424338 171586 424574
rect 171822 424338 171854 424574
rect 171234 388894 171854 424338
rect 171234 388658 171266 388894
rect 171502 388658 171586 388894
rect 171822 388658 171854 388894
rect 171234 388574 171854 388658
rect 171234 388338 171266 388574
rect 171502 388338 171586 388574
rect 171822 388338 171854 388574
rect 171234 352894 171854 388338
rect 171234 352658 171266 352894
rect 171502 352658 171586 352894
rect 171822 352658 171854 352894
rect 171234 352574 171854 352658
rect 171234 352338 171266 352574
rect 171502 352338 171586 352574
rect 171822 352338 171854 352574
rect 171234 316894 171854 352338
rect 171234 316658 171266 316894
rect 171502 316658 171586 316894
rect 171822 316658 171854 316894
rect 171234 316574 171854 316658
rect 171234 316338 171266 316574
rect 171502 316338 171586 316574
rect 171822 316338 171854 316574
rect 171234 280894 171854 316338
rect 171234 280658 171266 280894
rect 171502 280658 171586 280894
rect 171822 280658 171854 280894
rect 171234 280574 171854 280658
rect 171234 280338 171266 280574
rect 171502 280338 171586 280574
rect 171822 280338 171854 280574
rect 171234 244894 171854 280338
rect 171234 244658 171266 244894
rect 171502 244658 171586 244894
rect 171822 244658 171854 244894
rect 171234 244574 171854 244658
rect 171234 244338 171266 244574
rect 171502 244338 171586 244574
rect 171822 244338 171854 244574
rect 171234 208894 171854 244338
rect 171234 208658 171266 208894
rect 171502 208658 171586 208894
rect 171822 208658 171854 208894
rect 171234 208574 171854 208658
rect 171234 208338 171266 208574
rect 171502 208338 171586 208574
rect 171822 208338 171854 208574
rect 171234 192000 171854 208338
rect 174954 680614 175574 711002
rect 192954 710598 193574 711590
rect 192954 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 193574 710598
rect 192954 710278 193574 710362
rect 192954 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 193574 710278
rect 189234 708678 189854 709670
rect 189234 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 189854 708678
rect 189234 708358 189854 708442
rect 189234 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 189854 708358
rect 185514 706758 186134 707750
rect 185514 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 186134 706758
rect 185514 706438 186134 706522
rect 185514 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 186134 706438
rect 174954 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 175574 680614
rect 174954 680294 175574 680378
rect 174954 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 175574 680294
rect 174954 644614 175574 680058
rect 174954 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 175574 644614
rect 174954 644294 175574 644378
rect 174954 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 175574 644294
rect 174954 608614 175574 644058
rect 174954 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 175574 608614
rect 174954 608294 175574 608378
rect 174954 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 175574 608294
rect 174954 572614 175574 608058
rect 174954 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 175574 572614
rect 174954 572294 175574 572378
rect 174954 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 175574 572294
rect 174954 536614 175574 572058
rect 174954 536378 174986 536614
rect 175222 536378 175306 536614
rect 175542 536378 175574 536614
rect 174954 536294 175574 536378
rect 174954 536058 174986 536294
rect 175222 536058 175306 536294
rect 175542 536058 175574 536294
rect 174954 500614 175574 536058
rect 174954 500378 174986 500614
rect 175222 500378 175306 500614
rect 175542 500378 175574 500614
rect 174954 500294 175574 500378
rect 174954 500058 174986 500294
rect 175222 500058 175306 500294
rect 175542 500058 175574 500294
rect 174954 464614 175574 500058
rect 174954 464378 174986 464614
rect 175222 464378 175306 464614
rect 175542 464378 175574 464614
rect 174954 464294 175574 464378
rect 174954 464058 174986 464294
rect 175222 464058 175306 464294
rect 175542 464058 175574 464294
rect 174954 428614 175574 464058
rect 174954 428378 174986 428614
rect 175222 428378 175306 428614
rect 175542 428378 175574 428614
rect 174954 428294 175574 428378
rect 174954 428058 174986 428294
rect 175222 428058 175306 428294
rect 175542 428058 175574 428294
rect 174954 392614 175574 428058
rect 174954 392378 174986 392614
rect 175222 392378 175306 392614
rect 175542 392378 175574 392614
rect 174954 392294 175574 392378
rect 174954 392058 174986 392294
rect 175222 392058 175306 392294
rect 175542 392058 175574 392294
rect 174954 356614 175574 392058
rect 174954 356378 174986 356614
rect 175222 356378 175306 356614
rect 175542 356378 175574 356614
rect 174954 356294 175574 356378
rect 174954 356058 174986 356294
rect 175222 356058 175306 356294
rect 175542 356058 175574 356294
rect 174954 320614 175574 356058
rect 174954 320378 174986 320614
rect 175222 320378 175306 320614
rect 175542 320378 175574 320614
rect 174954 320294 175574 320378
rect 174954 320058 174986 320294
rect 175222 320058 175306 320294
rect 175542 320058 175574 320294
rect 174954 284614 175574 320058
rect 174954 284378 174986 284614
rect 175222 284378 175306 284614
rect 175542 284378 175574 284614
rect 174954 284294 175574 284378
rect 174954 284058 174986 284294
rect 175222 284058 175306 284294
rect 175542 284058 175574 284294
rect 174954 248614 175574 284058
rect 174954 248378 174986 248614
rect 175222 248378 175306 248614
rect 175542 248378 175574 248614
rect 174954 248294 175574 248378
rect 174954 248058 174986 248294
rect 175222 248058 175306 248294
rect 175542 248058 175574 248294
rect 174954 212614 175574 248058
rect 174954 212378 174986 212614
rect 175222 212378 175306 212614
rect 175542 212378 175574 212614
rect 174954 212294 175574 212378
rect 174954 212058 174986 212294
rect 175222 212058 175306 212294
rect 175542 212058 175574 212294
rect 162243 183454 162563 183486
rect 162243 183218 162285 183454
rect 162521 183218 162563 183454
rect 162243 183134 162563 183218
rect 162243 182898 162285 183134
rect 162521 182898 162563 183134
rect 162243 182866 162563 182898
rect 164840 183454 165160 183486
rect 164840 183218 164882 183454
rect 165118 183218 165160 183454
rect 164840 183134 165160 183218
rect 164840 182898 164882 183134
rect 165118 182898 165160 183134
rect 164840 182866 165160 182898
rect 167437 183454 167757 183486
rect 167437 183218 167479 183454
rect 167715 183218 167757 183454
rect 167437 183134 167757 183218
rect 167437 182898 167479 183134
rect 167715 182898 167757 183134
rect 167437 182866 167757 182898
rect 174954 176614 175574 212058
rect 174954 176378 174986 176614
rect 175222 176378 175306 176614
rect 175542 176378 175574 176614
rect 174954 176294 175574 176378
rect 174954 176058 174986 176294
rect 175222 176058 175306 176294
rect 175542 176058 175574 176294
rect 163541 165454 163861 165486
rect 163541 165218 163583 165454
rect 163819 165218 163861 165454
rect 163541 165134 163861 165218
rect 163541 164898 163583 165134
rect 163819 164898 163861 165134
rect 163541 164866 163861 164898
rect 166138 165454 166458 165486
rect 166138 165218 166180 165454
rect 166416 165218 166458 165454
rect 166138 165134 166458 165218
rect 166138 164898 166180 165134
rect 166416 164898 166458 165134
rect 166138 164866 166458 164898
rect 156954 158378 156986 158614
rect 157222 158378 157306 158614
rect 157542 158378 157574 158614
rect 156954 158294 157574 158378
rect 156954 158058 156986 158294
rect 157222 158058 157306 158294
rect 157542 158058 157574 158294
rect 156954 122614 157574 158058
rect 163794 156000 164414 158000
rect 167514 156000 168134 158000
rect 171234 156000 171854 158000
rect 162243 147454 162563 147486
rect 162243 147218 162285 147454
rect 162521 147218 162563 147454
rect 162243 147134 162563 147218
rect 162243 146898 162285 147134
rect 162521 146898 162563 147134
rect 162243 146866 162563 146898
rect 164840 147454 165160 147486
rect 164840 147218 164882 147454
rect 165118 147218 165160 147454
rect 164840 147134 165160 147218
rect 164840 146898 164882 147134
rect 165118 146898 165160 147134
rect 164840 146866 165160 146898
rect 167437 147454 167757 147486
rect 167437 147218 167479 147454
rect 167715 147218 167757 147454
rect 167437 147134 167757 147218
rect 167437 146898 167479 147134
rect 167715 146898 167757 147134
rect 167437 146866 167757 146898
rect 174954 140614 175574 176058
rect 174954 140378 174986 140614
rect 175222 140378 175306 140614
rect 175542 140378 175574 140614
rect 174954 140294 175574 140378
rect 174954 140058 174986 140294
rect 175222 140058 175306 140294
rect 175542 140058 175574 140294
rect 163541 129454 163861 129486
rect 163541 129218 163583 129454
rect 163819 129218 163861 129454
rect 163541 129134 163861 129218
rect 163541 128898 163583 129134
rect 163819 128898 163861 129134
rect 163541 128866 163861 128898
rect 166138 129454 166458 129486
rect 166138 129218 166180 129454
rect 166416 129218 166458 129454
rect 166138 129134 166458 129218
rect 166138 128898 166180 129134
rect 166416 128898 166458 129134
rect 166138 128866 166458 128898
rect 156954 122378 156986 122614
rect 157222 122378 157306 122614
rect 157542 122378 157574 122614
rect 156954 122294 157574 122378
rect 156954 122058 156986 122294
rect 157222 122058 157306 122294
rect 157542 122058 157574 122294
rect 156954 86614 157574 122058
rect 156954 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 157574 86614
rect 156954 86294 157574 86378
rect 156954 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 157574 86294
rect 156954 50614 157574 86058
rect 156954 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 157574 50614
rect 156954 50294 157574 50378
rect 156954 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 157574 50294
rect 156954 14614 157574 50058
rect 156954 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 157574 14614
rect 156954 14294 157574 14378
rect 156954 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 157574 14294
rect 138954 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 139574 -7066
rect 138954 -7386 139574 -7302
rect 138954 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 139574 -7386
rect 138954 -7654 139574 -7622
rect 156954 -6106 157574 14058
rect 163794 93454 164414 122000
rect 163794 93218 163826 93454
rect 164062 93218 164146 93454
rect 164382 93218 164414 93454
rect 163794 93134 164414 93218
rect 163794 92898 163826 93134
rect 164062 92898 164146 93134
rect 164382 92898 164414 93134
rect 163794 57454 164414 92898
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -1306 164414 20898
rect 163794 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 164414 -1306
rect 163794 -1626 164414 -1542
rect 163794 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 164414 -1626
rect 163794 -1894 164414 -1862
rect 167514 97174 168134 122000
rect 167514 96938 167546 97174
rect 167782 96938 167866 97174
rect 168102 96938 168134 97174
rect 167514 96854 168134 96938
rect 167514 96618 167546 96854
rect 167782 96618 167866 96854
rect 168102 96618 168134 96854
rect 167514 61174 168134 96618
rect 167514 60938 167546 61174
rect 167782 60938 167866 61174
rect 168102 60938 168134 61174
rect 167514 60854 168134 60938
rect 167514 60618 167546 60854
rect 167782 60618 167866 60854
rect 168102 60618 168134 60854
rect 167514 25174 168134 60618
rect 167514 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 168134 25174
rect 167514 24854 168134 24938
rect 167514 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 168134 24854
rect 167514 -3226 168134 24618
rect 167514 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 168134 -3226
rect 167514 -3546 168134 -3462
rect 167514 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 168134 -3546
rect 167514 -3814 168134 -3782
rect 171234 100894 171854 122000
rect 171234 100658 171266 100894
rect 171502 100658 171586 100894
rect 171822 100658 171854 100894
rect 171234 100574 171854 100658
rect 171234 100338 171266 100574
rect 171502 100338 171586 100574
rect 171822 100338 171854 100574
rect 171234 64894 171854 100338
rect 171234 64658 171266 64894
rect 171502 64658 171586 64894
rect 171822 64658 171854 64894
rect 171234 64574 171854 64658
rect 171234 64338 171266 64574
rect 171502 64338 171586 64574
rect 171822 64338 171854 64574
rect 171234 28894 171854 64338
rect 171234 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 171854 28894
rect 171234 28574 171854 28658
rect 171234 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 171854 28574
rect 171234 -5146 171854 28338
rect 171234 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 171854 -5146
rect 171234 -5466 171854 -5382
rect 171234 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 171854 -5466
rect 171234 -5734 171854 -5702
rect 174954 104614 175574 140058
rect 174954 104378 174986 104614
rect 175222 104378 175306 104614
rect 175542 104378 175574 104614
rect 174954 104294 175574 104378
rect 174954 104058 174986 104294
rect 175222 104058 175306 104294
rect 175542 104058 175574 104294
rect 174954 68614 175574 104058
rect 174954 68378 174986 68614
rect 175222 68378 175306 68614
rect 175542 68378 175574 68614
rect 174954 68294 175574 68378
rect 174954 68058 174986 68294
rect 175222 68058 175306 68294
rect 175542 68058 175574 68294
rect 174954 32614 175574 68058
rect 174954 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 175574 32614
rect 174954 32294 175574 32378
rect 174954 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 175574 32294
rect 156954 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 157574 -6106
rect 156954 -6426 157574 -6342
rect 156954 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 157574 -6426
rect 156954 -7654 157574 -6662
rect 174954 -7066 175574 32058
rect 181794 704838 182414 705830
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 543454 182414 578898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 507454 182414 542898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 181794 471454 182414 506898
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 181794 435454 182414 470898
rect 181794 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 182414 435454
rect 181794 435134 182414 435218
rect 181794 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 182414 435134
rect 181794 399454 182414 434898
rect 181794 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 182414 399454
rect 181794 399134 182414 399218
rect 181794 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 182414 399134
rect 181794 363454 182414 398898
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 181794 327454 182414 362898
rect 181794 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 182414 327454
rect 181794 327134 182414 327218
rect 181794 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 182414 327134
rect 181794 291454 182414 326898
rect 181794 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 182414 291454
rect 181794 291134 182414 291218
rect 181794 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 182414 291134
rect 181794 255454 182414 290898
rect 181794 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 182414 255454
rect 181794 255134 182414 255218
rect 181794 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 182414 255134
rect 181794 219454 182414 254898
rect 181794 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 182414 219454
rect 181794 219134 182414 219218
rect 181794 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 182414 219134
rect 181794 183454 182414 218898
rect 181794 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 182414 183454
rect 181794 183134 182414 183218
rect 181794 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 182414 183134
rect 181794 147454 182414 182898
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 111454 182414 146898
rect 181794 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 182414 111454
rect 181794 111134 182414 111218
rect 181794 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 182414 111134
rect 181794 75454 182414 110898
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 181794 39454 182414 74898
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -1894 182414 -902
rect 185514 691174 186134 706202
rect 185514 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 186134 691174
rect 185514 690854 186134 690938
rect 185514 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 186134 690854
rect 185514 655174 186134 690618
rect 185514 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 186134 655174
rect 185514 654854 186134 654938
rect 185514 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 186134 654854
rect 185514 619174 186134 654618
rect 185514 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 186134 619174
rect 185514 618854 186134 618938
rect 185514 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 186134 618854
rect 185514 583174 186134 618618
rect 185514 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 186134 583174
rect 185514 582854 186134 582938
rect 185514 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 186134 582854
rect 185514 547174 186134 582618
rect 185514 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 186134 547174
rect 185514 546854 186134 546938
rect 185514 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 186134 546854
rect 185514 511174 186134 546618
rect 185514 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 186134 511174
rect 185514 510854 186134 510938
rect 185514 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 186134 510854
rect 185514 475174 186134 510618
rect 185514 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 186134 475174
rect 185514 474854 186134 474938
rect 185514 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 186134 474854
rect 185514 439174 186134 474618
rect 185514 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 186134 439174
rect 185514 438854 186134 438938
rect 185514 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 186134 438854
rect 185514 403174 186134 438618
rect 185514 402938 185546 403174
rect 185782 402938 185866 403174
rect 186102 402938 186134 403174
rect 185514 402854 186134 402938
rect 185514 402618 185546 402854
rect 185782 402618 185866 402854
rect 186102 402618 186134 402854
rect 185514 367174 186134 402618
rect 185514 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 186134 367174
rect 185514 366854 186134 366938
rect 185514 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 186134 366854
rect 185514 331174 186134 366618
rect 185514 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 186134 331174
rect 185514 330854 186134 330938
rect 185514 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 186134 330854
rect 185514 295174 186134 330618
rect 185514 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 186134 295174
rect 185514 294854 186134 294938
rect 185514 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 186134 294854
rect 185514 259174 186134 294618
rect 185514 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 186134 259174
rect 185514 258854 186134 258938
rect 185514 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 186134 258854
rect 185514 223174 186134 258618
rect 185514 222938 185546 223174
rect 185782 222938 185866 223174
rect 186102 222938 186134 223174
rect 185514 222854 186134 222938
rect 185514 222618 185546 222854
rect 185782 222618 185866 222854
rect 186102 222618 186134 222854
rect 185514 187174 186134 222618
rect 185514 186938 185546 187174
rect 185782 186938 185866 187174
rect 186102 186938 186134 187174
rect 185514 186854 186134 186938
rect 185514 186618 185546 186854
rect 185782 186618 185866 186854
rect 186102 186618 186134 186854
rect 185514 151174 186134 186618
rect 185514 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 186134 151174
rect 185514 150854 186134 150938
rect 185514 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 186134 150854
rect 185514 115174 186134 150618
rect 185514 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 186134 115174
rect 185514 114854 186134 114938
rect 185514 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 186134 114854
rect 185514 79174 186134 114618
rect 185514 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 186134 79174
rect 185514 78854 186134 78938
rect 185514 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 186134 78854
rect 185514 43174 186134 78618
rect 185514 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 186134 43174
rect 185514 42854 186134 42938
rect 185514 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 186134 42854
rect 185514 7174 186134 42618
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 185514 -2266 186134 6618
rect 185514 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 186134 -2266
rect 185514 -2586 186134 -2502
rect 185514 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 186134 -2586
rect 185514 -3814 186134 -2822
rect 189234 694894 189854 708122
rect 189234 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 189854 694894
rect 189234 694574 189854 694658
rect 189234 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 189854 694574
rect 189234 658894 189854 694338
rect 189234 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 189854 658894
rect 189234 658574 189854 658658
rect 189234 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 189854 658574
rect 189234 622894 189854 658338
rect 189234 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 189854 622894
rect 189234 622574 189854 622658
rect 189234 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 189854 622574
rect 189234 586894 189854 622338
rect 189234 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 189854 586894
rect 189234 586574 189854 586658
rect 189234 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 189854 586574
rect 189234 550894 189854 586338
rect 189234 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 189854 550894
rect 189234 550574 189854 550658
rect 189234 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 189854 550574
rect 189234 514894 189854 550338
rect 189234 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 189854 514894
rect 189234 514574 189854 514658
rect 189234 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 189854 514574
rect 189234 478894 189854 514338
rect 189234 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 189854 478894
rect 189234 478574 189854 478658
rect 189234 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 189854 478574
rect 189234 442894 189854 478338
rect 189234 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 189854 442894
rect 189234 442574 189854 442658
rect 189234 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 189854 442574
rect 189234 406894 189854 442338
rect 189234 406658 189266 406894
rect 189502 406658 189586 406894
rect 189822 406658 189854 406894
rect 189234 406574 189854 406658
rect 189234 406338 189266 406574
rect 189502 406338 189586 406574
rect 189822 406338 189854 406574
rect 189234 370894 189854 406338
rect 189234 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 189854 370894
rect 189234 370574 189854 370658
rect 189234 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 189854 370574
rect 189234 334894 189854 370338
rect 189234 334658 189266 334894
rect 189502 334658 189586 334894
rect 189822 334658 189854 334894
rect 189234 334574 189854 334658
rect 189234 334338 189266 334574
rect 189502 334338 189586 334574
rect 189822 334338 189854 334574
rect 189234 298894 189854 334338
rect 189234 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 189854 298894
rect 189234 298574 189854 298658
rect 189234 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 189854 298574
rect 189234 262894 189854 298338
rect 189234 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 189854 262894
rect 189234 262574 189854 262658
rect 189234 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 189854 262574
rect 189234 226894 189854 262338
rect 189234 226658 189266 226894
rect 189502 226658 189586 226894
rect 189822 226658 189854 226894
rect 189234 226574 189854 226658
rect 189234 226338 189266 226574
rect 189502 226338 189586 226574
rect 189822 226338 189854 226574
rect 189234 190894 189854 226338
rect 189234 190658 189266 190894
rect 189502 190658 189586 190894
rect 189822 190658 189854 190894
rect 189234 190574 189854 190658
rect 189234 190338 189266 190574
rect 189502 190338 189586 190574
rect 189822 190338 189854 190574
rect 189234 154894 189854 190338
rect 189234 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 189854 154894
rect 189234 154574 189854 154658
rect 189234 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 189854 154574
rect 189234 118894 189854 154338
rect 189234 118658 189266 118894
rect 189502 118658 189586 118894
rect 189822 118658 189854 118894
rect 189234 118574 189854 118658
rect 189234 118338 189266 118574
rect 189502 118338 189586 118574
rect 189822 118338 189854 118574
rect 189234 82894 189854 118338
rect 189234 82658 189266 82894
rect 189502 82658 189586 82894
rect 189822 82658 189854 82894
rect 189234 82574 189854 82658
rect 189234 82338 189266 82574
rect 189502 82338 189586 82574
rect 189822 82338 189854 82574
rect 189234 46894 189854 82338
rect 189234 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 189854 46894
rect 189234 46574 189854 46658
rect 189234 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 189854 46574
rect 189234 10894 189854 46338
rect 189234 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 189854 10894
rect 189234 10574 189854 10658
rect 189234 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 189854 10574
rect 189234 -4186 189854 10338
rect 189234 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 189854 -4186
rect 189234 -4506 189854 -4422
rect 189234 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 189854 -4506
rect 189234 -5734 189854 -4742
rect 192954 698614 193574 710042
rect 210954 711558 211574 711590
rect 210954 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 211574 711558
rect 210954 711238 211574 711322
rect 210954 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 211574 711238
rect 207234 709638 207854 709670
rect 207234 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 207854 709638
rect 207234 709318 207854 709402
rect 207234 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 207854 709318
rect 203514 707718 204134 707750
rect 203514 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 204134 707718
rect 203514 707398 204134 707482
rect 203514 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 204134 707398
rect 192954 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 193574 698614
rect 192954 698294 193574 698378
rect 192954 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 193574 698294
rect 192954 662614 193574 698058
rect 192954 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 193574 662614
rect 192954 662294 193574 662378
rect 192954 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 193574 662294
rect 192954 626614 193574 662058
rect 192954 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 193574 626614
rect 192954 626294 193574 626378
rect 192954 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 193574 626294
rect 192954 590614 193574 626058
rect 192954 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 193574 590614
rect 192954 590294 193574 590378
rect 192954 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 193574 590294
rect 192954 554614 193574 590058
rect 192954 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 193574 554614
rect 192954 554294 193574 554378
rect 192954 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 193574 554294
rect 192954 518614 193574 554058
rect 192954 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 193574 518614
rect 192954 518294 193574 518378
rect 192954 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 193574 518294
rect 192954 482614 193574 518058
rect 192954 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 193574 482614
rect 192954 482294 193574 482378
rect 192954 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 193574 482294
rect 192954 446614 193574 482058
rect 192954 446378 192986 446614
rect 193222 446378 193306 446614
rect 193542 446378 193574 446614
rect 192954 446294 193574 446378
rect 192954 446058 192986 446294
rect 193222 446058 193306 446294
rect 193542 446058 193574 446294
rect 192954 410614 193574 446058
rect 192954 410378 192986 410614
rect 193222 410378 193306 410614
rect 193542 410378 193574 410614
rect 192954 410294 193574 410378
rect 192954 410058 192986 410294
rect 193222 410058 193306 410294
rect 193542 410058 193574 410294
rect 192954 374614 193574 410058
rect 192954 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 193574 374614
rect 192954 374294 193574 374378
rect 192954 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 193574 374294
rect 192954 338614 193574 374058
rect 192954 338378 192986 338614
rect 193222 338378 193306 338614
rect 193542 338378 193574 338614
rect 192954 338294 193574 338378
rect 192954 338058 192986 338294
rect 193222 338058 193306 338294
rect 193542 338058 193574 338294
rect 192954 302614 193574 338058
rect 192954 302378 192986 302614
rect 193222 302378 193306 302614
rect 193542 302378 193574 302614
rect 192954 302294 193574 302378
rect 192954 302058 192986 302294
rect 193222 302058 193306 302294
rect 193542 302058 193574 302294
rect 192954 266614 193574 302058
rect 199794 705798 200414 705830
rect 199794 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 200414 705798
rect 199794 705478 200414 705562
rect 199794 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 200414 705478
rect 199794 669454 200414 705242
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 561454 200414 596898
rect 199794 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 200414 561454
rect 199794 561134 200414 561218
rect 199794 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 200414 561134
rect 199794 525454 200414 560898
rect 199794 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 200414 525454
rect 199794 525134 200414 525218
rect 199794 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 200414 525134
rect 199794 489454 200414 524898
rect 199794 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 200414 489454
rect 199794 489134 200414 489218
rect 199794 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 200414 489134
rect 199794 453454 200414 488898
rect 199794 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 200414 453454
rect 199794 453134 200414 453218
rect 199794 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 200414 453134
rect 199794 417454 200414 452898
rect 199794 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 200414 417454
rect 199794 417134 200414 417218
rect 199794 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 200414 417134
rect 199794 381454 200414 416898
rect 199794 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 200414 381454
rect 199794 381134 200414 381218
rect 199794 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 200414 381134
rect 199794 345454 200414 380898
rect 199794 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 200414 345454
rect 199794 345134 200414 345218
rect 199794 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 200414 345134
rect 199794 309454 200414 344898
rect 199794 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 200414 309454
rect 199794 309134 200414 309218
rect 199794 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 200414 309134
rect 199794 302000 200414 308898
rect 203514 673174 204134 707162
rect 203514 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 204134 673174
rect 203514 672854 204134 672938
rect 203514 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 204134 672854
rect 203514 637174 204134 672618
rect 203514 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 204134 637174
rect 203514 636854 204134 636938
rect 203514 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 204134 636854
rect 203514 601174 204134 636618
rect 203514 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 204134 601174
rect 203514 600854 204134 600938
rect 203514 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 204134 600854
rect 203514 565174 204134 600618
rect 203514 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 204134 565174
rect 203514 564854 204134 564938
rect 203514 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 204134 564854
rect 203514 529174 204134 564618
rect 203514 528938 203546 529174
rect 203782 528938 203866 529174
rect 204102 528938 204134 529174
rect 203514 528854 204134 528938
rect 203514 528618 203546 528854
rect 203782 528618 203866 528854
rect 204102 528618 204134 528854
rect 203514 493174 204134 528618
rect 203514 492938 203546 493174
rect 203782 492938 203866 493174
rect 204102 492938 204134 493174
rect 203514 492854 204134 492938
rect 203514 492618 203546 492854
rect 203782 492618 203866 492854
rect 204102 492618 204134 492854
rect 203514 457174 204134 492618
rect 203514 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 204134 457174
rect 203514 456854 204134 456938
rect 203514 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 204134 456854
rect 203514 421174 204134 456618
rect 203514 420938 203546 421174
rect 203782 420938 203866 421174
rect 204102 420938 204134 421174
rect 203514 420854 204134 420938
rect 203514 420618 203546 420854
rect 203782 420618 203866 420854
rect 204102 420618 204134 420854
rect 203514 385174 204134 420618
rect 203514 384938 203546 385174
rect 203782 384938 203866 385174
rect 204102 384938 204134 385174
rect 203514 384854 204134 384938
rect 203514 384618 203546 384854
rect 203782 384618 203866 384854
rect 204102 384618 204134 384854
rect 203514 349174 204134 384618
rect 203514 348938 203546 349174
rect 203782 348938 203866 349174
rect 204102 348938 204134 349174
rect 203514 348854 204134 348938
rect 203514 348618 203546 348854
rect 203782 348618 203866 348854
rect 204102 348618 204134 348854
rect 203514 313174 204134 348618
rect 203514 312938 203546 313174
rect 203782 312938 203866 313174
rect 204102 312938 204134 313174
rect 203514 312854 204134 312938
rect 203514 312618 203546 312854
rect 203782 312618 203866 312854
rect 204102 312618 204134 312854
rect 203514 302000 204134 312618
rect 207234 676894 207854 709082
rect 207234 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 207854 676894
rect 207234 676574 207854 676658
rect 207234 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 207854 676574
rect 207234 640894 207854 676338
rect 207234 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 207854 640894
rect 207234 640574 207854 640658
rect 207234 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 207854 640574
rect 207234 604894 207854 640338
rect 207234 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 207854 604894
rect 207234 604574 207854 604658
rect 207234 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 207854 604574
rect 207234 568894 207854 604338
rect 207234 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 207854 568894
rect 207234 568574 207854 568658
rect 207234 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 207854 568574
rect 207234 532894 207854 568338
rect 207234 532658 207266 532894
rect 207502 532658 207586 532894
rect 207822 532658 207854 532894
rect 207234 532574 207854 532658
rect 207234 532338 207266 532574
rect 207502 532338 207586 532574
rect 207822 532338 207854 532574
rect 207234 496894 207854 532338
rect 207234 496658 207266 496894
rect 207502 496658 207586 496894
rect 207822 496658 207854 496894
rect 207234 496574 207854 496658
rect 207234 496338 207266 496574
rect 207502 496338 207586 496574
rect 207822 496338 207854 496574
rect 207234 460894 207854 496338
rect 207234 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 207854 460894
rect 207234 460574 207854 460658
rect 207234 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 207854 460574
rect 207234 424894 207854 460338
rect 207234 424658 207266 424894
rect 207502 424658 207586 424894
rect 207822 424658 207854 424894
rect 207234 424574 207854 424658
rect 207234 424338 207266 424574
rect 207502 424338 207586 424574
rect 207822 424338 207854 424574
rect 207234 388894 207854 424338
rect 207234 388658 207266 388894
rect 207502 388658 207586 388894
rect 207822 388658 207854 388894
rect 207234 388574 207854 388658
rect 207234 388338 207266 388574
rect 207502 388338 207586 388574
rect 207822 388338 207854 388574
rect 207234 352894 207854 388338
rect 207234 352658 207266 352894
rect 207502 352658 207586 352894
rect 207822 352658 207854 352894
rect 207234 352574 207854 352658
rect 207234 352338 207266 352574
rect 207502 352338 207586 352574
rect 207822 352338 207854 352574
rect 207234 316894 207854 352338
rect 207234 316658 207266 316894
rect 207502 316658 207586 316894
rect 207822 316658 207854 316894
rect 207234 316574 207854 316658
rect 207234 316338 207266 316574
rect 207502 316338 207586 316574
rect 207822 316338 207854 316574
rect 207234 302000 207854 316338
rect 210954 680614 211574 711002
rect 228954 710598 229574 711590
rect 228954 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 229574 710598
rect 228954 710278 229574 710362
rect 228954 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 229574 710278
rect 225234 708678 225854 709670
rect 225234 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 225854 708678
rect 225234 708358 225854 708442
rect 225234 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 225854 708358
rect 221514 706758 222134 707750
rect 221514 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 222134 706758
rect 221514 706438 222134 706522
rect 221514 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 222134 706438
rect 210954 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 211574 680614
rect 210954 680294 211574 680378
rect 210954 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 211574 680294
rect 210954 644614 211574 680058
rect 210954 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 211574 644614
rect 210954 644294 211574 644378
rect 210954 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 211574 644294
rect 210954 608614 211574 644058
rect 210954 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 211574 608614
rect 210954 608294 211574 608378
rect 210954 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 211574 608294
rect 210954 572614 211574 608058
rect 210954 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 211574 572614
rect 210954 572294 211574 572378
rect 210954 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 211574 572294
rect 210954 536614 211574 572058
rect 210954 536378 210986 536614
rect 211222 536378 211306 536614
rect 211542 536378 211574 536614
rect 210954 536294 211574 536378
rect 210954 536058 210986 536294
rect 211222 536058 211306 536294
rect 211542 536058 211574 536294
rect 210954 500614 211574 536058
rect 210954 500378 210986 500614
rect 211222 500378 211306 500614
rect 211542 500378 211574 500614
rect 210954 500294 211574 500378
rect 210954 500058 210986 500294
rect 211222 500058 211306 500294
rect 211542 500058 211574 500294
rect 210954 464614 211574 500058
rect 210954 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 211574 464614
rect 210954 464294 211574 464378
rect 210954 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 211574 464294
rect 210954 428614 211574 464058
rect 210954 428378 210986 428614
rect 211222 428378 211306 428614
rect 211542 428378 211574 428614
rect 210954 428294 211574 428378
rect 210954 428058 210986 428294
rect 211222 428058 211306 428294
rect 211542 428058 211574 428294
rect 210954 392614 211574 428058
rect 210954 392378 210986 392614
rect 211222 392378 211306 392614
rect 211542 392378 211574 392614
rect 210954 392294 211574 392378
rect 210954 392058 210986 392294
rect 211222 392058 211306 392294
rect 211542 392058 211574 392294
rect 210954 356614 211574 392058
rect 210954 356378 210986 356614
rect 211222 356378 211306 356614
rect 211542 356378 211574 356614
rect 210954 356294 211574 356378
rect 210954 356058 210986 356294
rect 211222 356058 211306 356294
rect 211542 356058 211574 356294
rect 210954 320614 211574 356058
rect 210954 320378 210986 320614
rect 211222 320378 211306 320614
rect 211542 320378 211574 320614
rect 210954 320294 211574 320378
rect 210954 320058 210986 320294
rect 211222 320058 211306 320294
rect 211542 320058 211574 320294
rect 210954 302000 211574 320058
rect 217794 704838 218414 705830
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 543454 218414 578898
rect 217794 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 218414 543454
rect 217794 543134 218414 543218
rect 217794 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 218414 543134
rect 217794 507454 218414 542898
rect 217794 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 218414 507454
rect 217794 507134 218414 507218
rect 217794 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 218414 507134
rect 217794 471454 218414 506898
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 217794 435454 218414 470898
rect 217794 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 218414 435454
rect 217794 435134 218414 435218
rect 217794 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 218414 435134
rect 217794 399454 218414 434898
rect 217794 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 218414 399454
rect 217794 399134 218414 399218
rect 217794 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 218414 399134
rect 217794 363454 218414 398898
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 217794 327454 218414 362898
rect 217794 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 218414 327454
rect 217794 327134 218414 327218
rect 217794 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 218414 327134
rect 217794 302000 218414 326898
rect 221514 691174 222134 706202
rect 221514 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 222134 691174
rect 221514 690854 222134 690938
rect 221514 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 222134 690854
rect 221514 655174 222134 690618
rect 221514 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 222134 655174
rect 221514 654854 222134 654938
rect 221514 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 222134 654854
rect 221514 619174 222134 654618
rect 221514 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 222134 619174
rect 221514 618854 222134 618938
rect 221514 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 222134 618854
rect 221514 583174 222134 618618
rect 221514 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 222134 583174
rect 221514 582854 222134 582938
rect 221514 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 222134 582854
rect 221514 547174 222134 582618
rect 221514 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 222134 547174
rect 221514 546854 222134 546938
rect 221514 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 222134 546854
rect 221514 511174 222134 546618
rect 221514 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 222134 511174
rect 221514 510854 222134 510938
rect 221514 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 222134 510854
rect 221514 475174 222134 510618
rect 221514 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 222134 475174
rect 221514 474854 222134 474938
rect 221514 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 222134 474854
rect 221514 439174 222134 474618
rect 221514 438938 221546 439174
rect 221782 438938 221866 439174
rect 222102 438938 222134 439174
rect 221514 438854 222134 438938
rect 221514 438618 221546 438854
rect 221782 438618 221866 438854
rect 222102 438618 222134 438854
rect 221514 403174 222134 438618
rect 221514 402938 221546 403174
rect 221782 402938 221866 403174
rect 222102 402938 222134 403174
rect 221514 402854 222134 402938
rect 221514 402618 221546 402854
rect 221782 402618 221866 402854
rect 222102 402618 222134 402854
rect 221514 367174 222134 402618
rect 221514 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 222134 367174
rect 221514 366854 222134 366938
rect 221514 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 222134 366854
rect 221514 331174 222134 366618
rect 221514 330938 221546 331174
rect 221782 330938 221866 331174
rect 222102 330938 222134 331174
rect 221514 330854 222134 330938
rect 221514 330618 221546 330854
rect 221782 330618 221866 330854
rect 222102 330618 222134 330854
rect 221514 302000 222134 330618
rect 225234 694894 225854 708122
rect 225234 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 225854 694894
rect 225234 694574 225854 694658
rect 225234 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 225854 694574
rect 225234 658894 225854 694338
rect 225234 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 225854 658894
rect 225234 658574 225854 658658
rect 225234 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 225854 658574
rect 225234 622894 225854 658338
rect 225234 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 225854 622894
rect 225234 622574 225854 622658
rect 225234 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 225854 622574
rect 225234 586894 225854 622338
rect 225234 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 225854 586894
rect 225234 586574 225854 586658
rect 225234 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 225854 586574
rect 225234 550894 225854 586338
rect 225234 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 225854 550894
rect 225234 550574 225854 550658
rect 225234 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 225854 550574
rect 225234 514894 225854 550338
rect 225234 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 225854 514894
rect 225234 514574 225854 514658
rect 225234 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 225854 514574
rect 225234 478894 225854 514338
rect 225234 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 225854 478894
rect 225234 478574 225854 478658
rect 225234 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 225854 478574
rect 225234 442894 225854 478338
rect 225234 442658 225266 442894
rect 225502 442658 225586 442894
rect 225822 442658 225854 442894
rect 225234 442574 225854 442658
rect 225234 442338 225266 442574
rect 225502 442338 225586 442574
rect 225822 442338 225854 442574
rect 225234 406894 225854 442338
rect 225234 406658 225266 406894
rect 225502 406658 225586 406894
rect 225822 406658 225854 406894
rect 225234 406574 225854 406658
rect 225234 406338 225266 406574
rect 225502 406338 225586 406574
rect 225822 406338 225854 406574
rect 225234 370894 225854 406338
rect 225234 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 225854 370894
rect 225234 370574 225854 370658
rect 225234 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 225854 370574
rect 225234 334894 225854 370338
rect 225234 334658 225266 334894
rect 225502 334658 225586 334894
rect 225822 334658 225854 334894
rect 225234 334574 225854 334658
rect 225234 334338 225266 334574
rect 225502 334338 225586 334574
rect 225822 334338 225854 334574
rect 225234 302000 225854 334338
rect 228954 698614 229574 710042
rect 246954 711558 247574 711590
rect 246954 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 247574 711558
rect 246954 711238 247574 711322
rect 246954 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 247574 711238
rect 243234 709638 243854 709670
rect 243234 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 243854 709638
rect 243234 709318 243854 709402
rect 243234 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 243854 709318
rect 239514 707718 240134 707750
rect 239514 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 240134 707718
rect 239514 707398 240134 707482
rect 239514 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 240134 707398
rect 228954 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 229574 698614
rect 228954 698294 229574 698378
rect 228954 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 229574 698294
rect 228954 662614 229574 698058
rect 228954 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 229574 662614
rect 228954 662294 229574 662378
rect 228954 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 229574 662294
rect 228954 626614 229574 662058
rect 228954 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 229574 626614
rect 228954 626294 229574 626378
rect 228954 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 229574 626294
rect 228954 590614 229574 626058
rect 228954 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 229574 590614
rect 228954 590294 229574 590378
rect 228954 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 229574 590294
rect 228954 554614 229574 590058
rect 228954 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 229574 554614
rect 228954 554294 229574 554378
rect 228954 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 229574 554294
rect 228954 518614 229574 554058
rect 228954 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 229574 518614
rect 228954 518294 229574 518378
rect 228954 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 229574 518294
rect 228954 482614 229574 518058
rect 228954 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 229574 482614
rect 228954 482294 229574 482378
rect 228954 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 229574 482294
rect 228954 446614 229574 482058
rect 228954 446378 228986 446614
rect 229222 446378 229306 446614
rect 229542 446378 229574 446614
rect 228954 446294 229574 446378
rect 228954 446058 228986 446294
rect 229222 446058 229306 446294
rect 229542 446058 229574 446294
rect 228954 410614 229574 446058
rect 228954 410378 228986 410614
rect 229222 410378 229306 410614
rect 229542 410378 229574 410614
rect 228954 410294 229574 410378
rect 228954 410058 228986 410294
rect 229222 410058 229306 410294
rect 229542 410058 229574 410294
rect 228954 374614 229574 410058
rect 228954 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 229574 374614
rect 228954 374294 229574 374378
rect 228954 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 229574 374294
rect 228954 338614 229574 374058
rect 228954 338378 228986 338614
rect 229222 338378 229306 338614
rect 229542 338378 229574 338614
rect 228954 338294 229574 338378
rect 228954 338058 228986 338294
rect 229222 338058 229306 338294
rect 229542 338058 229574 338294
rect 228954 302614 229574 338058
rect 228954 302378 228986 302614
rect 229222 302378 229306 302614
rect 229542 302378 229574 302614
rect 228954 302294 229574 302378
rect 228954 302058 228986 302294
rect 229222 302058 229306 302294
rect 229542 302058 229574 302294
rect 228954 302000 229574 302058
rect 235794 705798 236414 705830
rect 235794 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 236414 705798
rect 235794 705478 236414 705562
rect 235794 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 236414 705478
rect 235794 669454 236414 705242
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 597454 236414 632898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 561454 236414 596898
rect 235794 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 236414 561454
rect 235794 561134 236414 561218
rect 235794 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 236414 561134
rect 235794 525454 236414 560898
rect 235794 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 236414 525454
rect 235794 525134 236414 525218
rect 235794 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 236414 525134
rect 235794 489454 236414 524898
rect 235794 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 236414 489454
rect 235794 489134 236414 489218
rect 235794 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 236414 489134
rect 235794 453454 236414 488898
rect 235794 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 236414 453454
rect 235794 453134 236414 453218
rect 235794 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 236414 453134
rect 235794 417454 236414 452898
rect 235794 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 236414 417454
rect 235794 417134 236414 417218
rect 235794 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 236414 417134
rect 235794 381454 236414 416898
rect 235794 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 236414 381454
rect 235794 381134 236414 381218
rect 235794 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 236414 381134
rect 235794 345454 236414 380898
rect 235794 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 236414 345454
rect 235794 345134 236414 345218
rect 235794 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 236414 345134
rect 235794 309454 236414 344898
rect 235794 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 236414 309454
rect 235794 309134 236414 309218
rect 235794 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 236414 309134
rect 235794 302000 236414 308898
rect 239514 673174 240134 707162
rect 239514 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 240134 673174
rect 239514 672854 240134 672938
rect 239514 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 240134 672854
rect 239514 637174 240134 672618
rect 239514 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 240134 637174
rect 239514 636854 240134 636938
rect 239514 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 240134 636854
rect 239514 601174 240134 636618
rect 239514 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 240134 601174
rect 239514 600854 240134 600938
rect 239514 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 240134 600854
rect 239514 565174 240134 600618
rect 239514 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 240134 565174
rect 239514 564854 240134 564938
rect 239514 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 240134 564854
rect 239514 529174 240134 564618
rect 239514 528938 239546 529174
rect 239782 528938 239866 529174
rect 240102 528938 240134 529174
rect 239514 528854 240134 528938
rect 239514 528618 239546 528854
rect 239782 528618 239866 528854
rect 240102 528618 240134 528854
rect 239514 493174 240134 528618
rect 239514 492938 239546 493174
rect 239782 492938 239866 493174
rect 240102 492938 240134 493174
rect 239514 492854 240134 492938
rect 239514 492618 239546 492854
rect 239782 492618 239866 492854
rect 240102 492618 240134 492854
rect 239514 457174 240134 492618
rect 239514 456938 239546 457174
rect 239782 456938 239866 457174
rect 240102 456938 240134 457174
rect 239514 456854 240134 456938
rect 239514 456618 239546 456854
rect 239782 456618 239866 456854
rect 240102 456618 240134 456854
rect 239514 421174 240134 456618
rect 239514 420938 239546 421174
rect 239782 420938 239866 421174
rect 240102 420938 240134 421174
rect 239514 420854 240134 420938
rect 239514 420618 239546 420854
rect 239782 420618 239866 420854
rect 240102 420618 240134 420854
rect 239514 385174 240134 420618
rect 239514 384938 239546 385174
rect 239782 384938 239866 385174
rect 240102 384938 240134 385174
rect 239514 384854 240134 384938
rect 239514 384618 239546 384854
rect 239782 384618 239866 384854
rect 240102 384618 240134 384854
rect 239514 349174 240134 384618
rect 239514 348938 239546 349174
rect 239782 348938 239866 349174
rect 240102 348938 240134 349174
rect 239514 348854 240134 348938
rect 239514 348618 239546 348854
rect 239782 348618 239866 348854
rect 240102 348618 240134 348854
rect 239514 313174 240134 348618
rect 239514 312938 239546 313174
rect 239782 312938 239866 313174
rect 240102 312938 240134 313174
rect 239514 312854 240134 312938
rect 239514 312618 239546 312854
rect 239782 312618 239866 312854
rect 240102 312618 240134 312854
rect 239514 302000 240134 312618
rect 243234 676894 243854 709082
rect 243234 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 243854 676894
rect 243234 676574 243854 676658
rect 243234 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 243854 676574
rect 243234 640894 243854 676338
rect 243234 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 243854 640894
rect 243234 640574 243854 640658
rect 243234 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 243854 640574
rect 243234 604894 243854 640338
rect 243234 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 243854 604894
rect 243234 604574 243854 604658
rect 243234 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 243854 604574
rect 243234 568894 243854 604338
rect 243234 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 243854 568894
rect 243234 568574 243854 568658
rect 243234 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 243854 568574
rect 243234 532894 243854 568338
rect 243234 532658 243266 532894
rect 243502 532658 243586 532894
rect 243822 532658 243854 532894
rect 243234 532574 243854 532658
rect 243234 532338 243266 532574
rect 243502 532338 243586 532574
rect 243822 532338 243854 532574
rect 243234 496894 243854 532338
rect 243234 496658 243266 496894
rect 243502 496658 243586 496894
rect 243822 496658 243854 496894
rect 243234 496574 243854 496658
rect 243234 496338 243266 496574
rect 243502 496338 243586 496574
rect 243822 496338 243854 496574
rect 243234 460894 243854 496338
rect 243234 460658 243266 460894
rect 243502 460658 243586 460894
rect 243822 460658 243854 460894
rect 243234 460574 243854 460658
rect 243234 460338 243266 460574
rect 243502 460338 243586 460574
rect 243822 460338 243854 460574
rect 243234 424894 243854 460338
rect 243234 424658 243266 424894
rect 243502 424658 243586 424894
rect 243822 424658 243854 424894
rect 243234 424574 243854 424658
rect 243234 424338 243266 424574
rect 243502 424338 243586 424574
rect 243822 424338 243854 424574
rect 243234 388894 243854 424338
rect 243234 388658 243266 388894
rect 243502 388658 243586 388894
rect 243822 388658 243854 388894
rect 243234 388574 243854 388658
rect 243234 388338 243266 388574
rect 243502 388338 243586 388574
rect 243822 388338 243854 388574
rect 243234 352894 243854 388338
rect 243234 352658 243266 352894
rect 243502 352658 243586 352894
rect 243822 352658 243854 352894
rect 243234 352574 243854 352658
rect 243234 352338 243266 352574
rect 243502 352338 243586 352574
rect 243822 352338 243854 352574
rect 243234 316894 243854 352338
rect 243234 316658 243266 316894
rect 243502 316658 243586 316894
rect 243822 316658 243854 316894
rect 243234 316574 243854 316658
rect 243234 316338 243266 316574
rect 243502 316338 243586 316574
rect 243822 316338 243854 316574
rect 243234 302000 243854 316338
rect 246954 680614 247574 711002
rect 264954 710598 265574 711590
rect 264954 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 265574 710598
rect 264954 710278 265574 710362
rect 264954 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 265574 710278
rect 261234 708678 261854 709670
rect 261234 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 261854 708678
rect 261234 708358 261854 708442
rect 261234 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 261854 708358
rect 257514 706758 258134 707750
rect 257514 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 258134 706758
rect 257514 706438 258134 706522
rect 257514 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 258134 706438
rect 246954 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 247574 680614
rect 246954 680294 247574 680378
rect 246954 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 247574 680294
rect 246954 644614 247574 680058
rect 246954 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 247574 644614
rect 246954 644294 247574 644378
rect 246954 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 247574 644294
rect 246954 608614 247574 644058
rect 246954 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 247574 608614
rect 246954 608294 247574 608378
rect 246954 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 247574 608294
rect 246954 572614 247574 608058
rect 246954 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 247574 572614
rect 246954 572294 247574 572378
rect 246954 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 247574 572294
rect 246954 536614 247574 572058
rect 246954 536378 246986 536614
rect 247222 536378 247306 536614
rect 247542 536378 247574 536614
rect 246954 536294 247574 536378
rect 246954 536058 246986 536294
rect 247222 536058 247306 536294
rect 247542 536058 247574 536294
rect 246954 500614 247574 536058
rect 246954 500378 246986 500614
rect 247222 500378 247306 500614
rect 247542 500378 247574 500614
rect 246954 500294 247574 500378
rect 246954 500058 246986 500294
rect 247222 500058 247306 500294
rect 247542 500058 247574 500294
rect 246954 464614 247574 500058
rect 246954 464378 246986 464614
rect 247222 464378 247306 464614
rect 247542 464378 247574 464614
rect 246954 464294 247574 464378
rect 246954 464058 246986 464294
rect 247222 464058 247306 464294
rect 247542 464058 247574 464294
rect 246954 428614 247574 464058
rect 246954 428378 246986 428614
rect 247222 428378 247306 428614
rect 247542 428378 247574 428614
rect 246954 428294 247574 428378
rect 246954 428058 246986 428294
rect 247222 428058 247306 428294
rect 247542 428058 247574 428294
rect 246954 392614 247574 428058
rect 246954 392378 246986 392614
rect 247222 392378 247306 392614
rect 247542 392378 247574 392614
rect 246954 392294 247574 392378
rect 246954 392058 246986 392294
rect 247222 392058 247306 392294
rect 247542 392058 247574 392294
rect 246954 356614 247574 392058
rect 246954 356378 246986 356614
rect 247222 356378 247306 356614
rect 247542 356378 247574 356614
rect 246954 356294 247574 356378
rect 246954 356058 246986 356294
rect 247222 356058 247306 356294
rect 247542 356058 247574 356294
rect 246954 320614 247574 356058
rect 246954 320378 246986 320614
rect 247222 320378 247306 320614
rect 247542 320378 247574 320614
rect 246954 320294 247574 320378
rect 246954 320058 246986 320294
rect 247222 320058 247306 320294
rect 247542 320058 247574 320294
rect 246954 302000 247574 320058
rect 253794 704838 254414 705830
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 543454 254414 578898
rect 253794 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 254414 543454
rect 253794 543134 254414 543218
rect 253794 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 254414 543134
rect 253794 507454 254414 542898
rect 253794 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 254414 507454
rect 253794 507134 254414 507218
rect 253794 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 254414 507134
rect 253794 471454 254414 506898
rect 253794 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 254414 471454
rect 253794 471134 254414 471218
rect 253794 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 254414 471134
rect 253794 435454 254414 470898
rect 253794 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 254414 435454
rect 253794 435134 254414 435218
rect 253794 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 254414 435134
rect 253794 399454 254414 434898
rect 253794 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 254414 399454
rect 253794 399134 254414 399218
rect 253794 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 254414 399134
rect 253794 363454 254414 398898
rect 253794 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 254414 363454
rect 253794 363134 254414 363218
rect 253794 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 254414 363134
rect 253794 327454 254414 362898
rect 253794 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 254414 327454
rect 253794 327134 254414 327218
rect 253794 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 254414 327134
rect 253794 302000 254414 326898
rect 257514 691174 258134 706202
rect 257514 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 258134 691174
rect 257514 690854 258134 690938
rect 257514 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 258134 690854
rect 257514 655174 258134 690618
rect 257514 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 258134 655174
rect 257514 654854 258134 654938
rect 257514 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 258134 654854
rect 257514 619174 258134 654618
rect 257514 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 258134 619174
rect 257514 618854 258134 618938
rect 257514 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 258134 618854
rect 257514 583174 258134 618618
rect 257514 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 258134 583174
rect 257514 582854 258134 582938
rect 257514 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 258134 582854
rect 257514 547174 258134 582618
rect 257514 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 258134 547174
rect 257514 546854 258134 546938
rect 257514 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 258134 546854
rect 257514 511174 258134 546618
rect 257514 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 258134 511174
rect 257514 510854 258134 510938
rect 257514 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 258134 510854
rect 257514 475174 258134 510618
rect 257514 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 258134 475174
rect 257514 474854 258134 474938
rect 257514 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 258134 474854
rect 257514 439174 258134 474618
rect 257514 438938 257546 439174
rect 257782 438938 257866 439174
rect 258102 438938 258134 439174
rect 257514 438854 258134 438938
rect 257514 438618 257546 438854
rect 257782 438618 257866 438854
rect 258102 438618 258134 438854
rect 257514 403174 258134 438618
rect 257514 402938 257546 403174
rect 257782 402938 257866 403174
rect 258102 402938 258134 403174
rect 257514 402854 258134 402938
rect 257514 402618 257546 402854
rect 257782 402618 257866 402854
rect 258102 402618 258134 402854
rect 257514 367174 258134 402618
rect 257514 366938 257546 367174
rect 257782 366938 257866 367174
rect 258102 366938 258134 367174
rect 257514 366854 258134 366938
rect 257514 366618 257546 366854
rect 257782 366618 257866 366854
rect 258102 366618 258134 366854
rect 257514 331174 258134 366618
rect 257514 330938 257546 331174
rect 257782 330938 257866 331174
rect 258102 330938 258134 331174
rect 257514 330854 258134 330938
rect 257514 330618 257546 330854
rect 257782 330618 257866 330854
rect 258102 330618 258134 330854
rect 257514 302000 258134 330618
rect 261234 694894 261854 708122
rect 261234 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 261854 694894
rect 261234 694574 261854 694658
rect 261234 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 261854 694574
rect 261234 658894 261854 694338
rect 261234 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 261854 658894
rect 261234 658574 261854 658658
rect 261234 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 261854 658574
rect 261234 622894 261854 658338
rect 261234 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 261854 622894
rect 261234 622574 261854 622658
rect 261234 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 261854 622574
rect 261234 586894 261854 622338
rect 261234 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 261854 586894
rect 261234 586574 261854 586658
rect 261234 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 261854 586574
rect 261234 550894 261854 586338
rect 261234 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 261854 550894
rect 261234 550574 261854 550658
rect 261234 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 261854 550574
rect 261234 514894 261854 550338
rect 261234 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 261854 514894
rect 261234 514574 261854 514658
rect 261234 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 261854 514574
rect 261234 478894 261854 514338
rect 261234 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 261854 478894
rect 261234 478574 261854 478658
rect 261234 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 261854 478574
rect 261234 442894 261854 478338
rect 261234 442658 261266 442894
rect 261502 442658 261586 442894
rect 261822 442658 261854 442894
rect 261234 442574 261854 442658
rect 261234 442338 261266 442574
rect 261502 442338 261586 442574
rect 261822 442338 261854 442574
rect 261234 406894 261854 442338
rect 261234 406658 261266 406894
rect 261502 406658 261586 406894
rect 261822 406658 261854 406894
rect 261234 406574 261854 406658
rect 261234 406338 261266 406574
rect 261502 406338 261586 406574
rect 261822 406338 261854 406574
rect 261234 370894 261854 406338
rect 261234 370658 261266 370894
rect 261502 370658 261586 370894
rect 261822 370658 261854 370894
rect 261234 370574 261854 370658
rect 261234 370338 261266 370574
rect 261502 370338 261586 370574
rect 261822 370338 261854 370574
rect 261234 334894 261854 370338
rect 261234 334658 261266 334894
rect 261502 334658 261586 334894
rect 261822 334658 261854 334894
rect 261234 334574 261854 334658
rect 261234 334338 261266 334574
rect 261502 334338 261586 334574
rect 261822 334338 261854 334574
rect 261234 302000 261854 334338
rect 264954 698614 265574 710042
rect 282954 711558 283574 711590
rect 282954 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 283574 711558
rect 282954 711238 283574 711322
rect 282954 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 283574 711238
rect 279234 709638 279854 709670
rect 279234 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 279854 709638
rect 279234 709318 279854 709402
rect 279234 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 279854 709318
rect 275514 707718 276134 707750
rect 275514 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 276134 707718
rect 275514 707398 276134 707482
rect 275514 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 276134 707398
rect 264954 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 265574 698614
rect 264954 698294 265574 698378
rect 264954 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 265574 698294
rect 264954 662614 265574 698058
rect 264954 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 265574 662614
rect 264954 662294 265574 662378
rect 264954 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 265574 662294
rect 264954 626614 265574 662058
rect 264954 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 265574 626614
rect 264954 626294 265574 626378
rect 264954 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 265574 626294
rect 264954 590614 265574 626058
rect 264954 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 265574 590614
rect 264954 590294 265574 590378
rect 264954 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 265574 590294
rect 264954 554614 265574 590058
rect 264954 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 265574 554614
rect 264954 554294 265574 554378
rect 264954 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 265574 554294
rect 264954 518614 265574 554058
rect 264954 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 265574 518614
rect 264954 518294 265574 518378
rect 264954 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 265574 518294
rect 264954 482614 265574 518058
rect 264954 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 265574 482614
rect 264954 482294 265574 482378
rect 264954 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 265574 482294
rect 264954 446614 265574 482058
rect 264954 446378 264986 446614
rect 265222 446378 265306 446614
rect 265542 446378 265574 446614
rect 264954 446294 265574 446378
rect 264954 446058 264986 446294
rect 265222 446058 265306 446294
rect 265542 446058 265574 446294
rect 264954 410614 265574 446058
rect 264954 410378 264986 410614
rect 265222 410378 265306 410614
rect 265542 410378 265574 410614
rect 264954 410294 265574 410378
rect 264954 410058 264986 410294
rect 265222 410058 265306 410294
rect 265542 410058 265574 410294
rect 264954 374614 265574 410058
rect 264954 374378 264986 374614
rect 265222 374378 265306 374614
rect 265542 374378 265574 374614
rect 264954 374294 265574 374378
rect 264954 374058 264986 374294
rect 265222 374058 265306 374294
rect 265542 374058 265574 374294
rect 264954 338614 265574 374058
rect 264954 338378 264986 338614
rect 265222 338378 265306 338614
rect 265542 338378 265574 338614
rect 264954 338294 265574 338378
rect 264954 338058 264986 338294
rect 265222 338058 265306 338294
rect 265542 338058 265574 338294
rect 264954 302614 265574 338058
rect 264954 302378 264986 302614
rect 265222 302378 265306 302614
rect 265542 302378 265574 302614
rect 264954 302294 265574 302378
rect 264954 302058 264986 302294
rect 265222 302058 265306 302294
rect 265542 302058 265574 302294
rect 264954 302000 265574 302058
rect 271794 705798 272414 705830
rect 271794 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 272414 705798
rect 271794 705478 272414 705562
rect 271794 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 272414 705478
rect 271794 669454 272414 705242
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 561454 272414 596898
rect 271794 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 272414 561454
rect 271794 561134 272414 561218
rect 271794 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 272414 561134
rect 271794 525454 272414 560898
rect 271794 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 272414 525454
rect 271794 525134 272414 525218
rect 271794 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 272414 525134
rect 271794 489454 272414 524898
rect 271794 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 272414 489454
rect 271794 489134 272414 489218
rect 271794 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 272414 489134
rect 271794 453454 272414 488898
rect 271794 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 272414 453454
rect 271794 453134 272414 453218
rect 271794 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 272414 453134
rect 271794 417454 272414 452898
rect 271794 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 272414 417454
rect 271794 417134 272414 417218
rect 271794 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 272414 417134
rect 271794 381454 272414 416898
rect 271794 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 272414 381454
rect 271794 381134 272414 381218
rect 271794 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 272414 381134
rect 271794 345454 272414 380898
rect 271794 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 272414 345454
rect 271794 345134 272414 345218
rect 271794 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 272414 345134
rect 271794 309454 272414 344898
rect 271794 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 272414 309454
rect 271794 309134 272414 309218
rect 271794 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 272414 309134
rect 271794 302000 272414 308898
rect 275514 673174 276134 707162
rect 275514 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 276134 673174
rect 275514 672854 276134 672938
rect 275514 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 276134 672854
rect 275514 637174 276134 672618
rect 275514 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 276134 637174
rect 275514 636854 276134 636938
rect 275514 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 276134 636854
rect 275514 601174 276134 636618
rect 275514 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 276134 601174
rect 275514 600854 276134 600938
rect 275514 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 276134 600854
rect 275514 565174 276134 600618
rect 275514 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 276134 565174
rect 275514 564854 276134 564938
rect 275514 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 276134 564854
rect 275514 529174 276134 564618
rect 275514 528938 275546 529174
rect 275782 528938 275866 529174
rect 276102 528938 276134 529174
rect 275514 528854 276134 528938
rect 275514 528618 275546 528854
rect 275782 528618 275866 528854
rect 276102 528618 276134 528854
rect 275514 493174 276134 528618
rect 275514 492938 275546 493174
rect 275782 492938 275866 493174
rect 276102 492938 276134 493174
rect 275514 492854 276134 492938
rect 275514 492618 275546 492854
rect 275782 492618 275866 492854
rect 276102 492618 276134 492854
rect 275514 457174 276134 492618
rect 275514 456938 275546 457174
rect 275782 456938 275866 457174
rect 276102 456938 276134 457174
rect 275514 456854 276134 456938
rect 275514 456618 275546 456854
rect 275782 456618 275866 456854
rect 276102 456618 276134 456854
rect 275514 421174 276134 456618
rect 275514 420938 275546 421174
rect 275782 420938 275866 421174
rect 276102 420938 276134 421174
rect 275514 420854 276134 420938
rect 275514 420618 275546 420854
rect 275782 420618 275866 420854
rect 276102 420618 276134 420854
rect 275514 385174 276134 420618
rect 275514 384938 275546 385174
rect 275782 384938 275866 385174
rect 276102 384938 276134 385174
rect 275514 384854 276134 384938
rect 275514 384618 275546 384854
rect 275782 384618 275866 384854
rect 276102 384618 276134 384854
rect 275514 349174 276134 384618
rect 275514 348938 275546 349174
rect 275782 348938 275866 349174
rect 276102 348938 276134 349174
rect 275514 348854 276134 348938
rect 275514 348618 275546 348854
rect 275782 348618 275866 348854
rect 276102 348618 276134 348854
rect 275514 313174 276134 348618
rect 275514 312938 275546 313174
rect 275782 312938 275866 313174
rect 276102 312938 276134 313174
rect 275514 312854 276134 312938
rect 275514 312618 275546 312854
rect 275782 312618 275866 312854
rect 276102 312618 276134 312854
rect 275514 302000 276134 312618
rect 279234 676894 279854 709082
rect 279234 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 279854 676894
rect 279234 676574 279854 676658
rect 279234 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 279854 676574
rect 279234 640894 279854 676338
rect 279234 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 279854 640894
rect 279234 640574 279854 640658
rect 279234 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 279854 640574
rect 279234 604894 279854 640338
rect 279234 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 279854 604894
rect 279234 604574 279854 604658
rect 279234 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 279854 604574
rect 279234 568894 279854 604338
rect 279234 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 279854 568894
rect 279234 568574 279854 568658
rect 279234 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 279854 568574
rect 279234 532894 279854 568338
rect 279234 532658 279266 532894
rect 279502 532658 279586 532894
rect 279822 532658 279854 532894
rect 279234 532574 279854 532658
rect 279234 532338 279266 532574
rect 279502 532338 279586 532574
rect 279822 532338 279854 532574
rect 279234 496894 279854 532338
rect 279234 496658 279266 496894
rect 279502 496658 279586 496894
rect 279822 496658 279854 496894
rect 279234 496574 279854 496658
rect 279234 496338 279266 496574
rect 279502 496338 279586 496574
rect 279822 496338 279854 496574
rect 279234 460894 279854 496338
rect 279234 460658 279266 460894
rect 279502 460658 279586 460894
rect 279822 460658 279854 460894
rect 279234 460574 279854 460658
rect 279234 460338 279266 460574
rect 279502 460338 279586 460574
rect 279822 460338 279854 460574
rect 279234 424894 279854 460338
rect 279234 424658 279266 424894
rect 279502 424658 279586 424894
rect 279822 424658 279854 424894
rect 279234 424574 279854 424658
rect 279234 424338 279266 424574
rect 279502 424338 279586 424574
rect 279822 424338 279854 424574
rect 279234 388894 279854 424338
rect 279234 388658 279266 388894
rect 279502 388658 279586 388894
rect 279822 388658 279854 388894
rect 279234 388574 279854 388658
rect 279234 388338 279266 388574
rect 279502 388338 279586 388574
rect 279822 388338 279854 388574
rect 279234 352894 279854 388338
rect 279234 352658 279266 352894
rect 279502 352658 279586 352894
rect 279822 352658 279854 352894
rect 279234 352574 279854 352658
rect 279234 352338 279266 352574
rect 279502 352338 279586 352574
rect 279822 352338 279854 352574
rect 279234 316894 279854 352338
rect 279234 316658 279266 316894
rect 279502 316658 279586 316894
rect 279822 316658 279854 316894
rect 279234 316574 279854 316658
rect 279234 316338 279266 316574
rect 279502 316338 279586 316574
rect 279822 316338 279854 316574
rect 279234 302000 279854 316338
rect 282954 680614 283574 711002
rect 300954 710598 301574 711590
rect 300954 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 301574 710598
rect 300954 710278 301574 710362
rect 300954 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 301574 710278
rect 297234 708678 297854 709670
rect 297234 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 297854 708678
rect 297234 708358 297854 708442
rect 297234 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 297854 708358
rect 293514 706758 294134 707750
rect 293514 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 294134 706758
rect 293514 706438 294134 706522
rect 293514 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 294134 706438
rect 282954 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 283574 680614
rect 282954 680294 283574 680378
rect 282954 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 283574 680294
rect 282954 644614 283574 680058
rect 282954 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 283574 644614
rect 282954 644294 283574 644378
rect 282954 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 283574 644294
rect 282954 608614 283574 644058
rect 282954 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 283574 608614
rect 282954 608294 283574 608378
rect 282954 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 283574 608294
rect 282954 572614 283574 608058
rect 282954 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 283574 572614
rect 282954 572294 283574 572378
rect 282954 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 283574 572294
rect 282954 536614 283574 572058
rect 282954 536378 282986 536614
rect 283222 536378 283306 536614
rect 283542 536378 283574 536614
rect 282954 536294 283574 536378
rect 282954 536058 282986 536294
rect 283222 536058 283306 536294
rect 283542 536058 283574 536294
rect 282954 500614 283574 536058
rect 282954 500378 282986 500614
rect 283222 500378 283306 500614
rect 283542 500378 283574 500614
rect 282954 500294 283574 500378
rect 282954 500058 282986 500294
rect 283222 500058 283306 500294
rect 283542 500058 283574 500294
rect 282954 464614 283574 500058
rect 282954 464378 282986 464614
rect 283222 464378 283306 464614
rect 283542 464378 283574 464614
rect 282954 464294 283574 464378
rect 282954 464058 282986 464294
rect 283222 464058 283306 464294
rect 283542 464058 283574 464294
rect 282954 428614 283574 464058
rect 282954 428378 282986 428614
rect 283222 428378 283306 428614
rect 283542 428378 283574 428614
rect 282954 428294 283574 428378
rect 282954 428058 282986 428294
rect 283222 428058 283306 428294
rect 283542 428058 283574 428294
rect 282954 392614 283574 428058
rect 282954 392378 282986 392614
rect 283222 392378 283306 392614
rect 283542 392378 283574 392614
rect 282954 392294 283574 392378
rect 282954 392058 282986 392294
rect 283222 392058 283306 392294
rect 283542 392058 283574 392294
rect 282954 356614 283574 392058
rect 282954 356378 282986 356614
rect 283222 356378 283306 356614
rect 283542 356378 283574 356614
rect 282954 356294 283574 356378
rect 282954 356058 282986 356294
rect 283222 356058 283306 356294
rect 283542 356058 283574 356294
rect 282954 320614 283574 356058
rect 282954 320378 282986 320614
rect 283222 320378 283306 320614
rect 283542 320378 283574 320614
rect 282954 320294 283574 320378
rect 282954 320058 282986 320294
rect 283222 320058 283306 320294
rect 283542 320058 283574 320294
rect 282954 302000 283574 320058
rect 289794 704838 290414 705830
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 543454 290414 578898
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289794 507454 290414 542898
rect 289794 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 290414 507454
rect 289794 507134 290414 507218
rect 289794 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 290414 507134
rect 289794 471454 290414 506898
rect 289794 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 290414 471454
rect 289794 471134 290414 471218
rect 289794 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 290414 471134
rect 289794 435454 290414 470898
rect 289794 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 290414 435454
rect 289794 435134 290414 435218
rect 289794 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 290414 435134
rect 289794 399454 290414 434898
rect 289794 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 290414 399454
rect 289794 399134 290414 399218
rect 289794 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 290414 399134
rect 289794 363454 290414 398898
rect 289794 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 290414 363454
rect 289794 363134 290414 363218
rect 289794 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 290414 363134
rect 289794 327454 290414 362898
rect 289794 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 290414 327454
rect 289794 327134 290414 327218
rect 289794 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 290414 327134
rect 289794 302000 290414 326898
rect 293514 691174 294134 706202
rect 293514 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 294134 691174
rect 293514 690854 294134 690938
rect 293514 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 294134 690854
rect 293514 655174 294134 690618
rect 293514 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 294134 655174
rect 293514 654854 294134 654938
rect 293514 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 294134 654854
rect 293514 619174 294134 654618
rect 293514 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 294134 619174
rect 293514 618854 294134 618938
rect 293514 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 294134 618854
rect 293514 583174 294134 618618
rect 293514 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 294134 583174
rect 293514 582854 294134 582938
rect 293514 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 294134 582854
rect 293514 547174 294134 582618
rect 293514 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 294134 547174
rect 293514 546854 294134 546938
rect 293514 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 294134 546854
rect 293514 511174 294134 546618
rect 293514 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 294134 511174
rect 293514 510854 294134 510938
rect 293514 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 294134 510854
rect 293514 475174 294134 510618
rect 293514 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 294134 475174
rect 293514 474854 294134 474938
rect 293514 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 294134 474854
rect 293514 439174 294134 474618
rect 293514 438938 293546 439174
rect 293782 438938 293866 439174
rect 294102 438938 294134 439174
rect 293514 438854 294134 438938
rect 293514 438618 293546 438854
rect 293782 438618 293866 438854
rect 294102 438618 294134 438854
rect 293514 403174 294134 438618
rect 293514 402938 293546 403174
rect 293782 402938 293866 403174
rect 294102 402938 294134 403174
rect 293514 402854 294134 402938
rect 293514 402618 293546 402854
rect 293782 402618 293866 402854
rect 294102 402618 294134 402854
rect 293514 367174 294134 402618
rect 293514 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 294134 367174
rect 293514 366854 294134 366938
rect 293514 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 294134 366854
rect 293514 331174 294134 366618
rect 293514 330938 293546 331174
rect 293782 330938 293866 331174
rect 294102 330938 294134 331174
rect 293514 330854 294134 330938
rect 293514 330618 293546 330854
rect 293782 330618 293866 330854
rect 294102 330618 294134 330854
rect 293514 302000 294134 330618
rect 297234 694894 297854 708122
rect 297234 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 297854 694894
rect 297234 694574 297854 694658
rect 297234 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 297854 694574
rect 297234 658894 297854 694338
rect 297234 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 297854 658894
rect 297234 658574 297854 658658
rect 297234 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 297854 658574
rect 297234 622894 297854 658338
rect 297234 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 297854 622894
rect 297234 622574 297854 622658
rect 297234 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 297854 622574
rect 297234 586894 297854 622338
rect 297234 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 297854 586894
rect 297234 586574 297854 586658
rect 297234 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 297854 586574
rect 297234 550894 297854 586338
rect 297234 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 297854 550894
rect 297234 550574 297854 550658
rect 297234 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 297854 550574
rect 297234 514894 297854 550338
rect 297234 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 297854 514894
rect 297234 514574 297854 514658
rect 297234 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 297854 514574
rect 297234 478894 297854 514338
rect 297234 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 297854 478894
rect 297234 478574 297854 478658
rect 297234 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 297854 478574
rect 297234 442894 297854 478338
rect 297234 442658 297266 442894
rect 297502 442658 297586 442894
rect 297822 442658 297854 442894
rect 297234 442574 297854 442658
rect 297234 442338 297266 442574
rect 297502 442338 297586 442574
rect 297822 442338 297854 442574
rect 297234 406894 297854 442338
rect 297234 406658 297266 406894
rect 297502 406658 297586 406894
rect 297822 406658 297854 406894
rect 297234 406574 297854 406658
rect 297234 406338 297266 406574
rect 297502 406338 297586 406574
rect 297822 406338 297854 406574
rect 297234 370894 297854 406338
rect 297234 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 297854 370894
rect 297234 370574 297854 370658
rect 297234 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 297854 370574
rect 297234 334894 297854 370338
rect 297234 334658 297266 334894
rect 297502 334658 297586 334894
rect 297822 334658 297854 334894
rect 297234 334574 297854 334658
rect 297234 334338 297266 334574
rect 297502 334338 297586 334574
rect 297822 334338 297854 334574
rect 297234 302000 297854 334338
rect 300954 698614 301574 710042
rect 318954 711558 319574 711590
rect 318954 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 319574 711558
rect 318954 711238 319574 711322
rect 318954 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 319574 711238
rect 315234 709638 315854 709670
rect 315234 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 315854 709638
rect 315234 709318 315854 709402
rect 315234 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 315854 709318
rect 311514 707718 312134 707750
rect 311514 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 312134 707718
rect 311514 707398 312134 707482
rect 311514 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 312134 707398
rect 300954 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 301574 698614
rect 300954 698294 301574 698378
rect 300954 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 301574 698294
rect 300954 662614 301574 698058
rect 300954 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 301574 662614
rect 300954 662294 301574 662378
rect 300954 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 301574 662294
rect 300954 626614 301574 662058
rect 300954 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 301574 626614
rect 300954 626294 301574 626378
rect 300954 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 301574 626294
rect 300954 590614 301574 626058
rect 300954 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 301574 590614
rect 300954 590294 301574 590378
rect 300954 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 301574 590294
rect 300954 554614 301574 590058
rect 300954 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 301574 554614
rect 300954 554294 301574 554378
rect 300954 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 301574 554294
rect 300954 518614 301574 554058
rect 300954 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 301574 518614
rect 300954 518294 301574 518378
rect 300954 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 301574 518294
rect 300954 482614 301574 518058
rect 300954 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 301574 482614
rect 300954 482294 301574 482378
rect 300954 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 301574 482294
rect 300954 446614 301574 482058
rect 300954 446378 300986 446614
rect 301222 446378 301306 446614
rect 301542 446378 301574 446614
rect 300954 446294 301574 446378
rect 300954 446058 300986 446294
rect 301222 446058 301306 446294
rect 301542 446058 301574 446294
rect 300954 410614 301574 446058
rect 300954 410378 300986 410614
rect 301222 410378 301306 410614
rect 301542 410378 301574 410614
rect 300954 410294 301574 410378
rect 300954 410058 300986 410294
rect 301222 410058 301306 410294
rect 301542 410058 301574 410294
rect 300954 374614 301574 410058
rect 300954 374378 300986 374614
rect 301222 374378 301306 374614
rect 301542 374378 301574 374614
rect 300954 374294 301574 374378
rect 300954 374058 300986 374294
rect 301222 374058 301306 374294
rect 301542 374058 301574 374294
rect 300954 338614 301574 374058
rect 300954 338378 300986 338614
rect 301222 338378 301306 338614
rect 301542 338378 301574 338614
rect 300954 338294 301574 338378
rect 300954 338058 300986 338294
rect 301222 338058 301306 338294
rect 301542 338058 301574 338294
rect 300954 302614 301574 338058
rect 300954 302378 300986 302614
rect 301222 302378 301306 302614
rect 301542 302378 301574 302614
rect 300954 302294 301574 302378
rect 300954 302058 300986 302294
rect 301222 302058 301306 302294
rect 301542 302058 301574 302294
rect 300954 302000 301574 302058
rect 307794 705798 308414 705830
rect 307794 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 308414 705798
rect 307794 705478 308414 705562
rect 307794 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 308414 705478
rect 307794 669454 308414 705242
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 561454 308414 596898
rect 307794 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 308414 561454
rect 307794 561134 308414 561218
rect 307794 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 308414 561134
rect 307794 525454 308414 560898
rect 307794 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 308414 525454
rect 307794 525134 308414 525218
rect 307794 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 308414 525134
rect 307794 489454 308414 524898
rect 307794 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 308414 489454
rect 307794 489134 308414 489218
rect 307794 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 308414 489134
rect 307794 453454 308414 488898
rect 307794 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 308414 453454
rect 307794 453134 308414 453218
rect 307794 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 308414 453134
rect 307794 417454 308414 452898
rect 307794 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 308414 417454
rect 307794 417134 308414 417218
rect 307794 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 308414 417134
rect 307794 381454 308414 416898
rect 307794 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 308414 381454
rect 307794 381134 308414 381218
rect 307794 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 308414 381134
rect 307794 345454 308414 380898
rect 307794 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 308414 345454
rect 307794 345134 308414 345218
rect 307794 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 308414 345134
rect 307794 309454 308414 344898
rect 307794 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 308414 309454
rect 307794 309134 308414 309218
rect 307794 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 308414 309134
rect 204208 291454 204528 291486
rect 204208 291218 204250 291454
rect 204486 291218 204528 291454
rect 204208 291134 204528 291218
rect 204208 290898 204250 291134
rect 204486 290898 204528 291134
rect 204208 290866 204528 290898
rect 234928 291454 235248 291486
rect 234928 291218 234970 291454
rect 235206 291218 235248 291454
rect 234928 291134 235248 291218
rect 234928 290898 234970 291134
rect 235206 290898 235248 291134
rect 234928 290866 235248 290898
rect 265648 291454 265968 291486
rect 265648 291218 265690 291454
rect 265926 291218 265968 291454
rect 265648 291134 265968 291218
rect 265648 290898 265690 291134
rect 265926 290898 265968 291134
rect 265648 290866 265968 290898
rect 296368 291454 296688 291486
rect 296368 291218 296410 291454
rect 296646 291218 296688 291454
rect 296368 291134 296688 291218
rect 296368 290898 296410 291134
rect 296646 290898 296688 291134
rect 296368 290866 296688 290898
rect 219568 273454 219888 273486
rect 219568 273218 219610 273454
rect 219846 273218 219888 273454
rect 219568 273134 219888 273218
rect 219568 272898 219610 273134
rect 219846 272898 219888 273134
rect 219568 272866 219888 272898
rect 250288 273454 250608 273486
rect 250288 273218 250330 273454
rect 250566 273218 250608 273454
rect 250288 273134 250608 273218
rect 250288 272898 250330 273134
rect 250566 272898 250608 273134
rect 250288 272866 250608 272898
rect 281008 273454 281328 273486
rect 281008 273218 281050 273454
rect 281286 273218 281328 273454
rect 281008 273134 281328 273218
rect 281008 272898 281050 273134
rect 281286 272898 281328 273134
rect 281008 272866 281328 272898
rect 307794 273454 308414 308898
rect 307794 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 308414 273454
rect 307794 273134 308414 273218
rect 307794 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 308414 273134
rect 192954 266378 192986 266614
rect 193222 266378 193306 266614
rect 193542 266378 193574 266614
rect 192954 266294 193574 266378
rect 192954 266058 192986 266294
rect 193222 266058 193306 266294
rect 193542 266058 193574 266294
rect 192954 230614 193574 266058
rect 204208 255454 204528 255486
rect 204208 255218 204250 255454
rect 204486 255218 204528 255454
rect 204208 255134 204528 255218
rect 204208 254898 204250 255134
rect 204486 254898 204528 255134
rect 204208 254866 204528 254898
rect 234928 255454 235248 255486
rect 234928 255218 234970 255454
rect 235206 255218 235248 255454
rect 234928 255134 235248 255218
rect 234928 254898 234970 255134
rect 235206 254898 235248 255134
rect 234928 254866 235248 254898
rect 265648 255454 265968 255486
rect 265648 255218 265690 255454
rect 265926 255218 265968 255454
rect 265648 255134 265968 255218
rect 265648 254898 265690 255134
rect 265926 254898 265968 255134
rect 265648 254866 265968 254898
rect 296368 255454 296688 255486
rect 296368 255218 296410 255454
rect 296646 255218 296688 255454
rect 296368 255134 296688 255218
rect 296368 254898 296410 255134
rect 296646 254898 296688 255134
rect 296368 254866 296688 254898
rect 219568 237454 219888 237486
rect 219568 237218 219610 237454
rect 219846 237218 219888 237454
rect 219568 237134 219888 237218
rect 219568 236898 219610 237134
rect 219846 236898 219888 237134
rect 219568 236866 219888 236898
rect 250288 237454 250608 237486
rect 250288 237218 250330 237454
rect 250566 237218 250608 237454
rect 250288 237134 250608 237218
rect 250288 236898 250330 237134
rect 250566 236898 250608 237134
rect 250288 236866 250608 236898
rect 281008 237454 281328 237486
rect 281008 237218 281050 237454
rect 281286 237218 281328 237454
rect 281008 237134 281328 237218
rect 281008 236898 281050 237134
rect 281286 236898 281328 237134
rect 281008 236866 281328 236898
rect 307794 237454 308414 272898
rect 307794 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 308414 237454
rect 307794 237134 308414 237218
rect 307794 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 308414 237134
rect 192954 230378 192986 230614
rect 193222 230378 193306 230614
rect 193542 230378 193574 230614
rect 192954 230294 193574 230378
rect 192954 230058 192986 230294
rect 193222 230058 193306 230294
rect 193542 230058 193574 230294
rect 192954 194614 193574 230058
rect 204208 219454 204528 219486
rect 204208 219218 204250 219454
rect 204486 219218 204528 219454
rect 204208 219134 204528 219218
rect 204208 218898 204250 219134
rect 204486 218898 204528 219134
rect 204208 218866 204528 218898
rect 234928 219454 235248 219486
rect 234928 219218 234970 219454
rect 235206 219218 235248 219454
rect 234928 219134 235248 219218
rect 234928 218898 234970 219134
rect 235206 218898 235248 219134
rect 234928 218866 235248 218898
rect 265648 219454 265968 219486
rect 265648 219218 265690 219454
rect 265926 219218 265968 219454
rect 265648 219134 265968 219218
rect 265648 218898 265690 219134
rect 265926 218898 265968 219134
rect 265648 218866 265968 218898
rect 296368 219454 296688 219486
rect 296368 219218 296410 219454
rect 296646 219218 296688 219454
rect 296368 219134 296688 219218
rect 296368 218898 296410 219134
rect 296646 218898 296688 219134
rect 296368 218866 296688 218898
rect 219568 201454 219888 201486
rect 219568 201218 219610 201454
rect 219846 201218 219888 201454
rect 219568 201134 219888 201218
rect 219568 200898 219610 201134
rect 219846 200898 219888 201134
rect 219568 200866 219888 200898
rect 250288 201454 250608 201486
rect 250288 201218 250330 201454
rect 250566 201218 250608 201454
rect 250288 201134 250608 201218
rect 250288 200898 250330 201134
rect 250566 200898 250608 201134
rect 250288 200866 250608 200898
rect 281008 201454 281328 201486
rect 281008 201218 281050 201454
rect 281286 201218 281328 201454
rect 281008 201134 281328 201218
rect 281008 200898 281050 201134
rect 281286 200898 281328 201134
rect 281008 200866 281328 200898
rect 307794 201454 308414 236898
rect 307794 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 308414 201454
rect 307794 201134 308414 201218
rect 307794 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 308414 201134
rect 192954 194378 192986 194614
rect 193222 194378 193306 194614
rect 193542 194378 193574 194614
rect 192954 194294 193574 194378
rect 192954 194058 192986 194294
rect 193222 194058 193306 194294
rect 193542 194058 193574 194294
rect 192954 158614 193574 194058
rect 204208 183454 204528 183486
rect 204208 183218 204250 183454
rect 204486 183218 204528 183454
rect 204208 183134 204528 183218
rect 204208 182898 204250 183134
rect 204486 182898 204528 183134
rect 204208 182866 204528 182898
rect 234928 183454 235248 183486
rect 234928 183218 234970 183454
rect 235206 183218 235248 183454
rect 234928 183134 235248 183218
rect 234928 182898 234970 183134
rect 235206 182898 235248 183134
rect 234928 182866 235248 182898
rect 265648 183454 265968 183486
rect 265648 183218 265690 183454
rect 265926 183218 265968 183454
rect 265648 183134 265968 183218
rect 265648 182898 265690 183134
rect 265926 182898 265968 183134
rect 265648 182866 265968 182898
rect 296368 183454 296688 183486
rect 296368 183218 296410 183454
rect 296646 183218 296688 183454
rect 296368 183134 296688 183218
rect 296368 182898 296410 183134
rect 296646 182898 296688 183134
rect 296368 182866 296688 182898
rect 219568 165454 219888 165486
rect 219568 165218 219610 165454
rect 219846 165218 219888 165454
rect 219568 165134 219888 165218
rect 219568 164898 219610 165134
rect 219846 164898 219888 165134
rect 219568 164866 219888 164898
rect 250288 165454 250608 165486
rect 250288 165218 250330 165454
rect 250566 165218 250608 165454
rect 250288 165134 250608 165218
rect 250288 164898 250330 165134
rect 250566 164898 250608 165134
rect 250288 164866 250608 164898
rect 281008 165454 281328 165486
rect 281008 165218 281050 165454
rect 281286 165218 281328 165454
rect 281008 165134 281328 165218
rect 281008 164898 281050 165134
rect 281286 164898 281328 165134
rect 281008 164866 281328 164898
rect 307794 165454 308414 200898
rect 307794 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 308414 165454
rect 307794 165134 308414 165218
rect 307794 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 308414 165134
rect 192954 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 193574 158614
rect 192954 158294 193574 158378
rect 192954 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 193574 158294
rect 192954 122614 193574 158058
rect 204208 147454 204528 147486
rect 204208 147218 204250 147454
rect 204486 147218 204528 147454
rect 204208 147134 204528 147218
rect 204208 146898 204250 147134
rect 204486 146898 204528 147134
rect 204208 146866 204528 146898
rect 234928 147454 235248 147486
rect 234928 147218 234970 147454
rect 235206 147218 235248 147454
rect 234928 147134 235248 147218
rect 234928 146898 234970 147134
rect 235206 146898 235248 147134
rect 234928 146866 235248 146898
rect 265648 147454 265968 147486
rect 265648 147218 265690 147454
rect 265926 147218 265968 147454
rect 265648 147134 265968 147218
rect 265648 146898 265690 147134
rect 265926 146898 265968 147134
rect 265648 146866 265968 146898
rect 296368 147454 296688 147486
rect 296368 147218 296410 147454
rect 296646 147218 296688 147454
rect 296368 147134 296688 147218
rect 296368 146898 296410 147134
rect 296646 146898 296688 147134
rect 296368 146866 296688 146898
rect 219568 129454 219888 129486
rect 219568 129218 219610 129454
rect 219846 129218 219888 129454
rect 219568 129134 219888 129218
rect 219568 128898 219610 129134
rect 219846 128898 219888 129134
rect 219568 128866 219888 128898
rect 250288 129454 250608 129486
rect 250288 129218 250330 129454
rect 250566 129218 250608 129454
rect 250288 129134 250608 129218
rect 250288 128898 250330 129134
rect 250566 128898 250608 129134
rect 250288 128866 250608 128898
rect 281008 129454 281328 129486
rect 281008 129218 281050 129454
rect 281286 129218 281328 129454
rect 281008 129134 281328 129218
rect 281008 128898 281050 129134
rect 281286 128898 281328 129134
rect 281008 128866 281328 128898
rect 307794 129454 308414 164898
rect 307794 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 308414 129454
rect 307794 129134 308414 129218
rect 307794 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 308414 129134
rect 192954 122378 192986 122614
rect 193222 122378 193306 122614
rect 193542 122378 193574 122614
rect 192954 122294 193574 122378
rect 192954 122058 192986 122294
rect 193222 122058 193306 122294
rect 193542 122058 193574 122294
rect 192954 86614 193574 122058
rect 204208 111454 204528 111486
rect 204208 111218 204250 111454
rect 204486 111218 204528 111454
rect 204208 111134 204528 111218
rect 204208 110898 204250 111134
rect 204486 110898 204528 111134
rect 204208 110866 204528 110898
rect 234928 111454 235248 111486
rect 234928 111218 234970 111454
rect 235206 111218 235248 111454
rect 234928 111134 235248 111218
rect 234928 110898 234970 111134
rect 235206 110898 235248 111134
rect 234928 110866 235248 110898
rect 265648 111454 265968 111486
rect 265648 111218 265690 111454
rect 265926 111218 265968 111454
rect 265648 111134 265968 111218
rect 265648 110898 265690 111134
rect 265926 110898 265968 111134
rect 265648 110866 265968 110898
rect 296368 111454 296688 111486
rect 296368 111218 296410 111454
rect 296646 111218 296688 111454
rect 296368 111134 296688 111218
rect 296368 110898 296410 111134
rect 296646 110898 296688 111134
rect 296368 110866 296688 110898
rect 192954 86378 192986 86614
rect 193222 86378 193306 86614
rect 193542 86378 193574 86614
rect 192954 86294 193574 86378
rect 192954 86058 192986 86294
rect 193222 86058 193306 86294
rect 193542 86058 193574 86294
rect 192954 50614 193574 86058
rect 192954 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 193574 50614
rect 192954 50294 193574 50378
rect 192954 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 193574 50294
rect 192954 14614 193574 50058
rect 192954 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 193574 14614
rect 192954 14294 193574 14378
rect 192954 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 193574 14294
rect 174954 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 175574 -7066
rect 174954 -7386 175574 -7302
rect 174954 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 175574 -7386
rect 174954 -7654 175574 -7622
rect 192954 -6106 193574 14058
rect 199794 93454 200414 98000
rect 199794 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 200414 93454
rect 199794 93134 200414 93218
rect 199794 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 200414 93134
rect 199794 57454 200414 92898
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 21454 200414 56898
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -1306 200414 20898
rect 199794 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 200414 -1306
rect 199794 -1626 200414 -1542
rect 199794 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 200414 -1626
rect 199794 -1894 200414 -1862
rect 203514 97174 204134 98000
rect 203514 96938 203546 97174
rect 203782 96938 203866 97174
rect 204102 96938 204134 97174
rect 203514 96854 204134 96938
rect 203514 96618 203546 96854
rect 203782 96618 203866 96854
rect 204102 96618 204134 96854
rect 203514 61174 204134 96618
rect 203514 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 204134 61174
rect 203514 60854 204134 60938
rect 203514 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 204134 60854
rect 203514 25174 204134 60618
rect 203514 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 204134 25174
rect 203514 24854 204134 24938
rect 203514 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 204134 24854
rect 203514 -3226 204134 24618
rect 203514 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 204134 -3226
rect 203514 -3546 204134 -3462
rect 203514 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 204134 -3546
rect 203514 -3814 204134 -3782
rect 207234 64894 207854 98000
rect 207234 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 207854 64894
rect 207234 64574 207854 64658
rect 207234 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 207854 64574
rect 207234 28894 207854 64338
rect 207234 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 207854 28894
rect 207234 28574 207854 28658
rect 207234 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 207854 28574
rect 207234 -5146 207854 28338
rect 207234 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 207854 -5146
rect 207234 -5466 207854 -5382
rect 207234 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 207854 -5466
rect 207234 -5734 207854 -5702
rect 210954 68614 211574 98000
rect 210954 68378 210986 68614
rect 211222 68378 211306 68614
rect 211542 68378 211574 68614
rect 210954 68294 211574 68378
rect 210954 68058 210986 68294
rect 211222 68058 211306 68294
rect 211542 68058 211574 68294
rect 210954 32614 211574 68058
rect 210954 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 211574 32614
rect 210954 32294 211574 32378
rect 210954 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 211574 32294
rect 192954 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 193574 -6106
rect 192954 -6426 193574 -6342
rect 192954 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 193574 -6426
rect 192954 -7654 193574 -6662
rect 210954 -7066 211574 32058
rect 217794 75454 218414 98000
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 217794 39454 218414 74898
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -1894 218414 -902
rect 221514 79174 222134 98000
rect 221514 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 222134 79174
rect 221514 78854 222134 78938
rect 221514 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 222134 78854
rect 221514 43174 222134 78618
rect 221514 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 222134 43174
rect 221514 42854 222134 42938
rect 221514 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 222134 42854
rect 221514 7174 222134 42618
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -2266 222134 6618
rect 221514 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 222134 -2266
rect 221514 -2586 222134 -2502
rect 221514 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 222134 -2586
rect 221514 -3814 222134 -2822
rect 225234 82894 225854 98000
rect 225234 82658 225266 82894
rect 225502 82658 225586 82894
rect 225822 82658 225854 82894
rect 225234 82574 225854 82658
rect 225234 82338 225266 82574
rect 225502 82338 225586 82574
rect 225822 82338 225854 82574
rect 225234 46894 225854 82338
rect 225234 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 225854 46894
rect 225234 46574 225854 46658
rect 225234 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 225854 46574
rect 225234 10894 225854 46338
rect 225234 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 225854 10894
rect 225234 10574 225854 10658
rect 225234 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 225854 10574
rect 225234 -4186 225854 10338
rect 225234 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 225854 -4186
rect 225234 -4506 225854 -4422
rect 225234 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 225854 -4506
rect 225234 -5734 225854 -4742
rect 228954 86614 229574 98000
rect 228954 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 229574 86614
rect 228954 86294 229574 86378
rect 228954 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 229574 86294
rect 228954 50614 229574 86058
rect 228954 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 229574 50614
rect 228954 50294 229574 50378
rect 228954 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 229574 50294
rect 228954 14614 229574 50058
rect 228954 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 229574 14614
rect 228954 14294 229574 14378
rect 228954 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 229574 14294
rect 210954 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 211574 -7066
rect 210954 -7386 211574 -7302
rect 210954 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 211574 -7386
rect 210954 -7654 211574 -7622
rect 228954 -6106 229574 14058
rect 235794 93454 236414 98000
rect 235794 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 236414 93454
rect 235794 93134 236414 93218
rect 235794 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 236414 93134
rect 235794 57454 236414 92898
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -1306 236414 20898
rect 235794 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 236414 -1306
rect 235794 -1626 236414 -1542
rect 235794 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 236414 -1626
rect 235794 -1894 236414 -1862
rect 239514 97174 240134 98000
rect 239514 96938 239546 97174
rect 239782 96938 239866 97174
rect 240102 96938 240134 97174
rect 239514 96854 240134 96938
rect 239514 96618 239546 96854
rect 239782 96618 239866 96854
rect 240102 96618 240134 96854
rect 239514 61174 240134 96618
rect 239514 60938 239546 61174
rect 239782 60938 239866 61174
rect 240102 60938 240134 61174
rect 239514 60854 240134 60938
rect 239514 60618 239546 60854
rect 239782 60618 239866 60854
rect 240102 60618 240134 60854
rect 239514 25174 240134 60618
rect 239514 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 240134 25174
rect 239514 24854 240134 24938
rect 239514 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 240134 24854
rect 239514 -3226 240134 24618
rect 239514 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 240134 -3226
rect 239514 -3546 240134 -3462
rect 239514 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 240134 -3546
rect 239514 -3814 240134 -3782
rect 243234 64894 243854 98000
rect 243234 64658 243266 64894
rect 243502 64658 243586 64894
rect 243822 64658 243854 64894
rect 243234 64574 243854 64658
rect 243234 64338 243266 64574
rect 243502 64338 243586 64574
rect 243822 64338 243854 64574
rect 243234 28894 243854 64338
rect 243234 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 243854 28894
rect 243234 28574 243854 28658
rect 243234 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 243854 28574
rect 243234 -5146 243854 28338
rect 243234 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 243854 -5146
rect 243234 -5466 243854 -5382
rect 243234 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 243854 -5466
rect 243234 -5734 243854 -5702
rect 246954 68614 247574 98000
rect 246954 68378 246986 68614
rect 247222 68378 247306 68614
rect 247542 68378 247574 68614
rect 246954 68294 247574 68378
rect 246954 68058 246986 68294
rect 247222 68058 247306 68294
rect 247542 68058 247574 68294
rect 246954 32614 247574 68058
rect 246954 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 247574 32614
rect 246954 32294 247574 32378
rect 246954 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 247574 32294
rect 228954 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 229574 -6106
rect 228954 -6426 229574 -6342
rect 228954 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 229574 -6426
rect 228954 -7654 229574 -6662
rect 246954 -7066 247574 32058
rect 253794 75454 254414 98000
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253794 39454 254414 74898
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -1894 254414 -902
rect 257514 79174 258134 98000
rect 257514 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 258134 79174
rect 257514 78854 258134 78938
rect 257514 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 258134 78854
rect 257514 43174 258134 78618
rect 257514 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 258134 43174
rect 257514 42854 258134 42938
rect 257514 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 258134 42854
rect 257514 7174 258134 42618
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 257514 -2266 258134 6618
rect 257514 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 258134 -2266
rect 257514 -2586 258134 -2502
rect 257514 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 258134 -2586
rect 257514 -3814 258134 -2822
rect 261234 82894 261854 98000
rect 261234 82658 261266 82894
rect 261502 82658 261586 82894
rect 261822 82658 261854 82894
rect 261234 82574 261854 82658
rect 261234 82338 261266 82574
rect 261502 82338 261586 82574
rect 261822 82338 261854 82574
rect 261234 46894 261854 82338
rect 261234 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 261854 46894
rect 261234 46574 261854 46658
rect 261234 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 261854 46574
rect 261234 10894 261854 46338
rect 261234 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 261854 10894
rect 261234 10574 261854 10658
rect 261234 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 261854 10574
rect 261234 -4186 261854 10338
rect 261234 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 261854 -4186
rect 261234 -4506 261854 -4422
rect 261234 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 261854 -4506
rect 261234 -5734 261854 -4742
rect 264954 86614 265574 98000
rect 264954 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 265574 86614
rect 264954 86294 265574 86378
rect 264954 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 265574 86294
rect 264954 50614 265574 86058
rect 264954 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 265574 50614
rect 264954 50294 265574 50378
rect 264954 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 265574 50294
rect 264954 14614 265574 50058
rect 264954 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 265574 14614
rect 264954 14294 265574 14378
rect 264954 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 265574 14294
rect 246954 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 247574 -7066
rect 246954 -7386 247574 -7302
rect 246954 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 247574 -7386
rect 246954 -7654 247574 -7622
rect 264954 -6106 265574 14058
rect 271794 93454 272414 98000
rect 271794 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 272414 93454
rect 271794 93134 272414 93218
rect 271794 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 272414 93134
rect 271794 57454 272414 92898
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -1306 272414 20898
rect 271794 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 272414 -1306
rect 271794 -1626 272414 -1542
rect 271794 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 272414 -1626
rect 271794 -1894 272414 -1862
rect 275514 97174 276134 98000
rect 275514 96938 275546 97174
rect 275782 96938 275866 97174
rect 276102 96938 276134 97174
rect 275514 96854 276134 96938
rect 275514 96618 275546 96854
rect 275782 96618 275866 96854
rect 276102 96618 276134 96854
rect 275514 61174 276134 96618
rect 275514 60938 275546 61174
rect 275782 60938 275866 61174
rect 276102 60938 276134 61174
rect 275514 60854 276134 60938
rect 275514 60618 275546 60854
rect 275782 60618 275866 60854
rect 276102 60618 276134 60854
rect 275514 25174 276134 60618
rect 275514 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 276134 25174
rect 275514 24854 276134 24938
rect 275514 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 276134 24854
rect 275514 -3226 276134 24618
rect 275514 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 276134 -3226
rect 275514 -3546 276134 -3462
rect 275514 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 276134 -3546
rect 275514 -3814 276134 -3782
rect 279234 64894 279854 98000
rect 279234 64658 279266 64894
rect 279502 64658 279586 64894
rect 279822 64658 279854 64894
rect 279234 64574 279854 64658
rect 279234 64338 279266 64574
rect 279502 64338 279586 64574
rect 279822 64338 279854 64574
rect 279234 28894 279854 64338
rect 279234 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 279854 28894
rect 279234 28574 279854 28658
rect 279234 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 279854 28574
rect 279234 -5146 279854 28338
rect 279234 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 279854 -5146
rect 279234 -5466 279854 -5382
rect 279234 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 279854 -5466
rect 279234 -5734 279854 -5702
rect 282954 68614 283574 98000
rect 282954 68378 282986 68614
rect 283222 68378 283306 68614
rect 283542 68378 283574 68614
rect 282954 68294 283574 68378
rect 282954 68058 282986 68294
rect 283222 68058 283306 68294
rect 283542 68058 283574 68294
rect 282954 32614 283574 68058
rect 282954 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 283574 32614
rect 282954 32294 283574 32378
rect 282954 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 283574 32294
rect 264954 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 265574 -6106
rect 264954 -6426 265574 -6342
rect 264954 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 265574 -6426
rect 264954 -7654 265574 -6662
rect 282954 -7066 283574 32058
rect 289794 75454 290414 98000
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 289794 39454 290414 74898
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -1894 290414 -902
rect 293514 79174 294134 98000
rect 293514 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 294134 79174
rect 293514 78854 294134 78938
rect 293514 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 294134 78854
rect 293514 43174 294134 78618
rect 293514 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 294134 43174
rect 293514 42854 294134 42938
rect 293514 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 294134 42854
rect 293514 7174 294134 42618
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 293514 -2266 294134 6618
rect 293514 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 294134 -2266
rect 293514 -2586 294134 -2502
rect 293514 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 294134 -2586
rect 293514 -3814 294134 -2822
rect 297234 82894 297854 98000
rect 297234 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 297854 82894
rect 297234 82574 297854 82658
rect 297234 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 297854 82574
rect 297234 46894 297854 82338
rect 297234 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 297854 46894
rect 297234 46574 297854 46658
rect 297234 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 297854 46574
rect 297234 10894 297854 46338
rect 297234 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 297854 10894
rect 297234 10574 297854 10658
rect 297234 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 297854 10574
rect 297234 -4186 297854 10338
rect 297234 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 297854 -4186
rect 297234 -4506 297854 -4422
rect 297234 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 297854 -4506
rect 297234 -5734 297854 -4742
rect 300954 86614 301574 98000
rect 300954 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 301574 86614
rect 300954 86294 301574 86378
rect 300954 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 301574 86294
rect 300954 50614 301574 86058
rect 300954 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 301574 50614
rect 300954 50294 301574 50378
rect 300954 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 301574 50294
rect 300954 14614 301574 50058
rect 300954 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 301574 14614
rect 300954 14294 301574 14378
rect 300954 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 301574 14294
rect 282954 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 283574 -7066
rect 282954 -7386 283574 -7302
rect 282954 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 283574 -7386
rect 282954 -7654 283574 -7622
rect 300954 -6106 301574 14058
rect 307794 93454 308414 128898
rect 307794 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 308414 93454
rect 307794 93134 308414 93218
rect 307794 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 308414 93134
rect 307794 57454 308414 92898
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -1306 308414 20898
rect 307794 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 308414 -1306
rect 307794 -1626 308414 -1542
rect 307794 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 308414 -1626
rect 307794 -1894 308414 -1862
rect 311514 673174 312134 707162
rect 311514 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 312134 673174
rect 311514 672854 312134 672938
rect 311514 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 312134 672854
rect 311514 637174 312134 672618
rect 311514 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 312134 637174
rect 311514 636854 312134 636938
rect 311514 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 312134 636854
rect 311514 601174 312134 636618
rect 311514 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 312134 601174
rect 311514 600854 312134 600938
rect 311514 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 312134 600854
rect 311514 565174 312134 600618
rect 311514 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 312134 565174
rect 311514 564854 312134 564938
rect 311514 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 312134 564854
rect 311514 529174 312134 564618
rect 311514 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 312134 529174
rect 311514 528854 312134 528938
rect 311514 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 312134 528854
rect 311514 493174 312134 528618
rect 311514 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 312134 493174
rect 311514 492854 312134 492938
rect 311514 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 312134 492854
rect 311514 457174 312134 492618
rect 311514 456938 311546 457174
rect 311782 456938 311866 457174
rect 312102 456938 312134 457174
rect 311514 456854 312134 456938
rect 311514 456618 311546 456854
rect 311782 456618 311866 456854
rect 312102 456618 312134 456854
rect 311514 421174 312134 456618
rect 311514 420938 311546 421174
rect 311782 420938 311866 421174
rect 312102 420938 312134 421174
rect 311514 420854 312134 420938
rect 311514 420618 311546 420854
rect 311782 420618 311866 420854
rect 312102 420618 312134 420854
rect 311514 385174 312134 420618
rect 311514 384938 311546 385174
rect 311782 384938 311866 385174
rect 312102 384938 312134 385174
rect 311514 384854 312134 384938
rect 311514 384618 311546 384854
rect 311782 384618 311866 384854
rect 312102 384618 312134 384854
rect 311514 349174 312134 384618
rect 311514 348938 311546 349174
rect 311782 348938 311866 349174
rect 312102 348938 312134 349174
rect 311514 348854 312134 348938
rect 311514 348618 311546 348854
rect 311782 348618 311866 348854
rect 312102 348618 312134 348854
rect 311514 313174 312134 348618
rect 311514 312938 311546 313174
rect 311782 312938 311866 313174
rect 312102 312938 312134 313174
rect 311514 312854 312134 312938
rect 311514 312618 311546 312854
rect 311782 312618 311866 312854
rect 312102 312618 312134 312854
rect 311514 277174 312134 312618
rect 311514 276938 311546 277174
rect 311782 276938 311866 277174
rect 312102 276938 312134 277174
rect 311514 276854 312134 276938
rect 311514 276618 311546 276854
rect 311782 276618 311866 276854
rect 312102 276618 312134 276854
rect 311514 241174 312134 276618
rect 311514 240938 311546 241174
rect 311782 240938 311866 241174
rect 312102 240938 312134 241174
rect 311514 240854 312134 240938
rect 311514 240618 311546 240854
rect 311782 240618 311866 240854
rect 312102 240618 312134 240854
rect 311514 205174 312134 240618
rect 311514 204938 311546 205174
rect 311782 204938 311866 205174
rect 312102 204938 312134 205174
rect 311514 204854 312134 204938
rect 311514 204618 311546 204854
rect 311782 204618 311866 204854
rect 312102 204618 312134 204854
rect 311514 169174 312134 204618
rect 311514 168938 311546 169174
rect 311782 168938 311866 169174
rect 312102 168938 312134 169174
rect 311514 168854 312134 168938
rect 311514 168618 311546 168854
rect 311782 168618 311866 168854
rect 312102 168618 312134 168854
rect 311514 133174 312134 168618
rect 311514 132938 311546 133174
rect 311782 132938 311866 133174
rect 312102 132938 312134 133174
rect 311514 132854 312134 132938
rect 311514 132618 311546 132854
rect 311782 132618 311866 132854
rect 312102 132618 312134 132854
rect 311514 97174 312134 132618
rect 311514 96938 311546 97174
rect 311782 96938 311866 97174
rect 312102 96938 312134 97174
rect 311514 96854 312134 96938
rect 311514 96618 311546 96854
rect 311782 96618 311866 96854
rect 312102 96618 312134 96854
rect 311514 61174 312134 96618
rect 311514 60938 311546 61174
rect 311782 60938 311866 61174
rect 312102 60938 312134 61174
rect 311514 60854 312134 60938
rect 311514 60618 311546 60854
rect 311782 60618 311866 60854
rect 312102 60618 312134 60854
rect 311514 25174 312134 60618
rect 311514 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 312134 25174
rect 311514 24854 312134 24938
rect 311514 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 312134 24854
rect 311514 -3226 312134 24618
rect 311514 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 312134 -3226
rect 311514 -3546 312134 -3462
rect 311514 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 312134 -3546
rect 311514 -3814 312134 -3782
rect 315234 676894 315854 709082
rect 315234 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 315854 676894
rect 315234 676574 315854 676658
rect 315234 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 315854 676574
rect 315234 640894 315854 676338
rect 315234 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 315854 640894
rect 315234 640574 315854 640658
rect 315234 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 315854 640574
rect 315234 604894 315854 640338
rect 315234 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 315854 604894
rect 315234 604574 315854 604658
rect 315234 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 315854 604574
rect 315234 568894 315854 604338
rect 315234 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 315854 568894
rect 315234 568574 315854 568658
rect 315234 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 315854 568574
rect 315234 532894 315854 568338
rect 315234 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 315854 532894
rect 315234 532574 315854 532658
rect 315234 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 315854 532574
rect 315234 496894 315854 532338
rect 315234 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 315854 496894
rect 315234 496574 315854 496658
rect 315234 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 315854 496574
rect 315234 460894 315854 496338
rect 315234 460658 315266 460894
rect 315502 460658 315586 460894
rect 315822 460658 315854 460894
rect 315234 460574 315854 460658
rect 315234 460338 315266 460574
rect 315502 460338 315586 460574
rect 315822 460338 315854 460574
rect 315234 424894 315854 460338
rect 315234 424658 315266 424894
rect 315502 424658 315586 424894
rect 315822 424658 315854 424894
rect 315234 424574 315854 424658
rect 315234 424338 315266 424574
rect 315502 424338 315586 424574
rect 315822 424338 315854 424574
rect 315234 388894 315854 424338
rect 315234 388658 315266 388894
rect 315502 388658 315586 388894
rect 315822 388658 315854 388894
rect 315234 388574 315854 388658
rect 315234 388338 315266 388574
rect 315502 388338 315586 388574
rect 315822 388338 315854 388574
rect 315234 352894 315854 388338
rect 315234 352658 315266 352894
rect 315502 352658 315586 352894
rect 315822 352658 315854 352894
rect 315234 352574 315854 352658
rect 315234 352338 315266 352574
rect 315502 352338 315586 352574
rect 315822 352338 315854 352574
rect 315234 316894 315854 352338
rect 315234 316658 315266 316894
rect 315502 316658 315586 316894
rect 315822 316658 315854 316894
rect 315234 316574 315854 316658
rect 315234 316338 315266 316574
rect 315502 316338 315586 316574
rect 315822 316338 315854 316574
rect 315234 280894 315854 316338
rect 315234 280658 315266 280894
rect 315502 280658 315586 280894
rect 315822 280658 315854 280894
rect 315234 280574 315854 280658
rect 315234 280338 315266 280574
rect 315502 280338 315586 280574
rect 315822 280338 315854 280574
rect 315234 244894 315854 280338
rect 315234 244658 315266 244894
rect 315502 244658 315586 244894
rect 315822 244658 315854 244894
rect 315234 244574 315854 244658
rect 315234 244338 315266 244574
rect 315502 244338 315586 244574
rect 315822 244338 315854 244574
rect 315234 208894 315854 244338
rect 315234 208658 315266 208894
rect 315502 208658 315586 208894
rect 315822 208658 315854 208894
rect 315234 208574 315854 208658
rect 315234 208338 315266 208574
rect 315502 208338 315586 208574
rect 315822 208338 315854 208574
rect 315234 172894 315854 208338
rect 315234 172658 315266 172894
rect 315502 172658 315586 172894
rect 315822 172658 315854 172894
rect 315234 172574 315854 172658
rect 315234 172338 315266 172574
rect 315502 172338 315586 172574
rect 315822 172338 315854 172574
rect 315234 136894 315854 172338
rect 315234 136658 315266 136894
rect 315502 136658 315586 136894
rect 315822 136658 315854 136894
rect 315234 136574 315854 136658
rect 315234 136338 315266 136574
rect 315502 136338 315586 136574
rect 315822 136338 315854 136574
rect 315234 100894 315854 136338
rect 315234 100658 315266 100894
rect 315502 100658 315586 100894
rect 315822 100658 315854 100894
rect 315234 100574 315854 100658
rect 315234 100338 315266 100574
rect 315502 100338 315586 100574
rect 315822 100338 315854 100574
rect 315234 64894 315854 100338
rect 315234 64658 315266 64894
rect 315502 64658 315586 64894
rect 315822 64658 315854 64894
rect 315234 64574 315854 64658
rect 315234 64338 315266 64574
rect 315502 64338 315586 64574
rect 315822 64338 315854 64574
rect 315234 28894 315854 64338
rect 315234 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 315854 28894
rect 315234 28574 315854 28658
rect 315234 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 315854 28574
rect 315234 -5146 315854 28338
rect 315234 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 315854 -5146
rect 315234 -5466 315854 -5382
rect 315234 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 315854 -5466
rect 315234 -5734 315854 -5702
rect 318954 680614 319574 711002
rect 336954 710598 337574 711590
rect 336954 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 337574 710598
rect 336954 710278 337574 710362
rect 336954 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 337574 710278
rect 333234 708678 333854 709670
rect 333234 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 333854 708678
rect 333234 708358 333854 708442
rect 333234 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 333854 708358
rect 329514 706758 330134 707750
rect 329514 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 330134 706758
rect 329514 706438 330134 706522
rect 329514 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 330134 706438
rect 318954 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 319574 680614
rect 318954 680294 319574 680378
rect 318954 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 319574 680294
rect 318954 644614 319574 680058
rect 318954 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 319574 644614
rect 318954 644294 319574 644378
rect 318954 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 319574 644294
rect 318954 608614 319574 644058
rect 318954 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 319574 608614
rect 318954 608294 319574 608378
rect 318954 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 319574 608294
rect 318954 572614 319574 608058
rect 318954 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 319574 572614
rect 318954 572294 319574 572378
rect 318954 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 319574 572294
rect 318954 536614 319574 572058
rect 318954 536378 318986 536614
rect 319222 536378 319306 536614
rect 319542 536378 319574 536614
rect 318954 536294 319574 536378
rect 318954 536058 318986 536294
rect 319222 536058 319306 536294
rect 319542 536058 319574 536294
rect 318954 500614 319574 536058
rect 318954 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 319574 500614
rect 318954 500294 319574 500378
rect 318954 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 319574 500294
rect 318954 464614 319574 500058
rect 318954 464378 318986 464614
rect 319222 464378 319306 464614
rect 319542 464378 319574 464614
rect 318954 464294 319574 464378
rect 318954 464058 318986 464294
rect 319222 464058 319306 464294
rect 319542 464058 319574 464294
rect 318954 428614 319574 464058
rect 318954 428378 318986 428614
rect 319222 428378 319306 428614
rect 319542 428378 319574 428614
rect 318954 428294 319574 428378
rect 318954 428058 318986 428294
rect 319222 428058 319306 428294
rect 319542 428058 319574 428294
rect 318954 392614 319574 428058
rect 318954 392378 318986 392614
rect 319222 392378 319306 392614
rect 319542 392378 319574 392614
rect 318954 392294 319574 392378
rect 318954 392058 318986 392294
rect 319222 392058 319306 392294
rect 319542 392058 319574 392294
rect 318954 356614 319574 392058
rect 318954 356378 318986 356614
rect 319222 356378 319306 356614
rect 319542 356378 319574 356614
rect 318954 356294 319574 356378
rect 318954 356058 318986 356294
rect 319222 356058 319306 356294
rect 319542 356058 319574 356294
rect 318954 320614 319574 356058
rect 318954 320378 318986 320614
rect 319222 320378 319306 320614
rect 319542 320378 319574 320614
rect 318954 320294 319574 320378
rect 318954 320058 318986 320294
rect 319222 320058 319306 320294
rect 319542 320058 319574 320294
rect 318954 284614 319574 320058
rect 318954 284378 318986 284614
rect 319222 284378 319306 284614
rect 319542 284378 319574 284614
rect 318954 284294 319574 284378
rect 318954 284058 318986 284294
rect 319222 284058 319306 284294
rect 319542 284058 319574 284294
rect 318954 248614 319574 284058
rect 318954 248378 318986 248614
rect 319222 248378 319306 248614
rect 319542 248378 319574 248614
rect 318954 248294 319574 248378
rect 318954 248058 318986 248294
rect 319222 248058 319306 248294
rect 319542 248058 319574 248294
rect 318954 212614 319574 248058
rect 318954 212378 318986 212614
rect 319222 212378 319306 212614
rect 319542 212378 319574 212614
rect 318954 212294 319574 212378
rect 318954 212058 318986 212294
rect 319222 212058 319306 212294
rect 319542 212058 319574 212294
rect 318954 176614 319574 212058
rect 318954 176378 318986 176614
rect 319222 176378 319306 176614
rect 319542 176378 319574 176614
rect 318954 176294 319574 176378
rect 318954 176058 318986 176294
rect 319222 176058 319306 176294
rect 319542 176058 319574 176294
rect 318954 140614 319574 176058
rect 318954 140378 318986 140614
rect 319222 140378 319306 140614
rect 319542 140378 319574 140614
rect 318954 140294 319574 140378
rect 318954 140058 318986 140294
rect 319222 140058 319306 140294
rect 319542 140058 319574 140294
rect 318954 104614 319574 140058
rect 318954 104378 318986 104614
rect 319222 104378 319306 104614
rect 319542 104378 319574 104614
rect 318954 104294 319574 104378
rect 318954 104058 318986 104294
rect 319222 104058 319306 104294
rect 319542 104058 319574 104294
rect 318954 68614 319574 104058
rect 318954 68378 318986 68614
rect 319222 68378 319306 68614
rect 319542 68378 319574 68614
rect 318954 68294 319574 68378
rect 318954 68058 318986 68294
rect 319222 68058 319306 68294
rect 319542 68058 319574 68294
rect 318954 32614 319574 68058
rect 318954 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 319574 32614
rect 318954 32294 319574 32378
rect 318954 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 319574 32294
rect 300954 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 301574 -6106
rect 300954 -6426 301574 -6342
rect 300954 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 301574 -6426
rect 300954 -7654 301574 -6662
rect 318954 -7066 319574 32058
rect 325794 704838 326414 705830
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 543454 326414 578898
rect 325794 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 326414 543454
rect 325794 543134 326414 543218
rect 325794 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 326414 543134
rect 325794 507454 326414 542898
rect 325794 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 326414 507454
rect 325794 507134 326414 507218
rect 325794 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 326414 507134
rect 325794 471454 326414 506898
rect 325794 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 326414 471454
rect 325794 471134 326414 471218
rect 325794 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 326414 471134
rect 325794 435454 326414 470898
rect 325794 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 326414 435454
rect 325794 435134 326414 435218
rect 325794 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 326414 435134
rect 325794 399454 326414 434898
rect 325794 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 326414 399454
rect 325794 399134 326414 399218
rect 325794 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 326414 399134
rect 325794 363454 326414 398898
rect 325794 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 326414 363454
rect 325794 363134 326414 363218
rect 325794 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 326414 363134
rect 325794 327454 326414 362898
rect 325794 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 326414 327454
rect 325794 327134 326414 327218
rect 325794 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 326414 327134
rect 325794 291454 326414 326898
rect 325794 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 326414 291454
rect 325794 291134 326414 291218
rect 325794 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 326414 291134
rect 325794 255454 326414 290898
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 325794 219454 326414 254898
rect 325794 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 326414 219454
rect 325794 219134 326414 219218
rect 325794 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 326414 219134
rect 325794 183454 326414 218898
rect 325794 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 326414 183454
rect 325794 183134 326414 183218
rect 325794 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 326414 183134
rect 325794 147454 326414 182898
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 325794 111454 326414 146898
rect 325794 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 326414 111454
rect 325794 111134 326414 111218
rect 325794 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 326414 111134
rect 325794 75454 326414 110898
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -1894 326414 -902
rect 329514 691174 330134 706202
rect 329514 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 330134 691174
rect 329514 690854 330134 690938
rect 329514 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 330134 690854
rect 329514 655174 330134 690618
rect 329514 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 330134 655174
rect 329514 654854 330134 654938
rect 329514 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 330134 654854
rect 329514 619174 330134 654618
rect 329514 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 330134 619174
rect 329514 618854 330134 618938
rect 329514 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 330134 618854
rect 329514 583174 330134 618618
rect 329514 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 330134 583174
rect 329514 582854 330134 582938
rect 329514 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 330134 582854
rect 329514 547174 330134 582618
rect 329514 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 330134 547174
rect 329514 546854 330134 546938
rect 329514 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 330134 546854
rect 329514 511174 330134 546618
rect 329514 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 330134 511174
rect 329514 510854 330134 510938
rect 329514 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 330134 510854
rect 329514 475174 330134 510618
rect 329514 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 330134 475174
rect 329514 474854 330134 474938
rect 329514 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 330134 474854
rect 329514 439174 330134 474618
rect 329514 438938 329546 439174
rect 329782 438938 329866 439174
rect 330102 438938 330134 439174
rect 329514 438854 330134 438938
rect 329514 438618 329546 438854
rect 329782 438618 329866 438854
rect 330102 438618 330134 438854
rect 329514 403174 330134 438618
rect 329514 402938 329546 403174
rect 329782 402938 329866 403174
rect 330102 402938 330134 403174
rect 329514 402854 330134 402938
rect 329514 402618 329546 402854
rect 329782 402618 329866 402854
rect 330102 402618 330134 402854
rect 329514 367174 330134 402618
rect 329514 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 330134 367174
rect 329514 366854 330134 366938
rect 329514 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 330134 366854
rect 329514 331174 330134 366618
rect 329514 330938 329546 331174
rect 329782 330938 329866 331174
rect 330102 330938 330134 331174
rect 329514 330854 330134 330938
rect 329514 330618 329546 330854
rect 329782 330618 329866 330854
rect 330102 330618 330134 330854
rect 329514 295174 330134 330618
rect 329514 294938 329546 295174
rect 329782 294938 329866 295174
rect 330102 294938 330134 295174
rect 329514 294854 330134 294938
rect 329514 294618 329546 294854
rect 329782 294618 329866 294854
rect 330102 294618 330134 294854
rect 329514 259174 330134 294618
rect 329514 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 330134 259174
rect 329514 258854 330134 258938
rect 329514 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 330134 258854
rect 329514 223174 330134 258618
rect 329514 222938 329546 223174
rect 329782 222938 329866 223174
rect 330102 222938 330134 223174
rect 329514 222854 330134 222938
rect 329514 222618 329546 222854
rect 329782 222618 329866 222854
rect 330102 222618 330134 222854
rect 329514 187174 330134 222618
rect 329514 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 330134 187174
rect 329514 186854 330134 186938
rect 329514 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 330134 186854
rect 329514 151174 330134 186618
rect 329514 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 330134 151174
rect 329514 150854 330134 150938
rect 329514 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 330134 150854
rect 329514 115174 330134 150618
rect 329514 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 330134 115174
rect 329514 114854 330134 114938
rect 329514 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 330134 114854
rect 329514 79174 330134 114618
rect 329514 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 330134 79174
rect 329514 78854 330134 78938
rect 329514 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 330134 78854
rect 329514 43174 330134 78618
rect 329514 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 330134 43174
rect 329514 42854 330134 42938
rect 329514 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 330134 42854
rect 329514 7174 330134 42618
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 329514 -2266 330134 6618
rect 329514 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 330134 -2266
rect 329514 -2586 330134 -2502
rect 329514 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 330134 -2586
rect 329514 -3814 330134 -2822
rect 333234 694894 333854 708122
rect 333234 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 333854 694894
rect 333234 694574 333854 694658
rect 333234 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 333854 694574
rect 333234 658894 333854 694338
rect 333234 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 333854 658894
rect 333234 658574 333854 658658
rect 333234 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 333854 658574
rect 333234 622894 333854 658338
rect 333234 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 333854 622894
rect 333234 622574 333854 622658
rect 333234 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 333854 622574
rect 333234 586894 333854 622338
rect 333234 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 333854 586894
rect 333234 586574 333854 586658
rect 333234 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 333854 586574
rect 333234 550894 333854 586338
rect 333234 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 333854 550894
rect 333234 550574 333854 550658
rect 333234 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 333854 550574
rect 333234 514894 333854 550338
rect 333234 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 333854 514894
rect 333234 514574 333854 514658
rect 333234 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 333854 514574
rect 333234 478894 333854 514338
rect 333234 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 333854 478894
rect 333234 478574 333854 478658
rect 333234 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 333854 478574
rect 333234 442894 333854 478338
rect 333234 442658 333266 442894
rect 333502 442658 333586 442894
rect 333822 442658 333854 442894
rect 333234 442574 333854 442658
rect 333234 442338 333266 442574
rect 333502 442338 333586 442574
rect 333822 442338 333854 442574
rect 333234 406894 333854 442338
rect 333234 406658 333266 406894
rect 333502 406658 333586 406894
rect 333822 406658 333854 406894
rect 333234 406574 333854 406658
rect 333234 406338 333266 406574
rect 333502 406338 333586 406574
rect 333822 406338 333854 406574
rect 333234 370894 333854 406338
rect 333234 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 333854 370894
rect 333234 370574 333854 370658
rect 333234 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 333854 370574
rect 333234 334894 333854 370338
rect 333234 334658 333266 334894
rect 333502 334658 333586 334894
rect 333822 334658 333854 334894
rect 333234 334574 333854 334658
rect 333234 334338 333266 334574
rect 333502 334338 333586 334574
rect 333822 334338 333854 334574
rect 333234 298894 333854 334338
rect 333234 298658 333266 298894
rect 333502 298658 333586 298894
rect 333822 298658 333854 298894
rect 333234 298574 333854 298658
rect 333234 298338 333266 298574
rect 333502 298338 333586 298574
rect 333822 298338 333854 298574
rect 333234 262894 333854 298338
rect 333234 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 333854 262894
rect 333234 262574 333854 262658
rect 333234 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 333854 262574
rect 333234 226894 333854 262338
rect 333234 226658 333266 226894
rect 333502 226658 333586 226894
rect 333822 226658 333854 226894
rect 333234 226574 333854 226658
rect 333234 226338 333266 226574
rect 333502 226338 333586 226574
rect 333822 226338 333854 226574
rect 333234 190894 333854 226338
rect 333234 190658 333266 190894
rect 333502 190658 333586 190894
rect 333822 190658 333854 190894
rect 333234 190574 333854 190658
rect 333234 190338 333266 190574
rect 333502 190338 333586 190574
rect 333822 190338 333854 190574
rect 333234 154894 333854 190338
rect 333234 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 333854 154894
rect 333234 154574 333854 154658
rect 333234 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 333854 154574
rect 333234 118894 333854 154338
rect 333234 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 333854 118894
rect 333234 118574 333854 118658
rect 333234 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 333854 118574
rect 333234 82894 333854 118338
rect 333234 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 333854 82894
rect 333234 82574 333854 82658
rect 333234 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 333854 82574
rect 333234 46894 333854 82338
rect 333234 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 333854 46894
rect 333234 46574 333854 46658
rect 333234 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 333854 46574
rect 333234 10894 333854 46338
rect 333234 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 333854 10894
rect 333234 10574 333854 10658
rect 333234 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 333854 10574
rect 333234 -4186 333854 10338
rect 333234 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 333854 -4186
rect 333234 -4506 333854 -4422
rect 333234 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 333854 -4506
rect 333234 -5734 333854 -4742
rect 336954 698614 337574 710042
rect 354954 711558 355574 711590
rect 354954 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 355574 711558
rect 354954 711238 355574 711322
rect 354954 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 355574 711238
rect 351234 709638 351854 709670
rect 351234 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 351854 709638
rect 351234 709318 351854 709402
rect 351234 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 351854 709318
rect 347514 707718 348134 707750
rect 347514 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 348134 707718
rect 347514 707398 348134 707482
rect 347514 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 348134 707398
rect 336954 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 337574 698614
rect 336954 698294 337574 698378
rect 336954 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 337574 698294
rect 336954 662614 337574 698058
rect 336954 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 337574 662614
rect 336954 662294 337574 662378
rect 336954 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 337574 662294
rect 336954 626614 337574 662058
rect 336954 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 337574 626614
rect 336954 626294 337574 626378
rect 336954 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 337574 626294
rect 336954 590614 337574 626058
rect 336954 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 337574 590614
rect 336954 590294 337574 590378
rect 336954 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 337574 590294
rect 336954 554614 337574 590058
rect 336954 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 337574 554614
rect 336954 554294 337574 554378
rect 336954 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 337574 554294
rect 336954 518614 337574 554058
rect 336954 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 337574 518614
rect 336954 518294 337574 518378
rect 336954 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 337574 518294
rect 336954 482614 337574 518058
rect 336954 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 337574 482614
rect 336954 482294 337574 482378
rect 336954 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 337574 482294
rect 336954 446614 337574 482058
rect 336954 446378 336986 446614
rect 337222 446378 337306 446614
rect 337542 446378 337574 446614
rect 336954 446294 337574 446378
rect 336954 446058 336986 446294
rect 337222 446058 337306 446294
rect 337542 446058 337574 446294
rect 336954 410614 337574 446058
rect 336954 410378 336986 410614
rect 337222 410378 337306 410614
rect 337542 410378 337574 410614
rect 336954 410294 337574 410378
rect 336954 410058 336986 410294
rect 337222 410058 337306 410294
rect 337542 410058 337574 410294
rect 336954 374614 337574 410058
rect 336954 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 337574 374614
rect 336954 374294 337574 374378
rect 336954 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 337574 374294
rect 336954 338614 337574 374058
rect 336954 338378 336986 338614
rect 337222 338378 337306 338614
rect 337542 338378 337574 338614
rect 336954 338294 337574 338378
rect 336954 338058 336986 338294
rect 337222 338058 337306 338294
rect 337542 338058 337574 338294
rect 336954 302614 337574 338058
rect 336954 302378 336986 302614
rect 337222 302378 337306 302614
rect 337542 302378 337574 302614
rect 336954 302294 337574 302378
rect 336954 302058 336986 302294
rect 337222 302058 337306 302294
rect 337542 302058 337574 302294
rect 336954 266614 337574 302058
rect 336954 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 337574 266614
rect 336954 266294 337574 266378
rect 336954 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 337574 266294
rect 336954 230614 337574 266058
rect 336954 230378 336986 230614
rect 337222 230378 337306 230614
rect 337542 230378 337574 230614
rect 336954 230294 337574 230378
rect 336954 230058 336986 230294
rect 337222 230058 337306 230294
rect 337542 230058 337574 230294
rect 336954 194614 337574 230058
rect 336954 194378 336986 194614
rect 337222 194378 337306 194614
rect 337542 194378 337574 194614
rect 336954 194294 337574 194378
rect 336954 194058 336986 194294
rect 337222 194058 337306 194294
rect 337542 194058 337574 194294
rect 336954 158614 337574 194058
rect 336954 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 337574 158614
rect 336954 158294 337574 158378
rect 336954 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 337574 158294
rect 336954 122614 337574 158058
rect 336954 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 337574 122614
rect 336954 122294 337574 122378
rect 336954 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 337574 122294
rect 336954 86614 337574 122058
rect 336954 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 337574 86614
rect 336954 86294 337574 86378
rect 336954 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 337574 86294
rect 336954 50614 337574 86058
rect 336954 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 337574 50614
rect 336954 50294 337574 50378
rect 336954 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 337574 50294
rect 336954 14614 337574 50058
rect 336954 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 337574 14614
rect 336954 14294 337574 14378
rect 336954 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 337574 14294
rect 318954 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 319574 -7066
rect 318954 -7386 319574 -7302
rect 318954 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 319574 -7386
rect 318954 -7654 319574 -7622
rect 336954 -6106 337574 14058
rect 343794 705798 344414 705830
rect 343794 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 344414 705798
rect 343794 705478 344414 705562
rect 343794 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 344414 705478
rect 343794 669454 344414 705242
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 561454 344414 596898
rect 343794 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 344414 561454
rect 343794 561134 344414 561218
rect 343794 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 344414 561134
rect 343794 525454 344414 560898
rect 343794 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 344414 525454
rect 343794 525134 344414 525218
rect 343794 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 344414 525134
rect 343794 489454 344414 524898
rect 343794 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 344414 489454
rect 343794 489134 344414 489218
rect 343794 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 344414 489134
rect 343794 453454 344414 488898
rect 343794 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 344414 453454
rect 343794 453134 344414 453218
rect 343794 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 344414 453134
rect 343794 417454 344414 452898
rect 343794 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 344414 417454
rect 343794 417134 344414 417218
rect 343794 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 344414 417134
rect 343794 381454 344414 416898
rect 343794 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 344414 381454
rect 343794 381134 344414 381218
rect 343794 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 344414 381134
rect 343794 345454 344414 380898
rect 343794 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 344414 345454
rect 343794 345134 344414 345218
rect 343794 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 344414 345134
rect 343794 309454 344414 344898
rect 343794 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 344414 309454
rect 343794 309134 344414 309218
rect 343794 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 344414 309134
rect 343794 273454 344414 308898
rect 343794 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 344414 273454
rect 343794 273134 344414 273218
rect 343794 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 344414 273134
rect 343794 237454 344414 272898
rect 343794 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 344414 237454
rect 343794 237134 344414 237218
rect 343794 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 344414 237134
rect 343794 201454 344414 236898
rect 343794 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 344414 201454
rect 343794 201134 344414 201218
rect 343794 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 344414 201134
rect 343794 165454 344414 200898
rect 343794 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 344414 165454
rect 343794 165134 344414 165218
rect 343794 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 344414 165134
rect 343794 129454 344414 164898
rect 343794 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 344414 129454
rect 343794 129134 344414 129218
rect 343794 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 344414 129134
rect 343794 93454 344414 128898
rect 343794 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 344414 93454
rect 343794 93134 344414 93218
rect 343794 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 344414 93134
rect 343794 57454 344414 92898
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -1306 344414 20898
rect 343794 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 344414 -1306
rect 343794 -1626 344414 -1542
rect 343794 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 344414 -1626
rect 343794 -1894 344414 -1862
rect 347514 673174 348134 707162
rect 347514 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 348134 673174
rect 347514 672854 348134 672938
rect 347514 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 348134 672854
rect 347514 637174 348134 672618
rect 347514 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 348134 637174
rect 347514 636854 348134 636938
rect 347514 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 348134 636854
rect 347514 601174 348134 636618
rect 347514 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 348134 601174
rect 347514 600854 348134 600938
rect 347514 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 348134 600854
rect 347514 565174 348134 600618
rect 347514 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 348134 565174
rect 347514 564854 348134 564938
rect 347514 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 348134 564854
rect 347514 529174 348134 564618
rect 347514 528938 347546 529174
rect 347782 528938 347866 529174
rect 348102 528938 348134 529174
rect 347514 528854 348134 528938
rect 347514 528618 347546 528854
rect 347782 528618 347866 528854
rect 348102 528618 348134 528854
rect 347514 493174 348134 528618
rect 347514 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 348134 493174
rect 347514 492854 348134 492938
rect 347514 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 348134 492854
rect 347514 457174 348134 492618
rect 347514 456938 347546 457174
rect 347782 456938 347866 457174
rect 348102 456938 348134 457174
rect 347514 456854 348134 456938
rect 347514 456618 347546 456854
rect 347782 456618 347866 456854
rect 348102 456618 348134 456854
rect 347514 421174 348134 456618
rect 347514 420938 347546 421174
rect 347782 420938 347866 421174
rect 348102 420938 348134 421174
rect 347514 420854 348134 420938
rect 347514 420618 347546 420854
rect 347782 420618 347866 420854
rect 348102 420618 348134 420854
rect 347514 385174 348134 420618
rect 347514 384938 347546 385174
rect 347782 384938 347866 385174
rect 348102 384938 348134 385174
rect 347514 384854 348134 384938
rect 347514 384618 347546 384854
rect 347782 384618 347866 384854
rect 348102 384618 348134 384854
rect 347514 349174 348134 384618
rect 347514 348938 347546 349174
rect 347782 348938 347866 349174
rect 348102 348938 348134 349174
rect 347514 348854 348134 348938
rect 347514 348618 347546 348854
rect 347782 348618 347866 348854
rect 348102 348618 348134 348854
rect 347514 313174 348134 348618
rect 347514 312938 347546 313174
rect 347782 312938 347866 313174
rect 348102 312938 348134 313174
rect 347514 312854 348134 312938
rect 347514 312618 347546 312854
rect 347782 312618 347866 312854
rect 348102 312618 348134 312854
rect 347514 277174 348134 312618
rect 347514 276938 347546 277174
rect 347782 276938 347866 277174
rect 348102 276938 348134 277174
rect 347514 276854 348134 276938
rect 347514 276618 347546 276854
rect 347782 276618 347866 276854
rect 348102 276618 348134 276854
rect 347514 241174 348134 276618
rect 347514 240938 347546 241174
rect 347782 240938 347866 241174
rect 348102 240938 348134 241174
rect 347514 240854 348134 240938
rect 347514 240618 347546 240854
rect 347782 240618 347866 240854
rect 348102 240618 348134 240854
rect 347514 205174 348134 240618
rect 347514 204938 347546 205174
rect 347782 204938 347866 205174
rect 348102 204938 348134 205174
rect 347514 204854 348134 204938
rect 347514 204618 347546 204854
rect 347782 204618 347866 204854
rect 348102 204618 348134 204854
rect 347514 169174 348134 204618
rect 347514 168938 347546 169174
rect 347782 168938 347866 169174
rect 348102 168938 348134 169174
rect 347514 168854 348134 168938
rect 347514 168618 347546 168854
rect 347782 168618 347866 168854
rect 348102 168618 348134 168854
rect 347514 133174 348134 168618
rect 347514 132938 347546 133174
rect 347782 132938 347866 133174
rect 348102 132938 348134 133174
rect 347514 132854 348134 132938
rect 347514 132618 347546 132854
rect 347782 132618 347866 132854
rect 348102 132618 348134 132854
rect 347514 97174 348134 132618
rect 347514 96938 347546 97174
rect 347782 96938 347866 97174
rect 348102 96938 348134 97174
rect 347514 96854 348134 96938
rect 347514 96618 347546 96854
rect 347782 96618 347866 96854
rect 348102 96618 348134 96854
rect 347514 61174 348134 96618
rect 347514 60938 347546 61174
rect 347782 60938 347866 61174
rect 348102 60938 348134 61174
rect 347514 60854 348134 60938
rect 347514 60618 347546 60854
rect 347782 60618 347866 60854
rect 348102 60618 348134 60854
rect 347514 25174 348134 60618
rect 347514 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 348134 25174
rect 347514 24854 348134 24938
rect 347514 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 348134 24854
rect 347514 -3226 348134 24618
rect 347514 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 348134 -3226
rect 347514 -3546 348134 -3462
rect 347514 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 348134 -3546
rect 347514 -3814 348134 -3782
rect 351234 676894 351854 709082
rect 351234 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 351854 676894
rect 351234 676574 351854 676658
rect 351234 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 351854 676574
rect 351234 640894 351854 676338
rect 351234 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 351854 640894
rect 351234 640574 351854 640658
rect 351234 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 351854 640574
rect 351234 604894 351854 640338
rect 351234 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 351854 604894
rect 351234 604574 351854 604658
rect 351234 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 351854 604574
rect 351234 568894 351854 604338
rect 351234 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 351854 568894
rect 351234 568574 351854 568658
rect 351234 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 351854 568574
rect 351234 532894 351854 568338
rect 351234 532658 351266 532894
rect 351502 532658 351586 532894
rect 351822 532658 351854 532894
rect 351234 532574 351854 532658
rect 351234 532338 351266 532574
rect 351502 532338 351586 532574
rect 351822 532338 351854 532574
rect 351234 496894 351854 532338
rect 351234 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 351854 496894
rect 351234 496574 351854 496658
rect 351234 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 351854 496574
rect 351234 460894 351854 496338
rect 351234 460658 351266 460894
rect 351502 460658 351586 460894
rect 351822 460658 351854 460894
rect 351234 460574 351854 460658
rect 351234 460338 351266 460574
rect 351502 460338 351586 460574
rect 351822 460338 351854 460574
rect 351234 424894 351854 460338
rect 351234 424658 351266 424894
rect 351502 424658 351586 424894
rect 351822 424658 351854 424894
rect 351234 424574 351854 424658
rect 351234 424338 351266 424574
rect 351502 424338 351586 424574
rect 351822 424338 351854 424574
rect 351234 388894 351854 424338
rect 351234 388658 351266 388894
rect 351502 388658 351586 388894
rect 351822 388658 351854 388894
rect 351234 388574 351854 388658
rect 351234 388338 351266 388574
rect 351502 388338 351586 388574
rect 351822 388338 351854 388574
rect 351234 352894 351854 388338
rect 351234 352658 351266 352894
rect 351502 352658 351586 352894
rect 351822 352658 351854 352894
rect 351234 352574 351854 352658
rect 351234 352338 351266 352574
rect 351502 352338 351586 352574
rect 351822 352338 351854 352574
rect 351234 316894 351854 352338
rect 351234 316658 351266 316894
rect 351502 316658 351586 316894
rect 351822 316658 351854 316894
rect 351234 316574 351854 316658
rect 351234 316338 351266 316574
rect 351502 316338 351586 316574
rect 351822 316338 351854 316574
rect 351234 280894 351854 316338
rect 351234 280658 351266 280894
rect 351502 280658 351586 280894
rect 351822 280658 351854 280894
rect 351234 280574 351854 280658
rect 351234 280338 351266 280574
rect 351502 280338 351586 280574
rect 351822 280338 351854 280574
rect 351234 244894 351854 280338
rect 351234 244658 351266 244894
rect 351502 244658 351586 244894
rect 351822 244658 351854 244894
rect 351234 244574 351854 244658
rect 351234 244338 351266 244574
rect 351502 244338 351586 244574
rect 351822 244338 351854 244574
rect 351234 208894 351854 244338
rect 351234 208658 351266 208894
rect 351502 208658 351586 208894
rect 351822 208658 351854 208894
rect 351234 208574 351854 208658
rect 351234 208338 351266 208574
rect 351502 208338 351586 208574
rect 351822 208338 351854 208574
rect 351234 172894 351854 208338
rect 351234 172658 351266 172894
rect 351502 172658 351586 172894
rect 351822 172658 351854 172894
rect 351234 172574 351854 172658
rect 351234 172338 351266 172574
rect 351502 172338 351586 172574
rect 351822 172338 351854 172574
rect 351234 136894 351854 172338
rect 351234 136658 351266 136894
rect 351502 136658 351586 136894
rect 351822 136658 351854 136894
rect 351234 136574 351854 136658
rect 351234 136338 351266 136574
rect 351502 136338 351586 136574
rect 351822 136338 351854 136574
rect 351234 100894 351854 136338
rect 351234 100658 351266 100894
rect 351502 100658 351586 100894
rect 351822 100658 351854 100894
rect 351234 100574 351854 100658
rect 351234 100338 351266 100574
rect 351502 100338 351586 100574
rect 351822 100338 351854 100574
rect 351234 64894 351854 100338
rect 351234 64658 351266 64894
rect 351502 64658 351586 64894
rect 351822 64658 351854 64894
rect 351234 64574 351854 64658
rect 351234 64338 351266 64574
rect 351502 64338 351586 64574
rect 351822 64338 351854 64574
rect 351234 28894 351854 64338
rect 351234 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 351854 28894
rect 351234 28574 351854 28658
rect 351234 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 351854 28574
rect 351234 -5146 351854 28338
rect 351234 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 351854 -5146
rect 351234 -5466 351854 -5382
rect 351234 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 351854 -5466
rect 351234 -5734 351854 -5702
rect 354954 680614 355574 711002
rect 372954 710598 373574 711590
rect 372954 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 373574 710598
rect 372954 710278 373574 710362
rect 372954 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 373574 710278
rect 369234 708678 369854 709670
rect 369234 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 369854 708678
rect 369234 708358 369854 708442
rect 369234 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 369854 708358
rect 365514 706758 366134 707750
rect 365514 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 366134 706758
rect 365514 706438 366134 706522
rect 365514 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 366134 706438
rect 354954 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 355574 680614
rect 354954 680294 355574 680378
rect 354954 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 355574 680294
rect 354954 644614 355574 680058
rect 354954 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 355574 644614
rect 354954 644294 355574 644378
rect 354954 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 355574 644294
rect 354954 608614 355574 644058
rect 354954 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 355574 608614
rect 354954 608294 355574 608378
rect 354954 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 355574 608294
rect 354954 572614 355574 608058
rect 354954 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 355574 572614
rect 354954 572294 355574 572378
rect 354954 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 355574 572294
rect 354954 536614 355574 572058
rect 354954 536378 354986 536614
rect 355222 536378 355306 536614
rect 355542 536378 355574 536614
rect 354954 536294 355574 536378
rect 354954 536058 354986 536294
rect 355222 536058 355306 536294
rect 355542 536058 355574 536294
rect 354954 500614 355574 536058
rect 354954 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 355574 500614
rect 354954 500294 355574 500378
rect 354954 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 355574 500294
rect 354954 464614 355574 500058
rect 354954 464378 354986 464614
rect 355222 464378 355306 464614
rect 355542 464378 355574 464614
rect 354954 464294 355574 464378
rect 354954 464058 354986 464294
rect 355222 464058 355306 464294
rect 355542 464058 355574 464294
rect 354954 428614 355574 464058
rect 354954 428378 354986 428614
rect 355222 428378 355306 428614
rect 355542 428378 355574 428614
rect 354954 428294 355574 428378
rect 354954 428058 354986 428294
rect 355222 428058 355306 428294
rect 355542 428058 355574 428294
rect 354954 392614 355574 428058
rect 354954 392378 354986 392614
rect 355222 392378 355306 392614
rect 355542 392378 355574 392614
rect 354954 392294 355574 392378
rect 354954 392058 354986 392294
rect 355222 392058 355306 392294
rect 355542 392058 355574 392294
rect 354954 356614 355574 392058
rect 361794 704838 362414 705830
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 435454 362414 470898
rect 361794 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 362414 435454
rect 361794 435134 362414 435218
rect 361794 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 362414 435134
rect 361794 399454 362414 434898
rect 361794 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 362414 399454
rect 361794 399134 362414 399218
rect 361794 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 362414 399134
rect 361794 372000 362414 398898
rect 365514 691174 366134 706202
rect 365514 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 366134 691174
rect 365514 690854 366134 690938
rect 365514 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 366134 690854
rect 365514 655174 366134 690618
rect 365514 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 366134 655174
rect 365514 654854 366134 654938
rect 365514 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 366134 654854
rect 365514 619174 366134 654618
rect 365514 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 366134 619174
rect 365514 618854 366134 618938
rect 365514 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 366134 618854
rect 365514 583174 366134 618618
rect 365514 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 366134 583174
rect 365514 582854 366134 582938
rect 365514 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 366134 582854
rect 365514 547174 366134 582618
rect 365514 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 366134 547174
rect 365514 546854 366134 546938
rect 365514 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 366134 546854
rect 365514 511174 366134 546618
rect 365514 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 366134 511174
rect 365514 510854 366134 510938
rect 365514 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 366134 510854
rect 365514 475174 366134 510618
rect 365514 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 366134 475174
rect 365514 474854 366134 474938
rect 365514 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 366134 474854
rect 365514 439174 366134 474618
rect 365514 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 366134 439174
rect 365514 438854 366134 438938
rect 365514 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 366134 438854
rect 365514 403174 366134 438618
rect 365514 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 366134 403174
rect 365514 402854 366134 402938
rect 365514 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 366134 402854
rect 365514 372000 366134 402618
rect 369234 694894 369854 708122
rect 369234 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 369854 694894
rect 369234 694574 369854 694658
rect 369234 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 369854 694574
rect 369234 658894 369854 694338
rect 369234 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 369854 658894
rect 369234 658574 369854 658658
rect 369234 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 369854 658574
rect 369234 622894 369854 658338
rect 369234 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 369854 622894
rect 369234 622574 369854 622658
rect 369234 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 369854 622574
rect 369234 586894 369854 622338
rect 369234 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 369854 586894
rect 369234 586574 369854 586658
rect 369234 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 369854 586574
rect 369234 550894 369854 586338
rect 369234 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 369854 550894
rect 369234 550574 369854 550658
rect 369234 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 369854 550574
rect 369234 514894 369854 550338
rect 369234 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 369854 514894
rect 369234 514574 369854 514658
rect 369234 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 369854 514574
rect 369234 478894 369854 514338
rect 369234 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 369854 478894
rect 369234 478574 369854 478658
rect 369234 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 369854 478574
rect 369234 442894 369854 478338
rect 369234 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 369854 442894
rect 369234 442574 369854 442658
rect 369234 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 369854 442574
rect 369234 406894 369854 442338
rect 369234 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 369854 406894
rect 369234 406574 369854 406658
rect 369234 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 369854 406574
rect 369234 372000 369854 406338
rect 372954 698614 373574 710042
rect 390954 711558 391574 711590
rect 390954 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 391574 711558
rect 390954 711238 391574 711322
rect 390954 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 391574 711238
rect 387234 709638 387854 709670
rect 387234 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 387854 709638
rect 387234 709318 387854 709402
rect 387234 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 387854 709318
rect 383514 707718 384134 707750
rect 383514 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 384134 707718
rect 383514 707398 384134 707482
rect 383514 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 384134 707398
rect 372954 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 373574 698614
rect 372954 698294 373574 698378
rect 372954 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 373574 698294
rect 372954 662614 373574 698058
rect 372954 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 373574 662614
rect 372954 662294 373574 662378
rect 372954 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 373574 662294
rect 372954 626614 373574 662058
rect 372954 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 373574 626614
rect 372954 626294 373574 626378
rect 372954 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 373574 626294
rect 372954 590614 373574 626058
rect 372954 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 373574 590614
rect 372954 590294 373574 590378
rect 372954 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 373574 590294
rect 372954 554614 373574 590058
rect 372954 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 373574 554614
rect 372954 554294 373574 554378
rect 372954 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 373574 554294
rect 372954 518614 373574 554058
rect 372954 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 373574 518614
rect 372954 518294 373574 518378
rect 372954 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 373574 518294
rect 372954 482614 373574 518058
rect 372954 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 373574 482614
rect 372954 482294 373574 482378
rect 372954 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 373574 482294
rect 372954 446614 373574 482058
rect 372954 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 373574 446614
rect 372954 446294 373574 446378
rect 372954 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 373574 446294
rect 372954 410614 373574 446058
rect 372954 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 373574 410614
rect 372954 410294 373574 410378
rect 372954 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 373574 410294
rect 372954 374614 373574 410058
rect 372954 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 373574 374614
rect 372954 374294 373574 374378
rect 372954 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 373574 374294
rect 362243 363454 362563 363486
rect 362243 363218 362285 363454
rect 362521 363218 362563 363454
rect 362243 363134 362563 363218
rect 362243 362898 362285 363134
rect 362521 362898 362563 363134
rect 362243 362866 362563 362898
rect 364840 363454 365160 363486
rect 364840 363218 364882 363454
rect 365118 363218 365160 363454
rect 364840 363134 365160 363218
rect 364840 362898 364882 363134
rect 365118 362898 365160 363134
rect 364840 362866 365160 362898
rect 367437 363454 367757 363486
rect 367437 363218 367479 363454
rect 367715 363218 367757 363454
rect 367437 363134 367757 363218
rect 367437 362898 367479 363134
rect 367715 362898 367757 363134
rect 367437 362866 367757 362898
rect 354954 356378 354986 356614
rect 355222 356378 355306 356614
rect 355542 356378 355574 356614
rect 354954 356294 355574 356378
rect 354954 356058 354986 356294
rect 355222 356058 355306 356294
rect 355542 356058 355574 356294
rect 354954 320614 355574 356058
rect 372107 352476 372173 352477
rect 372107 352412 372108 352476
rect 372172 352412 372173 352476
rect 372107 352411 372173 352412
rect 371739 351388 371805 351389
rect 371739 351324 371740 351388
rect 371804 351324 371805 351388
rect 371739 351323 371805 351324
rect 371371 350844 371437 350845
rect 371371 350780 371372 350844
rect 371436 350780 371437 350844
rect 371371 350779 371437 350780
rect 363541 345454 363861 345486
rect 363541 345218 363583 345454
rect 363819 345218 363861 345454
rect 363541 345134 363861 345218
rect 363541 344898 363583 345134
rect 363819 344898 363861 345134
rect 363541 344866 363861 344898
rect 366138 345454 366458 345486
rect 366138 345218 366180 345454
rect 366416 345218 366458 345454
rect 366138 345134 366458 345218
rect 366138 344898 366180 345134
rect 366416 344898 366458 345134
rect 366138 344866 366458 344898
rect 371187 343364 371253 343365
rect 371187 343300 371188 343364
rect 371252 343300 371253 343364
rect 371187 343299 371253 343300
rect 361619 337788 361685 337789
rect 361619 337724 361620 337788
rect 361684 337724 361685 337788
rect 361619 337723 361685 337724
rect 354954 320378 354986 320614
rect 355222 320378 355306 320614
rect 355542 320378 355574 320614
rect 354954 320294 355574 320378
rect 354954 320058 354986 320294
rect 355222 320058 355306 320294
rect 355542 320058 355574 320294
rect 354954 284614 355574 320058
rect 354954 284378 354986 284614
rect 355222 284378 355306 284614
rect 355542 284378 355574 284614
rect 354954 284294 355574 284378
rect 354954 284058 354986 284294
rect 355222 284058 355306 284294
rect 355542 284058 355574 284294
rect 354954 248614 355574 284058
rect 361622 266117 361682 337723
rect 361794 327454 362414 338000
rect 364379 337788 364445 337789
rect 364379 337724 364380 337788
rect 364444 337724 364445 337788
rect 364379 337723 364445 337724
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 361794 300000 362414 326898
rect 362243 291454 362563 291486
rect 362243 291218 362285 291454
rect 362521 291218 362563 291454
rect 362243 291134 362563 291218
rect 362243 290898 362285 291134
rect 362521 290898 362563 291134
rect 362243 290866 362563 290898
rect 363541 273454 363861 273486
rect 363541 273218 363583 273454
rect 363819 273218 363861 273454
rect 363541 273134 363861 273218
rect 363541 272898 363583 273134
rect 363819 272898 363861 273134
rect 363541 272866 363861 272898
rect 364382 266117 364442 337723
rect 365514 331174 366134 338000
rect 365514 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 366134 331174
rect 365514 330854 366134 330938
rect 365514 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 366134 330854
rect 365514 300000 366134 330618
rect 369234 334894 369854 338000
rect 369234 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 369854 334894
rect 369234 334574 369854 334658
rect 369234 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 369854 334574
rect 369234 300000 369854 334338
rect 364840 291454 365160 291486
rect 364840 291218 364882 291454
rect 365118 291218 365160 291454
rect 364840 291134 365160 291218
rect 364840 290898 364882 291134
rect 365118 290898 365160 291134
rect 364840 290866 365160 290898
rect 367437 291454 367757 291486
rect 367437 291218 367479 291454
rect 367715 291218 367757 291454
rect 367437 291134 367757 291218
rect 367437 290898 367479 291134
rect 367715 290898 367757 291134
rect 367437 290866 367757 290898
rect 370267 274820 370333 274821
rect 370267 274756 370268 274820
rect 370332 274756 370333 274820
rect 370267 274755 370333 274756
rect 366138 273454 366458 273486
rect 366138 273218 366180 273454
rect 366416 273218 366458 273454
rect 366138 273134 366458 273218
rect 366138 272898 366180 273134
rect 366416 272898 366458 273134
rect 366138 272866 366458 272898
rect 370083 268428 370149 268429
rect 370083 268364 370084 268428
rect 370148 268364 370149 268428
rect 370083 268363 370149 268364
rect 361619 266116 361685 266117
rect 361619 266052 361620 266116
rect 361684 266052 361685 266116
rect 361619 266051 361685 266052
rect 364379 266116 364445 266117
rect 364379 266052 364380 266116
rect 364444 266052 364445 266116
rect 364379 266051 364445 266052
rect 354954 248378 354986 248614
rect 355222 248378 355306 248614
rect 355542 248378 355574 248614
rect 354954 248294 355574 248378
rect 354954 248058 354986 248294
rect 355222 248058 355306 248294
rect 355542 248058 355574 248294
rect 354954 212614 355574 248058
rect 354954 212378 354986 212614
rect 355222 212378 355306 212614
rect 355542 212378 355574 212614
rect 354954 212294 355574 212378
rect 354954 212058 354986 212294
rect 355222 212058 355306 212294
rect 355542 212058 355574 212294
rect 354954 176614 355574 212058
rect 361622 194581 361682 266051
rect 361794 255454 362414 266000
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 228000 362414 254898
rect 362243 219454 362563 219486
rect 362243 219218 362285 219454
rect 362521 219218 362563 219454
rect 362243 219134 362563 219218
rect 362243 218898 362285 219134
rect 362521 218898 362563 219134
rect 362243 218866 362563 218898
rect 363541 201454 363861 201486
rect 363541 201218 363583 201454
rect 363819 201218 363861 201454
rect 363541 201134 363861 201218
rect 363541 200898 363583 201134
rect 363819 200898 363861 201134
rect 363541 200866 363861 200898
rect 364382 196077 364442 266051
rect 365514 259174 366134 266000
rect 365514 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 366134 259174
rect 365514 258854 366134 258938
rect 365514 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 366134 258854
rect 365514 228000 366134 258618
rect 369234 262894 369854 266000
rect 369234 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 369854 262894
rect 369234 262574 369854 262658
rect 369234 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 369854 262574
rect 369234 228000 369854 262338
rect 364840 219454 365160 219486
rect 364840 219218 364882 219454
rect 365118 219218 365160 219454
rect 364840 219134 365160 219218
rect 364840 218898 364882 219134
rect 365118 218898 365160 219134
rect 364840 218866 365160 218898
rect 367437 219454 367757 219486
rect 367437 219218 367479 219454
rect 367715 219218 367757 219454
rect 367437 219134 367757 219218
rect 367437 218898 367479 219134
rect 367715 218898 367757 219134
rect 367437 218866 367757 218898
rect 366138 201454 366458 201486
rect 366138 201218 366180 201454
rect 366416 201218 366458 201454
rect 366138 201134 366458 201218
rect 366138 200898 366180 201134
rect 366416 200898 366458 201134
rect 366138 200866 366458 200898
rect 370086 196621 370146 268363
rect 370270 203149 370330 274755
rect 371190 271421 371250 343299
rect 371374 278901 371434 350779
rect 371742 279445 371802 351323
rect 372110 280533 372170 352411
rect 372954 338614 373574 374058
rect 372954 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 373574 338614
rect 372954 338294 373574 338378
rect 372954 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 373574 338294
rect 372954 302614 373574 338058
rect 372954 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 373574 302614
rect 372954 302294 373574 302378
rect 372954 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 373574 302294
rect 372107 280532 372173 280533
rect 372107 280468 372108 280532
rect 372172 280468 372173 280532
rect 372107 280467 372173 280468
rect 371923 279988 371989 279989
rect 371923 279924 371924 279988
rect 371988 279924 371989 279988
rect 371923 279923 371989 279924
rect 371739 279444 371805 279445
rect 371739 279380 371740 279444
rect 371804 279380 371805 279444
rect 371739 279379 371805 279380
rect 371371 278900 371437 278901
rect 371371 278836 371372 278900
rect 371436 278836 371437 278900
rect 371371 278835 371437 278836
rect 371187 271420 371253 271421
rect 371187 271356 371188 271420
rect 371252 271356 371253 271420
rect 371187 271355 371253 271356
rect 371190 267750 371250 271355
rect 371190 267690 371434 267750
rect 370267 203148 370333 203149
rect 370267 203084 370268 203148
rect 370332 203084 370333 203148
rect 370267 203083 370333 203084
rect 371374 199341 371434 267690
rect 371926 208453 371986 279923
rect 372110 225045 372170 280467
rect 372954 266614 373574 302058
rect 372954 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 373574 266614
rect 372954 266294 373574 266378
rect 372954 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 373574 266294
rect 372954 230614 373574 266058
rect 372954 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 373574 230614
rect 372954 230294 373574 230378
rect 372954 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 373574 230294
rect 372107 225044 372173 225045
rect 372107 224980 372108 225044
rect 372172 224980 372173 225044
rect 372107 224979 372173 224980
rect 371923 208452 371989 208453
rect 371923 208388 371924 208452
rect 371988 208388 371989 208452
rect 371923 208387 371989 208388
rect 371371 199340 371437 199341
rect 371371 199276 371372 199340
rect 371436 199276 371437 199340
rect 371371 199275 371437 199276
rect 370083 196620 370149 196621
rect 370083 196556 370084 196620
rect 370148 196556 370149 196620
rect 370083 196555 370149 196556
rect 364379 196076 364445 196077
rect 364379 196012 364380 196076
rect 364444 196012 364445 196076
rect 364379 196011 364445 196012
rect 372954 194614 373574 230058
rect 361619 194580 361685 194581
rect 361619 194516 361620 194580
rect 361684 194516 361685 194580
rect 361619 194515 361685 194516
rect 362723 194580 362789 194581
rect 362723 194516 362724 194580
rect 362788 194516 362789 194580
rect 362723 194515 362789 194516
rect 365299 194580 365365 194581
rect 365299 194516 365300 194580
rect 365364 194516 365365 194580
rect 365299 194515 365365 194516
rect 354954 176378 354986 176614
rect 355222 176378 355306 176614
rect 355542 176378 355574 176614
rect 354954 176294 355574 176378
rect 354954 176058 354986 176294
rect 355222 176058 355306 176294
rect 355542 176058 355574 176294
rect 354954 140614 355574 176058
rect 361794 183454 362414 194000
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 361794 156000 362414 182898
rect 362243 147454 362563 147486
rect 362243 147218 362285 147454
rect 362521 147218 362563 147454
rect 362243 147134 362563 147218
rect 362243 146898 362285 147134
rect 362521 146898 362563 147134
rect 362243 146866 362563 146898
rect 354954 140378 354986 140614
rect 355222 140378 355306 140614
rect 355542 140378 355574 140614
rect 354954 140294 355574 140378
rect 354954 140058 354986 140294
rect 355222 140058 355306 140294
rect 355542 140058 355574 140294
rect 354954 104614 355574 140058
rect 362726 123997 362786 194515
rect 364840 147454 365160 147486
rect 364840 147218 364882 147454
rect 365118 147218 365160 147454
rect 364840 147134 365160 147218
rect 364840 146898 364882 147134
rect 365118 146898 365160 147134
rect 364840 146866 365160 146898
rect 363541 129454 363861 129486
rect 363541 129218 363583 129454
rect 363819 129218 363861 129454
rect 363541 129134 363861 129218
rect 363541 128898 363583 129134
rect 363819 128898 363861 129134
rect 363541 128866 363861 128898
rect 365302 123997 365362 194515
rect 372954 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 373574 194614
rect 372954 194294 373574 194378
rect 372954 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 373574 194294
rect 365514 187174 366134 194000
rect 365514 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 366134 187174
rect 365514 186854 366134 186938
rect 365514 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 366134 186854
rect 365514 156000 366134 186618
rect 369234 190894 369854 194000
rect 369234 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 369854 190894
rect 369234 190574 369854 190658
rect 369234 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 369854 190574
rect 369234 156000 369854 190338
rect 371739 159356 371805 159357
rect 371739 159292 371740 159356
rect 371804 159292 371805 159356
rect 371739 159291 371805 159292
rect 370083 153100 370149 153101
rect 370083 153036 370084 153100
rect 370148 153036 370149 153100
rect 370083 153035 370149 153036
rect 367437 147454 367757 147486
rect 367437 147218 367479 147454
rect 367715 147218 367757 147454
rect 367437 147134 367757 147218
rect 367437 146898 367479 147134
rect 367715 146898 367757 147134
rect 367437 146866 367757 146898
rect 370086 142170 370146 153035
rect 369902 142110 370146 142170
rect 369902 134061 369962 142110
rect 369899 134060 369965 134061
rect 369899 133996 369900 134060
rect 369964 133996 369965 134060
rect 369899 133995 369965 133996
rect 366138 129454 366458 129486
rect 366138 129218 366180 129454
rect 366416 129218 366458 129454
rect 366138 129134 366458 129218
rect 366138 128898 366180 129134
rect 366416 128898 366458 129134
rect 366138 128866 366458 128898
rect 371742 127397 371802 159291
rect 372954 158614 373574 194058
rect 372954 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 373574 158614
rect 372954 158294 373574 158378
rect 372954 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 373574 158294
rect 371739 127396 371805 127397
rect 371739 127332 371740 127396
rect 371804 127332 371805 127396
rect 371739 127331 371805 127332
rect 362723 123996 362789 123997
rect 362723 123932 362724 123996
rect 362788 123932 362789 123996
rect 362723 123931 362789 123932
rect 365299 123996 365365 123997
rect 365299 123932 365300 123996
rect 365364 123932 365365 123996
rect 365299 123931 365365 123932
rect 372954 122614 373574 158058
rect 372954 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 373574 122614
rect 372954 122294 373574 122378
rect 372954 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 373574 122294
rect 354954 104378 354986 104614
rect 355222 104378 355306 104614
rect 355542 104378 355574 104614
rect 354954 104294 355574 104378
rect 354954 104058 354986 104294
rect 355222 104058 355306 104294
rect 355542 104058 355574 104294
rect 354954 68614 355574 104058
rect 354954 68378 354986 68614
rect 355222 68378 355306 68614
rect 355542 68378 355574 68614
rect 354954 68294 355574 68378
rect 354954 68058 354986 68294
rect 355222 68058 355306 68294
rect 355542 68058 355574 68294
rect 354954 32614 355574 68058
rect 354954 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 355574 32614
rect 354954 32294 355574 32378
rect 354954 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 355574 32294
rect 336954 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 337574 -6106
rect 336954 -6426 337574 -6342
rect 336954 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 337574 -6426
rect 336954 -7654 337574 -6662
rect 354954 -7066 355574 32058
rect 361794 111454 362414 122000
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -1894 362414 -902
rect 365514 115174 366134 122000
rect 365514 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 366134 115174
rect 365514 114854 366134 114938
rect 365514 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 366134 114854
rect 365514 79174 366134 114618
rect 365514 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 366134 79174
rect 365514 78854 366134 78938
rect 365514 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 366134 78854
rect 365514 43174 366134 78618
rect 365514 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 366134 43174
rect 365514 42854 366134 42938
rect 365514 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 366134 42854
rect 365514 7174 366134 42618
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 365514 -2266 366134 6618
rect 365514 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 366134 -2266
rect 365514 -2586 366134 -2502
rect 365514 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 366134 -2586
rect 365514 -3814 366134 -2822
rect 369234 118894 369854 122000
rect 369234 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 369854 118894
rect 369234 118574 369854 118658
rect 369234 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 369854 118574
rect 369234 82894 369854 118338
rect 369234 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 369854 82894
rect 369234 82574 369854 82658
rect 369234 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 369854 82574
rect 369234 46894 369854 82338
rect 369234 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 369854 46894
rect 369234 46574 369854 46658
rect 369234 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 369854 46574
rect 369234 10894 369854 46338
rect 369234 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 369854 10894
rect 369234 10574 369854 10658
rect 369234 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 369854 10574
rect 369234 -4186 369854 10338
rect 369234 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 369854 -4186
rect 369234 -4506 369854 -4422
rect 369234 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 369854 -4506
rect 369234 -5734 369854 -4742
rect 372954 86614 373574 122058
rect 372954 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 373574 86614
rect 372954 86294 373574 86378
rect 372954 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 373574 86294
rect 372954 50614 373574 86058
rect 372954 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 373574 50614
rect 372954 50294 373574 50378
rect 372954 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 373574 50294
rect 372954 14614 373574 50058
rect 372954 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 373574 14614
rect 372954 14294 373574 14378
rect 372954 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 373574 14294
rect 354954 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 355574 -7066
rect 354954 -7386 355574 -7302
rect 354954 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 355574 -7386
rect 354954 -7654 355574 -7622
rect 372954 -6106 373574 14058
rect 379794 705798 380414 705830
rect 379794 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 380414 705798
rect 379794 705478 380414 705562
rect 379794 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 380414 705478
rect 379794 669454 380414 705242
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 561454 380414 596898
rect 379794 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 380414 561454
rect 379794 561134 380414 561218
rect 379794 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 380414 561134
rect 379794 525454 380414 560898
rect 379794 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 380414 525454
rect 379794 525134 380414 525218
rect 379794 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 380414 525134
rect 379794 489454 380414 524898
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 379794 489134 380414 489218
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 379794 453454 380414 488898
rect 379794 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 380414 453454
rect 379794 453134 380414 453218
rect 379794 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 380414 453134
rect 379794 417454 380414 452898
rect 379794 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 380414 417454
rect 379794 417134 380414 417218
rect 379794 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 380414 417134
rect 379794 381454 380414 416898
rect 379794 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 380414 381454
rect 379794 381134 380414 381218
rect 379794 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 380414 381134
rect 379794 345454 380414 380898
rect 379794 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 380414 345454
rect 379794 345134 380414 345218
rect 379794 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 380414 345134
rect 379794 309454 380414 344898
rect 379794 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 380414 309454
rect 379794 309134 380414 309218
rect 379794 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 380414 309134
rect 379794 273454 380414 308898
rect 379794 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 380414 273454
rect 379794 273134 380414 273218
rect 379794 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 380414 273134
rect 379794 237454 380414 272898
rect 379794 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 380414 237454
rect 379794 237134 380414 237218
rect 379794 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 380414 237134
rect 379794 201454 380414 236898
rect 379794 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 380414 201454
rect 379794 201134 380414 201218
rect 379794 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 380414 201134
rect 379794 165454 380414 200898
rect 379794 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 380414 165454
rect 379794 165134 380414 165218
rect 379794 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 380414 165134
rect 379794 129454 380414 164898
rect 379794 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 380414 129454
rect 379794 129134 380414 129218
rect 379794 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 380414 129134
rect 379794 93454 380414 128898
rect 379794 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 380414 93454
rect 379794 93134 380414 93218
rect 379794 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 380414 93134
rect 379794 57454 380414 92898
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -1306 380414 20898
rect 379794 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 380414 -1306
rect 379794 -1626 380414 -1542
rect 379794 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 380414 -1626
rect 379794 -1894 380414 -1862
rect 383514 673174 384134 707162
rect 383514 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 384134 673174
rect 383514 672854 384134 672938
rect 383514 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 384134 672854
rect 383514 637174 384134 672618
rect 383514 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 384134 637174
rect 383514 636854 384134 636938
rect 383514 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 384134 636854
rect 383514 601174 384134 636618
rect 383514 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 384134 601174
rect 383514 600854 384134 600938
rect 383514 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 384134 600854
rect 383514 565174 384134 600618
rect 383514 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 384134 565174
rect 383514 564854 384134 564938
rect 383514 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 384134 564854
rect 383514 529174 384134 564618
rect 383514 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 384134 529174
rect 383514 528854 384134 528938
rect 383514 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 384134 528854
rect 383514 493174 384134 528618
rect 383514 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 384134 493174
rect 383514 492854 384134 492938
rect 383514 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 384134 492854
rect 383514 457174 384134 492618
rect 383514 456938 383546 457174
rect 383782 456938 383866 457174
rect 384102 456938 384134 457174
rect 383514 456854 384134 456938
rect 383514 456618 383546 456854
rect 383782 456618 383866 456854
rect 384102 456618 384134 456854
rect 383514 421174 384134 456618
rect 383514 420938 383546 421174
rect 383782 420938 383866 421174
rect 384102 420938 384134 421174
rect 383514 420854 384134 420938
rect 383514 420618 383546 420854
rect 383782 420618 383866 420854
rect 384102 420618 384134 420854
rect 383514 385174 384134 420618
rect 383514 384938 383546 385174
rect 383782 384938 383866 385174
rect 384102 384938 384134 385174
rect 383514 384854 384134 384938
rect 383514 384618 383546 384854
rect 383782 384618 383866 384854
rect 384102 384618 384134 384854
rect 383514 349174 384134 384618
rect 383514 348938 383546 349174
rect 383782 348938 383866 349174
rect 384102 348938 384134 349174
rect 383514 348854 384134 348938
rect 383514 348618 383546 348854
rect 383782 348618 383866 348854
rect 384102 348618 384134 348854
rect 383514 313174 384134 348618
rect 383514 312938 383546 313174
rect 383782 312938 383866 313174
rect 384102 312938 384134 313174
rect 383514 312854 384134 312938
rect 383514 312618 383546 312854
rect 383782 312618 383866 312854
rect 384102 312618 384134 312854
rect 383514 277174 384134 312618
rect 383514 276938 383546 277174
rect 383782 276938 383866 277174
rect 384102 276938 384134 277174
rect 383514 276854 384134 276938
rect 383514 276618 383546 276854
rect 383782 276618 383866 276854
rect 384102 276618 384134 276854
rect 383514 241174 384134 276618
rect 383514 240938 383546 241174
rect 383782 240938 383866 241174
rect 384102 240938 384134 241174
rect 383514 240854 384134 240938
rect 383514 240618 383546 240854
rect 383782 240618 383866 240854
rect 384102 240618 384134 240854
rect 383514 205174 384134 240618
rect 383514 204938 383546 205174
rect 383782 204938 383866 205174
rect 384102 204938 384134 205174
rect 383514 204854 384134 204938
rect 383514 204618 383546 204854
rect 383782 204618 383866 204854
rect 384102 204618 384134 204854
rect 383514 169174 384134 204618
rect 383514 168938 383546 169174
rect 383782 168938 383866 169174
rect 384102 168938 384134 169174
rect 383514 168854 384134 168938
rect 383514 168618 383546 168854
rect 383782 168618 383866 168854
rect 384102 168618 384134 168854
rect 383514 133174 384134 168618
rect 383514 132938 383546 133174
rect 383782 132938 383866 133174
rect 384102 132938 384134 133174
rect 383514 132854 384134 132938
rect 383514 132618 383546 132854
rect 383782 132618 383866 132854
rect 384102 132618 384134 132854
rect 383514 97174 384134 132618
rect 383514 96938 383546 97174
rect 383782 96938 383866 97174
rect 384102 96938 384134 97174
rect 383514 96854 384134 96938
rect 383514 96618 383546 96854
rect 383782 96618 383866 96854
rect 384102 96618 384134 96854
rect 383514 61174 384134 96618
rect 383514 60938 383546 61174
rect 383782 60938 383866 61174
rect 384102 60938 384134 61174
rect 383514 60854 384134 60938
rect 383514 60618 383546 60854
rect 383782 60618 383866 60854
rect 384102 60618 384134 60854
rect 383514 25174 384134 60618
rect 383514 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 384134 25174
rect 383514 24854 384134 24938
rect 383514 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 384134 24854
rect 383514 -3226 384134 24618
rect 383514 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 384134 -3226
rect 383514 -3546 384134 -3462
rect 383514 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 384134 -3546
rect 383514 -3814 384134 -3782
rect 387234 676894 387854 709082
rect 387234 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 387854 676894
rect 387234 676574 387854 676658
rect 387234 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 387854 676574
rect 387234 640894 387854 676338
rect 387234 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 387854 640894
rect 387234 640574 387854 640658
rect 387234 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 387854 640574
rect 387234 604894 387854 640338
rect 387234 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 387854 604894
rect 387234 604574 387854 604658
rect 387234 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 387854 604574
rect 387234 568894 387854 604338
rect 387234 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 387854 568894
rect 387234 568574 387854 568658
rect 387234 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 387854 568574
rect 387234 532894 387854 568338
rect 387234 532658 387266 532894
rect 387502 532658 387586 532894
rect 387822 532658 387854 532894
rect 387234 532574 387854 532658
rect 387234 532338 387266 532574
rect 387502 532338 387586 532574
rect 387822 532338 387854 532574
rect 387234 496894 387854 532338
rect 387234 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 387854 496894
rect 387234 496574 387854 496658
rect 387234 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 387854 496574
rect 387234 460894 387854 496338
rect 387234 460658 387266 460894
rect 387502 460658 387586 460894
rect 387822 460658 387854 460894
rect 387234 460574 387854 460658
rect 387234 460338 387266 460574
rect 387502 460338 387586 460574
rect 387822 460338 387854 460574
rect 387234 424894 387854 460338
rect 387234 424658 387266 424894
rect 387502 424658 387586 424894
rect 387822 424658 387854 424894
rect 387234 424574 387854 424658
rect 387234 424338 387266 424574
rect 387502 424338 387586 424574
rect 387822 424338 387854 424574
rect 387234 388894 387854 424338
rect 387234 388658 387266 388894
rect 387502 388658 387586 388894
rect 387822 388658 387854 388894
rect 387234 388574 387854 388658
rect 387234 388338 387266 388574
rect 387502 388338 387586 388574
rect 387822 388338 387854 388574
rect 387234 352894 387854 388338
rect 387234 352658 387266 352894
rect 387502 352658 387586 352894
rect 387822 352658 387854 352894
rect 387234 352574 387854 352658
rect 387234 352338 387266 352574
rect 387502 352338 387586 352574
rect 387822 352338 387854 352574
rect 387234 316894 387854 352338
rect 387234 316658 387266 316894
rect 387502 316658 387586 316894
rect 387822 316658 387854 316894
rect 387234 316574 387854 316658
rect 387234 316338 387266 316574
rect 387502 316338 387586 316574
rect 387822 316338 387854 316574
rect 387234 280894 387854 316338
rect 387234 280658 387266 280894
rect 387502 280658 387586 280894
rect 387822 280658 387854 280894
rect 387234 280574 387854 280658
rect 387234 280338 387266 280574
rect 387502 280338 387586 280574
rect 387822 280338 387854 280574
rect 387234 244894 387854 280338
rect 387234 244658 387266 244894
rect 387502 244658 387586 244894
rect 387822 244658 387854 244894
rect 387234 244574 387854 244658
rect 387234 244338 387266 244574
rect 387502 244338 387586 244574
rect 387822 244338 387854 244574
rect 387234 208894 387854 244338
rect 387234 208658 387266 208894
rect 387502 208658 387586 208894
rect 387822 208658 387854 208894
rect 387234 208574 387854 208658
rect 387234 208338 387266 208574
rect 387502 208338 387586 208574
rect 387822 208338 387854 208574
rect 387234 172894 387854 208338
rect 387234 172658 387266 172894
rect 387502 172658 387586 172894
rect 387822 172658 387854 172894
rect 387234 172574 387854 172658
rect 387234 172338 387266 172574
rect 387502 172338 387586 172574
rect 387822 172338 387854 172574
rect 387234 136894 387854 172338
rect 387234 136658 387266 136894
rect 387502 136658 387586 136894
rect 387822 136658 387854 136894
rect 387234 136574 387854 136658
rect 387234 136338 387266 136574
rect 387502 136338 387586 136574
rect 387822 136338 387854 136574
rect 387234 100894 387854 136338
rect 387234 100658 387266 100894
rect 387502 100658 387586 100894
rect 387822 100658 387854 100894
rect 387234 100574 387854 100658
rect 387234 100338 387266 100574
rect 387502 100338 387586 100574
rect 387822 100338 387854 100574
rect 387234 64894 387854 100338
rect 387234 64658 387266 64894
rect 387502 64658 387586 64894
rect 387822 64658 387854 64894
rect 387234 64574 387854 64658
rect 387234 64338 387266 64574
rect 387502 64338 387586 64574
rect 387822 64338 387854 64574
rect 387234 28894 387854 64338
rect 387234 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 387854 28894
rect 387234 28574 387854 28658
rect 387234 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 387854 28574
rect 387234 -5146 387854 28338
rect 387234 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 387854 -5146
rect 387234 -5466 387854 -5382
rect 387234 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 387854 -5466
rect 387234 -5734 387854 -5702
rect 390954 680614 391574 711002
rect 408954 710598 409574 711590
rect 408954 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 409574 710598
rect 408954 710278 409574 710362
rect 408954 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 409574 710278
rect 405234 708678 405854 709670
rect 405234 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 405854 708678
rect 405234 708358 405854 708442
rect 405234 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 405854 708358
rect 401514 706758 402134 707750
rect 401514 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 402134 706758
rect 401514 706438 402134 706522
rect 401514 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 402134 706438
rect 390954 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 391574 680614
rect 390954 680294 391574 680378
rect 390954 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 391574 680294
rect 390954 644614 391574 680058
rect 390954 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 391574 644614
rect 390954 644294 391574 644378
rect 390954 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 391574 644294
rect 390954 608614 391574 644058
rect 390954 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 391574 608614
rect 390954 608294 391574 608378
rect 390954 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 391574 608294
rect 390954 572614 391574 608058
rect 390954 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 391574 572614
rect 390954 572294 391574 572378
rect 390954 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 391574 572294
rect 390954 536614 391574 572058
rect 390954 536378 390986 536614
rect 391222 536378 391306 536614
rect 391542 536378 391574 536614
rect 390954 536294 391574 536378
rect 390954 536058 390986 536294
rect 391222 536058 391306 536294
rect 391542 536058 391574 536294
rect 390954 500614 391574 536058
rect 390954 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 391574 500614
rect 390954 500294 391574 500378
rect 390954 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 391574 500294
rect 390954 464614 391574 500058
rect 390954 464378 390986 464614
rect 391222 464378 391306 464614
rect 391542 464378 391574 464614
rect 390954 464294 391574 464378
rect 390954 464058 390986 464294
rect 391222 464058 391306 464294
rect 391542 464058 391574 464294
rect 390954 428614 391574 464058
rect 390954 428378 390986 428614
rect 391222 428378 391306 428614
rect 391542 428378 391574 428614
rect 390954 428294 391574 428378
rect 390954 428058 390986 428294
rect 391222 428058 391306 428294
rect 391542 428058 391574 428294
rect 390954 392614 391574 428058
rect 390954 392378 390986 392614
rect 391222 392378 391306 392614
rect 391542 392378 391574 392614
rect 390954 392294 391574 392378
rect 390954 392058 390986 392294
rect 391222 392058 391306 392294
rect 391542 392058 391574 392294
rect 390954 356614 391574 392058
rect 390954 356378 390986 356614
rect 391222 356378 391306 356614
rect 391542 356378 391574 356614
rect 390954 356294 391574 356378
rect 390954 356058 390986 356294
rect 391222 356058 391306 356294
rect 391542 356058 391574 356294
rect 390954 320614 391574 356058
rect 390954 320378 390986 320614
rect 391222 320378 391306 320614
rect 391542 320378 391574 320614
rect 390954 320294 391574 320378
rect 390954 320058 390986 320294
rect 391222 320058 391306 320294
rect 391542 320058 391574 320294
rect 390954 284614 391574 320058
rect 390954 284378 390986 284614
rect 391222 284378 391306 284614
rect 391542 284378 391574 284614
rect 390954 284294 391574 284378
rect 390954 284058 390986 284294
rect 391222 284058 391306 284294
rect 391542 284058 391574 284294
rect 390954 248614 391574 284058
rect 390954 248378 390986 248614
rect 391222 248378 391306 248614
rect 391542 248378 391574 248614
rect 390954 248294 391574 248378
rect 390954 248058 390986 248294
rect 391222 248058 391306 248294
rect 391542 248058 391574 248294
rect 390954 212614 391574 248058
rect 390954 212378 390986 212614
rect 391222 212378 391306 212614
rect 391542 212378 391574 212614
rect 390954 212294 391574 212378
rect 390954 212058 390986 212294
rect 391222 212058 391306 212294
rect 391542 212058 391574 212294
rect 390954 176614 391574 212058
rect 390954 176378 390986 176614
rect 391222 176378 391306 176614
rect 391542 176378 391574 176614
rect 390954 176294 391574 176378
rect 390954 176058 390986 176294
rect 391222 176058 391306 176294
rect 391542 176058 391574 176294
rect 390954 140614 391574 176058
rect 390954 140378 390986 140614
rect 391222 140378 391306 140614
rect 391542 140378 391574 140614
rect 390954 140294 391574 140378
rect 390954 140058 390986 140294
rect 391222 140058 391306 140294
rect 391542 140058 391574 140294
rect 390954 104614 391574 140058
rect 390954 104378 390986 104614
rect 391222 104378 391306 104614
rect 391542 104378 391574 104614
rect 390954 104294 391574 104378
rect 390954 104058 390986 104294
rect 391222 104058 391306 104294
rect 391542 104058 391574 104294
rect 390954 68614 391574 104058
rect 390954 68378 390986 68614
rect 391222 68378 391306 68614
rect 391542 68378 391574 68614
rect 390954 68294 391574 68378
rect 390954 68058 390986 68294
rect 391222 68058 391306 68294
rect 391542 68058 391574 68294
rect 390954 32614 391574 68058
rect 390954 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 391574 32614
rect 390954 32294 391574 32378
rect 390954 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 391574 32294
rect 372954 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 373574 -6106
rect 372954 -6426 373574 -6342
rect 372954 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 373574 -6426
rect 372954 -7654 373574 -6662
rect 390954 -7066 391574 32058
rect 397794 704838 398414 705830
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 397794 363454 398414 398898
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 219454 398414 254898
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397794 147454 398414 182898
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -1894 398414 -902
rect 401514 691174 402134 706202
rect 401514 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 402134 691174
rect 401514 690854 402134 690938
rect 401514 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 402134 690854
rect 401514 655174 402134 690618
rect 401514 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 402134 655174
rect 401514 654854 402134 654938
rect 401514 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 402134 654854
rect 401514 619174 402134 654618
rect 401514 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 402134 619174
rect 401514 618854 402134 618938
rect 401514 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 402134 618854
rect 401514 583174 402134 618618
rect 401514 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 402134 583174
rect 401514 582854 402134 582938
rect 401514 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 402134 582854
rect 401514 547174 402134 582618
rect 401514 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 402134 547174
rect 401514 546854 402134 546938
rect 401514 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 402134 546854
rect 401514 511174 402134 546618
rect 401514 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 402134 511174
rect 401514 510854 402134 510938
rect 401514 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 402134 510854
rect 401514 475174 402134 510618
rect 401514 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 402134 475174
rect 401514 474854 402134 474938
rect 401514 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 402134 474854
rect 401514 439174 402134 474618
rect 401514 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 402134 439174
rect 401514 438854 402134 438938
rect 401514 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 402134 438854
rect 401514 403174 402134 438618
rect 401514 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 402134 403174
rect 401514 402854 402134 402938
rect 401514 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 402134 402854
rect 401514 367174 402134 402618
rect 401514 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 402134 367174
rect 401514 366854 402134 366938
rect 401514 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 402134 366854
rect 401514 331174 402134 366618
rect 401514 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 402134 331174
rect 401514 330854 402134 330938
rect 401514 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 402134 330854
rect 401514 295174 402134 330618
rect 401514 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 402134 295174
rect 401514 294854 402134 294938
rect 401514 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 402134 294854
rect 401514 259174 402134 294618
rect 401514 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 402134 259174
rect 401514 258854 402134 258938
rect 401514 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 402134 258854
rect 401514 223174 402134 258618
rect 401514 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 402134 223174
rect 401514 222854 402134 222938
rect 401514 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 402134 222854
rect 401514 187174 402134 222618
rect 401514 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 402134 187174
rect 401514 186854 402134 186938
rect 401514 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 402134 186854
rect 401514 151174 402134 186618
rect 401514 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 402134 151174
rect 401514 150854 402134 150938
rect 401514 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 402134 150854
rect 401514 115174 402134 150618
rect 401514 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 402134 115174
rect 401514 114854 402134 114938
rect 401514 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 402134 114854
rect 401514 79174 402134 114618
rect 401514 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 402134 79174
rect 401514 78854 402134 78938
rect 401514 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 402134 78854
rect 401514 43174 402134 78618
rect 401514 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 402134 43174
rect 401514 42854 402134 42938
rect 401514 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 402134 42854
rect 401514 7174 402134 42618
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 401514 -2266 402134 6618
rect 401514 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 402134 -2266
rect 401514 -2586 402134 -2502
rect 401514 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 402134 -2586
rect 401514 -3814 402134 -2822
rect 405234 694894 405854 708122
rect 405234 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 405854 694894
rect 405234 694574 405854 694658
rect 405234 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 405854 694574
rect 405234 658894 405854 694338
rect 405234 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 405854 658894
rect 405234 658574 405854 658658
rect 405234 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 405854 658574
rect 405234 622894 405854 658338
rect 405234 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 405854 622894
rect 405234 622574 405854 622658
rect 405234 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 405854 622574
rect 405234 586894 405854 622338
rect 405234 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 405854 586894
rect 405234 586574 405854 586658
rect 405234 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 405854 586574
rect 405234 550894 405854 586338
rect 405234 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 405854 550894
rect 405234 550574 405854 550658
rect 405234 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 405854 550574
rect 405234 514894 405854 550338
rect 405234 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 405854 514894
rect 405234 514574 405854 514658
rect 405234 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 405854 514574
rect 405234 478894 405854 514338
rect 405234 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 405854 478894
rect 405234 478574 405854 478658
rect 405234 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 405854 478574
rect 405234 442894 405854 478338
rect 405234 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 405854 442894
rect 405234 442574 405854 442658
rect 405234 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 405854 442574
rect 405234 406894 405854 442338
rect 405234 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 405854 406894
rect 405234 406574 405854 406658
rect 405234 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 405854 406574
rect 405234 370894 405854 406338
rect 405234 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 405854 370894
rect 405234 370574 405854 370658
rect 405234 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 405854 370574
rect 405234 334894 405854 370338
rect 405234 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 405854 334894
rect 405234 334574 405854 334658
rect 405234 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 405854 334574
rect 405234 298894 405854 334338
rect 405234 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 405854 298894
rect 405234 298574 405854 298658
rect 405234 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 405854 298574
rect 405234 262894 405854 298338
rect 405234 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 405854 262894
rect 405234 262574 405854 262658
rect 405234 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 405854 262574
rect 405234 226894 405854 262338
rect 405234 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 405854 226894
rect 405234 226574 405854 226658
rect 405234 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 405854 226574
rect 405234 190894 405854 226338
rect 405234 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 405854 190894
rect 405234 190574 405854 190658
rect 405234 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 405854 190574
rect 405234 154894 405854 190338
rect 405234 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 405854 154894
rect 405234 154574 405854 154658
rect 405234 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 405854 154574
rect 405234 118894 405854 154338
rect 405234 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 405854 118894
rect 405234 118574 405854 118658
rect 405234 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 405854 118574
rect 405234 82894 405854 118338
rect 405234 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 405854 82894
rect 405234 82574 405854 82658
rect 405234 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 405854 82574
rect 405234 46894 405854 82338
rect 405234 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 405854 46894
rect 405234 46574 405854 46658
rect 405234 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 405854 46574
rect 405234 10894 405854 46338
rect 405234 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 405854 10894
rect 405234 10574 405854 10658
rect 405234 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 405854 10574
rect 405234 -4186 405854 10338
rect 405234 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 405854 -4186
rect 405234 -4506 405854 -4422
rect 405234 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 405854 -4506
rect 405234 -5734 405854 -4742
rect 408954 698614 409574 710042
rect 426954 711558 427574 711590
rect 426954 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 427574 711558
rect 426954 711238 427574 711322
rect 426954 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 427574 711238
rect 423234 709638 423854 709670
rect 423234 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 423854 709638
rect 423234 709318 423854 709402
rect 423234 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 423854 709318
rect 419514 707718 420134 707750
rect 419514 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 420134 707718
rect 419514 707398 420134 707482
rect 419514 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 420134 707398
rect 408954 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 409574 698614
rect 408954 698294 409574 698378
rect 408954 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 409574 698294
rect 408954 662614 409574 698058
rect 408954 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 409574 662614
rect 408954 662294 409574 662378
rect 408954 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 409574 662294
rect 408954 626614 409574 662058
rect 408954 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 409574 626614
rect 408954 626294 409574 626378
rect 408954 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 409574 626294
rect 408954 590614 409574 626058
rect 408954 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 409574 590614
rect 408954 590294 409574 590378
rect 408954 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 409574 590294
rect 408954 554614 409574 590058
rect 408954 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 409574 554614
rect 408954 554294 409574 554378
rect 408954 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 409574 554294
rect 408954 518614 409574 554058
rect 408954 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 409574 518614
rect 408954 518294 409574 518378
rect 408954 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 409574 518294
rect 408954 482614 409574 518058
rect 408954 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 409574 482614
rect 408954 482294 409574 482378
rect 408954 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 409574 482294
rect 408954 446614 409574 482058
rect 408954 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 409574 446614
rect 408954 446294 409574 446378
rect 408954 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 409574 446294
rect 408954 410614 409574 446058
rect 408954 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 409574 410614
rect 408954 410294 409574 410378
rect 408954 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 409574 410294
rect 408954 374614 409574 410058
rect 408954 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 409574 374614
rect 408954 374294 409574 374378
rect 408954 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 409574 374294
rect 408954 338614 409574 374058
rect 408954 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 409574 338614
rect 408954 338294 409574 338378
rect 408954 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 409574 338294
rect 408954 302614 409574 338058
rect 408954 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 409574 302614
rect 408954 302294 409574 302378
rect 408954 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 409574 302294
rect 408954 266614 409574 302058
rect 408954 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 409574 266614
rect 408954 266294 409574 266378
rect 408954 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 409574 266294
rect 408954 230614 409574 266058
rect 408954 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 409574 230614
rect 408954 230294 409574 230378
rect 408954 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 409574 230294
rect 408954 194614 409574 230058
rect 408954 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 409574 194614
rect 408954 194294 409574 194378
rect 408954 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 409574 194294
rect 408954 158614 409574 194058
rect 408954 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 409574 158614
rect 408954 158294 409574 158378
rect 408954 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 409574 158294
rect 408954 122614 409574 158058
rect 408954 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 409574 122614
rect 408954 122294 409574 122378
rect 408954 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 409574 122294
rect 408954 86614 409574 122058
rect 408954 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 409574 86614
rect 408954 86294 409574 86378
rect 408954 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 409574 86294
rect 408954 50614 409574 86058
rect 408954 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 409574 50614
rect 408954 50294 409574 50378
rect 408954 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 409574 50294
rect 408954 14614 409574 50058
rect 408954 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 409574 14614
rect 408954 14294 409574 14378
rect 408954 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 409574 14294
rect 390954 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 391574 -7066
rect 390954 -7386 391574 -7302
rect 390954 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 391574 -7386
rect 390954 -7654 391574 -7622
rect 408954 -6106 409574 14058
rect 415794 705798 416414 705830
rect 415794 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 416414 705798
rect 415794 705478 416414 705562
rect 415794 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 416414 705478
rect 415794 669454 416414 705242
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 561454 416414 596898
rect 415794 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 416414 561454
rect 415794 561134 416414 561218
rect 415794 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 416414 561134
rect 415794 525454 416414 560898
rect 415794 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 416414 525454
rect 415794 525134 416414 525218
rect 415794 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 416414 525134
rect 415794 489454 416414 524898
rect 415794 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 416414 489454
rect 415794 489134 416414 489218
rect 415794 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 416414 489134
rect 415794 453454 416414 488898
rect 415794 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 416414 453454
rect 415794 453134 416414 453218
rect 415794 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 416414 453134
rect 415794 417454 416414 452898
rect 415794 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 416414 417454
rect 415794 417134 416414 417218
rect 415794 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 416414 417134
rect 415794 381454 416414 416898
rect 415794 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 416414 381454
rect 415794 381134 416414 381218
rect 415794 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 416414 381134
rect 415794 345454 416414 380898
rect 415794 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 416414 345454
rect 415794 345134 416414 345218
rect 415794 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 416414 345134
rect 415794 309454 416414 344898
rect 415794 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 416414 309454
rect 415794 309134 416414 309218
rect 415794 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 416414 309134
rect 415794 273454 416414 308898
rect 415794 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 416414 273454
rect 415794 273134 416414 273218
rect 415794 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 416414 273134
rect 415794 237454 416414 272898
rect 415794 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 416414 237454
rect 415794 237134 416414 237218
rect 415794 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 416414 237134
rect 415794 201454 416414 236898
rect 415794 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 416414 201454
rect 415794 201134 416414 201218
rect 415794 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 416414 201134
rect 415794 165454 416414 200898
rect 415794 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 416414 165454
rect 415794 165134 416414 165218
rect 415794 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 416414 165134
rect 415794 129454 416414 164898
rect 415794 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 416414 129454
rect 415794 129134 416414 129218
rect 415794 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 416414 129134
rect 415794 93454 416414 128898
rect 415794 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 416414 93454
rect 415794 93134 416414 93218
rect 415794 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 416414 93134
rect 415794 57454 416414 92898
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -1306 416414 20898
rect 415794 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 416414 -1306
rect 415794 -1626 416414 -1542
rect 415794 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 416414 -1626
rect 415794 -1894 416414 -1862
rect 419514 673174 420134 707162
rect 419514 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 420134 673174
rect 419514 672854 420134 672938
rect 419514 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 420134 672854
rect 419514 637174 420134 672618
rect 419514 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 420134 637174
rect 419514 636854 420134 636938
rect 419514 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 420134 636854
rect 419514 601174 420134 636618
rect 419514 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 420134 601174
rect 419514 600854 420134 600938
rect 419514 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 420134 600854
rect 419514 565174 420134 600618
rect 419514 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 420134 565174
rect 419514 564854 420134 564938
rect 419514 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 420134 564854
rect 419514 529174 420134 564618
rect 419514 528938 419546 529174
rect 419782 528938 419866 529174
rect 420102 528938 420134 529174
rect 419514 528854 420134 528938
rect 419514 528618 419546 528854
rect 419782 528618 419866 528854
rect 420102 528618 420134 528854
rect 419514 493174 420134 528618
rect 419514 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 420134 493174
rect 419514 492854 420134 492938
rect 419514 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 420134 492854
rect 419514 457174 420134 492618
rect 419514 456938 419546 457174
rect 419782 456938 419866 457174
rect 420102 456938 420134 457174
rect 419514 456854 420134 456938
rect 419514 456618 419546 456854
rect 419782 456618 419866 456854
rect 420102 456618 420134 456854
rect 419514 421174 420134 456618
rect 419514 420938 419546 421174
rect 419782 420938 419866 421174
rect 420102 420938 420134 421174
rect 419514 420854 420134 420938
rect 419514 420618 419546 420854
rect 419782 420618 419866 420854
rect 420102 420618 420134 420854
rect 419514 385174 420134 420618
rect 419514 384938 419546 385174
rect 419782 384938 419866 385174
rect 420102 384938 420134 385174
rect 419514 384854 420134 384938
rect 419514 384618 419546 384854
rect 419782 384618 419866 384854
rect 420102 384618 420134 384854
rect 419514 349174 420134 384618
rect 419514 348938 419546 349174
rect 419782 348938 419866 349174
rect 420102 348938 420134 349174
rect 419514 348854 420134 348938
rect 419514 348618 419546 348854
rect 419782 348618 419866 348854
rect 420102 348618 420134 348854
rect 419514 313174 420134 348618
rect 419514 312938 419546 313174
rect 419782 312938 419866 313174
rect 420102 312938 420134 313174
rect 419514 312854 420134 312938
rect 419514 312618 419546 312854
rect 419782 312618 419866 312854
rect 420102 312618 420134 312854
rect 419514 277174 420134 312618
rect 419514 276938 419546 277174
rect 419782 276938 419866 277174
rect 420102 276938 420134 277174
rect 419514 276854 420134 276938
rect 419514 276618 419546 276854
rect 419782 276618 419866 276854
rect 420102 276618 420134 276854
rect 419514 241174 420134 276618
rect 419514 240938 419546 241174
rect 419782 240938 419866 241174
rect 420102 240938 420134 241174
rect 419514 240854 420134 240938
rect 419514 240618 419546 240854
rect 419782 240618 419866 240854
rect 420102 240618 420134 240854
rect 419514 205174 420134 240618
rect 419514 204938 419546 205174
rect 419782 204938 419866 205174
rect 420102 204938 420134 205174
rect 419514 204854 420134 204938
rect 419514 204618 419546 204854
rect 419782 204618 419866 204854
rect 420102 204618 420134 204854
rect 419514 169174 420134 204618
rect 419514 168938 419546 169174
rect 419782 168938 419866 169174
rect 420102 168938 420134 169174
rect 419514 168854 420134 168938
rect 419514 168618 419546 168854
rect 419782 168618 419866 168854
rect 420102 168618 420134 168854
rect 419514 133174 420134 168618
rect 419514 132938 419546 133174
rect 419782 132938 419866 133174
rect 420102 132938 420134 133174
rect 419514 132854 420134 132938
rect 419514 132618 419546 132854
rect 419782 132618 419866 132854
rect 420102 132618 420134 132854
rect 419514 97174 420134 132618
rect 419514 96938 419546 97174
rect 419782 96938 419866 97174
rect 420102 96938 420134 97174
rect 419514 96854 420134 96938
rect 419514 96618 419546 96854
rect 419782 96618 419866 96854
rect 420102 96618 420134 96854
rect 419514 61174 420134 96618
rect 419514 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 420134 61174
rect 419514 60854 420134 60938
rect 419514 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 420134 60854
rect 419514 25174 420134 60618
rect 419514 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 420134 25174
rect 419514 24854 420134 24938
rect 419514 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 420134 24854
rect 419514 -3226 420134 24618
rect 419514 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 420134 -3226
rect 419514 -3546 420134 -3462
rect 419514 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 420134 -3546
rect 419514 -3814 420134 -3782
rect 423234 676894 423854 709082
rect 423234 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 423854 676894
rect 423234 676574 423854 676658
rect 423234 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 423854 676574
rect 423234 640894 423854 676338
rect 423234 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 423854 640894
rect 423234 640574 423854 640658
rect 423234 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 423854 640574
rect 423234 604894 423854 640338
rect 423234 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 423854 604894
rect 423234 604574 423854 604658
rect 423234 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 423854 604574
rect 423234 568894 423854 604338
rect 423234 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 423854 568894
rect 423234 568574 423854 568658
rect 423234 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 423854 568574
rect 423234 532894 423854 568338
rect 423234 532658 423266 532894
rect 423502 532658 423586 532894
rect 423822 532658 423854 532894
rect 423234 532574 423854 532658
rect 423234 532338 423266 532574
rect 423502 532338 423586 532574
rect 423822 532338 423854 532574
rect 423234 496894 423854 532338
rect 423234 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 423854 496894
rect 423234 496574 423854 496658
rect 423234 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 423854 496574
rect 423234 460894 423854 496338
rect 423234 460658 423266 460894
rect 423502 460658 423586 460894
rect 423822 460658 423854 460894
rect 423234 460574 423854 460658
rect 423234 460338 423266 460574
rect 423502 460338 423586 460574
rect 423822 460338 423854 460574
rect 423234 424894 423854 460338
rect 423234 424658 423266 424894
rect 423502 424658 423586 424894
rect 423822 424658 423854 424894
rect 423234 424574 423854 424658
rect 423234 424338 423266 424574
rect 423502 424338 423586 424574
rect 423822 424338 423854 424574
rect 423234 388894 423854 424338
rect 423234 388658 423266 388894
rect 423502 388658 423586 388894
rect 423822 388658 423854 388894
rect 423234 388574 423854 388658
rect 423234 388338 423266 388574
rect 423502 388338 423586 388574
rect 423822 388338 423854 388574
rect 423234 352894 423854 388338
rect 423234 352658 423266 352894
rect 423502 352658 423586 352894
rect 423822 352658 423854 352894
rect 423234 352574 423854 352658
rect 423234 352338 423266 352574
rect 423502 352338 423586 352574
rect 423822 352338 423854 352574
rect 423234 316894 423854 352338
rect 423234 316658 423266 316894
rect 423502 316658 423586 316894
rect 423822 316658 423854 316894
rect 423234 316574 423854 316658
rect 423234 316338 423266 316574
rect 423502 316338 423586 316574
rect 423822 316338 423854 316574
rect 423234 280894 423854 316338
rect 423234 280658 423266 280894
rect 423502 280658 423586 280894
rect 423822 280658 423854 280894
rect 423234 280574 423854 280658
rect 423234 280338 423266 280574
rect 423502 280338 423586 280574
rect 423822 280338 423854 280574
rect 423234 244894 423854 280338
rect 423234 244658 423266 244894
rect 423502 244658 423586 244894
rect 423822 244658 423854 244894
rect 423234 244574 423854 244658
rect 423234 244338 423266 244574
rect 423502 244338 423586 244574
rect 423822 244338 423854 244574
rect 423234 208894 423854 244338
rect 423234 208658 423266 208894
rect 423502 208658 423586 208894
rect 423822 208658 423854 208894
rect 423234 208574 423854 208658
rect 423234 208338 423266 208574
rect 423502 208338 423586 208574
rect 423822 208338 423854 208574
rect 423234 172894 423854 208338
rect 423234 172658 423266 172894
rect 423502 172658 423586 172894
rect 423822 172658 423854 172894
rect 423234 172574 423854 172658
rect 423234 172338 423266 172574
rect 423502 172338 423586 172574
rect 423822 172338 423854 172574
rect 423234 136894 423854 172338
rect 423234 136658 423266 136894
rect 423502 136658 423586 136894
rect 423822 136658 423854 136894
rect 423234 136574 423854 136658
rect 423234 136338 423266 136574
rect 423502 136338 423586 136574
rect 423822 136338 423854 136574
rect 423234 100894 423854 136338
rect 423234 100658 423266 100894
rect 423502 100658 423586 100894
rect 423822 100658 423854 100894
rect 423234 100574 423854 100658
rect 423234 100338 423266 100574
rect 423502 100338 423586 100574
rect 423822 100338 423854 100574
rect 423234 64894 423854 100338
rect 423234 64658 423266 64894
rect 423502 64658 423586 64894
rect 423822 64658 423854 64894
rect 423234 64574 423854 64658
rect 423234 64338 423266 64574
rect 423502 64338 423586 64574
rect 423822 64338 423854 64574
rect 423234 28894 423854 64338
rect 423234 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 423854 28894
rect 423234 28574 423854 28658
rect 423234 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 423854 28574
rect 423234 -5146 423854 28338
rect 423234 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 423854 -5146
rect 423234 -5466 423854 -5382
rect 423234 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 423854 -5466
rect 423234 -5734 423854 -5702
rect 426954 680614 427574 711002
rect 444954 710598 445574 711590
rect 444954 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 445574 710598
rect 444954 710278 445574 710362
rect 444954 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 445574 710278
rect 441234 708678 441854 709670
rect 441234 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 441854 708678
rect 441234 708358 441854 708442
rect 441234 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 441854 708358
rect 437514 706758 438134 707750
rect 437514 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 438134 706758
rect 437514 706438 438134 706522
rect 437514 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 438134 706438
rect 426954 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 427574 680614
rect 426954 680294 427574 680378
rect 426954 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 427574 680294
rect 426954 644614 427574 680058
rect 426954 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 427574 644614
rect 426954 644294 427574 644378
rect 426954 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 427574 644294
rect 426954 608614 427574 644058
rect 426954 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 427574 608614
rect 426954 608294 427574 608378
rect 426954 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 427574 608294
rect 426954 572614 427574 608058
rect 426954 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 427574 572614
rect 426954 572294 427574 572378
rect 426954 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 427574 572294
rect 426954 536614 427574 572058
rect 426954 536378 426986 536614
rect 427222 536378 427306 536614
rect 427542 536378 427574 536614
rect 426954 536294 427574 536378
rect 426954 536058 426986 536294
rect 427222 536058 427306 536294
rect 427542 536058 427574 536294
rect 426954 500614 427574 536058
rect 426954 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 427574 500614
rect 426954 500294 427574 500378
rect 426954 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 427574 500294
rect 426954 464614 427574 500058
rect 426954 464378 426986 464614
rect 427222 464378 427306 464614
rect 427542 464378 427574 464614
rect 426954 464294 427574 464378
rect 426954 464058 426986 464294
rect 427222 464058 427306 464294
rect 427542 464058 427574 464294
rect 426954 428614 427574 464058
rect 426954 428378 426986 428614
rect 427222 428378 427306 428614
rect 427542 428378 427574 428614
rect 426954 428294 427574 428378
rect 426954 428058 426986 428294
rect 427222 428058 427306 428294
rect 427542 428058 427574 428294
rect 426954 392614 427574 428058
rect 426954 392378 426986 392614
rect 427222 392378 427306 392614
rect 427542 392378 427574 392614
rect 426954 392294 427574 392378
rect 426954 392058 426986 392294
rect 427222 392058 427306 392294
rect 427542 392058 427574 392294
rect 426954 356614 427574 392058
rect 433794 704838 434414 705830
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 435454 434414 470898
rect 433794 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 434414 435454
rect 433794 435134 434414 435218
rect 433794 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 434414 435134
rect 433794 399454 434414 434898
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 372000 434414 398898
rect 437514 691174 438134 706202
rect 437514 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 438134 691174
rect 437514 690854 438134 690938
rect 437514 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 438134 690854
rect 437514 655174 438134 690618
rect 437514 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 438134 655174
rect 437514 654854 438134 654938
rect 437514 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 438134 654854
rect 437514 619174 438134 654618
rect 437514 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 438134 619174
rect 437514 618854 438134 618938
rect 437514 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 438134 618854
rect 437514 583174 438134 618618
rect 437514 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 438134 583174
rect 437514 582854 438134 582938
rect 437514 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 438134 582854
rect 437514 547174 438134 582618
rect 437514 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 438134 547174
rect 437514 546854 438134 546938
rect 437514 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 438134 546854
rect 437514 511174 438134 546618
rect 437514 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 438134 511174
rect 437514 510854 438134 510938
rect 437514 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 438134 510854
rect 437514 475174 438134 510618
rect 437514 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 438134 475174
rect 437514 474854 438134 474938
rect 437514 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 438134 474854
rect 437514 439174 438134 474618
rect 437514 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 438134 439174
rect 437514 438854 438134 438938
rect 437514 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 438134 438854
rect 437514 403174 438134 438618
rect 437514 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 438134 403174
rect 437514 402854 438134 402938
rect 437514 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 438134 402854
rect 437514 372000 438134 402618
rect 441234 694894 441854 708122
rect 441234 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 441854 694894
rect 441234 694574 441854 694658
rect 441234 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 441854 694574
rect 441234 658894 441854 694338
rect 441234 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 441854 658894
rect 441234 658574 441854 658658
rect 441234 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 441854 658574
rect 441234 622894 441854 658338
rect 441234 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 441854 622894
rect 441234 622574 441854 622658
rect 441234 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 441854 622574
rect 441234 586894 441854 622338
rect 441234 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 441854 586894
rect 441234 586574 441854 586658
rect 441234 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 441854 586574
rect 441234 550894 441854 586338
rect 441234 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 441854 550894
rect 441234 550574 441854 550658
rect 441234 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 441854 550574
rect 441234 514894 441854 550338
rect 441234 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 441854 514894
rect 441234 514574 441854 514658
rect 441234 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 441854 514574
rect 441234 478894 441854 514338
rect 441234 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 441854 478894
rect 441234 478574 441854 478658
rect 441234 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 441854 478574
rect 441234 442894 441854 478338
rect 441234 442658 441266 442894
rect 441502 442658 441586 442894
rect 441822 442658 441854 442894
rect 441234 442574 441854 442658
rect 441234 442338 441266 442574
rect 441502 442338 441586 442574
rect 441822 442338 441854 442574
rect 441234 406894 441854 442338
rect 441234 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 441854 406894
rect 441234 406574 441854 406658
rect 441234 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 441854 406574
rect 441234 372000 441854 406338
rect 444954 698614 445574 710042
rect 462954 711558 463574 711590
rect 462954 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 463574 711558
rect 462954 711238 463574 711322
rect 462954 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 463574 711238
rect 459234 709638 459854 709670
rect 459234 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 459854 709638
rect 459234 709318 459854 709402
rect 459234 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 459854 709318
rect 455514 707718 456134 707750
rect 455514 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 456134 707718
rect 455514 707398 456134 707482
rect 455514 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 456134 707398
rect 444954 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 445574 698614
rect 444954 698294 445574 698378
rect 444954 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 445574 698294
rect 444954 662614 445574 698058
rect 444954 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 445574 662614
rect 444954 662294 445574 662378
rect 444954 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 445574 662294
rect 444954 626614 445574 662058
rect 444954 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 445574 626614
rect 444954 626294 445574 626378
rect 444954 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 445574 626294
rect 444954 590614 445574 626058
rect 444954 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 445574 590614
rect 444954 590294 445574 590378
rect 444954 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 445574 590294
rect 444954 554614 445574 590058
rect 444954 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 445574 554614
rect 444954 554294 445574 554378
rect 444954 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 445574 554294
rect 444954 518614 445574 554058
rect 444954 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 445574 518614
rect 444954 518294 445574 518378
rect 444954 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 445574 518294
rect 444954 482614 445574 518058
rect 444954 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 445574 482614
rect 444954 482294 445574 482378
rect 444954 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 445574 482294
rect 444954 446614 445574 482058
rect 444954 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 445574 446614
rect 444954 446294 445574 446378
rect 444954 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 445574 446294
rect 444954 410614 445574 446058
rect 444954 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 445574 410614
rect 444954 410294 445574 410378
rect 444954 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 445574 410294
rect 444954 374614 445574 410058
rect 444954 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 445574 374614
rect 444954 374294 445574 374378
rect 444954 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 445574 374294
rect 434243 363454 434563 363486
rect 434243 363218 434285 363454
rect 434521 363218 434563 363454
rect 434243 363134 434563 363218
rect 434243 362898 434285 363134
rect 434521 362898 434563 363134
rect 434243 362866 434563 362898
rect 436840 363454 437160 363486
rect 436840 363218 436882 363454
rect 437118 363218 437160 363454
rect 436840 363134 437160 363218
rect 436840 362898 436882 363134
rect 437118 362898 437160 363134
rect 436840 362866 437160 362898
rect 439437 363454 439757 363486
rect 439437 363218 439479 363454
rect 439715 363218 439757 363454
rect 439437 363134 439757 363218
rect 439437 362898 439479 363134
rect 439715 362898 439757 363134
rect 439437 362866 439757 362898
rect 426954 356378 426986 356614
rect 427222 356378 427306 356614
rect 427542 356378 427574 356614
rect 426954 356294 427574 356378
rect 426954 356058 426986 356294
rect 427222 356058 427306 356294
rect 427542 356058 427574 356294
rect 426954 320614 427574 356058
rect 435541 345454 435861 345486
rect 435541 345218 435583 345454
rect 435819 345218 435861 345454
rect 435541 345134 435861 345218
rect 435541 344898 435583 345134
rect 435819 344898 435861 345134
rect 435541 344866 435861 344898
rect 438138 345454 438458 345486
rect 438138 345218 438180 345454
rect 438416 345218 438458 345454
rect 438138 345134 438458 345218
rect 438138 344898 438180 345134
rect 438416 344898 438458 345134
rect 438138 344866 438458 344898
rect 444954 338614 445574 374058
rect 444954 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 445574 338614
rect 444954 338294 445574 338378
rect 444954 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 445574 338294
rect 426954 320378 426986 320614
rect 427222 320378 427306 320614
rect 427542 320378 427574 320614
rect 426954 320294 427574 320378
rect 426954 320058 426986 320294
rect 427222 320058 427306 320294
rect 427542 320058 427574 320294
rect 426954 284614 427574 320058
rect 433794 327454 434414 338000
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 300000 434414 326898
rect 437514 331174 438134 338000
rect 437514 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 438134 331174
rect 437514 330854 438134 330938
rect 437514 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 438134 330854
rect 437514 300000 438134 330618
rect 441234 334894 441854 338000
rect 441234 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 441854 334894
rect 441234 334574 441854 334658
rect 441234 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 441854 334574
rect 441234 300000 441854 334338
rect 444954 302614 445574 338058
rect 444954 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 445574 302614
rect 444954 302294 445574 302378
rect 444954 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 445574 302294
rect 434243 291454 434563 291486
rect 434243 291218 434285 291454
rect 434521 291218 434563 291454
rect 434243 291134 434563 291218
rect 434243 290898 434285 291134
rect 434521 290898 434563 291134
rect 434243 290866 434563 290898
rect 436840 291454 437160 291486
rect 436840 291218 436882 291454
rect 437118 291218 437160 291454
rect 436840 291134 437160 291218
rect 436840 290898 436882 291134
rect 437118 290898 437160 291134
rect 436840 290866 437160 290898
rect 439437 291454 439757 291486
rect 439437 291218 439479 291454
rect 439715 291218 439757 291454
rect 439437 291134 439757 291218
rect 439437 290898 439479 291134
rect 439715 290898 439757 291134
rect 439437 290866 439757 290898
rect 426954 284378 426986 284614
rect 427222 284378 427306 284614
rect 427542 284378 427574 284614
rect 426954 284294 427574 284378
rect 426954 284058 426986 284294
rect 427222 284058 427306 284294
rect 427542 284058 427574 284294
rect 426954 248614 427574 284058
rect 435541 273454 435861 273486
rect 435541 273218 435583 273454
rect 435819 273218 435861 273454
rect 435541 273134 435861 273218
rect 435541 272898 435583 273134
rect 435819 272898 435861 273134
rect 435541 272866 435861 272898
rect 438138 273454 438458 273486
rect 438138 273218 438180 273454
rect 438416 273218 438458 273454
rect 438138 273134 438458 273218
rect 438138 272898 438180 273134
rect 438416 272898 438458 273134
rect 438138 272866 438458 272898
rect 444954 266614 445574 302058
rect 444954 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 445574 266614
rect 444954 266294 445574 266378
rect 444954 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 445574 266294
rect 426954 248378 426986 248614
rect 427222 248378 427306 248614
rect 427542 248378 427574 248614
rect 426954 248294 427574 248378
rect 426954 248058 426986 248294
rect 427222 248058 427306 248294
rect 427542 248058 427574 248294
rect 426954 212614 427574 248058
rect 433794 255454 434414 266000
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 228000 434414 254898
rect 437514 259174 438134 266000
rect 437514 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 438134 259174
rect 437514 258854 438134 258938
rect 437514 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 438134 258854
rect 437514 228000 438134 258618
rect 441234 262894 441854 266000
rect 441234 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 441854 262894
rect 441234 262574 441854 262658
rect 441234 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 441854 262574
rect 441234 228000 441854 262338
rect 444954 230614 445574 266058
rect 444954 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 445574 230614
rect 444954 230294 445574 230378
rect 444954 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 445574 230294
rect 434243 219454 434563 219486
rect 434243 219218 434285 219454
rect 434521 219218 434563 219454
rect 434243 219134 434563 219218
rect 434243 218898 434285 219134
rect 434521 218898 434563 219134
rect 434243 218866 434563 218898
rect 436840 219454 437160 219486
rect 436840 219218 436882 219454
rect 437118 219218 437160 219454
rect 436840 219134 437160 219218
rect 436840 218898 436882 219134
rect 437118 218898 437160 219134
rect 436840 218866 437160 218898
rect 439437 219454 439757 219486
rect 439437 219218 439479 219454
rect 439715 219218 439757 219454
rect 439437 219134 439757 219218
rect 439437 218898 439479 219134
rect 439715 218898 439757 219134
rect 439437 218866 439757 218898
rect 426954 212378 426986 212614
rect 427222 212378 427306 212614
rect 427542 212378 427574 212614
rect 426954 212294 427574 212378
rect 426954 212058 426986 212294
rect 427222 212058 427306 212294
rect 427542 212058 427574 212294
rect 426954 176614 427574 212058
rect 435541 201454 435861 201486
rect 435541 201218 435583 201454
rect 435819 201218 435861 201454
rect 435541 201134 435861 201218
rect 435541 200898 435583 201134
rect 435819 200898 435861 201134
rect 435541 200866 435861 200898
rect 438138 201454 438458 201486
rect 438138 201218 438180 201454
rect 438416 201218 438458 201454
rect 438138 201134 438458 201218
rect 438138 200898 438180 201134
rect 438416 200898 438458 201134
rect 438138 200866 438458 200898
rect 444954 194614 445574 230058
rect 444954 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 445574 194614
rect 444954 194294 445574 194378
rect 444954 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 445574 194294
rect 426954 176378 426986 176614
rect 427222 176378 427306 176614
rect 427542 176378 427574 176614
rect 426954 176294 427574 176378
rect 426954 176058 426986 176294
rect 427222 176058 427306 176294
rect 427542 176058 427574 176294
rect 426954 140614 427574 176058
rect 433794 183454 434414 194000
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 433794 156000 434414 182898
rect 437514 187174 438134 194000
rect 437514 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 438134 187174
rect 437514 186854 438134 186938
rect 437514 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 438134 186854
rect 437514 156000 438134 186618
rect 441234 190894 441854 194000
rect 441234 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 441854 190894
rect 441234 190574 441854 190658
rect 441234 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 441854 190574
rect 441234 156000 441854 190338
rect 444954 158614 445574 194058
rect 444954 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 445574 158614
rect 444954 158294 445574 158378
rect 444954 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 445574 158294
rect 434243 147454 434563 147486
rect 434243 147218 434285 147454
rect 434521 147218 434563 147454
rect 434243 147134 434563 147218
rect 434243 146898 434285 147134
rect 434521 146898 434563 147134
rect 434243 146866 434563 146898
rect 436840 147454 437160 147486
rect 436840 147218 436882 147454
rect 437118 147218 437160 147454
rect 436840 147134 437160 147218
rect 436840 146898 436882 147134
rect 437118 146898 437160 147134
rect 436840 146866 437160 146898
rect 439437 147454 439757 147486
rect 439437 147218 439479 147454
rect 439715 147218 439757 147454
rect 439437 147134 439757 147218
rect 439437 146898 439479 147134
rect 439715 146898 439757 147134
rect 439437 146866 439757 146898
rect 426954 140378 426986 140614
rect 427222 140378 427306 140614
rect 427542 140378 427574 140614
rect 426954 140294 427574 140378
rect 426954 140058 426986 140294
rect 427222 140058 427306 140294
rect 427542 140058 427574 140294
rect 426954 104614 427574 140058
rect 435541 129454 435861 129486
rect 435541 129218 435583 129454
rect 435819 129218 435861 129454
rect 435541 129134 435861 129218
rect 435541 128898 435583 129134
rect 435819 128898 435861 129134
rect 435541 128866 435861 128898
rect 438138 129454 438458 129486
rect 438138 129218 438180 129454
rect 438416 129218 438458 129454
rect 438138 129134 438458 129218
rect 438138 128898 438180 129134
rect 438416 128898 438458 129134
rect 438138 128866 438458 128898
rect 444954 122614 445574 158058
rect 444954 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 445574 122614
rect 444954 122294 445574 122378
rect 444954 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 445574 122294
rect 426954 104378 426986 104614
rect 427222 104378 427306 104614
rect 427542 104378 427574 104614
rect 426954 104294 427574 104378
rect 426954 104058 426986 104294
rect 427222 104058 427306 104294
rect 427542 104058 427574 104294
rect 426954 68614 427574 104058
rect 426954 68378 426986 68614
rect 427222 68378 427306 68614
rect 427542 68378 427574 68614
rect 426954 68294 427574 68378
rect 426954 68058 426986 68294
rect 427222 68058 427306 68294
rect 427542 68058 427574 68294
rect 426954 32614 427574 68058
rect 426954 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 427574 32614
rect 426954 32294 427574 32378
rect 426954 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 427574 32294
rect 408954 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 409574 -6106
rect 408954 -6426 409574 -6342
rect 408954 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 409574 -6426
rect 408954 -7654 409574 -6662
rect 426954 -7066 427574 32058
rect 433794 111454 434414 122000
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -1894 434414 -902
rect 437514 115174 438134 122000
rect 437514 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 438134 115174
rect 437514 114854 438134 114938
rect 437514 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 438134 114854
rect 437514 79174 438134 114618
rect 437514 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 438134 79174
rect 437514 78854 438134 78938
rect 437514 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 438134 78854
rect 437514 43174 438134 78618
rect 437514 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 438134 43174
rect 437514 42854 438134 42938
rect 437514 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 438134 42854
rect 437514 7174 438134 42618
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -2266 438134 6618
rect 437514 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 438134 -2266
rect 437514 -2586 438134 -2502
rect 437514 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 438134 -2586
rect 437514 -3814 438134 -2822
rect 441234 118894 441854 122000
rect 441234 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 441854 118894
rect 441234 118574 441854 118658
rect 441234 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 441854 118574
rect 441234 82894 441854 118338
rect 441234 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 441854 82894
rect 441234 82574 441854 82658
rect 441234 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 441854 82574
rect 441234 46894 441854 82338
rect 441234 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 441854 46894
rect 441234 46574 441854 46658
rect 441234 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 441854 46574
rect 441234 10894 441854 46338
rect 441234 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 441854 10894
rect 441234 10574 441854 10658
rect 441234 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 441854 10574
rect 441234 -4186 441854 10338
rect 441234 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 441854 -4186
rect 441234 -4506 441854 -4422
rect 441234 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 441854 -4506
rect 441234 -5734 441854 -4742
rect 444954 86614 445574 122058
rect 444954 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 445574 86614
rect 444954 86294 445574 86378
rect 444954 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 445574 86294
rect 444954 50614 445574 86058
rect 444954 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 445574 50614
rect 444954 50294 445574 50378
rect 444954 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 445574 50294
rect 444954 14614 445574 50058
rect 444954 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 445574 14614
rect 444954 14294 445574 14378
rect 444954 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 445574 14294
rect 426954 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 427574 -7066
rect 426954 -7386 427574 -7302
rect 426954 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 427574 -7386
rect 426954 -7654 427574 -7622
rect 444954 -6106 445574 14058
rect 451794 705798 452414 705830
rect 451794 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 452414 705798
rect 451794 705478 452414 705562
rect 451794 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 452414 705478
rect 451794 669454 452414 705242
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 453454 452414 488898
rect 451794 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 452414 453454
rect 451794 453134 452414 453218
rect 451794 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 452414 453134
rect 451794 417454 452414 452898
rect 451794 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 452414 417454
rect 451794 417134 452414 417218
rect 451794 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 452414 417134
rect 451794 381454 452414 416898
rect 451794 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 452414 381454
rect 451794 381134 452414 381218
rect 451794 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 452414 381134
rect 451794 345454 452414 380898
rect 451794 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 452414 345454
rect 451794 345134 452414 345218
rect 451794 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 452414 345134
rect 451794 309454 452414 344898
rect 451794 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 452414 309454
rect 451794 309134 452414 309218
rect 451794 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 452414 309134
rect 451794 273454 452414 308898
rect 451794 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 452414 273454
rect 451794 273134 452414 273218
rect 451794 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 452414 273134
rect 451794 237454 452414 272898
rect 451794 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 452414 237454
rect 451794 237134 452414 237218
rect 451794 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 452414 237134
rect 451794 201454 452414 236898
rect 451794 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 452414 201454
rect 451794 201134 452414 201218
rect 451794 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 452414 201134
rect 451794 165454 452414 200898
rect 451794 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 452414 165454
rect 451794 165134 452414 165218
rect 451794 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 452414 165134
rect 451794 129454 452414 164898
rect 451794 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 452414 129454
rect 451794 129134 452414 129218
rect 451794 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 452414 129134
rect 451794 93454 452414 128898
rect 451794 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 452414 93454
rect 451794 93134 452414 93218
rect 451794 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 452414 93134
rect 451794 57454 452414 92898
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -1306 452414 20898
rect 451794 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 452414 -1306
rect 451794 -1626 452414 -1542
rect 451794 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 452414 -1626
rect 451794 -1894 452414 -1862
rect 455514 673174 456134 707162
rect 455514 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 456134 673174
rect 455514 672854 456134 672938
rect 455514 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 456134 672854
rect 455514 637174 456134 672618
rect 455514 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 456134 637174
rect 455514 636854 456134 636938
rect 455514 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 456134 636854
rect 455514 601174 456134 636618
rect 455514 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 456134 601174
rect 455514 600854 456134 600938
rect 455514 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 456134 600854
rect 455514 565174 456134 600618
rect 455514 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 456134 565174
rect 455514 564854 456134 564938
rect 455514 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 456134 564854
rect 455514 529174 456134 564618
rect 455514 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 456134 529174
rect 455514 528854 456134 528938
rect 455514 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 456134 528854
rect 455514 493174 456134 528618
rect 455514 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 456134 493174
rect 455514 492854 456134 492938
rect 455514 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 456134 492854
rect 455514 457174 456134 492618
rect 455514 456938 455546 457174
rect 455782 456938 455866 457174
rect 456102 456938 456134 457174
rect 455514 456854 456134 456938
rect 455514 456618 455546 456854
rect 455782 456618 455866 456854
rect 456102 456618 456134 456854
rect 455514 421174 456134 456618
rect 455514 420938 455546 421174
rect 455782 420938 455866 421174
rect 456102 420938 456134 421174
rect 455514 420854 456134 420938
rect 455514 420618 455546 420854
rect 455782 420618 455866 420854
rect 456102 420618 456134 420854
rect 455514 385174 456134 420618
rect 455514 384938 455546 385174
rect 455782 384938 455866 385174
rect 456102 384938 456134 385174
rect 455514 384854 456134 384938
rect 455514 384618 455546 384854
rect 455782 384618 455866 384854
rect 456102 384618 456134 384854
rect 455514 349174 456134 384618
rect 455514 348938 455546 349174
rect 455782 348938 455866 349174
rect 456102 348938 456134 349174
rect 455514 348854 456134 348938
rect 455514 348618 455546 348854
rect 455782 348618 455866 348854
rect 456102 348618 456134 348854
rect 455514 313174 456134 348618
rect 455514 312938 455546 313174
rect 455782 312938 455866 313174
rect 456102 312938 456134 313174
rect 455514 312854 456134 312938
rect 455514 312618 455546 312854
rect 455782 312618 455866 312854
rect 456102 312618 456134 312854
rect 455514 277174 456134 312618
rect 455514 276938 455546 277174
rect 455782 276938 455866 277174
rect 456102 276938 456134 277174
rect 455514 276854 456134 276938
rect 455514 276618 455546 276854
rect 455782 276618 455866 276854
rect 456102 276618 456134 276854
rect 455514 241174 456134 276618
rect 455514 240938 455546 241174
rect 455782 240938 455866 241174
rect 456102 240938 456134 241174
rect 455514 240854 456134 240938
rect 455514 240618 455546 240854
rect 455782 240618 455866 240854
rect 456102 240618 456134 240854
rect 455514 205174 456134 240618
rect 455514 204938 455546 205174
rect 455782 204938 455866 205174
rect 456102 204938 456134 205174
rect 455514 204854 456134 204938
rect 455514 204618 455546 204854
rect 455782 204618 455866 204854
rect 456102 204618 456134 204854
rect 455514 169174 456134 204618
rect 455514 168938 455546 169174
rect 455782 168938 455866 169174
rect 456102 168938 456134 169174
rect 455514 168854 456134 168938
rect 455514 168618 455546 168854
rect 455782 168618 455866 168854
rect 456102 168618 456134 168854
rect 455514 133174 456134 168618
rect 455514 132938 455546 133174
rect 455782 132938 455866 133174
rect 456102 132938 456134 133174
rect 455514 132854 456134 132938
rect 455514 132618 455546 132854
rect 455782 132618 455866 132854
rect 456102 132618 456134 132854
rect 455514 97174 456134 132618
rect 455514 96938 455546 97174
rect 455782 96938 455866 97174
rect 456102 96938 456134 97174
rect 455514 96854 456134 96938
rect 455514 96618 455546 96854
rect 455782 96618 455866 96854
rect 456102 96618 456134 96854
rect 455514 61174 456134 96618
rect 455514 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 456134 61174
rect 455514 60854 456134 60938
rect 455514 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 456134 60854
rect 455514 25174 456134 60618
rect 455514 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 456134 25174
rect 455514 24854 456134 24938
rect 455514 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 456134 24854
rect 455514 -3226 456134 24618
rect 455514 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 456134 -3226
rect 455514 -3546 456134 -3462
rect 455514 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 456134 -3546
rect 455514 -3814 456134 -3782
rect 459234 676894 459854 709082
rect 459234 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 459854 676894
rect 459234 676574 459854 676658
rect 459234 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 459854 676574
rect 459234 640894 459854 676338
rect 459234 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 459854 640894
rect 459234 640574 459854 640658
rect 459234 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 459854 640574
rect 459234 604894 459854 640338
rect 459234 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 459854 604894
rect 459234 604574 459854 604658
rect 459234 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 459854 604574
rect 459234 568894 459854 604338
rect 459234 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 459854 568894
rect 459234 568574 459854 568658
rect 459234 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 459854 568574
rect 459234 532894 459854 568338
rect 459234 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 459854 532894
rect 459234 532574 459854 532658
rect 459234 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 459854 532574
rect 459234 496894 459854 532338
rect 459234 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 459854 496894
rect 459234 496574 459854 496658
rect 459234 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 459854 496574
rect 459234 460894 459854 496338
rect 459234 460658 459266 460894
rect 459502 460658 459586 460894
rect 459822 460658 459854 460894
rect 459234 460574 459854 460658
rect 459234 460338 459266 460574
rect 459502 460338 459586 460574
rect 459822 460338 459854 460574
rect 459234 424894 459854 460338
rect 459234 424658 459266 424894
rect 459502 424658 459586 424894
rect 459822 424658 459854 424894
rect 459234 424574 459854 424658
rect 459234 424338 459266 424574
rect 459502 424338 459586 424574
rect 459822 424338 459854 424574
rect 459234 388894 459854 424338
rect 459234 388658 459266 388894
rect 459502 388658 459586 388894
rect 459822 388658 459854 388894
rect 459234 388574 459854 388658
rect 459234 388338 459266 388574
rect 459502 388338 459586 388574
rect 459822 388338 459854 388574
rect 459234 352894 459854 388338
rect 459234 352658 459266 352894
rect 459502 352658 459586 352894
rect 459822 352658 459854 352894
rect 459234 352574 459854 352658
rect 459234 352338 459266 352574
rect 459502 352338 459586 352574
rect 459822 352338 459854 352574
rect 459234 316894 459854 352338
rect 459234 316658 459266 316894
rect 459502 316658 459586 316894
rect 459822 316658 459854 316894
rect 459234 316574 459854 316658
rect 459234 316338 459266 316574
rect 459502 316338 459586 316574
rect 459822 316338 459854 316574
rect 459234 280894 459854 316338
rect 459234 280658 459266 280894
rect 459502 280658 459586 280894
rect 459822 280658 459854 280894
rect 459234 280574 459854 280658
rect 459234 280338 459266 280574
rect 459502 280338 459586 280574
rect 459822 280338 459854 280574
rect 459234 244894 459854 280338
rect 459234 244658 459266 244894
rect 459502 244658 459586 244894
rect 459822 244658 459854 244894
rect 459234 244574 459854 244658
rect 459234 244338 459266 244574
rect 459502 244338 459586 244574
rect 459822 244338 459854 244574
rect 459234 208894 459854 244338
rect 459234 208658 459266 208894
rect 459502 208658 459586 208894
rect 459822 208658 459854 208894
rect 459234 208574 459854 208658
rect 459234 208338 459266 208574
rect 459502 208338 459586 208574
rect 459822 208338 459854 208574
rect 459234 172894 459854 208338
rect 459234 172658 459266 172894
rect 459502 172658 459586 172894
rect 459822 172658 459854 172894
rect 459234 172574 459854 172658
rect 459234 172338 459266 172574
rect 459502 172338 459586 172574
rect 459822 172338 459854 172574
rect 459234 136894 459854 172338
rect 459234 136658 459266 136894
rect 459502 136658 459586 136894
rect 459822 136658 459854 136894
rect 459234 136574 459854 136658
rect 459234 136338 459266 136574
rect 459502 136338 459586 136574
rect 459822 136338 459854 136574
rect 459234 100894 459854 136338
rect 459234 100658 459266 100894
rect 459502 100658 459586 100894
rect 459822 100658 459854 100894
rect 459234 100574 459854 100658
rect 459234 100338 459266 100574
rect 459502 100338 459586 100574
rect 459822 100338 459854 100574
rect 459234 64894 459854 100338
rect 459234 64658 459266 64894
rect 459502 64658 459586 64894
rect 459822 64658 459854 64894
rect 459234 64574 459854 64658
rect 459234 64338 459266 64574
rect 459502 64338 459586 64574
rect 459822 64338 459854 64574
rect 459234 28894 459854 64338
rect 459234 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 459854 28894
rect 459234 28574 459854 28658
rect 459234 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 459854 28574
rect 459234 -5146 459854 28338
rect 459234 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 459854 -5146
rect 459234 -5466 459854 -5382
rect 459234 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 459854 -5466
rect 459234 -5734 459854 -5702
rect 462954 680614 463574 711002
rect 480954 710598 481574 711590
rect 480954 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 481574 710598
rect 480954 710278 481574 710362
rect 480954 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 481574 710278
rect 477234 708678 477854 709670
rect 477234 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 477854 708678
rect 477234 708358 477854 708442
rect 477234 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 477854 708358
rect 473514 706758 474134 707750
rect 473514 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 474134 706758
rect 473514 706438 474134 706522
rect 473514 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 474134 706438
rect 462954 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 463574 680614
rect 462954 680294 463574 680378
rect 462954 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 463574 680294
rect 462954 644614 463574 680058
rect 462954 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 463574 644614
rect 462954 644294 463574 644378
rect 462954 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 463574 644294
rect 462954 608614 463574 644058
rect 462954 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 463574 608614
rect 462954 608294 463574 608378
rect 462954 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 463574 608294
rect 462954 572614 463574 608058
rect 462954 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 463574 572614
rect 462954 572294 463574 572378
rect 462954 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 463574 572294
rect 462954 536614 463574 572058
rect 462954 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 463574 536614
rect 462954 536294 463574 536378
rect 462954 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 463574 536294
rect 462954 500614 463574 536058
rect 462954 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 463574 500614
rect 462954 500294 463574 500378
rect 462954 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 463574 500294
rect 462954 464614 463574 500058
rect 462954 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 463574 464614
rect 462954 464294 463574 464378
rect 462954 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 463574 464294
rect 462954 428614 463574 464058
rect 462954 428378 462986 428614
rect 463222 428378 463306 428614
rect 463542 428378 463574 428614
rect 462954 428294 463574 428378
rect 462954 428058 462986 428294
rect 463222 428058 463306 428294
rect 463542 428058 463574 428294
rect 462954 392614 463574 428058
rect 462954 392378 462986 392614
rect 463222 392378 463306 392614
rect 463542 392378 463574 392614
rect 462954 392294 463574 392378
rect 462954 392058 462986 392294
rect 463222 392058 463306 392294
rect 463542 392058 463574 392294
rect 462954 356614 463574 392058
rect 462954 356378 462986 356614
rect 463222 356378 463306 356614
rect 463542 356378 463574 356614
rect 462954 356294 463574 356378
rect 462954 356058 462986 356294
rect 463222 356058 463306 356294
rect 463542 356058 463574 356294
rect 462954 320614 463574 356058
rect 462954 320378 462986 320614
rect 463222 320378 463306 320614
rect 463542 320378 463574 320614
rect 462954 320294 463574 320378
rect 462954 320058 462986 320294
rect 463222 320058 463306 320294
rect 463542 320058 463574 320294
rect 462954 284614 463574 320058
rect 462954 284378 462986 284614
rect 463222 284378 463306 284614
rect 463542 284378 463574 284614
rect 462954 284294 463574 284378
rect 462954 284058 462986 284294
rect 463222 284058 463306 284294
rect 463542 284058 463574 284294
rect 462954 248614 463574 284058
rect 462954 248378 462986 248614
rect 463222 248378 463306 248614
rect 463542 248378 463574 248614
rect 462954 248294 463574 248378
rect 462954 248058 462986 248294
rect 463222 248058 463306 248294
rect 463542 248058 463574 248294
rect 462954 212614 463574 248058
rect 462954 212378 462986 212614
rect 463222 212378 463306 212614
rect 463542 212378 463574 212614
rect 462954 212294 463574 212378
rect 462954 212058 462986 212294
rect 463222 212058 463306 212294
rect 463542 212058 463574 212294
rect 462954 176614 463574 212058
rect 462954 176378 462986 176614
rect 463222 176378 463306 176614
rect 463542 176378 463574 176614
rect 462954 176294 463574 176378
rect 462954 176058 462986 176294
rect 463222 176058 463306 176294
rect 463542 176058 463574 176294
rect 462954 140614 463574 176058
rect 462954 140378 462986 140614
rect 463222 140378 463306 140614
rect 463542 140378 463574 140614
rect 462954 140294 463574 140378
rect 462954 140058 462986 140294
rect 463222 140058 463306 140294
rect 463542 140058 463574 140294
rect 462954 104614 463574 140058
rect 462954 104378 462986 104614
rect 463222 104378 463306 104614
rect 463542 104378 463574 104614
rect 462954 104294 463574 104378
rect 462954 104058 462986 104294
rect 463222 104058 463306 104294
rect 463542 104058 463574 104294
rect 462954 68614 463574 104058
rect 462954 68378 462986 68614
rect 463222 68378 463306 68614
rect 463542 68378 463574 68614
rect 462954 68294 463574 68378
rect 462954 68058 462986 68294
rect 463222 68058 463306 68294
rect 463542 68058 463574 68294
rect 462954 32614 463574 68058
rect 462954 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 463574 32614
rect 462954 32294 463574 32378
rect 462954 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 463574 32294
rect 444954 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 445574 -6106
rect 444954 -6426 445574 -6342
rect 444954 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 445574 -6426
rect 444954 -7654 445574 -6662
rect 462954 -7066 463574 32058
rect 469794 704838 470414 705830
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 363454 470414 398898
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 291454 470414 326898
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -1894 470414 -902
rect 473514 691174 474134 706202
rect 473514 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 474134 691174
rect 473514 690854 474134 690938
rect 473514 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 474134 690854
rect 473514 655174 474134 690618
rect 473514 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 474134 655174
rect 473514 654854 474134 654938
rect 473514 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 474134 654854
rect 473514 619174 474134 654618
rect 473514 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 474134 619174
rect 473514 618854 474134 618938
rect 473514 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 474134 618854
rect 473514 583174 474134 618618
rect 473514 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 474134 583174
rect 473514 582854 474134 582938
rect 473514 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 474134 582854
rect 473514 547174 474134 582618
rect 473514 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 474134 547174
rect 473514 546854 474134 546938
rect 473514 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 474134 546854
rect 473514 511174 474134 546618
rect 473514 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 474134 511174
rect 473514 510854 474134 510938
rect 473514 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 474134 510854
rect 473514 475174 474134 510618
rect 473514 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 474134 475174
rect 473514 474854 474134 474938
rect 473514 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 474134 474854
rect 473514 439174 474134 474618
rect 473514 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 474134 439174
rect 473514 438854 474134 438938
rect 473514 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 474134 438854
rect 473514 403174 474134 438618
rect 473514 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 474134 403174
rect 473514 402854 474134 402938
rect 473514 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 474134 402854
rect 473514 367174 474134 402618
rect 473514 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 474134 367174
rect 473514 366854 474134 366938
rect 473514 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 474134 366854
rect 473514 331174 474134 366618
rect 473514 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 474134 331174
rect 473514 330854 474134 330938
rect 473514 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 474134 330854
rect 473514 295174 474134 330618
rect 473514 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 474134 295174
rect 473514 294854 474134 294938
rect 473514 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 474134 294854
rect 473514 259174 474134 294618
rect 473514 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 474134 259174
rect 473514 258854 474134 258938
rect 473514 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 474134 258854
rect 473514 223174 474134 258618
rect 473514 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 474134 223174
rect 473514 222854 474134 222938
rect 473514 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 474134 222854
rect 473514 187174 474134 222618
rect 473514 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 474134 187174
rect 473514 186854 474134 186938
rect 473514 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 474134 186854
rect 473514 151174 474134 186618
rect 473514 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 474134 151174
rect 473514 150854 474134 150938
rect 473514 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 474134 150854
rect 473514 115174 474134 150618
rect 473514 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 474134 115174
rect 473514 114854 474134 114938
rect 473514 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 474134 114854
rect 473514 79174 474134 114618
rect 473514 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 474134 79174
rect 473514 78854 474134 78938
rect 473514 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 474134 78854
rect 473514 43174 474134 78618
rect 473514 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 474134 43174
rect 473514 42854 474134 42938
rect 473514 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 474134 42854
rect 473514 7174 474134 42618
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -2266 474134 6618
rect 473514 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 474134 -2266
rect 473514 -2586 474134 -2502
rect 473514 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 474134 -2586
rect 473514 -3814 474134 -2822
rect 477234 694894 477854 708122
rect 477234 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 477854 694894
rect 477234 694574 477854 694658
rect 477234 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 477854 694574
rect 477234 658894 477854 694338
rect 477234 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 477854 658894
rect 477234 658574 477854 658658
rect 477234 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 477854 658574
rect 477234 622894 477854 658338
rect 477234 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 477854 622894
rect 477234 622574 477854 622658
rect 477234 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 477854 622574
rect 477234 586894 477854 622338
rect 477234 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 477854 586894
rect 477234 586574 477854 586658
rect 477234 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 477854 586574
rect 477234 550894 477854 586338
rect 477234 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 477854 550894
rect 477234 550574 477854 550658
rect 477234 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 477854 550574
rect 477234 514894 477854 550338
rect 477234 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 477854 514894
rect 477234 514574 477854 514658
rect 477234 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 477854 514574
rect 477234 478894 477854 514338
rect 477234 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 477854 478894
rect 477234 478574 477854 478658
rect 477234 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 477854 478574
rect 477234 442894 477854 478338
rect 477234 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 477854 442894
rect 477234 442574 477854 442658
rect 477234 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 477854 442574
rect 477234 406894 477854 442338
rect 477234 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 477854 406894
rect 477234 406574 477854 406658
rect 477234 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 477854 406574
rect 477234 370894 477854 406338
rect 477234 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 477854 370894
rect 477234 370574 477854 370658
rect 477234 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 477854 370574
rect 477234 334894 477854 370338
rect 477234 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 477854 334894
rect 477234 334574 477854 334658
rect 477234 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 477854 334574
rect 477234 298894 477854 334338
rect 477234 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 477854 298894
rect 477234 298574 477854 298658
rect 477234 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 477854 298574
rect 477234 262894 477854 298338
rect 477234 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 477854 262894
rect 477234 262574 477854 262658
rect 477234 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 477854 262574
rect 477234 226894 477854 262338
rect 477234 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 477854 226894
rect 477234 226574 477854 226658
rect 477234 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 477854 226574
rect 477234 190894 477854 226338
rect 477234 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 477854 190894
rect 477234 190574 477854 190658
rect 477234 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 477854 190574
rect 477234 154894 477854 190338
rect 477234 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 477854 154894
rect 477234 154574 477854 154658
rect 477234 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 477854 154574
rect 477234 118894 477854 154338
rect 477234 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 477854 118894
rect 477234 118574 477854 118658
rect 477234 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 477854 118574
rect 477234 82894 477854 118338
rect 477234 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 477854 82894
rect 477234 82574 477854 82658
rect 477234 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 477854 82574
rect 477234 46894 477854 82338
rect 477234 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 477854 46894
rect 477234 46574 477854 46658
rect 477234 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 477854 46574
rect 477234 10894 477854 46338
rect 477234 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 477854 10894
rect 477234 10574 477854 10658
rect 477234 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 477854 10574
rect 477234 -4186 477854 10338
rect 477234 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 477854 -4186
rect 477234 -4506 477854 -4422
rect 477234 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 477854 -4506
rect 477234 -5734 477854 -4742
rect 480954 698614 481574 710042
rect 498954 711558 499574 711590
rect 498954 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 499574 711558
rect 498954 711238 499574 711322
rect 498954 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 499574 711238
rect 495234 709638 495854 709670
rect 495234 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 495854 709638
rect 495234 709318 495854 709402
rect 495234 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 495854 709318
rect 491514 707718 492134 707750
rect 491514 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 492134 707718
rect 491514 707398 492134 707482
rect 491514 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 492134 707398
rect 480954 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 481574 698614
rect 480954 698294 481574 698378
rect 480954 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 481574 698294
rect 480954 662614 481574 698058
rect 480954 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 481574 662614
rect 480954 662294 481574 662378
rect 480954 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 481574 662294
rect 480954 626614 481574 662058
rect 480954 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 481574 626614
rect 480954 626294 481574 626378
rect 480954 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 481574 626294
rect 480954 590614 481574 626058
rect 480954 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 481574 590614
rect 480954 590294 481574 590378
rect 480954 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 481574 590294
rect 480954 554614 481574 590058
rect 480954 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 481574 554614
rect 480954 554294 481574 554378
rect 480954 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 481574 554294
rect 480954 518614 481574 554058
rect 480954 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 481574 518614
rect 480954 518294 481574 518378
rect 480954 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 481574 518294
rect 480954 482614 481574 518058
rect 480954 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 481574 482614
rect 480954 482294 481574 482378
rect 480954 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 481574 482294
rect 480954 446614 481574 482058
rect 480954 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 481574 446614
rect 480954 446294 481574 446378
rect 480954 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 481574 446294
rect 480954 410614 481574 446058
rect 480954 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 481574 410614
rect 480954 410294 481574 410378
rect 480954 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 481574 410294
rect 480954 374614 481574 410058
rect 480954 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 481574 374614
rect 480954 374294 481574 374378
rect 480954 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 481574 374294
rect 480954 338614 481574 374058
rect 480954 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 481574 338614
rect 480954 338294 481574 338378
rect 480954 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 481574 338294
rect 480954 302614 481574 338058
rect 480954 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 481574 302614
rect 480954 302294 481574 302378
rect 480954 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 481574 302294
rect 480954 266614 481574 302058
rect 480954 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 481574 266614
rect 480954 266294 481574 266378
rect 480954 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 481574 266294
rect 480954 230614 481574 266058
rect 480954 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 481574 230614
rect 480954 230294 481574 230378
rect 480954 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 481574 230294
rect 480954 194614 481574 230058
rect 480954 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 481574 194614
rect 480954 194294 481574 194378
rect 480954 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 481574 194294
rect 480954 158614 481574 194058
rect 480954 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 481574 158614
rect 480954 158294 481574 158378
rect 480954 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 481574 158294
rect 480954 122614 481574 158058
rect 480954 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 481574 122614
rect 480954 122294 481574 122378
rect 480954 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 481574 122294
rect 480954 86614 481574 122058
rect 480954 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 481574 86614
rect 480954 86294 481574 86378
rect 480954 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 481574 86294
rect 480954 50614 481574 86058
rect 480954 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 481574 50614
rect 480954 50294 481574 50378
rect 480954 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 481574 50294
rect 480954 14614 481574 50058
rect 480954 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 481574 14614
rect 480954 14294 481574 14378
rect 480954 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 481574 14294
rect 462954 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 463574 -7066
rect 462954 -7386 463574 -7302
rect 462954 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 463574 -7386
rect 462954 -7654 463574 -7622
rect 480954 -6106 481574 14058
rect 487794 705798 488414 705830
rect 487794 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 488414 705798
rect 487794 705478 488414 705562
rect 487794 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 488414 705478
rect 487794 669454 488414 705242
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597454 488414 632898
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 561454 488414 596898
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 453454 488414 488898
rect 487794 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 488414 453454
rect 487794 453134 488414 453218
rect 487794 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 488414 453134
rect 487794 417454 488414 452898
rect 487794 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 488414 417454
rect 487794 417134 488414 417218
rect 487794 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 488414 417134
rect 487794 381454 488414 416898
rect 487794 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 488414 381454
rect 487794 381134 488414 381218
rect 487794 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 488414 381134
rect 487794 345454 488414 380898
rect 487794 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 488414 345454
rect 487794 345134 488414 345218
rect 487794 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 488414 345134
rect 487794 309454 488414 344898
rect 487794 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 488414 309454
rect 487794 309134 488414 309218
rect 487794 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 488414 309134
rect 487794 273454 488414 308898
rect 487794 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 488414 273454
rect 487794 273134 488414 273218
rect 487794 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 488414 273134
rect 487794 237454 488414 272898
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 487794 201454 488414 236898
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 165454 488414 200898
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 129454 488414 164898
rect 487794 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 488414 129454
rect 487794 129134 488414 129218
rect 487794 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 488414 129134
rect 487794 93454 488414 128898
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -1306 488414 20898
rect 487794 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 488414 -1306
rect 487794 -1626 488414 -1542
rect 487794 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 488414 -1626
rect 487794 -1894 488414 -1862
rect 491514 673174 492134 707162
rect 491514 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 492134 673174
rect 491514 672854 492134 672938
rect 491514 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 492134 672854
rect 491514 637174 492134 672618
rect 491514 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 492134 637174
rect 491514 636854 492134 636938
rect 491514 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 492134 636854
rect 491514 601174 492134 636618
rect 491514 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 492134 601174
rect 491514 600854 492134 600938
rect 491514 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 492134 600854
rect 491514 565174 492134 600618
rect 491514 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 492134 565174
rect 491514 564854 492134 564938
rect 491514 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 492134 564854
rect 491514 529174 492134 564618
rect 491514 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 492134 529174
rect 491514 528854 492134 528938
rect 491514 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 492134 528854
rect 491514 493174 492134 528618
rect 491514 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 492134 493174
rect 491514 492854 492134 492938
rect 491514 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 492134 492854
rect 491514 457174 492134 492618
rect 491514 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 492134 457174
rect 491514 456854 492134 456938
rect 491514 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 492134 456854
rect 491514 421174 492134 456618
rect 491514 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 492134 421174
rect 491514 420854 492134 420938
rect 491514 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 492134 420854
rect 491514 385174 492134 420618
rect 491514 384938 491546 385174
rect 491782 384938 491866 385174
rect 492102 384938 492134 385174
rect 491514 384854 492134 384938
rect 491514 384618 491546 384854
rect 491782 384618 491866 384854
rect 492102 384618 492134 384854
rect 491514 349174 492134 384618
rect 491514 348938 491546 349174
rect 491782 348938 491866 349174
rect 492102 348938 492134 349174
rect 491514 348854 492134 348938
rect 491514 348618 491546 348854
rect 491782 348618 491866 348854
rect 492102 348618 492134 348854
rect 491514 313174 492134 348618
rect 491514 312938 491546 313174
rect 491782 312938 491866 313174
rect 492102 312938 492134 313174
rect 491514 312854 492134 312938
rect 491514 312618 491546 312854
rect 491782 312618 491866 312854
rect 492102 312618 492134 312854
rect 491514 277174 492134 312618
rect 491514 276938 491546 277174
rect 491782 276938 491866 277174
rect 492102 276938 492134 277174
rect 491514 276854 492134 276938
rect 491514 276618 491546 276854
rect 491782 276618 491866 276854
rect 492102 276618 492134 276854
rect 491514 241174 492134 276618
rect 491514 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 492134 241174
rect 491514 240854 492134 240938
rect 491514 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 492134 240854
rect 491514 205174 492134 240618
rect 491514 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 492134 205174
rect 491514 204854 492134 204938
rect 491514 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 492134 204854
rect 491514 169174 492134 204618
rect 491514 168938 491546 169174
rect 491782 168938 491866 169174
rect 492102 168938 492134 169174
rect 491514 168854 492134 168938
rect 491514 168618 491546 168854
rect 491782 168618 491866 168854
rect 492102 168618 492134 168854
rect 491514 133174 492134 168618
rect 491514 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 492134 133174
rect 491514 132854 492134 132938
rect 491514 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 492134 132854
rect 491514 97174 492134 132618
rect 491514 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 492134 97174
rect 491514 96854 492134 96938
rect 491514 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 492134 96854
rect 491514 61174 492134 96618
rect 491514 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 492134 61174
rect 491514 60854 492134 60938
rect 491514 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 492134 60854
rect 491514 25174 492134 60618
rect 491514 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 492134 25174
rect 491514 24854 492134 24938
rect 491514 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 492134 24854
rect 491514 -3226 492134 24618
rect 491514 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 492134 -3226
rect 491514 -3546 492134 -3462
rect 491514 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 492134 -3546
rect 491514 -3814 492134 -3782
rect 495234 676894 495854 709082
rect 495234 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 495854 676894
rect 495234 676574 495854 676658
rect 495234 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 495854 676574
rect 495234 640894 495854 676338
rect 495234 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 495854 640894
rect 495234 640574 495854 640658
rect 495234 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 495854 640574
rect 495234 604894 495854 640338
rect 495234 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 495854 604894
rect 495234 604574 495854 604658
rect 495234 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 495854 604574
rect 495234 568894 495854 604338
rect 495234 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 495854 568894
rect 495234 568574 495854 568658
rect 495234 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 495854 568574
rect 495234 532894 495854 568338
rect 495234 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 495854 532894
rect 495234 532574 495854 532658
rect 495234 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 495854 532574
rect 495234 496894 495854 532338
rect 495234 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 495854 496894
rect 495234 496574 495854 496658
rect 495234 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 495854 496574
rect 495234 460894 495854 496338
rect 495234 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 495854 460894
rect 495234 460574 495854 460658
rect 495234 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 495854 460574
rect 495234 424894 495854 460338
rect 495234 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 495854 424894
rect 495234 424574 495854 424658
rect 495234 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 495854 424574
rect 495234 388894 495854 424338
rect 495234 388658 495266 388894
rect 495502 388658 495586 388894
rect 495822 388658 495854 388894
rect 495234 388574 495854 388658
rect 495234 388338 495266 388574
rect 495502 388338 495586 388574
rect 495822 388338 495854 388574
rect 495234 352894 495854 388338
rect 495234 352658 495266 352894
rect 495502 352658 495586 352894
rect 495822 352658 495854 352894
rect 495234 352574 495854 352658
rect 495234 352338 495266 352574
rect 495502 352338 495586 352574
rect 495822 352338 495854 352574
rect 495234 316894 495854 352338
rect 495234 316658 495266 316894
rect 495502 316658 495586 316894
rect 495822 316658 495854 316894
rect 495234 316574 495854 316658
rect 495234 316338 495266 316574
rect 495502 316338 495586 316574
rect 495822 316338 495854 316574
rect 495234 280894 495854 316338
rect 495234 280658 495266 280894
rect 495502 280658 495586 280894
rect 495822 280658 495854 280894
rect 495234 280574 495854 280658
rect 495234 280338 495266 280574
rect 495502 280338 495586 280574
rect 495822 280338 495854 280574
rect 495234 244894 495854 280338
rect 495234 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 495854 244894
rect 495234 244574 495854 244658
rect 495234 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 495854 244574
rect 495234 208894 495854 244338
rect 495234 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 495854 208894
rect 495234 208574 495854 208658
rect 495234 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 495854 208574
rect 495234 172894 495854 208338
rect 495234 172658 495266 172894
rect 495502 172658 495586 172894
rect 495822 172658 495854 172894
rect 495234 172574 495854 172658
rect 495234 172338 495266 172574
rect 495502 172338 495586 172574
rect 495822 172338 495854 172574
rect 495234 136894 495854 172338
rect 495234 136658 495266 136894
rect 495502 136658 495586 136894
rect 495822 136658 495854 136894
rect 495234 136574 495854 136658
rect 495234 136338 495266 136574
rect 495502 136338 495586 136574
rect 495822 136338 495854 136574
rect 495234 100894 495854 136338
rect 495234 100658 495266 100894
rect 495502 100658 495586 100894
rect 495822 100658 495854 100894
rect 495234 100574 495854 100658
rect 495234 100338 495266 100574
rect 495502 100338 495586 100574
rect 495822 100338 495854 100574
rect 495234 64894 495854 100338
rect 495234 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 495854 64894
rect 495234 64574 495854 64658
rect 495234 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 495854 64574
rect 495234 28894 495854 64338
rect 495234 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 495854 28894
rect 495234 28574 495854 28658
rect 495234 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 495854 28574
rect 495234 -5146 495854 28338
rect 495234 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 495854 -5146
rect 495234 -5466 495854 -5382
rect 495234 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 495854 -5466
rect 495234 -5734 495854 -5702
rect 498954 680614 499574 711002
rect 516954 710598 517574 711590
rect 516954 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 517574 710598
rect 516954 710278 517574 710362
rect 516954 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 517574 710278
rect 513234 708678 513854 709670
rect 513234 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 513854 708678
rect 513234 708358 513854 708442
rect 513234 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 513854 708358
rect 509514 706758 510134 707750
rect 509514 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 510134 706758
rect 509514 706438 510134 706522
rect 509514 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 510134 706438
rect 498954 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 499574 680614
rect 498954 680294 499574 680378
rect 498954 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 499574 680294
rect 498954 644614 499574 680058
rect 498954 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 499574 644614
rect 498954 644294 499574 644378
rect 498954 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 499574 644294
rect 498954 608614 499574 644058
rect 498954 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 499574 608614
rect 498954 608294 499574 608378
rect 498954 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 499574 608294
rect 498954 572614 499574 608058
rect 498954 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 499574 572614
rect 498954 572294 499574 572378
rect 498954 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 499574 572294
rect 498954 536614 499574 572058
rect 498954 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 499574 536614
rect 498954 536294 499574 536378
rect 498954 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 499574 536294
rect 498954 500614 499574 536058
rect 498954 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 499574 500614
rect 498954 500294 499574 500378
rect 498954 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 499574 500294
rect 498954 464614 499574 500058
rect 498954 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 499574 464614
rect 498954 464294 499574 464378
rect 498954 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 499574 464294
rect 498954 428614 499574 464058
rect 498954 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 499574 428614
rect 498954 428294 499574 428378
rect 498954 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 499574 428294
rect 498954 392614 499574 428058
rect 498954 392378 498986 392614
rect 499222 392378 499306 392614
rect 499542 392378 499574 392614
rect 498954 392294 499574 392378
rect 498954 392058 498986 392294
rect 499222 392058 499306 392294
rect 499542 392058 499574 392294
rect 498954 356614 499574 392058
rect 498954 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 499574 356614
rect 498954 356294 499574 356378
rect 498954 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 499574 356294
rect 498954 320614 499574 356058
rect 498954 320378 498986 320614
rect 499222 320378 499306 320614
rect 499542 320378 499574 320614
rect 498954 320294 499574 320378
rect 498954 320058 498986 320294
rect 499222 320058 499306 320294
rect 499542 320058 499574 320294
rect 498954 284614 499574 320058
rect 498954 284378 498986 284614
rect 499222 284378 499306 284614
rect 499542 284378 499574 284614
rect 498954 284294 499574 284378
rect 498954 284058 498986 284294
rect 499222 284058 499306 284294
rect 499542 284058 499574 284294
rect 498954 248614 499574 284058
rect 498954 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 499574 248614
rect 498954 248294 499574 248378
rect 498954 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 499574 248294
rect 498954 212614 499574 248058
rect 498954 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 499574 212614
rect 498954 212294 499574 212378
rect 498954 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 499574 212294
rect 498954 176614 499574 212058
rect 498954 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 499574 176614
rect 498954 176294 499574 176378
rect 498954 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 499574 176294
rect 498954 140614 499574 176058
rect 498954 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 499574 140614
rect 498954 140294 499574 140378
rect 498954 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 499574 140294
rect 498954 104614 499574 140058
rect 498954 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 499574 104614
rect 498954 104294 499574 104378
rect 498954 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 499574 104294
rect 498954 68614 499574 104058
rect 498954 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 499574 68614
rect 498954 68294 499574 68378
rect 498954 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 499574 68294
rect 498954 32614 499574 68058
rect 498954 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 499574 32614
rect 498954 32294 499574 32378
rect 498954 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 499574 32294
rect 480954 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 481574 -6106
rect 480954 -6426 481574 -6342
rect 480954 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 481574 -6426
rect 480954 -7654 481574 -6662
rect 498954 -7066 499574 32058
rect 505794 704838 506414 705830
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -1894 506414 -902
rect 509514 691174 510134 706202
rect 509514 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 510134 691174
rect 509514 690854 510134 690938
rect 509514 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 510134 690854
rect 509514 655174 510134 690618
rect 509514 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 510134 655174
rect 509514 654854 510134 654938
rect 509514 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 510134 654854
rect 509514 619174 510134 654618
rect 509514 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 510134 619174
rect 509514 618854 510134 618938
rect 509514 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 510134 618854
rect 509514 583174 510134 618618
rect 509514 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 510134 583174
rect 509514 582854 510134 582938
rect 509514 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 510134 582854
rect 509514 547174 510134 582618
rect 509514 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 510134 547174
rect 509514 546854 510134 546938
rect 509514 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 510134 546854
rect 509514 511174 510134 546618
rect 509514 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 510134 511174
rect 509514 510854 510134 510938
rect 509514 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 510134 510854
rect 509514 475174 510134 510618
rect 509514 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 510134 475174
rect 509514 474854 510134 474938
rect 509514 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 510134 474854
rect 509514 439174 510134 474618
rect 509514 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 510134 439174
rect 509514 438854 510134 438938
rect 509514 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 510134 438854
rect 509514 403174 510134 438618
rect 509514 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 510134 403174
rect 509514 402854 510134 402938
rect 509514 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 510134 402854
rect 509514 367174 510134 402618
rect 509514 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 510134 367174
rect 509514 366854 510134 366938
rect 509514 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 510134 366854
rect 509514 331174 510134 366618
rect 509514 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 510134 331174
rect 509514 330854 510134 330938
rect 509514 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 510134 330854
rect 509514 295174 510134 330618
rect 509514 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 510134 295174
rect 509514 294854 510134 294938
rect 509514 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 510134 294854
rect 509514 259174 510134 294618
rect 509514 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 510134 259174
rect 509514 258854 510134 258938
rect 509514 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 510134 258854
rect 509514 223174 510134 258618
rect 509514 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 510134 223174
rect 509514 222854 510134 222938
rect 509514 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 510134 222854
rect 509514 187174 510134 222618
rect 509514 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 510134 187174
rect 509514 186854 510134 186938
rect 509514 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 510134 186854
rect 509514 151174 510134 186618
rect 509514 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 510134 151174
rect 509514 150854 510134 150938
rect 509514 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 510134 150854
rect 509514 115174 510134 150618
rect 509514 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 510134 115174
rect 509514 114854 510134 114938
rect 509514 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 510134 114854
rect 509514 79174 510134 114618
rect 509514 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 510134 79174
rect 509514 78854 510134 78938
rect 509514 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 510134 78854
rect 509514 43174 510134 78618
rect 509514 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 510134 43174
rect 509514 42854 510134 42938
rect 509514 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 510134 42854
rect 509514 7174 510134 42618
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -2266 510134 6618
rect 509514 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 510134 -2266
rect 509514 -2586 510134 -2502
rect 509514 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 510134 -2586
rect 509514 -3814 510134 -2822
rect 513234 694894 513854 708122
rect 513234 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 513854 694894
rect 513234 694574 513854 694658
rect 513234 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 513854 694574
rect 513234 658894 513854 694338
rect 513234 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 513854 658894
rect 513234 658574 513854 658658
rect 513234 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 513854 658574
rect 513234 622894 513854 658338
rect 513234 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 513854 622894
rect 513234 622574 513854 622658
rect 513234 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 513854 622574
rect 513234 586894 513854 622338
rect 513234 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 513854 586894
rect 513234 586574 513854 586658
rect 513234 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 513854 586574
rect 513234 550894 513854 586338
rect 513234 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 513854 550894
rect 513234 550574 513854 550658
rect 513234 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 513854 550574
rect 513234 514894 513854 550338
rect 513234 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 513854 514894
rect 513234 514574 513854 514658
rect 513234 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 513854 514574
rect 513234 478894 513854 514338
rect 513234 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 513854 478894
rect 513234 478574 513854 478658
rect 513234 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 513854 478574
rect 513234 442894 513854 478338
rect 513234 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 513854 442894
rect 513234 442574 513854 442658
rect 513234 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 513854 442574
rect 513234 406894 513854 442338
rect 513234 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 513854 406894
rect 513234 406574 513854 406658
rect 513234 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 513854 406574
rect 513234 370894 513854 406338
rect 513234 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 513854 370894
rect 513234 370574 513854 370658
rect 513234 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 513854 370574
rect 513234 334894 513854 370338
rect 513234 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 513854 334894
rect 513234 334574 513854 334658
rect 513234 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 513854 334574
rect 513234 298894 513854 334338
rect 513234 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 513854 298894
rect 513234 298574 513854 298658
rect 513234 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 513854 298574
rect 513234 262894 513854 298338
rect 513234 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 513854 262894
rect 513234 262574 513854 262658
rect 513234 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 513854 262574
rect 513234 226894 513854 262338
rect 513234 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 513854 226894
rect 513234 226574 513854 226658
rect 513234 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 513854 226574
rect 513234 190894 513854 226338
rect 513234 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 513854 190894
rect 513234 190574 513854 190658
rect 513234 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 513854 190574
rect 513234 154894 513854 190338
rect 513234 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 513854 154894
rect 513234 154574 513854 154658
rect 513234 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 513854 154574
rect 513234 118894 513854 154338
rect 513234 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 513854 118894
rect 513234 118574 513854 118658
rect 513234 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 513854 118574
rect 513234 82894 513854 118338
rect 513234 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 513854 82894
rect 513234 82574 513854 82658
rect 513234 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 513854 82574
rect 513234 46894 513854 82338
rect 513234 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 513854 46894
rect 513234 46574 513854 46658
rect 513234 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 513854 46574
rect 513234 10894 513854 46338
rect 513234 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 513854 10894
rect 513234 10574 513854 10658
rect 513234 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 513854 10574
rect 513234 -4186 513854 10338
rect 513234 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 513854 -4186
rect 513234 -4506 513854 -4422
rect 513234 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 513854 -4506
rect 513234 -5734 513854 -4742
rect 516954 698614 517574 710042
rect 534954 711558 535574 711590
rect 534954 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 535574 711558
rect 534954 711238 535574 711322
rect 534954 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 535574 711238
rect 531234 709638 531854 709670
rect 531234 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 531854 709638
rect 531234 709318 531854 709402
rect 531234 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 531854 709318
rect 527514 707718 528134 707750
rect 527514 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 528134 707718
rect 527514 707398 528134 707482
rect 527514 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 528134 707398
rect 516954 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 517574 698614
rect 516954 698294 517574 698378
rect 516954 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 517574 698294
rect 516954 662614 517574 698058
rect 516954 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 517574 662614
rect 516954 662294 517574 662378
rect 516954 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 517574 662294
rect 516954 626614 517574 662058
rect 516954 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 517574 626614
rect 516954 626294 517574 626378
rect 516954 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 517574 626294
rect 516954 590614 517574 626058
rect 516954 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 517574 590614
rect 516954 590294 517574 590378
rect 516954 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 517574 590294
rect 516954 554614 517574 590058
rect 516954 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 517574 554614
rect 516954 554294 517574 554378
rect 516954 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 517574 554294
rect 516954 518614 517574 554058
rect 516954 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 517574 518614
rect 516954 518294 517574 518378
rect 516954 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 517574 518294
rect 516954 482614 517574 518058
rect 516954 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 517574 482614
rect 516954 482294 517574 482378
rect 516954 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 517574 482294
rect 516954 446614 517574 482058
rect 516954 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 517574 446614
rect 516954 446294 517574 446378
rect 516954 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 517574 446294
rect 516954 410614 517574 446058
rect 516954 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 517574 410614
rect 516954 410294 517574 410378
rect 516954 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 517574 410294
rect 516954 374614 517574 410058
rect 516954 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 517574 374614
rect 516954 374294 517574 374378
rect 516954 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 517574 374294
rect 516954 338614 517574 374058
rect 516954 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 517574 338614
rect 516954 338294 517574 338378
rect 516954 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 517574 338294
rect 516954 302614 517574 338058
rect 516954 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 517574 302614
rect 516954 302294 517574 302378
rect 516954 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 517574 302294
rect 516954 266614 517574 302058
rect 516954 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 517574 266614
rect 516954 266294 517574 266378
rect 516954 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 517574 266294
rect 516954 230614 517574 266058
rect 516954 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 517574 230614
rect 516954 230294 517574 230378
rect 516954 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 517574 230294
rect 516954 194614 517574 230058
rect 516954 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 517574 194614
rect 516954 194294 517574 194378
rect 516954 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 517574 194294
rect 516954 158614 517574 194058
rect 516954 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 517574 158614
rect 516954 158294 517574 158378
rect 516954 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 517574 158294
rect 516954 122614 517574 158058
rect 516954 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 517574 122614
rect 516954 122294 517574 122378
rect 516954 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 517574 122294
rect 516954 86614 517574 122058
rect 516954 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 517574 86614
rect 516954 86294 517574 86378
rect 516954 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 517574 86294
rect 516954 50614 517574 86058
rect 516954 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 517574 50614
rect 516954 50294 517574 50378
rect 516954 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 517574 50294
rect 516954 14614 517574 50058
rect 516954 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 517574 14614
rect 516954 14294 517574 14378
rect 516954 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 517574 14294
rect 498954 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 499574 -7066
rect 498954 -7386 499574 -7302
rect 498954 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 499574 -7386
rect 498954 -7654 499574 -7622
rect 516954 -6106 517574 14058
rect 523794 705798 524414 705830
rect 523794 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 524414 705798
rect 523794 705478 524414 705562
rect 523794 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 524414 705478
rect 523794 669454 524414 705242
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -1306 524414 20898
rect 523794 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 524414 -1306
rect 523794 -1626 524414 -1542
rect 523794 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 524414 -1626
rect 523794 -1894 524414 -1862
rect 527514 673174 528134 707162
rect 527514 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 528134 673174
rect 527514 672854 528134 672938
rect 527514 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 528134 672854
rect 527514 637174 528134 672618
rect 527514 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 528134 637174
rect 527514 636854 528134 636938
rect 527514 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 528134 636854
rect 527514 601174 528134 636618
rect 527514 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 528134 601174
rect 527514 600854 528134 600938
rect 527514 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 528134 600854
rect 527514 565174 528134 600618
rect 527514 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 528134 565174
rect 527514 564854 528134 564938
rect 527514 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 528134 564854
rect 527514 529174 528134 564618
rect 527514 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 528134 529174
rect 527514 528854 528134 528938
rect 527514 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 528134 528854
rect 527514 493174 528134 528618
rect 527514 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 528134 493174
rect 527514 492854 528134 492938
rect 527514 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 528134 492854
rect 527514 457174 528134 492618
rect 527514 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 528134 457174
rect 527514 456854 528134 456938
rect 527514 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 528134 456854
rect 527514 421174 528134 456618
rect 527514 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 528134 421174
rect 527514 420854 528134 420938
rect 527514 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 528134 420854
rect 527514 385174 528134 420618
rect 527514 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 528134 385174
rect 527514 384854 528134 384938
rect 527514 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 528134 384854
rect 527514 349174 528134 384618
rect 527514 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 528134 349174
rect 527514 348854 528134 348938
rect 527514 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 528134 348854
rect 527514 313174 528134 348618
rect 527514 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 528134 313174
rect 527514 312854 528134 312938
rect 527514 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 528134 312854
rect 527514 277174 528134 312618
rect 527514 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 528134 277174
rect 527514 276854 528134 276938
rect 527514 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 528134 276854
rect 527514 241174 528134 276618
rect 527514 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 528134 241174
rect 527514 240854 528134 240938
rect 527514 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 528134 240854
rect 527514 205174 528134 240618
rect 527514 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 528134 205174
rect 527514 204854 528134 204938
rect 527514 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 528134 204854
rect 527514 169174 528134 204618
rect 527514 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 528134 169174
rect 527514 168854 528134 168938
rect 527514 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 528134 168854
rect 527514 133174 528134 168618
rect 527514 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 528134 133174
rect 527514 132854 528134 132938
rect 527514 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 528134 132854
rect 527514 97174 528134 132618
rect 527514 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 528134 97174
rect 527514 96854 528134 96938
rect 527514 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 528134 96854
rect 527514 61174 528134 96618
rect 527514 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 528134 61174
rect 527514 60854 528134 60938
rect 527514 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 528134 60854
rect 527514 25174 528134 60618
rect 527514 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 528134 25174
rect 527514 24854 528134 24938
rect 527514 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 528134 24854
rect 527514 -3226 528134 24618
rect 527514 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 528134 -3226
rect 527514 -3546 528134 -3462
rect 527514 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 528134 -3546
rect 527514 -3814 528134 -3782
rect 531234 676894 531854 709082
rect 531234 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 531854 676894
rect 531234 676574 531854 676658
rect 531234 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 531854 676574
rect 531234 640894 531854 676338
rect 531234 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 531854 640894
rect 531234 640574 531854 640658
rect 531234 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 531854 640574
rect 531234 604894 531854 640338
rect 531234 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 531854 604894
rect 531234 604574 531854 604658
rect 531234 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 531854 604574
rect 531234 568894 531854 604338
rect 531234 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 531854 568894
rect 531234 568574 531854 568658
rect 531234 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 531854 568574
rect 531234 532894 531854 568338
rect 531234 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 531854 532894
rect 531234 532574 531854 532658
rect 531234 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 531854 532574
rect 531234 496894 531854 532338
rect 531234 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 531854 496894
rect 531234 496574 531854 496658
rect 531234 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 531854 496574
rect 531234 460894 531854 496338
rect 531234 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 531854 460894
rect 531234 460574 531854 460658
rect 531234 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 531854 460574
rect 531234 424894 531854 460338
rect 531234 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 531854 424894
rect 531234 424574 531854 424658
rect 531234 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 531854 424574
rect 531234 388894 531854 424338
rect 531234 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 531854 388894
rect 531234 388574 531854 388658
rect 531234 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 531854 388574
rect 531234 352894 531854 388338
rect 531234 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 531854 352894
rect 531234 352574 531854 352658
rect 531234 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 531854 352574
rect 531234 316894 531854 352338
rect 531234 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 531854 316894
rect 531234 316574 531854 316658
rect 531234 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 531854 316574
rect 531234 280894 531854 316338
rect 531234 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 531854 280894
rect 531234 280574 531854 280658
rect 531234 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 531854 280574
rect 531234 244894 531854 280338
rect 531234 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 531854 244894
rect 531234 244574 531854 244658
rect 531234 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 531854 244574
rect 531234 208894 531854 244338
rect 531234 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 531854 208894
rect 531234 208574 531854 208658
rect 531234 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 531854 208574
rect 531234 172894 531854 208338
rect 531234 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 531854 172894
rect 531234 172574 531854 172658
rect 531234 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 531854 172574
rect 531234 136894 531854 172338
rect 531234 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 531854 136894
rect 531234 136574 531854 136658
rect 531234 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 531854 136574
rect 531234 100894 531854 136338
rect 531234 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 531854 100894
rect 531234 100574 531854 100658
rect 531234 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 531854 100574
rect 531234 64894 531854 100338
rect 531234 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 531854 64894
rect 531234 64574 531854 64658
rect 531234 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 531854 64574
rect 531234 28894 531854 64338
rect 531234 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 531854 28894
rect 531234 28574 531854 28658
rect 531234 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 531854 28574
rect 531234 -5146 531854 28338
rect 531234 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 531854 -5146
rect 531234 -5466 531854 -5382
rect 531234 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 531854 -5466
rect 531234 -5734 531854 -5702
rect 534954 680614 535574 711002
rect 552954 710598 553574 711590
rect 552954 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 553574 710598
rect 552954 710278 553574 710362
rect 552954 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 553574 710278
rect 549234 708678 549854 709670
rect 549234 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 549854 708678
rect 549234 708358 549854 708442
rect 549234 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 549854 708358
rect 545514 706758 546134 707750
rect 545514 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 546134 706758
rect 545514 706438 546134 706522
rect 545514 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 546134 706438
rect 534954 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 535574 680614
rect 534954 680294 535574 680378
rect 534954 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 535574 680294
rect 534954 644614 535574 680058
rect 534954 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 535574 644614
rect 534954 644294 535574 644378
rect 534954 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 535574 644294
rect 534954 608614 535574 644058
rect 534954 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 535574 608614
rect 534954 608294 535574 608378
rect 534954 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 535574 608294
rect 534954 572614 535574 608058
rect 534954 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 535574 572614
rect 534954 572294 535574 572378
rect 534954 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 535574 572294
rect 534954 536614 535574 572058
rect 534954 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 535574 536614
rect 534954 536294 535574 536378
rect 534954 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 535574 536294
rect 534954 500614 535574 536058
rect 534954 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 535574 500614
rect 534954 500294 535574 500378
rect 534954 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 535574 500294
rect 534954 464614 535574 500058
rect 534954 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 535574 464614
rect 534954 464294 535574 464378
rect 534954 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 535574 464294
rect 534954 428614 535574 464058
rect 534954 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 535574 428614
rect 534954 428294 535574 428378
rect 534954 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 535574 428294
rect 534954 392614 535574 428058
rect 534954 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 535574 392614
rect 534954 392294 535574 392378
rect 534954 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 535574 392294
rect 534954 356614 535574 392058
rect 534954 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 535574 356614
rect 534954 356294 535574 356378
rect 534954 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 535574 356294
rect 534954 320614 535574 356058
rect 534954 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 535574 320614
rect 534954 320294 535574 320378
rect 534954 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 535574 320294
rect 534954 284614 535574 320058
rect 534954 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 535574 284614
rect 534954 284294 535574 284378
rect 534954 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 535574 284294
rect 534954 248614 535574 284058
rect 534954 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 535574 248614
rect 534954 248294 535574 248378
rect 534954 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 535574 248294
rect 534954 212614 535574 248058
rect 534954 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 535574 212614
rect 534954 212294 535574 212378
rect 534954 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 535574 212294
rect 534954 176614 535574 212058
rect 534954 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 535574 176614
rect 534954 176294 535574 176378
rect 534954 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 535574 176294
rect 534954 140614 535574 176058
rect 534954 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 535574 140614
rect 534954 140294 535574 140378
rect 534954 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 535574 140294
rect 534954 104614 535574 140058
rect 534954 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 535574 104614
rect 534954 104294 535574 104378
rect 534954 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 535574 104294
rect 534954 68614 535574 104058
rect 534954 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 535574 68614
rect 534954 68294 535574 68378
rect 534954 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 535574 68294
rect 534954 32614 535574 68058
rect 534954 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 535574 32614
rect 534954 32294 535574 32378
rect 534954 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 535574 32294
rect 516954 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 517574 -6106
rect 516954 -6426 517574 -6342
rect 516954 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 517574 -6426
rect 516954 -7654 517574 -6662
rect 534954 -7066 535574 32058
rect 541794 704838 542414 705830
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -1894 542414 -902
rect 545514 691174 546134 706202
rect 545514 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 546134 691174
rect 545514 690854 546134 690938
rect 545514 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 546134 690854
rect 545514 655174 546134 690618
rect 545514 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 546134 655174
rect 545514 654854 546134 654938
rect 545514 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 546134 654854
rect 545514 619174 546134 654618
rect 545514 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 546134 619174
rect 545514 618854 546134 618938
rect 545514 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 546134 618854
rect 545514 583174 546134 618618
rect 545514 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 546134 583174
rect 545514 582854 546134 582938
rect 545514 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 546134 582854
rect 545514 547174 546134 582618
rect 545514 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 546134 547174
rect 545514 546854 546134 546938
rect 545514 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 546134 546854
rect 545514 511174 546134 546618
rect 545514 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 546134 511174
rect 545514 510854 546134 510938
rect 545514 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 546134 510854
rect 545514 475174 546134 510618
rect 545514 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 546134 475174
rect 545514 474854 546134 474938
rect 545514 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 546134 474854
rect 545514 439174 546134 474618
rect 545514 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 546134 439174
rect 545514 438854 546134 438938
rect 545514 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 546134 438854
rect 545514 403174 546134 438618
rect 545514 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 546134 403174
rect 545514 402854 546134 402938
rect 545514 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 546134 402854
rect 545514 367174 546134 402618
rect 545514 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 546134 367174
rect 545514 366854 546134 366938
rect 545514 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 546134 366854
rect 545514 331174 546134 366618
rect 545514 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 546134 331174
rect 545514 330854 546134 330938
rect 545514 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 546134 330854
rect 545514 295174 546134 330618
rect 545514 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 546134 295174
rect 545514 294854 546134 294938
rect 545514 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 546134 294854
rect 545514 259174 546134 294618
rect 545514 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 546134 259174
rect 545514 258854 546134 258938
rect 545514 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 546134 258854
rect 545514 223174 546134 258618
rect 545514 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 546134 223174
rect 545514 222854 546134 222938
rect 545514 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 546134 222854
rect 545514 187174 546134 222618
rect 545514 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 546134 187174
rect 545514 186854 546134 186938
rect 545514 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 546134 186854
rect 545514 151174 546134 186618
rect 545514 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 546134 151174
rect 545514 150854 546134 150938
rect 545514 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 546134 150854
rect 545514 115174 546134 150618
rect 545514 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 546134 115174
rect 545514 114854 546134 114938
rect 545514 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 546134 114854
rect 545514 79174 546134 114618
rect 545514 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 546134 79174
rect 545514 78854 546134 78938
rect 545514 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 546134 78854
rect 545514 43174 546134 78618
rect 545514 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 546134 43174
rect 545514 42854 546134 42938
rect 545514 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 546134 42854
rect 545514 7174 546134 42618
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -2266 546134 6618
rect 545514 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 546134 -2266
rect 545514 -2586 546134 -2502
rect 545514 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 546134 -2586
rect 545514 -3814 546134 -2822
rect 549234 694894 549854 708122
rect 549234 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 549854 694894
rect 549234 694574 549854 694658
rect 549234 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 549854 694574
rect 549234 658894 549854 694338
rect 549234 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 549854 658894
rect 549234 658574 549854 658658
rect 549234 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 549854 658574
rect 549234 622894 549854 658338
rect 549234 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 549854 622894
rect 549234 622574 549854 622658
rect 549234 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 549854 622574
rect 549234 586894 549854 622338
rect 549234 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 549854 586894
rect 549234 586574 549854 586658
rect 549234 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 549854 586574
rect 549234 550894 549854 586338
rect 549234 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 549854 550894
rect 549234 550574 549854 550658
rect 549234 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 549854 550574
rect 549234 514894 549854 550338
rect 549234 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 549854 514894
rect 549234 514574 549854 514658
rect 549234 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 549854 514574
rect 549234 478894 549854 514338
rect 549234 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 549854 478894
rect 549234 478574 549854 478658
rect 549234 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 549854 478574
rect 549234 442894 549854 478338
rect 549234 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 549854 442894
rect 549234 442574 549854 442658
rect 549234 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 549854 442574
rect 549234 406894 549854 442338
rect 549234 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 549854 406894
rect 549234 406574 549854 406658
rect 549234 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 549854 406574
rect 549234 370894 549854 406338
rect 549234 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 549854 370894
rect 549234 370574 549854 370658
rect 549234 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 549854 370574
rect 549234 334894 549854 370338
rect 549234 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 549854 334894
rect 549234 334574 549854 334658
rect 549234 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 549854 334574
rect 549234 298894 549854 334338
rect 549234 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 549854 298894
rect 549234 298574 549854 298658
rect 549234 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 549854 298574
rect 549234 262894 549854 298338
rect 549234 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 549854 262894
rect 549234 262574 549854 262658
rect 549234 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 549854 262574
rect 549234 226894 549854 262338
rect 549234 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 549854 226894
rect 549234 226574 549854 226658
rect 549234 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 549854 226574
rect 549234 190894 549854 226338
rect 549234 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 549854 190894
rect 549234 190574 549854 190658
rect 549234 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 549854 190574
rect 549234 154894 549854 190338
rect 549234 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 549854 154894
rect 549234 154574 549854 154658
rect 549234 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 549854 154574
rect 549234 118894 549854 154338
rect 549234 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 549854 118894
rect 549234 118574 549854 118658
rect 549234 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 549854 118574
rect 549234 82894 549854 118338
rect 549234 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 549854 82894
rect 549234 82574 549854 82658
rect 549234 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 549854 82574
rect 549234 46894 549854 82338
rect 549234 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 549854 46894
rect 549234 46574 549854 46658
rect 549234 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 549854 46574
rect 549234 10894 549854 46338
rect 549234 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 549854 10894
rect 549234 10574 549854 10658
rect 549234 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 549854 10574
rect 549234 -4186 549854 10338
rect 549234 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 549854 -4186
rect 549234 -4506 549854 -4422
rect 549234 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 549854 -4506
rect 549234 -5734 549854 -4742
rect 552954 698614 553574 710042
rect 570954 711558 571574 711590
rect 570954 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 571574 711558
rect 570954 711238 571574 711322
rect 570954 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 571574 711238
rect 567234 709638 567854 709670
rect 567234 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 567854 709638
rect 567234 709318 567854 709402
rect 567234 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 567854 709318
rect 563514 707718 564134 707750
rect 563514 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 564134 707718
rect 563514 707398 564134 707482
rect 563514 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 564134 707398
rect 552954 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 553574 698614
rect 552954 698294 553574 698378
rect 552954 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 553574 698294
rect 552954 662614 553574 698058
rect 552954 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 553574 662614
rect 552954 662294 553574 662378
rect 552954 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 553574 662294
rect 552954 626614 553574 662058
rect 552954 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 553574 626614
rect 552954 626294 553574 626378
rect 552954 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 553574 626294
rect 552954 590614 553574 626058
rect 552954 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 553574 590614
rect 552954 590294 553574 590378
rect 552954 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 553574 590294
rect 552954 554614 553574 590058
rect 552954 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 553574 554614
rect 552954 554294 553574 554378
rect 552954 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 553574 554294
rect 552954 518614 553574 554058
rect 552954 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 553574 518614
rect 552954 518294 553574 518378
rect 552954 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 553574 518294
rect 552954 482614 553574 518058
rect 552954 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 553574 482614
rect 552954 482294 553574 482378
rect 552954 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 553574 482294
rect 552954 446614 553574 482058
rect 552954 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 553574 446614
rect 552954 446294 553574 446378
rect 552954 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 553574 446294
rect 552954 410614 553574 446058
rect 552954 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 553574 410614
rect 552954 410294 553574 410378
rect 552954 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 553574 410294
rect 552954 374614 553574 410058
rect 552954 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 553574 374614
rect 552954 374294 553574 374378
rect 552954 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 553574 374294
rect 552954 338614 553574 374058
rect 552954 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 553574 338614
rect 552954 338294 553574 338378
rect 552954 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 553574 338294
rect 552954 302614 553574 338058
rect 552954 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 553574 302614
rect 552954 302294 553574 302378
rect 552954 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 553574 302294
rect 552954 266614 553574 302058
rect 552954 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 553574 266614
rect 552954 266294 553574 266378
rect 552954 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 553574 266294
rect 552954 230614 553574 266058
rect 552954 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 553574 230614
rect 552954 230294 553574 230378
rect 552954 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 553574 230294
rect 552954 194614 553574 230058
rect 552954 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 553574 194614
rect 552954 194294 553574 194378
rect 552954 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 553574 194294
rect 552954 158614 553574 194058
rect 552954 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 553574 158614
rect 552954 158294 553574 158378
rect 552954 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 553574 158294
rect 552954 122614 553574 158058
rect 552954 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 553574 122614
rect 552954 122294 553574 122378
rect 552954 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 553574 122294
rect 552954 86614 553574 122058
rect 552954 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 553574 86614
rect 552954 86294 553574 86378
rect 552954 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 553574 86294
rect 552954 50614 553574 86058
rect 552954 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 553574 50614
rect 552954 50294 553574 50378
rect 552954 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 553574 50294
rect 552954 14614 553574 50058
rect 552954 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 553574 14614
rect 552954 14294 553574 14378
rect 552954 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 553574 14294
rect 534954 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 535574 -7066
rect 534954 -7386 535574 -7302
rect 534954 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 535574 -7386
rect 534954 -7654 535574 -7622
rect 552954 -6106 553574 14058
rect 559794 705798 560414 705830
rect 559794 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 560414 705798
rect 559794 705478 560414 705562
rect 559794 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 560414 705478
rect 559794 669454 560414 705242
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -1306 560414 20898
rect 559794 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 560414 -1306
rect 559794 -1626 560414 -1542
rect 559794 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 560414 -1626
rect 559794 -1894 560414 -1862
rect 563514 673174 564134 707162
rect 563514 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 564134 673174
rect 563514 672854 564134 672938
rect 563514 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 564134 672854
rect 563514 637174 564134 672618
rect 563514 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 564134 637174
rect 563514 636854 564134 636938
rect 563514 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 564134 636854
rect 563514 601174 564134 636618
rect 563514 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 564134 601174
rect 563514 600854 564134 600938
rect 563514 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 564134 600854
rect 563514 565174 564134 600618
rect 563514 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 564134 565174
rect 563514 564854 564134 564938
rect 563514 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 564134 564854
rect 563514 529174 564134 564618
rect 563514 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 564134 529174
rect 563514 528854 564134 528938
rect 563514 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 564134 528854
rect 563514 493174 564134 528618
rect 563514 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 564134 493174
rect 563514 492854 564134 492938
rect 563514 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 564134 492854
rect 563514 457174 564134 492618
rect 563514 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 564134 457174
rect 563514 456854 564134 456938
rect 563514 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 564134 456854
rect 563514 421174 564134 456618
rect 563514 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 564134 421174
rect 563514 420854 564134 420938
rect 563514 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 564134 420854
rect 563514 385174 564134 420618
rect 563514 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 564134 385174
rect 563514 384854 564134 384938
rect 563514 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 564134 384854
rect 563514 349174 564134 384618
rect 563514 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 564134 349174
rect 563514 348854 564134 348938
rect 563514 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 564134 348854
rect 563514 313174 564134 348618
rect 563514 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 564134 313174
rect 563514 312854 564134 312938
rect 563514 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 564134 312854
rect 563514 277174 564134 312618
rect 563514 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 564134 277174
rect 563514 276854 564134 276938
rect 563514 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 564134 276854
rect 563514 241174 564134 276618
rect 563514 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 564134 241174
rect 563514 240854 564134 240938
rect 563514 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 564134 240854
rect 563514 205174 564134 240618
rect 563514 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 564134 205174
rect 563514 204854 564134 204938
rect 563514 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 564134 204854
rect 563514 169174 564134 204618
rect 563514 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 564134 169174
rect 563514 168854 564134 168938
rect 563514 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 564134 168854
rect 563514 133174 564134 168618
rect 563514 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 564134 133174
rect 563514 132854 564134 132938
rect 563514 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 564134 132854
rect 563514 97174 564134 132618
rect 563514 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 564134 97174
rect 563514 96854 564134 96938
rect 563514 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 564134 96854
rect 563514 61174 564134 96618
rect 563514 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 564134 61174
rect 563514 60854 564134 60938
rect 563514 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 564134 60854
rect 563514 25174 564134 60618
rect 563514 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 564134 25174
rect 563514 24854 564134 24938
rect 563514 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 564134 24854
rect 563514 -3226 564134 24618
rect 563514 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 564134 -3226
rect 563514 -3546 564134 -3462
rect 563514 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 564134 -3546
rect 563514 -3814 564134 -3782
rect 567234 676894 567854 709082
rect 567234 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 567854 676894
rect 567234 676574 567854 676658
rect 567234 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 567854 676574
rect 567234 640894 567854 676338
rect 567234 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 567854 640894
rect 567234 640574 567854 640658
rect 567234 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 567854 640574
rect 567234 604894 567854 640338
rect 567234 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 567854 604894
rect 567234 604574 567854 604658
rect 567234 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 567854 604574
rect 567234 568894 567854 604338
rect 567234 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 567854 568894
rect 567234 568574 567854 568658
rect 567234 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 567854 568574
rect 567234 532894 567854 568338
rect 567234 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 567854 532894
rect 567234 532574 567854 532658
rect 567234 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 567854 532574
rect 567234 496894 567854 532338
rect 567234 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 567854 496894
rect 567234 496574 567854 496658
rect 567234 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 567854 496574
rect 567234 460894 567854 496338
rect 567234 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 567854 460894
rect 567234 460574 567854 460658
rect 567234 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 567854 460574
rect 567234 424894 567854 460338
rect 567234 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 567854 424894
rect 567234 424574 567854 424658
rect 567234 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 567854 424574
rect 567234 388894 567854 424338
rect 567234 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 567854 388894
rect 567234 388574 567854 388658
rect 567234 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 567854 388574
rect 567234 352894 567854 388338
rect 567234 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 567854 352894
rect 567234 352574 567854 352658
rect 567234 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 567854 352574
rect 567234 316894 567854 352338
rect 567234 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 567854 316894
rect 567234 316574 567854 316658
rect 567234 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 567854 316574
rect 567234 280894 567854 316338
rect 567234 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 567854 280894
rect 567234 280574 567854 280658
rect 567234 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 567854 280574
rect 567234 244894 567854 280338
rect 567234 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 567854 244894
rect 567234 244574 567854 244658
rect 567234 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 567854 244574
rect 567234 208894 567854 244338
rect 567234 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 567854 208894
rect 567234 208574 567854 208658
rect 567234 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 567854 208574
rect 567234 172894 567854 208338
rect 567234 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 567854 172894
rect 567234 172574 567854 172658
rect 567234 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 567854 172574
rect 567234 136894 567854 172338
rect 567234 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 567854 136894
rect 567234 136574 567854 136658
rect 567234 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 567854 136574
rect 567234 100894 567854 136338
rect 567234 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 567854 100894
rect 567234 100574 567854 100658
rect 567234 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 567854 100574
rect 567234 64894 567854 100338
rect 567234 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 567854 64894
rect 567234 64574 567854 64658
rect 567234 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 567854 64574
rect 567234 28894 567854 64338
rect 567234 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 567854 28894
rect 567234 28574 567854 28658
rect 567234 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 567854 28574
rect 567234 -5146 567854 28338
rect 567234 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 567854 -5146
rect 567234 -5466 567854 -5382
rect 567234 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 567854 -5466
rect 567234 -5734 567854 -5702
rect 570954 680614 571574 711002
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 581514 706758 582134 707750
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 581514 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 582134 706758
rect 581514 706438 582134 706522
rect 581514 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 582134 706438
rect 570954 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 571574 680614
rect 570954 680294 571574 680378
rect 570954 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 571574 680294
rect 570954 644614 571574 680058
rect 570954 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 571574 644614
rect 570954 644294 571574 644378
rect 570954 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 571574 644294
rect 570954 608614 571574 644058
rect 570954 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 571574 608614
rect 570954 608294 571574 608378
rect 570954 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 571574 608294
rect 570954 572614 571574 608058
rect 570954 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 571574 572614
rect 570954 572294 571574 572378
rect 570954 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 571574 572294
rect 570954 536614 571574 572058
rect 570954 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 571574 536614
rect 570954 536294 571574 536378
rect 570954 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 571574 536294
rect 570954 500614 571574 536058
rect 570954 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 571574 500614
rect 570954 500294 571574 500378
rect 570954 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 571574 500294
rect 570954 464614 571574 500058
rect 570954 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 571574 464614
rect 570954 464294 571574 464378
rect 570954 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 571574 464294
rect 570954 428614 571574 464058
rect 570954 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 571574 428614
rect 570954 428294 571574 428378
rect 570954 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 571574 428294
rect 570954 392614 571574 428058
rect 570954 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 571574 392614
rect 570954 392294 571574 392378
rect 570954 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 571574 392294
rect 570954 356614 571574 392058
rect 570954 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 571574 356614
rect 570954 356294 571574 356378
rect 570954 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 571574 356294
rect 570954 320614 571574 356058
rect 570954 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 571574 320614
rect 570954 320294 571574 320378
rect 570954 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 571574 320294
rect 570954 284614 571574 320058
rect 570954 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 571574 284614
rect 570954 284294 571574 284378
rect 570954 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 571574 284294
rect 570954 248614 571574 284058
rect 570954 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 571574 248614
rect 570954 248294 571574 248378
rect 570954 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 571574 248294
rect 570954 212614 571574 248058
rect 570954 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 571574 212614
rect 570954 212294 571574 212378
rect 570954 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 571574 212294
rect 570954 176614 571574 212058
rect 570954 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 571574 176614
rect 570954 176294 571574 176378
rect 570954 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 571574 176294
rect 570954 140614 571574 176058
rect 570954 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 571574 140614
rect 570954 140294 571574 140378
rect 570954 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 571574 140294
rect 570954 104614 571574 140058
rect 570954 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 571574 104614
rect 570954 104294 571574 104378
rect 570954 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 571574 104294
rect 570954 68614 571574 104058
rect 570954 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 571574 68614
rect 570954 68294 571574 68378
rect 570954 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 571574 68294
rect 570954 32614 571574 68058
rect 570954 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 571574 32614
rect 570954 32294 571574 32378
rect 570954 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 571574 32294
rect 552954 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 553574 -6106
rect 552954 -6426 553574 -6342
rect 552954 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 553574 -6426
rect 552954 -7654 553574 -6662
rect 570954 -7066 571574 32058
rect 577794 704838 578414 705830
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -1894 578414 -902
rect 581514 691174 582134 706202
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -2266 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 669454 586890 705242
rect 586270 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect 586270 669134 586890 669218
rect 586270 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect 586270 633454 586890 668898
rect 586270 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect 586270 633134 586890 633218
rect 586270 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect 586270 597454 586890 632898
rect 586270 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect 586270 597134 586890 597218
rect 586270 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect 586270 561454 586890 596898
rect 586270 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect 586270 561134 586890 561218
rect 586270 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect 586270 525454 586890 560898
rect 586270 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect 586270 525134 586890 525218
rect 586270 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect 586270 489454 586890 524898
rect 586270 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect 586270 489134 586890 489218
rect 586270 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect 586270 453454 586890 488898
rect 586270 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect 586270 453134 586890 453218
rect 586270 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect 586270 417454 586890 452898
rect 586270 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect 586270 417134 586890 417218
rect 586270 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect 586270 381454 586890 416898
rect 586270 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect 586270 381134 586890 381218
rect 586270 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect 586270 345454 586890 380898
rect 586270 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect 586270 345134 586890 345218
rect 586270 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect 586270 309454 586890 344898
rect 586270 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect 586270 309134 586890 309218
rect 586270 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect 586270 273454 586890 308898
rect 586270 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect 586270 273134 586890 273218
rect 586270 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect 586270 237454 586890 272898
rect 586270 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect 586270 237134 586890 237218
rect 586270 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect 586270 201454 586890 236898
rect 586270 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect 586270 201134 586890 201218
rect 586270 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect 586270 165454 586890 200898
rect 586270 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect 586270 165134 586890 165218
rect 586270 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect 586270 129454 586890 164898
rect 586270 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect 586270 129134 586890 129218
rect 586270 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect 586270 93454 586890 128898
rect 586270 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect 586270 93134 586890 93218
rect 586270 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect 586270 57454 586890 92898
rect 586270 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect 586270 57134 586890 57218
rect 586270 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect 586270 21454 586890 56898
rect 586270 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect 586270 21134 586890 21218
rect 586270 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect 586270 -1306 586890 20898
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 691174 587850 706202
rect 587230 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 587850 691174
rect 587230 690854 587850 690938
rect 587230 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 587850 690854
rect 587230 655174 587850 690618
rect 587230 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 587850 655174
rect 587230 654854 587850 654938
rect 587230 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 587850 654854
rect 587230 619174 587850 654618
rect 587230 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 587850 619174
rect 587230 618854 587850 618938
rect 587230 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 587850 618854
rect 587230 583174 587850 618618
rect 587230 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 587850 583174
rect 587230 582854 587850 582938
rect 587230 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 587850 582854
rect 587230 547174 587850 582618
rect 587230 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 587850 547174
rect 587230 546854 587850 546938
rect 587230 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 587850 546854
rect 587230 511174 587850 546618
rect 587230 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 587850 511174
rect 587230 510854 587850 510938
rect 587230 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 587850 510854
rect 587230 475174 587850 510618
rect 587230 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 587850 475174
rect 587230 474854 587850 474938
rect 587230 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 587850 474854
rect 587230 439174 587850 474618
rect 587230 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 587850 439174
rect 587230 438854 587850 438938
rect 587230 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 587850 438854
rect 587230 403174 587850 438618
rect 587230 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 587850 403174
rect 587230 402854 587850 402938
rect 587230 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 587850 402854
rect 587230 367174 587850 402618
rect 587230 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 587850 367174
rect 587230 366854 587850 366938
rect 587230 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 587850 366854
rect 587230 331174 587850 366618
rect 587230 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 587850 331174
rect 587230 330854 587850 330938
rect 587230 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 587850 330854
rect 587230 295174 587850 330618
rect 587230 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 587850 295174
rect 587230 294854 587850 294938
rect 587230 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 587850 294854
rect 587230 259174 587850 294618
rect 587230 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 587850 259174
rect 587230 258854 587850 258938
rect 587230 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 587850 258854
rect 587230 223174 587850 258618
rect 587230 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 587850 223174
rect 587230 222854 587850 222938
rect 587230 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 587850 222854
rect 587230 187174 587850 222618
rect 587230 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 587850 187174
rect 587230 186854 587850 186938
rect 587230 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 587850 186854
rect 587230 151174 587850 186618
rect 587230 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 587850 151174
rect 587230 150854 587850 150938
rect 587230 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 587850 150854
rect 587230 115174 587850 150618
rect 587230 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 587850 115174
rect 587230 114854 587850 114938
rect 587230 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 587850 114854
rect 587230 79174 587850 114618
rect 587230 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 587850 79174
rect 587230 78854 587850 78938
rect 587230 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 587850 78854
rect 587230 43174 587850 78618
rect 587230 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 587850 43174
rect 587230 42854 587850 42938
rect 587230 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 587850 42854
rect 587230 7174 587850 42618
rect 587230 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 587850 7174
rect 587230 6854 587850 6938
rect 587230 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 587850 6854
rect 581514 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 582134 -2266
rect 581514 -2586 582134 -2502
rect 581514 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 582134 -2586
rect 581514 -3814 582134 -2822
rect 587230 -2266 587850 6618
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 673174 588810 707162
rect 588190 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect 588190 672854 588810 672938
rect 588190 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect 588190 637174 588810 672618
rect 588190 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect 588190 636854 588810 636938
rect 588190 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect 588190 601174 588810 636618
rect 588190 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect 588190 600854 588810 600938
rect 588190 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect 588190 565174 588810 600618
rect 588190 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect 588190 564854 588810 564938
rect 588190 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect 588190 529174 588810 564618
rect 588190 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect 588190 528854 588810 528938
rect 588190 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect 588190 493174 588810 528618
rect 588190 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect 588190 492854 588810 492938
rect 588190 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect 588190 457174 588810 492618
rect 588190 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect 588190 456854 588810 456938
rect 588190 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect 588190 421174 588810 456618
rect 588190 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect 588190 420854 588810 420938
rect 588190 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect 588190 385174 588810 420618
rect 588190 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect 588190 384854 588810 384938
rect 588190 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect 588190 349174 588810 384618
rect 588190 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect 588190 348854 588810 348938
rect 588190 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect 588190 313174 588810 348618
rect 588190 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect 588190 312854 588810 312938
rect 588190 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect 588190 277174 588810 312618
rect 588190 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect 588190 276854 588810 276938
rect 588190 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect 588190 241174 588810 276618
rect 588190 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect 588190 240854 588810 240938
rect 588190 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect 588190 205174 588810 240618
rect 588190 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect 588190 204854 588810 204938
rect 588190 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect 588190 169174 588810 204618
rect 588190 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect 588190 168854 588810 168938
rect 588190 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect 588190 133174 588810 168618
rect 588190 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect 588190 132854 588810 132938
rect 588190 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect 588190 97174 588810 132618
rect 588190 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect 588190 96854 588810 96938
rect 588190 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect 588190 61174 588810 96618
rect 588190 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect 588190 60854 588810 60938
rect 588190 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect 588190 25174 588810 60618
rect 588190 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect 588190 24854 588810 24938
rect 588190 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect 588190 -3226 588810 24618
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 694894 589770 708122
rect 589150 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 589770 694894
rect 589150 694574 589770 694658
rect 589150 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 589770 694574
rect 589150 658894 589770 694338
rect 589150 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 589770 658894
rect 589150 658574 589770 658658
rect 589150 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 589770 658574
rect 589150 622894 589770 658338
rect 589150 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 589770 622894
rect 589150 622574 589770 622658
rect 589150 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 589770 622574
rect 589150 586894 589770 622338
rect 589150 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 589770 586894
rect 589150 586574 589770 586658
rect 589150 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 589770 586574
rect 589150 550894 589770 586338
rect 589150 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 589770 550894
rect 589150 550574 589770 550658
rect 589150 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 589770 550574
rect 589150 514894 589770 550338
rect 589150 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 589770 514894
rect 589150 514574 589770 514658
rect 589150 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 589770 514574
rect 589150 478894 589770 514338
rect 589150 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 589770 478894
rect 589150 478574 589770 478658
rect 589150 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 589770 478574
rect 589150 442894 589770 478338
rect 589150 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 589770 442894
rect 589150 442574 589770 442658
rect 589150 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 589770 442574
rect 589150 406894 589770 442338
rect 589150 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 589770 406894
rect 589150 406574 589770 406658
rect 589150 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 589770 406574
rect 589150 370894 589770 406338
rect 589150 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 589770 370894
rect 589150 370574 589770 370658
rect 589150 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 589770 370574
rect 589150 334894 589770 370338
rect 589150 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 589770 334894
rect 589150 334574 589770 334658
rect 589150 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 589770 334574
rect 589150 298894 589770 334338
rect 589150 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 589770 298894
rect 589150 298574 589770 298658
rect 589150 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 589770 298574
rect 589150 262894 589770 298338
rect 589150 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 589770 262894
rect 589150 262574 589770 262658
rect 589150 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 589770 262574
rect 589150 226894 589770 262338
rect 589150 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 589770 226894
rect 589150 226574 589770 226658
rect 589150 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 589770 226574
rect 589150 190894 589770 226338
rect 589150 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 589770 190894
rect 589150 190574 589770 190658
rect 589150 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 589770 190574
rect 589150 154894 589770 190338
rect 589150 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 589770 154894
rect 589150 154574 589770 154658
rect 589150 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 589770 154574
rect 589150 118894 589770 154338
rect 589150 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 589770 118894
rect 589150 118574 589770 118658
rect 589150 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 589770 118574
rect 589150 82894 589770 118338
rect 589150 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 589770 82894
rect 589150 82574 589770 82658
rect 589150 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 589770 82574
rect 589150 46894 589770 82338
rect 589150 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 589770 46894
rect 589150 46574 589770 46658
rect 589150 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 589770 46574
rect 589150 10894 589770 46338
rect 589150 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 589770 10894
rect 589150 10574 589770 10658
rect 589150 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 589770 10574
rect 589150 -4186 589770 10338
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 676894 590730 709082
rect 590110 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect 590110 676574 590730 676658
rect 590110 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect 590110 640894 590730 676338
rect 590110 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect 590110 640574 590730 640658
rect 590110 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect 590110 604894 590730 640338
rect 590110 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect 590110 604574 590730 604658
rect 590110 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect 590110 568894 590730 604338
rect 590110 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect 590110 568574 590730 568658
rect 590110 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect 590110 532894 590730 568338
rect 590110 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect 590110 532574 590730 532658
rect 590110 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect 590110 496894 590730 532338
rect 590110 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect 590110 496574 590730 496658
rect 590110 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect 590110 460894 590730 496338
rect 590110 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect 590110 460574 590730 460658
rect 590110 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect 590110 424894 590730 460338
rect 590110 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect 590110 424574 590730 424658
rect 590110 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect 590110 388894 590730 424338
rect 590110 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect 590110 388574 590730 388658
rect 590110 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect 590110 352894 590730 388338
rect 590110 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect 590110 352574 590730 352658
rect 590110 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect 590110 316894 590730 352338
rect 590110 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect 590110 316574 590730 316658
rect 590110 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect 590110 280894 590730 316338
rect 590110 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect 590110 280574 590730 280658
rect 590110 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect 590110 244894 590730 280338
rect 590110 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect 590110 244574 590730 244658
rect 590110 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect 590110 208894 590730 244338
rect 590110 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect 590110 208574 590730 208658
rect 590110 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect 590110 172894 590730 208338
rect 590110 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect 590110 172574 590730 172658
rect 590110 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect 590110 136894 590730 172338
rect 590110 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect 590110 136574 590730 136658
rect 590110 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect 590110 100894 590730 136338
rect 590110 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect 590110 100574 590730 100658
rect 590110 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect 590110 64894 590730 100338
rect 590110 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect 590110 64574 590730 64658
rect 590110 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect 590110 28894 590730 64338
rect 590110 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect 590110 28574 590730 28658
rect 590110 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect 590110 -5146 590730 28338
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 698614 591690 710042
rect 591070 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 591690 698614
rect 591070 698294 591690 698378
rect 591070 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 591690 698294
rect 591070 662614 591690 698058
rect 591070 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 591690 662614
rect 591070 662294 591690 662378
rect 591070 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 591690 662294
rect 591070 626614 591690 662058
rect 591070 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 591690 626614
rect 591070 626294 591690 626378
rect 591070 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 591690 626294
rect 591070 590614 591690 626058
rect 591070 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 591690 590614
rect 591070 590294 591690 590378
rect 591070 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 591690 590294
rect 591070 554614 591690 590058
rect 591070 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 591690 554614
rect 591070 554294 591690 554378
rect 591070 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 591690 554294
rect 591070 518614 591690 554058
rect 591070 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 591690 518614
rect 591070 518294 591690 518378
rect 591070 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 591690 518294
rect 591070 482614 591690 518058
rect 591070 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 591690 482614
rect 591070 482294 591690 482378
rect 591070 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 591690 482294
rect 591070 446614 591690 482058
rect 591070 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 591690 446614
rect 591070 446294 591690 446378
rect 591070 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 591690 446294
rect 591070 410614 591690 446058
rect 591070 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 591690 410614
rect 591070 410294 591690 410378
rect 591070 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 591690 410294
rect 591070 374614 591690 410058
rect 591070 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 591690 374614
rect 591070 374294 591690 374378
rect 591070 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 591690 374294
rect 591070 338614 591690 374058
rect 591070 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 591690 338614
rect 591070 338294 591690 338378
rect 591070 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 591690 338294
rect 591070 302614 591690 338058
rect 591070 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 591690 302614
rect 591070 302294 591690 302378
rect 591070 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 591690 302294
rect 591070 266614 591690 302058
rect 591070 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 591690 266614
rect 591070 266294 591690 266378
rect 591070 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 591690 266294
rect 591070 230614 591690 266058
rect 591070 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 591690 230614
rect 591070 230294 591690 230378
rect 591070 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 591690 230294
rect 591070 194614 591690 230058
rect 591070 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 591690 194614
rect 591070 194294 591690 194378
rect 591070 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 591690 194294
rect 591070 158614 591690 194058
rect 591070 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 591690 158614
rect 591070 158294 591690 158378
rect 591070 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 591690 158294
rect 591070 122614 591690 158058
rect 591070 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 591690 122614
rect 591070 122294 591690 122378
rect 591070 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 591690 122294
rect 591070 86614 591690 122058
rect 591070 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 591690 86614
rect 591070 86294 591690 86378
rect 591070 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 591690 86294
rect 591070 50614 591690 86058
rect 591070 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 591690 50614
rect 591070 50294 591690 50378
rect 591070 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 591690 50294
rect 591070 14614 591690 50058
rect 591070 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 591690 14614
rect 591070 14294 591690 14378
rect 591070 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 591690 14294
rect 591070 -6106 591690 14058
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 680614 592650 711002
rect 592030 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect 592030 680294 592650 680378
rect 592030 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect 592030 644614 592650 680058
rect 592030 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect 592030 644294 592650 644378
rect 592030 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect 592030 608614 592650 644058
rect 592030 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect 592030 608294 592650 608378
rect 592030 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect 592030 572614 592650 608058
rect 592030 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect 592030 572294 592650 572378
rect 592030 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect 592030 536614 592650 572058
rect 592030 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect 592030 536294 592650 536378
rect 592030 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect 592030 500614 592650 536058
rect 592030 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect 592030 500294 592650 500378
rect 592030 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect 592030 464614 592650 500058
rect 592030 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect 592030 464294 592650 464378
rect 592030 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect 592030 428614 592650 464058
rect 592030 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect 592030 428294 592650 428378
rect 592030 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect 592030 392614 592650 428058
rect 592030 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect 592030 392294 592650 392378
rect 592030 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect 592030 356614 592650 392058
rect 592030 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect 592030 356294 592650 356378
rect 592030 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect 592030 320614 592650 356058
rect 592030 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect 592030 320294 592650 320378
rect 592030 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect 592030 284614 592650 320058
rect 592030 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect 592030 284294 592650 284378
rect 592030 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect 592030 248614 592650 284058
rect 592030 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect 592030 248294 592650 248378
rect 592030 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect 592030 212614 592650 248058
rect 592030 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect 592030 212294 592650 212378
rect 592030 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect 592030 176614 592650 212058
rect 592030 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect 592030 176294 592650 176378
rect 592030 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect 592030 140614 592650 176058
rect 592030 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect 592030 140294 592650 140378
rect 592030 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect 592030 104614 592650 140058
rect 592030 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect 592030 104294 592650 104378
rect 592030 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect 592030 68614 592650 104058
rect 592030 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect 592030 68294 592650 68378
rect 592030 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect 592030 32614 592650 68058
rect 592030 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect 592030 32294 592650 32378
rect 592030 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect 570954 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 571574 -7066
rect 570954 -7386 571574 -7302
rect 570954 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 571574 -7386
rect 570954 -7654 571574 -7622
rect 592030 -7066 592650 32058
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 680378 -8458 680614
rect -8374 680378 -8138 680614
rect -8694 680058 -8458 680294
rect -8374 680058 -8138 680294
rect -8694 644378 -8458 644614
rect -8374 644378 -8138 644614
rect -8694 644058 -8458 644294
rect -8374 644058 -8138 644294
rect -8694 608378 -8458 608614
rect -8374 608378 -8138 608614
rect -8694 608058 -8458 608294
rect -8374 608058 -8138 608294
rect -8694 572378 -8458 572614
rect -8374 572378 -8138 572614
rect -8694 572058 -8458 572294
rect -8374 572058 -8138 572294
rect -8694 536378 -8458 536614
rect -8374 536378 -8138 536614
rect -8694 536058 -8458 536294
rect -8374 536058 -8138 536294
rect -8694 500378 -8458 500614
rect -8374 500378 -8138 500614
rect -8694 500058 -8458 500294
rect -8374 500058 -8138 500294
rect -8694 464378 -8458 464614
rect -8374 464378 -8138 464614
rect -8694 464058 -8458 464294
rect -8374 464058 -8138 464294
rect -8694 428378 -8458 428614
rect -8374 428378 -8138 428614
rect -8694 428058 -8458 428294
rect -8374 428058 -8138 428294
rect -8694 392378 -8458 392614
rect -8374 392378 -8138 392614
rect -8694 392058 -8458 392294
rect -8374 392058 -8138 392294
rect -8694 356378 -8458 356614
rect -8374 356378 -8138 356614
rect -8694 356058 -8458 356294
rect -8374 356058 -8138 356294
rect -8694 320378 -8458 320614
rect -8374 320378 -8138 320614
rect -8694 320058 -8458 320294
rect -8374 320058 -8138 320294
rect -8694 284378 -8458 284614
rect -8374 284378 -8138 284614
rect -8694 284058 -8458 284294
rect -8374 284058 -8138 284294
rect -8694 248378 -8458 248614
rect -8374 248378 -8138 248614
rect -8694 248058 -8458 248294
rect -8374 248058 -8138 248294
rect -8694 212378 -8458 212614
rect -8374 212378 -8138 212614
rect -8694 212058 -8458 212294
rect -8374 212058 -8138 212294
rect -8694 176378 -8458 176614
rect -8374 176378 -8138 176614
rect -8694 176058 -8458 176294
rect -8374 176058 -8138 176294
rect -8694 140378 -8458 140614
rect -8374 140378 -8138 140614
rect -8694 140058 -8458 140294
rect -8374 140058 -8138 140294
rect -8694 104378 -8458 104614
rect -8374 104378 -8138 104614
rect -8694 104058 -8458 104294
rect -8374 104058 -8138 104294
rect -8694 68378 -8458 68614
rect -8374 68378 -8138 68614
rect -8694 68058 -8458 68294
rect -8374 68058 -8138 68294
rect -8694 32378 -8458 32614
rect -8374 32378 -8138 32614
rect -8694 32058 -8458 32294
rect -8374 32058 -8138 32294
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect 12986 710362 13222 710598
rect 13306 710362 13542 710598
rect 12986 710042 13222 710278
rect 13306 710042 13542 710278
rect -7734 698378 -7498 698614
rect -7414 698378 -7178 698614
rect -7734 698058 -7498 698294
rect -7414 698058 -7178 698294
rect -7734 662378 -7498 662614
rect -7414 662378 -7178 662614
rect -7734 662058 -7498 662294
rect -7414 662058 -7178 662294
rect -7734 626378 -7498 626614
rect -7414 626378 -7178 626614
rect -7734 626058 -7498 626294
rect -7414 626058 -7178 626294
rect -7734 590378 -7498 590614
rect -7414 590378 -7178 590614
rect -7734 590058 -7498 590294
rect -7414 590058 -7178 590294
rect -7734 554378 -7498 554614
rect -7414 554378 -7178 554614
rect -7734 554058 -7498 554294
rect -7414 554058 -7178 554294
rect -7734 518378 -7498 518614
rect -7414 518378 -7178 518614
rect -7734 518058 -7498 518294
rect -7414 518058 -7178 518294
rect -7734 482378 -7498 482614
rect -7414 482378 -7178 482614
rect -7734 482058 -7498 482294
rect -7414 482058 -7178 482294
rect -7734 446378 -7498 446614
rect -7414 446378 -7178 446614
rect -7734 446058 -7498 446294
rect -7414 446058 -7178 446294
rect -7734 410378 -7498 410614
rect -7414 410378 -7178 410614
rect -7734 410058 -7498 410294
rect -7414 410058 -7178 410294
rect -7734 374378 -7498 374614
rect -7414 374378 -7178 374614
rect -7734 374058 -7498 374294
rect -7414 374058 -7178 374294
rect -7734 338378 -7498 338614
rect -7414 338378 -7178 338614
rect -7734 338058 -7498 338294
rect -7414 338058 -7178 338294
rect -7734 302378 -7498 302614
rect -7414 302378 -7178 302614
rect -7734 302058 -7498 302294
rect -7414 302058 -7178 302294
rect -7734 266378 -7498 266614
rect -7414 266378 -7178 266614
rect -7734 266058 -7498 266294
rect -7414 266058 -7178 266294
rect -7734 230378 -7498 230614
rect -7414 230378 -7178 230614
rect -7734 230058 -7498 230294
rect -7414 230058 -7178 230294
rect -7734 194378 -7498 194614
rect -7414 194378 -7178 194614
rect -7734 194058 -7498 194294
rect -7414 194058 -7178 194294
rect -7734 158378 -7498 158614
rect -7414 158378 -7178 158614
rect -7734 158058 -7498 158294
rect -7414 158058 -7178 158294
rect -7734 122378 -7498 122614
rect -7414 122378 -7178 122614
rect -7734 122058 -7498 122294
rect -7414 122058 -7178 122294
rect -7734 86378 -7498 86614
rect -7414 86378 -7178 86614
rect -7734 86058 -7498 86294
rect -7414 86058 -7178 86294
rect -7734 50378 -7498 50614
rect -7414 50378 -7178 50614
rect -7734 50058 -7498 50294
rect -7414 50058 -7178 50294
rect -7734 14378 -7498 14614
rect -7414 14378 -7178 14614
rect -7734 14058 -7498 14294
rect -7414 14058 -7178 14294
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 676658 -6538 676894
rect -6454 676658 -6218 676894
rect -6774 676338 -6538 676574
rect -6454 676338 -6218 676574
rect -6774 640658 -6538 640894
rect -6454 640658 -6218 640894
rect -6774 640338 -6538 640574
rect -6454 640338 -6218 640574
rect -6774 604658 -6538 604894
rect -6454 604658 -6218 604894
rect -6774 604338 -6538 604574
rect -6454 604338 -6218 604574
rect -6774 568658 -6538 568894
rect -6454 568658 -6218 568894
rect -6774 568338 -6538 568574
rect -6454 568338 -6218 568574
rect -6774 532658 -6538 532894
rect -6454 532658 -6218 532894
rect -6774 532338 -6538 532574
rect -6454 532338 -6218 532574
rect -6774 496658 -6538 496894
rect -6454 496658 -6218 496894
rect -6774 496338 -6538 496574
rect -6454 496338 -6218 496574
rect -6774 460658 -6538 460894
rect -6454 460658 -6218 460894
rect -6774 460338 -6538 460574
rect -6454 460338 -6218 460574
rect -6774 424658 -6538 424894
rect -6454 424658 -6218 424894
rect -6774 424338 -6538 424574
rect -6454 424338 -6218 424574
rect -6774 388658 -6538 388894
rect -6454 388658 -6218 388894
rect -6774 388338 -6538 388574
rect -6454 388338 -6218 388574
rect -6774 352658 -6538 352894
rect -6454 352658 -6218 352894
rect -6774 352338 -6538 352574
rect -6454 352338 -6218 352574
rect -6774 316658 -6538 316894
rect -6454 316658 -6218 316894
rect -6774 316338 -6538 316574
rect -6454 316338 -6218 316574
rect -6774 280658 -6538 280894
rect -6454 280658 -6218 280894
rect -6774 280338 -6538 280574
rect -6454 280338 -6218 280574
rect -6774 244658 -6538 244894
rect -6454 244658 -6218 244894
rect -6774 244338 -6538 244574
rect -6454 244338 -6218 244574
rect -6774 208658 -6538 208894
rect -6454 208658 -6218 208894
rect -6774 208338 -6538 208574
rect -6454 208338 -6218 208574
rect -6774 172658 -6538 172894
rect -6454 172658 -6218 172894
rect -6774 172338 -6538 172574
rect -6454 172338 -6218 172574
rect -6774 136658 -6538 136894
rect -6454 136658 -6218 136894
rect -6774 136338 -6538 136574
rect -6454 136338 -6218 136574
rect -6774 100658 -6538 100894
rect -6454 100658 -6218 100894
rect -6774 100338 -6538 100574
rect -6454 100338 -6218 100574
rect -6774 64658 -6538 64894
rect -6454 64658 -6218 64894
rect -6774 64338 -6538 64574
rect -6454 64338 -6218 64574
rect -6774 28658 -6538 28894
rect -6454 28658 -6218 28894
rect -6774 28338 -6538 28574
rect -6454 28338 -6218 28574
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect 9266 708442 9502 708678
rect 9586 708442 9822 708678
rect 9266 708122 9502 708358
rect 9586 708122 9822 708358
rect -5814 694658 -5578 694894
rect -5494 694658 -5258 694894
rect -5814 694338 -5578 694574
rect -5494 694338 -5258 694574
rect -5814 658658 -5578 658894
rect -5494 658658 -5258 658894
rect -5814 658338 -5578 658574
rect -5494 658338 -5258 658574
rect -5814 622658 -5578 622894
rect -5494 622658 -5258 622894
rect -5814 622338 -5578 622574
rect -5494 622338 -5258 622574
rect -5814 586658 -5578 586894
rect -5494 586658 -5258 586894
rect -5814 586338 -5578 586574
rect -5494 586338 -5258 586574
rect -5814 550658 -5578 550894
rect -5494 550658 -5258 550894
rect -5814 550338 -5578 550574
rect -5494 550338 -5258 550574
rect -5814 514658 -5578 514894
rect -5494 514658 -5258 514894
rect -5814 514338 -5578 514574
rect -5494 514338 -5258 514574
rect -5814 478658 -5578 478894
rect -5494 478658 -5258 478894
rect -5814 478338 -5578 478574
rect -5494 478338 -5258 478574
rect -5814 442658 -5578 442894
rect -5494 442658 -5258 442894
rect -5814 442338 -5578 442574
rect -5494 442338 -5258 442574
rect -5814 406658 -5578 406894
rect -5494 406658 -5258 406894
rect -5814 406338 -5578 406574
rect -5494 406338 -5258 406574
rect -5814 370658 -5578 370894
rect -5494 370658 -5258 370894
rect -5814 370338 -5578 370574
rect -5494 370338 -5258 370574
rect -5814 334658 -5578 334894
rect -5494 334658 -5258 334894
rect -5814 334338 -5578 334574
rect -5494 334338 -5258 334574
rect -5814 298658 -5578 298894
rect -5494 298658 -5258 298894
rect -5814 298338 -5578 298574
rect -5494 298338 -5258 298574
rect -5814 262658 -5578 262894
rect -5494 262658 -5258 262894
rect -5814 262338 -5578 262574
rect -5494 262338 -5258 262574
rect -5814 226658 -5578 226894
rect -5494 226658 -5258 226894
rect -5814 226338 -5578 226574
rect -5494 226338 -5258 226574
rect -5814 190658 -5578 190894
rect -5494 190658 -5258 190894
rect -5814 190338 -5578 190574
rect -5494 190338 -5258 190574
rect -5814 154658 -5578 154894
rect -5494 154658 -5258 154894
rect -5814 154338 -5578 154574
rect -5494 154338 -5258 154574
rect -5814 118658 -5578 118894
rect -5494 118658 -5258 118894
rect -5814 118338 -5578 118574
rect -5494 118338 -5258 118574
rect -5814 82658 -5578 82894
rect -5494 82658 -5258 82894
rect -5814 82338 -5578 82574
rect -5494 82338 -5258 82574
rect -5814 46658 -5578 46894
rect -5494 46658 -5258 46894
rect -5814 46338 -5578 46574
rect -5494 46338 -5258 46574
rect -5814 10658 -5578 10894
rect -5494 10658 -5258 10894
rect -5814 10338 -5578 10574
rect -5494 10338 -5258 10574
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 672938 -4618 673174
rect -4534 672938 -4298 673174
rect -4854 672618 -4618 672854
rect -4534 672618 -4298 672854
rect -4854 636938 -4618 637174
rect -4534 636938 -4298 637174
rect -4854 636618 -4618 636854
rect -4534 636618 -4298 636854
rect -4854 600938 -4618 601174
rect -4534 600938 -4298 601174
rect -4854 600618 -4618 600854
rect -4534 600618 -4298 600854
rect -4854 564938 -4618 565174
rect -4534 564938 -4298 565174
rect -4854 564618 -4618 564854
rect -4534 564618 -4298 564854
rect -4854 528938 -4618 529174
rect -4534 528938 -4298 529174
rect -4854 528618 -4618 528854
rect -4534 528618 -4298 528854
rect -4854 492938 -4618 493174
rect -4534 492938 -4298 493174
rect -4854 492618 -4618 492854
rect -4534 492618 -4298 492854
rect -4854 456938 -4618 457174
rect -4534 456938 -4298 457174
rect -4854 456618 -4618 456854
rect -4534 456618 -4298 456854
rect -4854 420938 -4618 421174
rect -4534 420938 -4298 421174
rect -4854 420618 -4618 420854
rect -4534 420618 -4298 420854
rect -4854 384938 -4618 385174
rect -4534 384938 -4298 385174
rect -4854 384618 -4618 384854
rect -4534 384618 -4298 384854
rect -4854 348938 -4618 349174
rect -4534 348938 -4298 349174
rect -4854 348618 -4618 348854
rect -4534 348618 -4298 348854
rect -4854 312938 -4618 313174
rect -4534 312938 -4298 313174
rect -4854 312618 -4618 312854
rect -4534 312618 -4298 312854
rect -4854 276938 -4618 277174
rect -4534 276938 -4298 277174
rect -4854 276618 -4618 276854
rect -4534 276618 -4298 276854
rect -4854 240938 -4618 241174
rect -4534 240938 -4298 241174
rect -4854 240618 -4618 240854
rect -4534 240618 -4298 240854
rect -4854 204938 -4618 205174
rect -4534 204938 -4298 205174
rect -4854 204618 -4618 204854
rect -4534 204618 -4298 204854
rect -4854 168938 -4618 169174
rect -4534 168938 -4298 169174
rect -4854 168618 -4618 168854
rect -4534 168618 -4298 168854
rect -4854 132938 -4618 133174
rect -4534 132938 -4298 133174
rect -4854 132618 -4618 132854
rect -4534 132618 -4298 132854
rect -4854 96938 -4618 97174
rect -4534 96938 -4298 97174
rect -4854 96618 -4618 96854
rect -4534 96618 -4298 96854
rect -4854 60938 -4618 61174
rect -4534 60938 -4298 61174
rect -4854 60618 -4618 60854
rect -4534 60618 -4298 60854
rect -4854 24938 -4618 25174
rect -4534 24938 -4298 25174
rect -4854 24618 -4618 24854
rect -4534 24618 -4298 24854
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect 5546 706522 5782 706758
rect 5866 706522 6102 706758
rect 5546 706202 5782 706438
rect 5866 706202 6102 706438
rect -3894 690938 -3658 691174
rect -3574 690938 -3338 691174
rect -3894 690618 -3658 690854
rect -3574 690618 -3338 690854
rect -3894 654938 -3658 655174
rect -3574 654938 -3338 655174
rect -3894 654618 -3658 654854
rect -3574 654618 -3338 654854
rect -3894 618938 -3658 619174
rect -3574 618938 -3338 619174
rect -3894 618618 -3658 618854
rect -3574 618618 -3338 618854
rect -3894 582938 -3658 583174
rect -3574 582938 -3338 583174
rect -3894 582618 -3658 582854
rect -3574 582618 -3338 582854
rect -3894 546938 -3658 547174
rect -3574 546938 -3338 547174
rect -3894 546618 -3658 546854
rect -3574 546618 -3338 546854
rect -3894 510938 -3658 511174
rect -3574 510938 -3338 511174
rect -3894 510618 -3658 510854
rect -3574 510618 -3338 510854
rect -3894 474938 -3658 475174
rect -3574 474938 -3338 475174
rect -3894 474618 -3658 474854
rect -3574 474618 -3338 474854
rect -3894 438938 -3658 439174
rect -3574 438938 -3338 439174
rect -3894 438618 -3658 438854
rect -3574 438618 -3338 438854
rect -3894 402938 -3658 403174
rect -3574 402938 -3338 403174
rect -3894 402618 -3658 402854
rect -3574 402618 -3338 402854
rect -3894 366938 -3658 367174
rect -3574 366938 -3338 367174
rect -3894 366618 -3658 366854
rect -3574 366618 -3338 366854
rect -3894 330938 -3658 331174
rect -3574 330938 -3338 331174
rect -3894 330618 -3658 330854
rect -3574 330618 -3338 330854
rect -3894 294938 -3658 295174
rect -3574 294938 -3338 295174
rect -3894 294618 -3658 294854
rect -3574 294618 -3338 294854
rect -3894 258938 -3658 259174
rect -3574 258938 -3338 259174
rect -3894 258618 -3658 258854
rect -3574 258618 -3338 258854
rect -3894 222938 -3658 223174
rect -3574 222938 -3338 223174
rect -3894 222618 -3658 222854
rect -3574 222618 -3338 222854
rect -3894 186938 -3658 187174
rect -3574 186938 -3338 187174
rect -3894 186618 -3658 186854
rect -3574 186618 -3338 186854
rect -3894 150938 -3658 151174
rect -3574 150938 -3338 151174
rect -3894 150618 -3658 150854
rect -3574 150618 -3338 150854
rect -3894 114938 -3658 115174
rect -3574 114938 -3338 115174
rect -3894 114618 -3658 114854
rect -3574 114618 -3338 114854
rect -3894 78938 -3658 79174
rect -3574 78938 -3338 79174
rect -3894 78618 -3658 78854
rect -3574 78618 -3338 78854
rect -3894 42938 -3658 43174
rect -3574 42938 -3338 43174
rect -3894 42618 -3658 42854
rect -3574 42618 -3338 42854
rect -3894 6938 -3658 7174
rect -3574 6938 -3338 7174
rect -3894 6618 -3658 6854
rect -3574 6618 -3338 6854
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 669218 -2698 669454
rect -2614 669218 -2378 669454
rect -2934 668898 -2698 669134
rect -2614 668898 -2378 669134
rect -2934 633218 -2698 633454
rect -2614 633218 -2378 633454
rect -2934 632898 -2698 633134
rect -2614 632898 -2378 633134
rect -2934 597218 -2698 597454
rect -2614 597218 -2378 597454
rect -2934 596898 -2698 597134
rect -2614 596898 -2378 597134
rect -2934 561218 -2698 561454
rect -2614 561218 -2378 561454
rect -2934 560898 -2698 561134
rect -2614 560898 -2378 561134
rect -2934 525218 -2698 525454
rect -2614 525218 -2378 525454
rect -2934 524898 -2698 525134
rect -2614 524898 -2378 525134
rect -2934 489218 -2698 489454
rect -2614 489218 -2378 489454
rect -2934 488898 -2698 489134
rect -2614 488898 -2378 489134
rect -2934 453218 -2698 453454
rect -2614 453218 -2378 453454
rect -2934 452898 -2698 453134
rect -2614 452898 -2378 453134
rect -2934 417218 -2698 417454
rect -2614 417218 -2378 417454
rect -2934 416898 -2698 417134
rect -2614 416898 -2378 417134
rect -2934 381218 -2698 381454
rect -2614 381218 -2378 381454
rect -2934 380898 -2698 381134
rect -2614 380898 -2378 381134
rect -2934 345218 -2698 345454
rect -2614 345218 -2378 345454
rect -2934 344898 -2698 345134
rect -2614 344898 -2378 345134
rect -2934 309218 -2698 309454
rect -2614 309218 -2378 309454
rect -2934 308898 -2698 309134
rect -2614 308898 -2378 309134
rect -2934 273218 -2698 273454
rect -2614 273218 -2378 273454
rect -2934 272898 -2698 273134
rect -2614 272898 -2378 273134
rect -2934 237218 -2698 237454
rect -2614 237218 -2378 237454
rect -2934 236898 -2698 237134
rect -2614 236898 -2378 237134
rect -2934 201218 -2698 201454
rect -2614 201218 -2378 201454
rect -2934 200898 -2698 201134
rect -2614 200898 -2378 201134
rect -2934 165218 -2698 165454
rect -2614 165218 -2378 165454
rect -2934 164898 -2698 165134
rect -2614 164898 -2378 165134
rect -2934 129218 -2698 129454
rect -2614 129218 -2378 129454
rect -2934 128898 -2698 129134
rect -2614 128898 -2378 129134
rect -2934 93218 -2698 93454
rect -2614 93218 -2378 93454
rect -2934 92898 -2698 93134
rect -2614 92898 -2378 93134
rect -2934 57218 -2698 57454
rect -2614 57218 -2378 57454
rect -2934 56898 -2698 57134
rect -2614 56898 -2378 57134
rect -2934 21218 -2698 21454
rect -2614 21218 -2378 21454
rect -2934 20898 -2698 21134
rect -2614 20898 -2378 21134
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect 5546 -2502 5782 -2266
rect 5866 -2502 6102 -2266
rect 5546 -2822 5782 -2586
rect 5866 -2822 6102 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect 9266 694658 9502 694894
rect 9586 694658 9822 694894
rect 9266 694338 9502 694574
rect 9586 694338 9822 694574
rect 9266 658658 9502 658894
rect 9586 658658 9822 658894
rect 9266 658338 9502 658574
rect 9586 658338 9822 658574
rect 9266 622658 9502 622894
rect 9586 622658 9822 622894
rect 9266 622338 9502 622574
rect 9586 622338 9822 622574
rect 9266 586658 9502 586894
rect 9586 586658 9822 586894
rect 9266 586338 9502 586574
rect 9586 586338 9822 586574
rect 9266 550658 9502 550894
rect 9586 550658 9822 550894
rect 9266 550338 9502 550574
rect 9586 550338 9822 550574
rect 9266 514658 9502 514894
rect 9586 514658 9822 514894
rect 9266 514338 9502 514574
rect 9586 514338 9822 514574
rect 9266 478658 9502 478894
rect 9586 478658 9822 478894
rect 9266 478338 9502 478574
rect 9586 478338 9822 478574
rect 9266 442658 9502 442894
rect 9586 442658 9822 442894
rect 9266 442338 9502 442574
rect 9586 442338 9822 442574
rect 9266 406658 9502 406894
rect 9586 406658 9822 406894
rect 9266 406338 9502 406574
rect 9586 406338 9822 406574
rect 9266 370658 9502 370894
rect 9586 370658 9822 370894
rect 9266 370338 9502 370574
rect 9586 370338 9822 370574
rect 9266 334658 9502 334894
rect 9586 334658 9822 334894
rect 9266 334338 9502 334574
rect 9586 334338 9822 334574
rect 9266 298658 9502 298894
rect 9586 298658 9822 298894
rect 9266 298338 9502 298574
rect 9586 298338 9822 298574
rect 9266 262658 9502 262894
rect 9586 262658 9822 262894
rect 9266 262338 9502 262574
rect 9586 262338 9822 262574
rect 9266 226658 9502 226894
rect 9586 226658 9822 226894
rect 9266 226338 9502 226574
rect 9586 226338 9822 226574
rect 9266 190658 9502 190894
rect 9586 190658 9822 190894
rect 9266 190338 9502 190574
rect 9586 190338 9822 190574
rect 9266 154658 9502 154894
rect 9586 154658 9822 154894
rect 9266 154338 9502 154574
rect 9586 154338 9822 154574
rect 9266 118658 9502 118894
rect 9586 118658 9822 118894
rect 9266 118338 9502 118574
rect 9586 118338 9822 118574
rect 9266 82658 9502 82894
rect 9586 82658 9822 82894
rect 9266 82338 9502 82574
rect 9586 82338 9822 82574
rect 9266 46658 9502 46894
rect 9586 46658 9822 46894
rect 9266 46338 9502 46574
rect 9586 46338 9822 46574
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect 9266 -4422 9502 -4186
rect 9586 -4422 9822 -4186
rect 9266 -4742 9502 -4506
rect 9586 -4742 9822 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect 30986 711322 31222 711558
rect 31306 711322 31542 711558
rect 30986 711002 31222 711238
rect 31306 711002 31542 711238
rect 27266 709402 27502 709638
rect 27586 709402 27822 709638
rect 27266 709082 27502 709318
rect 27586 709082 27822 709318
rect 23546 707482 23782 707718
rect 23866 707482 24102 707718
rect 23546 707162 23782 707398
rect 23866 707162 24102 707398
rect 12986 698378 13222 698614
rect 13306 698378 13542 698614
rect 12986 698058 13222 698294
rect 13306 698058 13542 698294
rect 12986 662378 13222 662614
rect 13306 662378 13542 662614
rect 12986 662058 13222 662294
rect 13306 662058 13542 662294
rect 12986 626378 13222 626614
rect 13306 626378 13542 626614
rect 12986 626058 13222 626294
rect 13306 626058 13542 626294
rect 12986 590378 13222 590614
rect 13306 590378 13542 590614
rect 12986 590058 13222 590294
rect 13306 590058 13542 590294
rect 12986 554378 13222 554614
rect 13306 554378 13542 554614
rect 12986 554058 13222 554294
rect 13306 554058 13542 554294
rect 12986 518378 13222 518614
rect 13306 518378 13542 518614
rect 12986 518058 13222 518294
rect 13306 518058 13542 518294
rect 12986 482378 13222 482614
rect 13306 482378 13542 482614
rect 12986 482058 13222 482294
rect 13306 482058 13542 482294
rect 12986 446378 13222 446614
rect 13306 446378 13542 446614
rect 12986 446058 13222 446294
rect 13306 446058 13542 446294
rect 12986 410378 13222 410614
rect 13306 410378 13542 410614
rect 12986 410058 13222 410294
rect 13306 410058 13542 410294
rect 12986 374378 13222 374614
rect 13306 374378 13542 374614
rect 12986 374058 13222 374294
rect 13306 374058 13542 374294
rect 12986 338378 13222 338614
rect 13306 338378 13542 338614
rect 12986 338058 13222 338294
rect 13306 338058 13542 338294
rect 12986 302378 13222 302614
rect 13306 302378 13542 302614
rect 12986 302058 13222 302294
rect 13306 302058 13542 302294
rect 12986 266378 13222 266614
rect 13306 266378 13542 266614
rect 12986 266058 13222 266294
rect 13306 266058 13542 266294
rect 12986 230378 13222 230614
rect 13306 230378 13542 230614
rect 12986 230058 13222 230294
rect 13306 230058 13542 230294
rect 12986 194378 13222 194614
rect 13306 194378 13542 194614
rect 12986 194058 13222 194294
rect 13306 194058 13542 194294
rect 12986 158378 13222 158614
rect 13306 158378 13542 158614
rect 12986 158058 13222 158294
rect 13306 158058 13542 158294
rect 12986 122378 13222 122614
rect 13306 122378 13542 122614
rect 12986 122058 13222 122294
rect 13306 122058 13542 122294
rect 12986 86378 13222 86614
rect 13306 86378 13542 86614
rect 12986 86058 13222 86294
rect 13306 86058 13542 86294
rect 12986 50378 13222 50614
rect 13306 50378 13542 50614
rect 12986 50058 13222 50294
rect 13306 50058 13542 50294
rect 12986 14378 13222 14614
rect 13306 14378 13542 14614
rect 12986 14058 13222 14294
rect 13306 14058 13542 14294
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect 19826 705562 20062 705798
rect 20146 705562 20382 705798
rect 19826 705242 20062 705478
rect 20146 705242 20382 705478
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -1542 20062 -1306
rect 20146 -1542 20382 -1306
rect 19826 -1862 20062 -1626
rect 20146 -1862 20382 -1626
rect 23546 672938 23782 673174
rect 23866 672938 24102 673174
rect 23546 672618 23782 672854
rect 23866 672618 24102 672854
rect 23546 636938 23782 637174
rect 23866 636938 24102 637174
rect 23546 636618 23782 636854
rect 23866 636618 24102 636854
rect 23546 600938 23782 601174
rect 23866 600938 24102 601174
rect 23546 600618 23782 600854
rect 23866 600618 24102 600854
rect 23546 564938 23782 565174
rect 23866 564938 24102 565174
rect 23546 564618 23782 564854
rect 23866 564618 24102 564854
rect 23546 528938 23782 529174
rect 23866 528938 24102 529174
rect 23546 528618 23782 528854
rect 23866 528618 24102 528854
rect 23546 492938 23782 493174
rect 23866 492938 24102 493174
rect 23546 492618 23782 492854
rect 23866 492618 24102 492854
rect 23546 456938 23782 457174
rect 23866 456938 24102 457174
rect 23546 456618 23782 456854
rect 23866 456618 24102 456854
rect 23546 420938 23782 421174
rect 23866 420938 24102 421174
rect 23546 420618 23782 420854
rect 23866 420618 24102 420854
rect 23546 384938 23782 385174
rect 23866 384938 24102 385174
rect 23546 384618 23782 384854
rect 23866 384618 24102 384854
rect 23546 348938 23782 349174
rect 23866 348938 24102 349174
rect 23546 348618 23782 348854
rect 23866 348618 24102 348854
rect 23546 312938 23782 313174
rect 23866 312938 24102 313174
rect 23546 312618 23782 312854
rect 23866 312618 24102 312854
rect 23546 276938 23782 277174
rect 23866 276938 24102 277174
rect 23546 276618 23782 276854
rect 23866 276618 24102 276854
rect 23546 240938 23782 241174
rect 23866 240938 24102 241174
rect 23546 240618 23782 240854
rect 23866 240618 24102 240854
rect 23546 204938 23782 205174
rect 23866 204938 24102 205174
rect 23546 204618 23782 204854
rect 23866 204618 24102 204854
rect 23546 168938 23782 169174
rect 23866 168938 24102 169174
rect 23546 168618 23782 168854
rect 23866 168618 24102 168854
rect 23546 132938 23782 133174
rect 23866 132938 24102 133174
rect 23546 132618 23782 132854
rect 23866 132618 24102 132854
rect 23546 96938 23782 97174
rect 23866 96938 24102 97174
rect 23546 96618 23782 96854
rect 23866 96618 24102 96854
rect 23546 60938 23782 61174
rect 23866 60938 24102 61174
rect 23546 60618 23782 60854
rect 23866 60618 24102 60854
rect 23546 24938 23782 25174
rect 23866 24938 24102 25174
rect 23546 24618 23782 24854
rect 23866 24618 24102 24854
rect 23546 -3462 23782 -3226
rect 23866 -3462 24102 -3226
rect 23546 -3782 23782 -3546
rect 23866 -3782 24102 -3546
rect 27266 676658 27502 676894
rect 27586 676658 27822 676894
rect 27266 676338 27502 676574
rect 27586 676338 27822 676574
rect 27266 640658 27502 640894
rect 27586 640658 27822 640894
rect 27266 640338 27502 640574
rect 27586 640338 27822 640574
rect 27266 604658 27502 604894
rect 27586 604658 27822 604894
rect 27266 604338 27502 604574
rect 27586 604338 27822 604574
rect 27266 568658 27502 568894
rect 27586 568658 27822 568894
rect 27266 568338 27502 568574
rect 27586 568338 27822 568574
rect 27266 532658 27502 532894
rect 27586 532658 27822 532894
rect 27266 532338 27502 532574
rect 27586 532338 27822 532574
rect 27266 496658 27502 496894
rect 27586 496658 27822 496894
rect 27266 496338 27502 496574
rect 27586 496338 27822 496574
rect 27266 460658 27502 460894
rect 27586 460658 27822 460894
rect 27266 460338 27502 460574
rect 27586 460338 27822 460574
rect 27266 424658 27502 424894
rect 27586 424658 27822 424894
rect 27266 424338 27502 424574
rect 27586 424338 27822 424574
rect 27266 388658 27502 388894
rect 27586 388658 27822 388894
rect 27266 388338 27502 388574
rect 27586 388338 27822 388574
rect 27266 352658 27502 352894
rect 27586 352658 27822 352894
rect 27266 352338 27502 352574
rect 27586 352338 27822 352574
rect 27266 316658 27502 316894
rect 27586 316658 27822 316894
rect 27266 316338 27502 316574
rect 27586 316338 27822 316574
rect 27266 280658 27502 280894
rect 27586 280658 27822 280894
rect 27266 280338 27502 280574
rect 27586 280338 27822 280574
rect 27266 244658 27502 244894
rect 27586 244658 27822 244894
rect 27266 244338 27502 244574
rect 27586 244338 27822 244574
rect 27266 208658 27502 208894
rect 27586 208658 27822 208894
rect 27266 208338 27502 208574
rect 27586 208338 27822 208574
rect 27266 172658 27502 172894
rect 27586 172658 27822 172894
rect 27266 172338 27502 172574
rect 27586 172338 27822 172574
rect 27266 136658 27502 136894
rect 27586 136658 27822 136894
rect 27266 136338 27502 136574
rect 27586 136338 27822 136574
rect 27266 100658 27502 100894
rect 27586 100658 27822 100894
rect 27266 100338 27502 100574
rect 27586 100338 27822 100574
rect 27266 64658 27502 64894
rect 27586 64658 27822 64894
rect 27266 64338 27502 64574
rect 27586 64338 27822 64574
rect 27266 28658 27502 28894
rect 27586 28658 27822 28894
rect 27266 28338 27502 28574
rect 27586 28338 27822 28574
rect 27266 -5382 27502 -5146
rect 27586 -5382 27822 -5146
rect 27266 -5702 27502 -5466
rect 27586 -5702 27822 -5466
rect 48986 710362 49222 710598
rect 49306 710362 49542 710598
rect 48986 710042 49222 710278
rect 49306 710042 49542 710278
rect 45266 708442 45502 708678
rect 45586 708442 45822 708678
rect 45266 708122 45502 708358
rect 45586 708122 45822 708358
rect 41546 706522 41782 706758
rect 41866 706522 42102 706758
rect 41546 706202 41782 706438
rect 41866 706202 42102 706438
rect 30986 680378 31222 680614
rect 31306 680378 31542 680614
rect 30986 680058 31222 680294
rect 31306 680058 31542 680294
rect 30986 644378 31222 644614
rect 31306 644378 31542 644614
rect 30986 644058 31222 644294
rect 31306 644058 31542 644294
rect 30986 608378 31222 608614
rect 31306 608378 31542 608614
rect 30986 608058 31222 608294
rect 31306 608058 31542 608294
rect 30986 572378 31222 572614
rect 31306 572378 31542 572614
rect 30986 572058 31222 572294
rect 31306 572058 31542 572294
rect 30986 536378 31222 536614
rect 31306 536378 31542 536614
rect 30986 536058 31222 536294
rect 31306 536058 31542 536294
rect 30986 500378 31222 500614
rect 31306 500378 31542 500614
rect 30986 500058 31222 500294
rect 31306 500058 31542 500294
rect 30986 464378 31222 464614
rect 31306 464378 31542 464614
rect 30986 464058 31222 464294
rect 31306 464058 31542 464294
rect 30986 428378 31222 428614
rect 31306 428378 31542 428614
rect 30986 428058 31222 428294
rect 31306 428058 31542 428294
rect 30986 392378 31222 392614
rect 31306 392378 31542 392614
rect 30986 392058 31222 392294
rect 31306 392058 31542 392294
rect 30986 356378 31222 356614
rect 31306 356378 31542 356614
rect 30986 356058 31222 356294
rect 31306 356058 31542 356294
rect 30986 320378 31222 320614
rect 31306 320378 31542 320614
rect 30986 320058 31222 320294
rect 31306 320058 31542 320294
rect 30986 284378 31222 284614
rect 31306 284378 31542 284614
rect 30986 284058 31222 284294
rect 31306 284058 31542 284294
rect 30986 248378 31222 248614
rect 31306 248378 31542 248614
rect 30986 248058 31222 248294
rect 31306 248058 31542 248294
rect 30986 212378 31222 212614
rect 31306 212378 31542 212614
rect 30986 212058 31222 212294
rect 31306 212058 31542 212294
rect 30986 176378 31222 176614
rect 31306 176378 31542 176614
rect 30986 176058 31222 176294
rect 31306 176058 31542 176294
rect 30986 140378 31222 140614
rect 31306 140378 31542 140614
rect 30986 140058 31222 140294
rect 31306 140058 31542 140294
rect 30986 104378 31222 104614
rect 31306 104378 31542 104614
rect 30986 104058 31222 104294
rect 31306 104058 31542 104294
rect 30986 68378 31222 68614
rect 31306 68378 31542 68614
rect 30986 68058 31222 68294
rect 31306 68058 31542 68294
rect 30986 32378 31222 32614
rect 31306 32378 31542 32614
rect 30986 32058 31222 32294
rect 31306 32058 31542 32294
rect 12986 -6342 13222 -6106
rect 13306 -6342 13542 -6106
rect 12986 -6662 13222 -6426
rect 13306 -6662 13542 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 41546 654938 41782 655174
rect 41866 654938 42102 655174
rect 41546 654618 41782 654854
rect 41866 654618 42102 654854
rect 41546 618938 41782 619174
rect 41866 618938 42102 619174
rect 41546 618618 41782 618854
rect 41866 618618 42102 618854
rect 41546 582938 41782 583174
rect 41866 582938 42102 583174
rect 41546 582618 41782 582854
rect 41866 582618 42102 582854
rect 41546 546938 41782 547174
rect 41866 546938 42102 547174
rect 41546 546618 41782 546854
rect 41866 546618 42102 546854
rect 41546 510938 41782 511174
rect 41866 510938 42102 511174
rect 41546 510618 41782 510854
rect 41866 510618 42102 510854
rect 41546 474938 41782 475174
rect 41866 474938 42102 475174
rect 41546 474618 41782 474854
rect 41866 474618 42102 474854
rect 41546 438938 41782 439174
rect 41866 438938 42102 439174
rect 41546 438618 41782 438854
rect 41866 438618 42102 438854
rect 41546 402938 41782 403174
rect 41866 402938 42102 403174
rect 41546 402618 41782 402854
rect 41866 402618 42102 402854
rect 41546 366938 41782 367174
rect 41866 366938 42102 367174
rect 41546 366618 41782 366854
rect 41866 366618 42102 366854
rect 41546 330938 41782 331174
rect 41866 330938 42102 331174
rect 41546 330618 41782 330854
rect 41866 330618 42102 330854
rect 41546 294938 41782 295174
rect 41866 294938 42102 295174
rect 41546 294618 41782 294854
rect 41866 294618 42102 294854
rect 41546 258938 41782 259174
rect 41866 258938 42102 259174
rect 41546 258618 41782 258854
rect 41866 258618 42102 258854
rect 41546 222938 41782 223174
rect 41866 222938 42102 223174
rect 41546 222618 41782 222854
rect 41866 222618 42102 222854
rect 41546 186938 41782 187174
rect 41866 186938 42102 187174
rect 41546 186618 41782 186854
rect 41866 186618 42102 186854
rect 41546 150938 41782 151174
rect 41866 150938 42102 151174
rect 41546 150618 41782 150854
rect 41866 150618 42102 150854
rect 41546 114938 41782 115174
rect 41866 114938 42102 115174
rect 41546 114618 41782 114854
rect 41866 114618 42102 114854
rect 41546 78938 41782 79174
rect 41866 78938 42102 79174
rect 41546 78618 41782 78854
rect 41866 78618 42102 78854
rect 41546 42938 41782 43174
rect 41866 42938 42102 43174
rect 41546 42618 41782 42854
rect 41866 42618 42102 42854
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 41546 -2502 41782 -2266
rect 41866 -2502 42102 -2266
rect 41546 -2822 41782 -2586
rect 41866 -2822 42102 -2586
rect 45266 694658 45502 694894
rect 45586 694658 45822 694894
rect 45266 694338 45502 694574
rect 45586 694338 45822 694574
rect 45266 658658 45502 658894
rect 45586 658658 45822 658894
rect 45266 658338 45502 658574
rect 45586 658338 45822 658574
rect 45266 622658 45502 622894
rect 45586 622658 45822 622894
rect 45266 622338 45502 622574
rect 45586 622338 45822 622574
rect 45266 586658 45502 586894
rect 45586 586658 45822 586894
rect 45266 586338 45502 586574
rect 45586 586338 45822 586574
rect 45266 550658 45502 550894
rect 45586 550658 45822 550894
rect 45266 550338 45502 550574
rect 45586 550338 45822 550574
rect 45266 514658 45502 514894
rect 45586 514658 45822 514894
rect 45266 514338 45502 514574
rect 45586 514338 45822 514574
rect 45266 478658 45502 478894
rect 45586 478658 45822 478894
rect 45266 478338 45502 478574
rect 45586 478338 45822 478574
rect 45266 442658 45502 442894
rect 45586 442658 45822 442894
rect 45266 442338 45502 442574
rect 45586 442338 45822 442574
rect 45266 406658 45502 406894
rect 45586 406658 45822 406894
rect 45266 406338 45502 406574
rect 45586 406338 45822 406574
rect 45266 370658 45502 370894
rect 45586 370658 45822 370894
rect 45266 370338 45502 370574
rect 45586 370338 45822 370574
rect 45266 334658 45502 334894
rect 45586 334658 45822 334894
rect 45266 334338 45502 334574
rect 45586 334338 45822 334574
rect 45266 298658 45502 298894
rect 45586 298658 45822 298894
rect 45266 298338 45502 298574
rect 45586 298338 45822 298574
rect 45266 262658 45502 262894
rect 45586 262658 45822 262894
rect 45266 262338 45502 262574
rect 45586 262338 45822 262574
rect 45266 226658 45502 226894
rect 45586 226658 45822 226894
rect 45266 226338 45502 226574
rect 45586 226338 45822 226574
rect 45266 190658 45502 190894
rect 45586 190658 45822 190894
rect 45266 190338 45502 190574
rect 45586 190338 45822 190574
rect 45266 154658 45502 154894
rect 45586 154658 45822 154894
rect 45266 154338 45502 154574
rect 45586 154338 45822 154574
rect 45266 118658 45502 118894
rect 45586 118658 45822 118894
rect 45266 118338 45502 118574
rect 45586 118338 45822 118574
rect 45266 82658 45502 82894
rect 45586 82658 45822 82894
rect 45266 82338 45502 82574
rect 45586 82338 45822 82574
rect 45266 46658 45502 46894
rect 45586 46658 45822 46894
rect 45266 46338 45502 46574
rect 45586 46338 45822 46574
rect 45266 10658 45502 10894
rect 45586 10658 45822 10894
rect 45266 10338 45502 10574
rect 45586 10338 45822 10574
rect 45266 -4422 45502 -4186
rect 45586 -4422 45822 -4186
rect 45266 -4742 45502 -4506
rect 45586 -4742 45822 -4506
rect 66986 711322 67222 711558
rect 67306 711322 67542 711558
rect 66986 711002 67222 711238
rect 67306 711002 67542 711238
rect 63266 709402 63502 709638
rect 63586 709402 63822 709638
rect 63266 709082 63502 709318
rect 63586 709082 63822 709318
rect 59546 707482 59782 707718
rect 59866 707482 60102 707718
rect 59546 707162 59782 707398
rect 59866 707162 60102 707398
rect 48986 698378 49222 698614
rect 49306 698378 49542 698614
rect 48986 698058 49222 698294
rect 49306 698058 49542 698294
rect 48986 662378 49222 662614
rect 49306 662378 49542 662614
rect 48986 662058 49222 662294
rect 49306 662058 49542 662294
rect 48986 626378 49222 626614
rect 49306 626378 49542 626614
rect 48986 626058 49222 626294
rect 49306 626058 49542 626294
rect 48986 590378 49222 590614
rect 49306 590378 49542 590614
rect 48986 590058 49222 590294
rect 49306 590058 49542 590294
rect 48986 554378 49222 554614
rect 49306 554378 49542 554614
rect 48986 554058 49222 554294
rect 49306 554058 49542 554294
rect 48986 518378 49222 518614
rect 49306 518378 49542 518614
rect 48986 518058 49222 518294
rect 49306 518058 49542 518294
rect 48986 482378 49222 482614
rect 49306 482378 49542 482614
rect 48986 482058 49222 482294
rect 49306 482058 49542 482294
rect 48986 446378 49222 446614
rect 49306 446378 49542 446614
rect 48986 446058 49222 446294
rect 49306 446058 49542 446294
rect 48986 410378 49222 410614
rect 49306 410378 49542 410614
rect 48986 410058 49222 410294
rect 49306 410058 49542 410294
rect 48986 374378 49222 374614
rect 49306 374378 49542 374614
rect 48986 374058 49222 374294
rect 49306 374058 49542 374294
rect 48986 338378 49222 338614
rect 49306 338378 49542 338614
rect 48986 338058 49222 338294
rect 49306 338058 49542 338294
rect 48986 302378 49222 302614
rect 49306 302378 49542 302614
rect 48986 302058 49222 302294
rect 49306 302058 49542 302294
rect 48986 266378 49222 266614
rect 49306 266378 49542 266614
rect 48986 266058 49222 266294
rect 49306 266058 49542 266294
rect 48986 230378 49222 230614
rect 49306 230378 49542 230614
rect 48986 230058 49222 230294
rect 49306 230058 49542 230294
rect 48986 194378 49222 194614
rect 49306 194378 49542 194614
rect 48986 194058 49222 194294
rect 49306 194058 49542 194294
rect 48986 158378 49222 158614
rect 49306 158378 49542 158614
rect 48986 158058 49222 158294
rect 49306 158058 49542 158294
rect 48986 122378 49222 122614
rect 49306 122378 49542 122614
rect 48986 122058 49222 122294
rect 49306 122058 49542 122294
rect 48986 86378 49222 86614
rect 49306 86378 49542 86614
rect 48986 86058 49222 86294
rect 49306 86058 49542 86294
rect 48986 50378 49222 50614
rect 49306 50378 49542 50614
rect 48986 50058 49222 50294
rect 49306 50058 49542 50294
rect 48986 14378 49222 14614
rect 49306 14378 49542 14614
rect 48986 14058 49222 14294
rect 49306 14058 49542 14294
rect 30986 -7302 31222 -7066
rect 31306 -7302 31542 -7066
rect 30986 -7622 31222 -7386
rect 31306 -7622 31542 -7386
rect 55826 705562 56062 705798
rect 56146 705562 56382 705798
rect 55826 705242 56062 705478
rect 56146 705242 56382 705478
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -1542 56062 -1306
rect 56146 -1542 56382 -1306
rect 55826 -1862 56062 -1626
rect 56146 -1862 56382 -1626
rect 59546 672938 59782 673174
rect 59866 672938 60102 673174
rect 59546 672618 59782 672854
rect 59866 672618 60102 672854
rect 59546 636938 59782 637174
rect 59866 636938 60102 637174
rect 59546 636618 59782 636854
rect 59866 636618 60102 636854
rect 59546 600938 59782 601174
rect 59866 600938 60102 601174
rect 59546 600618 59782 600854
rect 59866 600618 60102 600854
rect 59546 564938 59782 565174
rect 59866 564938 60102 565174
rect 59546 564618 59782 564854
rect 59866 564618 60102 564854
rect 59546 528938 59782 529174
rect 59866 528938 60102 529174
rect 59546 528618 59782 528854
rect 59866 528618 60102 528854
rect 59546 492938 59782 493174
rect 59866 492938 60102 493174
rect 59546 492618 59782 492854
rect 59866 492618 60102 492854
rect 59546 456938 59782 457174
rect 59866 456938 60102 457174
rect 59546 456618 59782 456854
rect 59866 456618 60102 456854
rect 59546 420938 59782 421174
rect 59866 420938 60102 421174
rect 59546 420618 59782 420854
rect 59866 420618 60102 420854
rect 59546 384938 59782 385174
rect 59866 384938 60102 385174
rect 59546 384618 59782 384854
rect 59866 384618 60102 384854
rect 59546 348938 59782 349174
rect 59866 348938 60102 349174
rect 59546 348618 59782 348854
rect 59866 348618 60102 348854
rect 59546 312938 59782 313174
rect 59866 312938 60102 313174
rect 59546 312618 59782 312854
rect 59866 312618 60102 312854
rect 59546 276938 59782 277174
rect 59866 276938 60102 277174
rect 59546 276618 59782 276854
rect 59866 276618 60102 276854
rect 59546 240938 59782 241174
rect 59866 240938 60102 241174
rect 59546 240618 59782 240854
rect 59866 240618 60102 240854
rect 59546 204938 59782 205174
rect 59866 204938 60102 205174
rect 59546 204618 59782 204854
rect 59866 204618 60102 204854
rect 59546 168938 59782 169174
rect 59866 168938 60102 169174
rect 59546 168618 59782 168854
rect 59866 168618 60102 168854
rect 59546 132938 59782 133174
rect 59866 132938 60102 133174
rect 59546 132618 59782 132854
rect 59866 132618 60102 132854
rect 59546 96938 59782 97174
rect 59866 96938 60102 97174
rect 59546 96618 59782 96854
rect 59866 96618 60102 96854
rect 59546 60938 59782 61174
rect 59866 60938 60102 61174
rect 59546 60618 59782 60854
rect 59866 60618 60102 60854
rect 59546 24938 59782 25174
rect 59866 24938 60102 25174
rect 59546 24618 59782 24854
rect 59866 24618 60102 24854
rect 59546 -3462 59782 -3226
rect 59866 -3462 60102 -3226
rect 59546 -3782 59782 -3546
rect 59866 -3782 60102 -3546
rect 63266 676658 63502 676894
rect 63586 676658 63822 676894
rect 63266 676338 63502 676574
rect 63586 676338 63822 676574
rect 63266 640658 63502 640894
rect 63586 640658 63822 640894
rect 63266 640338 63502 640574
rect 63586 640338 63822 640574
rect 63266 604658 63502 604894
rect 63586 604658 63822 604894
rect 63266 604338 63502 604574
rect 63586 604338 63822 604574
rect 63266 568658 63502 568894
rect 63586 568658 63822 568894
rect 63266 568338 63502 568574
rect 63586 568338 63822 568574
rect 63266 532658 63502 532894
rect 63586 532658 63822 532894
rect 63266 532338 63502 532574
rect 63586 532338 63822 532574
rect 63266 496658 63502 496894
rect 63586 496658 63822 496894
rect 63266 496338 63502 496574
rect 63586 496338 63822 496574
rect 63266 460658 63502 460894
rect 63586 460658 63822 460894
rect 63266 460338 63502 460574
rect 63586 460338 63822 460574
rect 63266 424658 63502 424894
rect 63586 424658 63822 424894
rect 63266 424338 63502 424574
rect 63586 424338 63822 424574
rect 63266 388658 63502 388894
rect 63586 388658 63822 388894
rect 63266 388338 63502 388574
rect 63586 388338 63822 388574
rect 63266 352658 63502 352894
rect 63586 352658 63822 352894
rect 63266 352338 63502 352574
rect 63586 352338 63822 352574
rect 63266 316658 63502 316894
rect 63586 316658 63822 316894
rect 63266 316338 63502 316574
rect 63586 316338 63822 316574
rect 63266 280658 63502 280894
rect 63586 280658 63822 280894
rect 63266 280338 63502 280574
rect 63586 280338 63822 280574
rect 63266 244658 63502 244894
rect 63586 244658 63822 244894
rect 63266 244338 63502 244574
rect 63586 244338 63822 244574
rect 63266 208658 63502 208894
rect 63586 208658 63822 208894
rect 63266 208338 63502 208574
rect 63586 208338 63822 208574
rect 63266 172658 63502 172894
rect 63586 172658 63822 172894
rect 63266 172338 63502 172574
rect 63586 172338 63822 172574
rect 63266 136658 63502 136894
rect 63586 136658 63822 136894
rect 63266 136338 63502 136574
rect 63586 136338 63822 136574
rect 63266 100658 63502 100894
rect 63586 100658 63822 100894
rect 63266 100338 63502 100574
rect 63586 100338 63822 100574
rect 63266 64658 63502 64894
rect 63586 64658 63822 64894
rect 63266 64338 63502 64574
rect 63586 64338 63822 64574
rect 63266 28658 63502 28894
rect 63586 28658 63822 28894
rect 63266 28338 63502 28574
rect 63586 28338 63822 28574
rect 63266 -5382 63502 -5146
rect 63586 -5382 63822 -5146
rect 63266 -5702 63502 -5466
rect 63586 -5702 63822 -5466
rect 84986 710362 85222 710598
rect 85306 710362 85542 710598
rect 84986 710042 85222 710278
rect 85306 710042 85542 710278
rect 81266 708442 81502 708678
rect 81586 708442 81822 708678
rect 81266 708122 81502 708358
rect 81586 708122 81822 708358
rect 77546 706522 77782 706758
rect 77866 706522 78102 706758
rect 77546 706202 77782 706438
rect 77866 706202 78102 706438
rect 66986 680378 67222 680614
rect 67306 680378 67542 680614
rect 66986 680058 67222 680294
rect 67306 680058 67542 680294
rect 66986 644378 67222 644614
rect 67306 644378 67542 644614
rect 66986 644058 67222 644294
rect 67306 644058 67542 644294
rect 66986 608378 67222 608614
rect 67306 608378 67542 608614
rect 66986 608058 67222 608294
rect 67306 608058 67542 608294
rect 66986 572378 67222 572614
rect 67306 572378 67542 572614
rect 66986 572058 67222 572294
rect 67306 572058 67542 572294
rect 66986 536378 67222 536614
rect 67306 536378 67542 536614
rect 66986 536058 67222 536294
rect 67306 536058 67542 536294
rect 66986 500378 67222 500614
rect 67306 500378 67542 500614
rect 66986 500058 67222 500294
rect 67306 500058 67542 500294
rect 66986 464378 67222 464614
rect 67306 464378 67542 464614
rect 66986 464058 67222 464294
rect 67306 464058 67542 464294
rect 66986 428378 67222 428614
rect 67306 428378 67542 428614
rect 66986 428058 67222 428294
rect 67306 428058 67542 428294
rect 66986 392378 67222 392614
rect 67306 392378 67542 392614
rect 66986 392058 67222 392294
rect 67306 392058 67542 392294
rect 66986 356378 67222 356614
rect 67306 356378 67542 356614
rect 66986 356058 67222 356294
rect 67306 356058 67542 356294
rect 66986 320378 67222 320614
rect 67306 320378 67542 320614
rect 66986 320058 67222 320294
rect 67306 320058 67542 320294
rect 66986 284378 67222 284614
rect 67306 284378 67542 284614
rect 66986 284058 67222 284294
rect 67306 284058 67542 284294
rect 66986 248378 67222 248614
rect 67306 248378 67542 248614
rect 66986 248058 67222 248294
rect 67306 248058 67542 248294
rect 66986 212378 67222 212614
rect 67306 212378 67542 212614
rect 66986 212058 67222 212294
rect 67306 212058 67542 212294
rect 66986 176378 67222 176614
rect 67306 176378 67542 176614
rect 66986 176058 67222 176294
rect 67306 176058 67542 176294
rect 66986 140378 67222 140614
rect 67306 140378 67542 140614
rect 66986 140058 67222 140294
rect 67306 140058 67542 140294
rect 66986 104378 67222 104614
rect 67306 104378 67542 104614
rect 66986 104058 67222 104294
rect 67306 104058 67542 104294
rect 66986 68378 67222 68614
rect 67306 68378 67542 68614
rect 66986 68058 67222 68294
rect 67306 68058 67542 68294
rect 66986 32378 67222 32614
rect 67306 32378 67542 32614
rect 66986 32058 67222 32294
rect 67306 32058 67542 32294
rect 48986 -6342 49222 -6106
rect 49306 -6342 49542 -6106
rect 48986 -6662 49222 -6426
rect 49306 -6662 49542 -6426
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 73826 579218 74062 579454
rect 74146 579218 74382 579454
rect 73826 578898 74062 579134
rect 74146 578898 74382 579134
rect 73826 543218 74062 543454
rect 74146 543218 74382 543454
rect 73826 542898 74062 543134
rect 74146 542898 74382 543134
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 73826 435218 74062 435454
rect 74146 435218 74382 435454
rect 73826 434898 74062 435134
rect 74146 434898 74382 435134
rect 73826 399218 74062 399454
rect 74146 399218 74382 399454
rect 73826 398898 74062 399134
rect 74146 398898 74382 399134
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 73826 327218 74062 327454
rect 74146 327218 74382 327454
rect 73826 326898 74062 327134
rect 74146 326898 74382 327134
rect 73826 291218 74062 291454
rect 74146 291218 74382 291454
rect 73826 290898 74062 291134
rect 74146 290898 74382 291134
rect 73826 255218 74062 255454
rect 74146 255218 74382 255454
rect 73826 254898 74062 255134
rect 74146 254898 74382 255134
rect 73826 219218 74062 219454
rect 74146 219218 74382 219454
rect 73826 218898 74062 219134
rect 74146 218898 74382 219134
rect 73826 183218 74062 183454
rect 74146 183218 74382 183454
rect 73826 182898 74062 183134
rect 74146 182898 74382 183134
rect 73826 147218 74062 147454
rect 74146 147218 74382 147454
rect 73826 146898 74062 147134
rect 74146 146898 74382 147134
rect 73826 111218 74062 111454
rect 74146 111218 74382 111454
rect 73826 110898 74062 111134
rect 74146 110898 74382 111134
rect 73826 75218 74062 75454
rect 74146 75218 74382 75454
rect 73826 74898 74062 75134
rect 74146 74898 74382 75134
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 77546 654938 77782 655174
rect 77866 654938 78102 655174
rect 77546 654618 77782 654854
rect 77866 654618 78102 654854
rect 77546 618938 77782 619174
rect 77866 618938 78102 619174
rect 77546 618618 77782 618854
rect 77866 618618 78102 618854
rect 77546 582938 77782 583174
rect 77866 582938 78102 583174
rect 77546 582618 77782 582854
rect 77866 582618 78102 582854
rect 77546 546938 77782 547174
rect 77866 546938 78102 547174
rect 77546 546618 77782 546854
rect 77866 546618 78102 546854
rect 77546 510938 77782 511174
rect 77866 510938 78102 511174
rect 77546 510618 77782 510854
rect 77866 510618 78102 510854
rect 77546 474938 77782 475174
rect 77866 474938 78102 475174
rect 77546 474618 77782 474854
rect 77866 474618 78102 474854
rect 77546 438938 77782 439174
rect 77866 438938 78102 439174
rect 77546 438618 77782 438854
rect 77866 438618 78102 438854
rect 77546 402938 77782 403174
rect 77866 402938 78102 403174
rect 77546 402618 77782 402854
rect 77866 402618 78102 402854
rect 77546 366938 77782 367174
rect 77866 366938 78102 367174
rect 77546 366618 77782 366854
rect 77866 366618 78102 366854
rect 77546 330938 77782 331174
rect 77866 330938 78102 331174
rect 77546 330618 77782 330854
rect 77866 330618 78102 330854
rect 77546 294938 77782 295174
rect 77866 294938 78102 295174
rect 77546 294618 77782 294854
rect 77866 294618 78102 294854
rect 77546 258938 77782 259174
rect 77866 258938 78102 259174
rect 77546 258618 77782 258854
rect 77866 258618 78102 258854
rect 77546 222938 77782 223174
rect 77866 222938 78102 223174
rect 77546 222618 77782 222854
rect 77866 222618 78102 222854
rect 77546 186938 77782 187174
rect 77866 186938 78102 187174
rect 77546 186618 77782 186854
rect 77866 186618 78102 186854
rect 77546 150938 77782 151174
rect 77866 150938 78102 151174
rect 77546 150618 77782 150854
rect 77866 150618 78102 150854
rect 77546 114938 77782 115174
rect 77866 114938 78102 115174
rect 77546 114618 77782 114854
rect 77866 114618 78102 114854
rect 77546 78938 77782 79174
rect 77866 78938 78102 79174
rect 77546 78618 77782 78854
rect 77866 78618 78102 78854
rect 77546 42938 77782 43174
rect 77866 42938 78102 43174
rect 77546 42618 77782 42854
rect 77866 42618 78102 42854
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 77546 -2502 77782 -2266
rect 77866 -2502 78102 -2266
rect 77546 -2822 77782 -2586
rect 77866 -2822 78102 -2586
rect 81266 694658 81502 694894
rect 81586 694658 81822 694894
rect 81266 694338 81502 694574
rect 81586 694338 81822 694574
rect 81266 658658 81502 658894
rect 81586 658658 81822 658894
rect 81266 658338 81502 658574
rect 81586 658338 81822 658574
rect 81266 622658 81502 622894
rect 81586 622658 81822 622894
rect 81266 622338 81502 622574
rect 81586 622338 81822 622574
rect 81266 586658 81502 586894
rect 81586 586658 81822 586894
rect 81266 586338 81502 586574
rect 81586 586338 81822 586574
rect 81266 550658 81502 550894
rect 81586 550658 81822 550894
rect 81266 550338 81502 550574
rect 81586 550338 81822 550574
rect 81266 514658 81502 514894
rect 81586 514658 81822 514894
rect 81266 514338 81502 514574
rect 81586 514338 81822 514574
rect 81266 478658 81502 478894
rect 81586 478658 81822 478894
rect 81266 478338 81502 478574
rect 81586 478338 81822 478574
rect 81266 442658 81502 442894
rect 81586 442658 81822 442894
rect 81266 442338 81502 442574
rect 81586 442338 81822 442574
rect 81266 406658 81502 406894
rect 81586 406658 81822 406894
rect 81266 406338 81502 406574
rect 81586 406338 81822 406574
rect 81266 370658 81502 370894
rect 81586 370658 81822 370894
rect 81266 370338 81502 370574
rect 81586 370338 81822 370574
rect 81266 334658 81502 334894
rect 81586 334658 81822 334894
rect 81266 334338 81502 334574
rect 81586 334338 81822 334574
rect 81266 298658 81502 298894
rect 81586 298658 81822 298894
rect 81266 298338 81502 298574
rect 81586 298338 81822 298574
rect 81266 262658 81502 262894
rect 81586 262658 81822 262894
rect 81266 262338 81502 262574
rect 81586 262338 81822 262574
rect 81266 226658 81502 226894
rect 81586 226658 81822 226894
rect 81266 226338 81502 226574
rect 81586 226338 81822 226574
rect 81266 190658 81502 190894
rect 81586 190658 81822 190894
rect 81266 190338 81502 190574
rect 81586 190338 81822 190574
rect 81266 154658 81502 154894
rect 81586 154658 81822 154894
rect 81266 154338 81502 154574
rect 81586 154338 81822 154574
rect 81266 118658 81502 118894
rect 81586 118658 81822 118894
rect 81266 118338 81502 118574
rect 81586 118338 81822 118574
rect 81266 82658 81502 82894
rect 81586 82658 81822 82894
rect 81266 82338 81502 82574
rect 81586 82338 81822 82574
rect 81266 46658 81502 46894
rect 81586 46658 81822 46894
rect 81266 46338 81502 46574
rect 81586 46338 81822 46574
rect 81266 10658 81502 10894
rect 81586 10658 81822 10894
rect 81266 10338 81502 10574
rect 81586 10338 81822 10574
rect 81266 -4422 81502 -4186
rect 81586 -4422 81822 -4186
rect 81266 -4742 81502 -4506
rect 81586 -4742 81822 -4506
rect 102986 711322 103222 711558
rect 103306 711322 103542 711558
rect 102986 711002 103222 711238
rect 103306 711002 103542 711238
rect 99266 709402 99502 709638
rect 99586 709402 99822 709638
rect 99266 709082 99502 709318
rect 99586 709082 99822 709318
rect 95546 707482 95782 707718
rect 95866 707482 96102 707718
rect 95546 707162 95782 707398
rect 95866 707162 96102 707398
rect 84986 698378 85222 698614
rect 85306 698378 85542 698614
rect 84986 698058 85222 698294
rect 85306 698058 85542 698294
rect 84986 662378 85222 662614
rect 85306 662378 85542 662614
rect 84986 662058 85222 662294
rect 85306 662058 85542 662294
rect 84986 626378 85222 626614
rect 85306 626378 85542 626614
rect 84986 626058 85222 626294
rect 85306 626058 85542 626294
rect 84986 590378 85222 590614
rect 85306 590378 85542 590614
rect 84986 590058 85222 590294
rect 85306 590058 85542 590294
rect 84986 554378 85222 554614
rect 85306 554378 85542 554614
rect 84986 554058 85222 554294
rect 85306 554058 85542 554294
rect 84986 518378 85222 518614
rect 85306 518378 85542 518614
rect 84986 518058 85222 518294
rect 85306 518058 85542 518294
rect 84986 482378 85222 482614
rect 85306 482378 85542 482614
rect 84986 482058 85222 482294
rect 85306 482058 85542 482294
rect 84986 446378 85222 446614
rect 85306 446378 85542 446614
rect 84986 446058 85222 446294
rect 85306 446058 85542 446294
rect 84986 410378 85222 410614
rect 85306 410378 85542 410614
rect 84986 410058 85222 410294
rect 85306 410058 85542 410294
rect 84986 374378 85222 374614
rect 85306 374378 85542 374614
rect 84986 374058 85222 374294
rect 85306 374058 85542 374294
rect 84986 338378 85222 338614
rect 85306 338378 85542 338614
rect 84986 338058 85222 338294
rect 85306 338058 85542 338294
rect 84986 302378 85222 302614
rect 85306 302378 85542 302614
rect 84986 302058 85222 302294
rect 85306 302058 85542 302294
rect 84986 266378 85222 266614
rect 85306 266378 85542 266614
rect 84986 266058 85222 266294
rect 85306 266058 85542 266294
rect 84986 230378 85222 230614
rect 85306 230378 85542 230614
rect 84986 230058 85222 230294
rect 85306 230058 85542 230294
rect 84986 194378 85222 194614
rect 85306 194378 85542 194614
rect 84986 194058 85222 194294
rect 85306 194058 85542 194294
rect 84986 158378 85222 158614
rect 85306 158378 85542 158614
rect 84986 158058 85222 158294
rect 85306 158058 85542 158294
rect 84986 122378 85222 122614
rect 85306 122378 85542 122614
rect 84986 122058 85222 122294
rect 85306 122058 85542 122294
rect 84986 86378 85222 86614
rect 85306 86378 85542 86614
rect 84986 86058 85222 86294
rect 85306 86058 85542 86294
rect 84986 50378 85222 50614
rect 85306 50378 85542 50614
rect 84986 50058 85222 50294
rect 85306 50058 85542 50294
rect 84986 14378 85222 14614
rect 85306 14378 85542 14614
rect 84986 14058 85222 14294
rect 85306 14058 85542 14294
rect 66986 -7302 67222 -7066
rect 67306 -7302 67542 -7066
rect 66986 -7622 67222 -7386
rect 67306 -7622 67542 -7386
rect 91826 705562 92062 705798
rect 92146 705562 92382 705798
rect 91826 705242 92062 705478
rect 92146 705242 92382 705478
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 91826 561218 92062 561454
rect 92146 561218 92382 561454
rect 91826 560898 92062 561134
rect 92146 560898 92382 561134
rect 91826 525218 92062 525454
rect 92146 525218 92382 525454
rect 91826 524898 92062 525134
rect 92146 524898 92382 525134
rect 91826 489218 92062 489454
rect 92146 489218 92382 489454
rect 91826 488898 92062 489134
rect 92146 488898 92382 489134
rect 91826 453218 92062 453454
rect 92146 453218 92382 453454
rect 91826 452898 92062 453134
rect 92146 452898 92382 453134
rect 91826 417218 92062 417454
rect 92146 417218 92382 417454
rect 91826 416898 92062 417134
rect 92146 416898 92382 417134
rect 91826 381218 92062 381454
rect 92146 381218 92382 381454
rect 91826 380898 92062 381134
rect 92146 380898 92382 381134
rect 91826 345218 92062 345454
rect 92146 345218 92382 345454
rect 91826 344898 92062 345134
rect 92146 344898 92382 345134
rect 91826 309218 92062 309454
rect 92146 309218 92382 309454
rect 91826 308898 92062 309134
rect 92146 308898 92382 309134
rect 91826 273218 92062 273454
rect 92146 273218 92382 273454
rect 91826 272898 92062 273134
rect 92146 272898 92382 273134
rect 91826 237218 92062 237454
rect 92146 237218 92382 237454
rect 91826 236898 92062 237134
rect 92146 236898 92382 237134
rect 91826 201218 92062 201454
rect 92146 201218 92382 201454
rect 91826 200898 92062 201134
rect 92146 200898 92382 201134
rect 91826 165218 92062 165454
rect 92146 165218 92382 165454
rect 91826 164898 92062 165134
rect 92146 164898 92382 165134
rect 91826 129218 92062 129454
rect 92146 129218 92382 129454
rect 91826 128898 92062 129134
rect 92146 128898 92382 129134
rect 91826 93218 92062 93454
rect 92146 93218 92382 93454
rect 91826 92898 92062 93134
rect 92146 92898 92382 93134
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -1542 92062 -1306
rect 92146 -1542 92382 -1306
rect 91826 -1862 92062 -1626
rect 92146 -1862 92382 -1626
rect 95546 672938 95782 673174
rect 95866 672938 96102 673174
rect 95546 672618 95782 672854
rect 95866 672618 96102 672854
rect 95546 636938 95782 637174
rect 95866 636938 96102 637174
rect 95546 636618 95782 636854
rect 95866 636618 96102 636854
rect 95546 600938 95782 601174
rect 95866 600938 96102 601174
rect 95546 600618 95782 600854
rect 95866 600618 96102 600854
rect 95546 564938 95782 565174
rect 95866 564938 96102 565174
rect 95546 564618 95782 564854
rect 95866 564618 96102 564854
rect 95546 528938 95782 529174
rect 95866 528938 96102 529174
rect 95546 528618 95782 528854
rect 95866 528618 96102 528854
rect 95546 492938 95782 493174
rect 95866 492938 96102 493174
rect 95546 492618 95782 492854
rect 95866 492618 96102 492854
rect 95546 456938 95782 457174
rect 95866 456938 96102 457174
rect 95546 456618 95782 456854
rect 95866 456618 96102 456854
rect 95546 420938 95782 421174
rect 95866 420938 96102 421174
rect 95546 420618 95782 420854
rect 95866 420618 96102 420854
rect 95546 384938 95782 385174
rect 95866 384938 96102 385174
rect 95546 384618 95782 384854
rect 95866 384618 96102 384854
rect 95546 348938 95782 349174
rect 95866 348938 96102 349174
rect 95546 348618 95782 348854
rect 95866 348618 96102 348854
rect 95546 312938 95782 313174
rect 95866 312938 96102 313174
rect 95546 312618 95782 312854
rect 95866 312618 96102 312854
rect 95546 276938 95782 277174
rect 95866 276938 96102 277174
rect 95546 276618 95782 276854
rect 95866 276618 96102 276854
rect 95546 240938 95782 241174
rect 95866 240938 96102 241174
rect 95546 240618 95782 240854
rect 95866 240618 96102 240854
rect 95546 204938 95782 205174
rect 95866 204938 96102 205174
rect 95546 204618 95782 204854
rect 95866 204618 96102 204854
rect 95546 168938 95782 169174
rect 95866 168938 96102 169174
rect 95546 168618 95782 168854
rect 95866 168618 96102 168854
rect 95546 132938 95782 133174
rect 95866 132938 96102 133174
rect 95546 132618 95782 132854
rect 95866 132618 96102 132854
rect 95546 96938 95782 97174
rect 95866 96938 96102 97174
rect 95546 96618 95782 96854
rect 95866 96618 96102 96854
rect 95546 60938 95782 61174
rect 95866 60938 96102 61174
rect 95546 60618 95782 60854
rect 95866 60618 96102 60854
rect 95546 24938 95782 25174
rect 95866 24938 96102 25174
rect 95546 24618 95782 24854
rect 95866 24618 96102 24854
rect 95546 -3462 95782 -3226
rect 95866 -3462 96102 -3226
rect 95546 -3782 95782 -3546
rect 95866 -3782 96102 -3546
rect 99266 676658 99502 676894
rect 99586 676658 99822 676894
rect 99266 676338 99502 676574
rect 99586 676338 99822 676574
rect 99266 640658 99502 640894
rect 99586 640658 99822 640894
rect 99266 640338 99502 640574
rect 99586 640338 99822 640574
rect 99266 604658 99502 604894
rect 99586 604658 99822 604894
rect 99266 604338 99502 604574
rect 99586 604338 99822 604574
rect 99266 568658 99502 568894
rect 99586 568658 99822 568894
rect 99266 568338 99502 568574
rect 99586 568338 99822 568574
rect 99266 532658 99502 532894
rect 99586 532658 99822 532894
rect 99266 532338 99502 532574
rect 99586 532338 99822 532574
rect 99266 496658 99502 496894
rect 99586 496658 99822 496894
rect 99266 496338 99502 496574
rect 99586 496338 99822 496574
rect 99266 460658 99502 460894
rect 99586 460658 99822 460894
rect 99266 460338 99502 460574
rect 99586 460338 99822 460574
rect 99266 424658 99502 424894
rect 99586 424658 99822 424894
rect 99266 424338 99502 424574
rect 99586 424338 99822 424574
rect 99266 388658 99502 388894
rect 99586 388658 99822 388894
rect 99266 388338 99502 388574
rect 99586 388338 99822 388574
rect 99266 352658 99502 352894
rect 99586 352658 99822 352894
rect 99266 352338 99502 352574
rect 99586 352338 99822 352574
rect 99266 316658 99502 316894
rect 99586 316658 99822 316894
rect 99266 316338 99502 316574
rect 99586 316338 99822 316574
rect 99266 280658 99502 280894
rect 99586 280658 99822 280894
rect 99266 280338 99502 280574
rect 99586 280338 99822 280574
rect 99266 244658 99502 244894
rect 99586 244658 99822 244894
rect 99266 244338 99502 244574
rect 99586 244338 99822 244574
rect 99266 208658 99502 208894
rect 99586 208658 99822 208894
rect 99266 208338 99502 208574
rect 99586 208338 99822 208574
rect 99266 172658 99502 172894
rect 99586 172658 99822 172894
rect 99266 172338 99502 172574
rect 99586 172338 99822 172574
rect 99266 136658 99502 136894
rect 99586 136658 99822 136894
rect 99266 136338 99502 136574
rect 99586 136338 99822 136574
rect 99266 100658 99502 100894
rect 99586 100658 99822 100894
rect 99266 100338 99502 100574
rect 99586 100338 99822 100574
rect 99266 64658 99502 64894
rect 99586 64658 99822 64894
rect 99266 64338 99502 64574
rect 99586 64338 99822 64574
rect 99266 28658 99502 28894
rect 99586 28658 99822 28894
rect 99266 28338 99502 28574
rect 99586 28338 99822 28574
rect 99266 -5382 99502 -5146
rect 99586 -5382 99822 -5146
rect 99266 -5702 99502 -5466
rect 99586 -5702 99822 -5466
rect 120986 710362 121222 710598
rect 121306 710362 121542 710598
rect 120986 710042 121222 710278
rect 121306 710042 121542 710278
rect 117266 708442 117502 708678
rect 117586 708442 117822 708678
rect 117266 708122 117502 708358
rect 117586 708122 117822 708358
rect 113546 706522 113782 706758
rect 113866 706522 114102 706758
rect 113546 706202 113782 706438
rect 113866 706202 114102 706438
rect 102986 680378 103222 680614
rect 103306 680378 103542 680614
rect 102986 680058 103222 680294
rect 103306 680058 103542 680294
rect 102986 644378 103222 644614
rect 103306 644378 103542 644614
rect 102986 644058 103222 644294
rect 103306 644058 103542 644294
rect 102986 608378 103222 608614
rect 103306 608378 103542 608614
rect 102986 608058 103222 608294
rect 103306 608058 103542 608294
rect 102986 572378 103222 572614
rect 103306 572378 103542 572614
rect 102986 572058 103222 572294
rect 103306 572058 103542 572294
rect 102986 536378 103222 536614
rect 103306 536378 103542 536614
rect 102986 536058 103222 536294
rect 103306 536058 103542 536294
rect 102986 500378 103222 500614
rect 103306 500378 103542 500614
rect 102986 500058 103222 500294
rect 103306 500058 103542 500294
rect 102986 464378 103222 464614
rect 103306 464378 103542 464614
rect 102986 464058 103222 464294
rect 103306 464058 103542 464294
rect 102986 428378 103222 428614
rect 103306 428378 103542 428614
rect 102986 428058 103222 428294
rect 103306 428058 103542 428294
rect 102986 392378 103222 392614
rect 103306 392378 103542 392614
rect 102986 392058 103222 392294
rect 103306 392058 103542 392294
rect 102986 356378 103222 356614
rect 103306 356378 103542 356614
rect 102986 356058 103222 356294
rect 103306 356058 103542 356294
rect 102986 320378 103222 320614
rect 103306 320378 103542 320614
rect 102986 320058 103222 320294
rect 103306 320058 103542 320294
rect 102986 284378 103222 284614
rect 103306 284378 103542 284614
rect 102986 284058 103222 284294
rect 103306 284058 103542 284294
rect 102986 248378 103222 248614
rect 103306 248378 103542 248614
rect 102986 248058 103222 248294
rect 103306 248058 103542 248294
rect 102986 212378 103222 212614
rect 103306 212378 103542 212614
rect 102986 212058 103222 212294
rect 103306 212058 103542 212294
rect 102986 176378 103222 176614
rect 103306 176378 103542 176614
rect 102986 176058 103222 176294
rect 103306 176058 103542 176294
rect 102986 140378 103222 140614
rect 103306 140378 103542 140614
rect 102986 140058 103222 140294
rect 103306 140058 103542 140294
rect 102986 104378 103222 104614
rect 103306 104378 103542 104614
rect 102986 104058 103222 104294
rect 103306 104058 103542 104294
rect 102986 68378 103222 68614
rect 103306 68378 103542 68614
rect 102986 68058 103222 68294
rect 103306 68058 103542 68294
rect 102986 32378 103222 32614
rect 103306 32378 103542 32614
rect 102986 32058 103222 32294
rect 103306 32058 103542 32294
rect 84986 -6342 85222 -6106
rect 85306 -6342 85542 -6106
rect 84986 -6662 85222 -6426
rect 85306 -6662 85542 -6426
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 109826 507218 110062 507454
rect 110146 507218 110382 507454
rect 109826 506898 110062 507134
rect 110146 506898 110382 507134
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 109826 435218 110062 435454
rect 110146 435218 110382 435454
rect 109826 434898 110062 435134
rect 110146 434898 110382 435134
rect 109826 399218 110062 399454
rect 110146 399218 110382 399454
rect 109826 398898 110062 399134
rect 110146 398898 110382 399134
rect 109826 363218 110062 363454
rect 110146 363218 110382 363454
rect 109826 362898 110062 363134
rect 110146 362898 110382 363134
rect 109826 327218 110062 327454
rect 110146 327218 110382 327454
rect 109826 326898 110062 327134
rect 110146 326898 110382 327134
rect 109826 291218 110062 291454
rect 110146 291218 110382 291454
rect 109826 290898 110062 291134
rect 110146 290898 110382 291134
rect 109826 255218 110062 255454
rect 110146 255218 110382 255454
rect 109826 254898 110062 255134
rect 110146 254898 110382 255134
rect 109826 219218 110062 219454
rect 110146 219218 110382 219454
rect 109826 218898 110062 219134
rect 110146 218898 110382 219134
rect 109826 183218 110062 183454
rect 110146 183218 110382 183454
rect 109826 182898 110062 183134
rect 110146 182898 110382 183134
rect 109826 147218 110062 147454
rect 110146 147218 110382 147454
rect 109826 146898 110062 147134
rect 110146 146898 110382 147134
rect 109826 111218 110062 111454
rect 110146 111218 110382 111454
rect 109826 110898 110062 111134
rect 110146 110898 110382 111134
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 690938 113782 691174
rect 113866 690938 114102 691174
rect 113546 690618 113782 690854
rect 113866 690618 114102 690854
rect 113546 654938 113782 655174
rect 113866 654938 114102 655174
rect 113546 654618 113782 654854
rect 113866 654618 114102 654854
rect 113546 618938 113782 619174
rect 113866 618938 114102 619174
rect 113546 618618 113782 618854
rect 113866 618618 114102 618854
rect 113546 582938 113782 583174
rect 113866 582938 114102 583174
rect 113546 582618 113782 582854
rect 113866 582618 114102 582854
rect 113546 546938 113782 547174
rect 113866 546938 114102 547174
rect 113546 546618 113782 546854
rect 113866 546618 114102 546854
rect 113546 510938 113782 511174
rect 113866 510938 114102 511174
rect 113546 510618 113782 510854
rect 113866 510618 114102 510854
rect 113546 474938 113782 475174
rect 113866 474938 114102 475174
rect 113546 474618 113782 474854
rect 113866 474618 114102 474854
rect 113546 438938 113782 439174
rect 113866 438938 114102 439174
rect 113546 438618 113782 438854
rect 113866 438618 114102 438854
rect 113546 402938 113782 403174
rect 113866 402938 114102 403174
rect 113546 402618 113782 402854
rect 113866 402618 114102 402854
rect 113546 366938 113782 367174
rect 113866 366938 114102 367174
rect 113546 366618 113782 366854
rect 113866 366618 114102 366854
rect 113546 330938 113782 331174
rect 113866 330938 114102 331174
rect 113546 330618 113782 330854
rect 113866 330618 114102 330854
rect 113546 294938 113782 295174
rect 113866 294938 114102 295174
rect 113546 294618 113782 294854
rect 113866 294618 114102 294854
rect 113546 258938 113782 259174
rect 113866 258938 114102 259174
rect 113546 258618 113782 258854
rect 113866 258618 114102 258854
rect 113546 222938 113782 223174
rect 113866 222938 114102 223174
rect 113546 222618 113782 222854
rect 113866 222618 114102 222854
rect 113546 186938 113782 187174
rect 113866 186938 114102 187174
rect 113546 186618 113782 186854
rect 113866 186618 114102 186854
rect 113546 150938 113782 151174
rect 113866 150938 114102 151174
rect 113546 150618 113782 150854
rect 113866 150618 114102 150854
rect 113546 114938 113782 115174
rect 113866 114938 114102 115174
rect 113546 114618 113782 114854
rect 113866 114618 114102 114854
rect 113546 78938 113782 79174
rect 113866 78938 114102 79174
rect 113546 78618 113782 78854
rect 113866 78618 114102 78854
rect 113546 42938 113782 43174
rect 113866 42938 114102 43174
rect 113546 42618 113782 42854
rect 113866 42618 114102 42854
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 113546 -2502 113782 -2266
rect 113866 -2502 114102 -2266
rect 113546 -2822 113782 -2586
rect 113866 -2822 114102 -2586
rect 117266 694658 117502 694894
rect 117586 694658 117822 694894
rect 117266 694338 117502 694574
rect 117586 694338 117822 694574
rect 117266 658658 117502 658894
rect 117586 658658 117822 658894
rect 117266 658338 117502 658574
rect 117586 658338 117822 658574
rect 117266 622658 117502 622894
rect 117586 622658 117822 622894
rect 117266 622338 117502 622574
rect 117586 622338 117822 622574
rect 117266 586658 117502 586894
rect 117586 586658 117822 586894
rect 117266 586338 117502 586574
rect 117586 586338 117822 586574
rect 117266 550658 117502 550894
rect 117586 550658 117822 550894
rect 117266 550338 117502 550574
rect 117586 550338 117822 550574
rect 117266 514658 117502 514894
rect 117586 514658 117822 514894
rect 117266 514338 117502 514574
rect 117586 514338 117822 514574
rect 117266 478658 117502 478894
rect 117586 478658 117822 478894
rect 117266 478338 117502 478574
rect 117586 478338 117822 478574
rect 117266 442658 117502 442894
rect 117586 442658 117822 442894
rect 117266 442338 117502 442574
rect 117586 442338 117822 442574
rect 117266 406658 117502 406894
rect 117586 406658 117822 406894
rect 117266 406338 117502 406574
rect 117586 406338 117822 406574
rect 117266 370658 117502 370894
rect 117586 370658 117822 370894
rect 117266 370338 117502 370574
rect 117586 370338 117822 370574
rect 117266 334658 117502 334894
rect 117586 334658 117822 334894
rect 117266 334338 117502 334574
rect 117586 334338 117822 334574
rect 117266 298658 117502 298894
rect 117586 298658 117822 298894
rect 117266 298338 117502 298574
rect 117586 298338 117822 298574
rect 117266 262658 117502 262894
rect 117586 262658 117822 262894
rect 117266 262338 117502 262574
rect 117586 262338 117822 262574
rect 117266 226658 117502 226894
rect 117586 226658 117822 226894
rect 117266 226338 117502 226574
rect 117586 226338 117822 226574
rect 117266 190658 117502 190894
rect 117586 190658 117822 190894
rect 117266 190338 117502 190574
rect 117586 190338 117822 190574
rect 117266 154658 117502 154894
rect 117586 154658 117822 154894
rect 117266 154338 117502 154574
rect 117586 154338 117822 154574
rect 117266 118658 117502 118894
rect 117586 118658 117822 118894
rect 117266 118338 117502 118574
rect 117586 118338 117822 118574
rect 117266 82658 117502 82894
rect 117586 82658 117822 82894
rect 117266 82338 117502 82574
rect 117586 82338 117822 82574
rect 117266 46658 117502 46894
rect 117586 46658 117822 46894
rect 117266 46338 117502 46574
rect 117586 46338 117822 46574
rect 117266 10658 117502 10894
rect 117586 10658 117822 10894
rect 117266 10338 117502 10574
rect 117586 10338 117822 10574
rect 117266 -4422 117502 -4186
rect 117586 -4422 117822 -4186
rect 117266 -4742 117502 -4506
rect 117586 -4742 117822 -4506
rect 138986 711322 139222 711558
rect 139306 711322 139542 711558
rect 138986 711002 139222 711238
rect 139306 711002 139542 711238
rect 135266 709402 135502 709638
rect 135586 709402 135822 709638
rect 135266 709082 135502 709318
rect 135586 709082 135822 709318
rect 131546 707482 131782 707718
rect 131866 707482 132102 707718
rect 131546 707162 131782 707398
rect 131866 707162 132102 707398
rect 120986 698378 121222 698614
rect 121306 698378 121542 698614
rect 120986 698058 121222 698294
rect 121306 698058 121542 698294
rect 120986 662378 121222 662614
rect 121306 662378 121542 662614
rect 120986 662058 121222 662294
rect 121306 662058 121542 662294
rect 120986 626378 121222 626614
rect 121306 626378 121542 626614
rect 120986 626058 121222 626294
rect 121306 626058 121542 626294
rect 120986 590378 121222 590614
rect 121306 590378 121542 590614
rect 120986 590058 121222 590294
rect 121306 590058 121542 590294
rect 120986 554378 121222 554614
rect 121306 554378 121542 554614
rect 120986 554058 121222 554294
rect 121306 554058 121542 554294
rect 120986 518378 121222 518614
rect 121306 518378 121542 518614
rect 120986 518058 121222 518294
rect 121306 518058 121542 518294
rect 120986 482378 121222 482614
rect 121306 482378 121542 482614
rect 120986 482058 121222 482294
rect 121306 482058 121542 482294
rect 120986 446378 121222 446614
rect 121306 446378 121542 446614
rect 120986 446058 121222 446294
rect 121306 446058 121542 446294
rect 120986 410378 121222 410614
rect 121306 410378 121542 410614
rect 120986 410058 121222 410294
rect 121306 410058 121542 410294
rect 120986 374378 121222 374614
rect 121306 374378 121542 374614
rect 120986 374058 121222 374294
rect 121306 374058 121542 374294
rect 120986 338378 121222 338614
rect 121306 338378 121542 338614
rect 120986 338058 121222 338294
rect 121306 338058 121542 338294
rect 120986 302378 121222 302614
rect 121306 302378 121542 302614
rect 120986 302058 121222 302294
rect 121306 302058 121542 302294
rect 120986 266378 121222 266614
rect 121306 266378 121542 266614
rect 120986 266058 121222 266294
rect 121306 266058 121542 266294
rect 120986 230378 121222 230614
rect 121306 230378 121542 230614
rect 120986 230058 121222 230294
rect 121306 230058 121542 230294
rect 120986 194378 121222 194614
rect 121306 194378 121542 194614
rect 120986 194058 121222 194294
rect 121306 194058 121542 194294
rect 120986 158378 121222 158614
rect 121306 158378 121542 158614
rect 120986 158058 121222 158294
rect 121306 158058 121542 158294
rect 120986 122378 121222 122614
rect 121306 122378 121542 122614
rect 120986 122058 121222 122294
rect 121306 122058 121542 122294
rect 120986 86378 121222 86614
rect 121306 86378 121542 86614
rect 120986 86058 121222 86294
rect 121306 86058 121542 86294
rect 120986 50378 121222 50614
rect 121306 50378 121542 50614
rect 120986 50058 121222 50294
rect 121306 50058 121542 50294
rect 120986 14378 121222 14614
rect 121306 14378 121542 14614
rect 120986 14058 121222 14294
rect 121306 14058 121542 14294
rect 102986 -7302 103222 -7066
rect 103306 -7302 103542 -7066
rect 102986 -7622 103222 -7386
rect 103306 -7622 103542 -7386
rect 127826 705562 128062 705798
rect 128146 705562 128382 705798
rect 127826 705242 128062 705478
rect 128146 705242 128382 705478
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 127826 561218 128062 561454
rect 128146 561218 128382 561454
rect 127826 560898 128062 561134
rect 128146 560898 128382 561134
rect 127826 525218 128062 525454
rect 128146 525218 128382 525454
rect 127826 524898 128062 525134
rect 128146 524898 128382 525134
rect 127826 489218 128062 489454
rect 128146 489218 128382 489454
rect 127826 488898 128062 489134
rect 128146 488898 128382 489134
rect 127826 453218 128062 453454
rect 128146 453218 128382 453454
rect 127826 452898 128062 453134
rect 128146 452898 128382 453134
rect 127826 417218 128062 417454
rect 128146 417218 128382 417454
rect 127826 416898 128062 417134
rect 128146 416898 128382 417134
rect 127826 381218 128062 381454
rect 128146 381218 128382 381454
rect 127826 380898 128062 381134
rect 128146 380898 128382 381134
rect 127826 345218 128062 345454
rect 128146 345218 128382 345454
rect 127826 344898 128062 345134
rect 128146 344898 128382 345134
rect 127826 309218 128062 309454
rect 128146 309218 128382 309454
rect 127826 308898 128062 309134
rect 128146 308898 128382 309134
rect 127826 273218 128062 273454
rect 128146 273218 128382 273454
rect 127826 272898 128062 273134
rect 128146 272898 128382 273134
rect 127826 237218 128062 237454
rect 128146 237218 128382 237454
rect 127826 236898 128062 237134
rect 128146 236898 128382 237134
rect 127826 201218 128062 201454
rect 128146 201218 128382 201454
rect 127826 200898 128062 201134
rect 128146 200898 128382 201134
rect 127826 165218 128062 165454
rect 128146 165218 128382 165454
rect 127826 164898 128062 165134
rect 128146 164898 128382 165134
rect 127826 129218 128062 129454
rect 128146 129218 128382 129454
rect 127826 128898 128062 129134
rect 128146 128898 128382 129134
rect 127826 93218 128062 93454
rect 128146 93218 128382 93454
rect 127826 92898 128062 93134
rect 128146 92898 128382 93134
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -1542 128062 -1306
rect 128146 -1542 128382 -1306
rect 127826 -1862 128062 -1626
rect 128146 -1862 128382 -1626
rect 131546 672938 131782 673174
rect 131866 672938 132102 673174
rect 131546 672618 131782 672854
rect 131866 672618 132102 672854
rect 131546 636938 131782 637174
rect 131866 636938 132102 637174
rect 131546 636618 131782 636854
rect 131866 636618 132102 636854
rect 131546 600938 131782 601174
rect 131866 600938 132102 601174
rect 131546 600618 131782 600854
rect 131866 600618 132102 600854
rect 131546 564938 131782 565174
rect 131866 564938 132102 565174
rect 131546 564618 131782 564854
rect 131866 564618 132102 564854
rect 131546 528938 131782 529174
rect 131866 528938 132102 529174
rect 131546 528618 131782 528854
rect 131866 528618 132102 528854
rect 131546 492938 131782 493174
rect 131866 492938 132102 493174
rect 131546 492618 131782 492854
rect 131866 492618 132102 492854
rect 131546 456938 131782 457174
rect 131866 456938 132102 457174
rect 131546 456618 131782 456854
rect 131866 456618 132102 456854
rect 131546 420938 131782 421174
rect 131866 420938 132102 421174
rect 131546 420618 131782 420854
rect 131866 420618 132102 420854
rect 131546 384938 131782 385174
rect 131866 384938 132102 385174
rect 131546 384618 131782 384854
rect 131866 384618 132102 384854
rect 131546 348938 131782 349174
rect 131866 348938 132102 349174
rect 131546 348618 131782 348854
rect 131866 348618 132102 348854
rect 131546 312938 131782 313174
rect 131866 312938 132102 313174
rect 131546 312618 131782 312854
rect 131866 312618 132102 312854
rect 131546 276938 131782 277174
rect 131866 276938 132102 277174
rect 131546 276618 131782 276854
rect 131866 276618 132102 276854
rect 131546 240938 131782 241174
rect 131866 240938 132102 241174
rect 131546 240618 131782 240854
rect 131866 240618 132102 240854
rect 131546 204938 131782 205174
rect 131866 204938 132102 205174
rect 131546 204618 131782 204854
rect 131866 204618 132102 204854
rect 131546 168938 131782 169174
rect 131866 168938 132102 169174
rect 131546 168618 131782 168854
rect 131866 168618 132102 168854
rect 131546 132938 131782 133174
rect 131866 132938 132102 133174
rect 131546 132618 131782 132854
rect 131866 132618 132102 132854
rect 131546 96938 131782 97174
rect 131866 96938 132102 97174
rect 131546 96618 131782 96854
rect 131866 96618 132102 96854
rect 131546 60938 131782 61174
rect 131866 60938 132102 61174
rect 131546 60618 131782 60854
rect 131866 60618 132102 60854
rect 131546 24938 131782 25174
rect 131866 24938 132102 25174
rect 131546 24618 131782 24854
rect 131866 24618 132102 24854
rect 131546 -3462 131782 -3226
rect 131866 -3462 132102 -3226
rect 131546 -3782 131782 -3546
rect 131866 -3782 132102 -3546
rect 135266 676658 135502 676894
rect 135586 676658 135822 676894
rect 135266 676338 135502 676574
rect 135586 676338 135822 676574
rect 135266 640658 135502 640894
rect 135586 640658 135822 640894
rect 135266 640338 135502 640574
rect 135586 640338 135822 640574
rect 135266 604658 135502 604894
rect 135586 604658 135822 604894
rect 135266 604338 135502 604574
rect 135586 604338 135822 604574
rect 135266 568658 135502 568894
rect 135586 568658 135822 568894
rect 135266 568338 135502 568574
rect 135586 568338 135822 568574
rect 135266 532658 135502 532894
rect 135586 532658 135822 532894
rect 135266 532338 135502 532574
rect 135586 532338 135822 532574
rect 135266 496658 135502 496894
rect 135586 496658 135822 496894
rect 135266 496338 135502 496574
rect 135586 496338 135822 496574
rect 135266 460658 135502 460894
rect 135586 460658 135822 460894
rect 135266 460338 135502 460574
rect 135586 460338 135822 460574
rect 135266 424658 135502 424894
rect 135586 424658 135822 424894
rect 135266 424338 135502 424574
rect 135586 424338 135822 424574
rect 135266 388658 135502 388894
rect 135586 388658 135822 388894
rect 135266 388338 135502 388574
rect 135586 388338 135822 388574
rect 135266 352658 135502 352894
rect 135586 352658 135822 352894
rect 135266 352338 135502 352574
rect 135586 352338 135822 352574
rect 135266 316658 135502 316894
rect 135586 316658 135822 316894
rect 135266 316338 135502 316574
rect 135586 316338 135822 316574
rect 135266 280658 135502 280894
rect 135586 280658 135822 280894
rect 135266 280338 135502 280574
rect 135586 280338 135822 280574
rect 135266 244658 135502 244894
rect 135586 244658 135822 244894
rect 135266 244338 135502 244574
rect 135586 244338 135822 244574
rect 135266 208658 135502 208894
rect 135586 208658 135822 208894
rect 135266 208338 135502 208574
rect 135586 208338 135822 208574
rect 135266 172658 135502 172894
rect 135586 172658 135822 172894
rect 135266 172338 135502 172574
rect 135586 172338 135822 172574
rect 135266 136658 135502 136894
rect 135586 136658 135822 136894
rect 135266 136338 135502 136574
rect 135586 136338 135822 136574
rect 135266 100658 135502 100894
rect 135586 100658 135822 100894
rect 135266 100338 135502 100574
rect 135586 100338 135822 100574
rect 135266 64658 135502 64894
rect 135586 64658 135822 64894
rect 135266 64338 135502 64574
rect 135586 64338 135822 64574
rect 135266 28658 135502 28894
rect 135586 28658 135822 28894
rect 135266 28338 135502 28574
rect 135586 28338 135822 28574
rect 135266 -5382 135502 -5146
rect 135586 -5382 135822 -5146
rect 135266 -5702 135502 -5466
rect 135586 -5702 135822 -5466
rect 156986 710362 157222 710598
rect 157306 710362 157542 710598
rect 156986 710042 157222 710278
rect 157306 710042 157542 710278
rect 153266 708442 153502 708678
rect 153586 708442 153822 708678
rect 153266 708122 153502 708358
rect 153586 708122 153822 708358
rect 149546 706522 149782 706758
rect 149866 706522 150102 706758
rect 149546 706202 149782 706438
rect 149866 706202 150102 706438
rect 138986 680378 139222 680614
rect 139306 680378 139542 680614
rect 138986 680058 139222 680294
rect 139306 680058 139542 680294
rect 138986 644378 139222 644614
rect 139306 644378 139542 644614
rect 138986 644058 139222 644294
rect 139306 644058 139542 644294
rect 138986 608378 139222 608614
rect 139306 608378 139542 608614
rect 138986 608058 139222 608294
rect 139306 608058 139542 608294
rect 138986 572378 139222 572614
rect 139306 572378 139542 572614
rect 138986 572058 139222 572294
rect 139306 572058 139542 572294
rect 138986 536378 139222 536614
rect 139306 536378 139542 536614
rect 138986 536058 139222 536294
rect 139306 536058 139542 536294
rect 138986 500378 139222 500614
rect 139306 500378 139542 500614
rect 138986 500058 139222 500294
rect 139306 500058 139542 500294
rect 138986 464378 139222 464614
rect 139306 464378 139542 464614
rect 138986 464058 139222 464294
rect 139306 464058 139542 464294
rect 138986 428378 139222 428614
rect 139306 428378 139542 428614
rect 138986 428058 139222 428294
rect 139306 428058 139542 428294
rect 138986 392378 139222 392614
rect 139306 392378 139542 392614
rect 138986 392058 139222 392294
rect 139306 392058 139542 392294
rect 138986 356378 139222 356614
rect 139306 356378 139542 356614
rect 138986 356058 139222 356294
rect 139306 356058 139542 356294
rect 138986 320378 139222 320614
rect 139306 320378 139542 320614
rect 138986 320058 139222 320294
rect 139306 320058 139542 320294
rect 138986 284378 139222 284614
rect 139306 284378 139542 284614
rect 138986 284058 139222 284294
rect 139306 284058 139542 284294
rect 138986 248378 139222 248614
rect 139306 248378 139542 248614
rect 138986 248058 139222 248294
rect 139306 248058 139542 248294
rect 138986 212378 139222 212614
rect 139306 212378 139542 212614
rect 138986 212058 139222 212294
rect 139306 212058 139542 212294
rect 138986 176378 139222 176614
rect 139306 176378 139542 176614
rect 138986 176058 139222 176294
rect 139306 176058 139542 176294
rect 138986 140378 139222 140614
rect 139306 140378 139542 140614
rect 138986 140058 139222 140294
rect 139306 140058 139542 140294
rect 138986 104378 139222 104614
rect 139306 104378 139542 104614
rect 138986 104058 139222 104294
rect 139306 104058 139542 104294
rect 138986 68378 139222 68614
rect 139306 68378 139542 68614
rect 138986 68058 139222 68294
rect 139306 68058 139542 68294
rect 138986 32378 139222 32614
rect 139306 32378 139542 32614
rect 138986 32058 139222 32294
rect 139306 32058 139542 32294
rect 120986 -6342 121222 -6106
rect 121306 -6342 121542 -6106
rect 120986 -6662 121222 -6426
rect 121306 -6662 121542 -6426
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 145826 507218 146062 507454
rect 146146 507218 146382 507454
rect 145826 506898 146062 507134
rect 146146 506898 146382 507134
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 145826 435218 146062 435454
rect 146146 435218 146382 435454
rect 145826 434898 146062 435134
rect 146146 434898 146382 435134
rect 145826 399218 146062 399454
rect 146146 399218 146382 399454
rect 145826 398898 146062 399134
rect 146146 398898 146382 399134
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 145826 327218 146062 327454
rect 146146 327218 146382 327454
rect 145826 326898 146062 327134
rect 146146 326898 146382 327134
rect 145826 291218 146062 291454
rect 146146 291218 146382 291454
rect 145826 290898 146062 291134
rect 146146 290898 146382 291134
rect 145826 255218 146062 255454
rect 146146 255218 146382 255454
rect 145826 254898 146062 255134
rect 146146 254898 146382 255134
rect 145826 219218 146062 219454
rect 146146 219218 146382 219454
rect 145826 218898 146062 219134
rect 146146 218898 146382 219134
rect 145826 183218 146062 183454
rect 146146 183218 146382 183454
rect 145826 182898 146062 183134
rect 146146 182898 146382 183134
rect 145826 147218 146062 147454
rect 146146 147218 146382 147454
rect 145826 146898 146062 147134
rect 146146 146898 146382 147134
rect 145826 111218 146062 111454
rect 146146 111218 146382 111454
rect 145826 110898 146062 111134
rect 146146 110898 146382 111134
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 149546 654938 149782 655174
rect 149866 654938 150102 655174
rect 149546 654618 149782 654854
rect 149866 654618 150102 654854
rect 149546 618938 149782 619174
rect 149866 618938 150102 619174
rect 149546 618618 149782 618854
rect 149866 618618 150102 618854
rect 149546 582938 149782 583174
rect 149866 582938 150102 583174
rect 149546 582618 149782 582854
rect 149866 582618 150102 582854
rect 149546 546938 149782 547174
rect 149866 546938 150102 547174
rect 149546 546618 149782 546854
rect 149866 546618 150102 546854
rect 149546 510938 149782 511174
rect 149866 510938 150102 511174
rect 149546 510618 149782 510854
rect 149866 510618 150102 510854
rect 149546 474938 149782 475174
rect 149866 474938 150102 475174
rect 149546 474618 149782 474854
rect 149866 474618 150102 474854
rect 149546 438938 149782 439174
rect 149866 438938 150102 439174
rect 149546 438618 149782 438854
rect 149866 438618 150102 438854
rect 149546 402938 149782 403174
rect 149866 402938 150102 403174
rect 149546 402618 149782 402854
rect 149866 402618 150102 402854
rect 149546 366938 149782 367174
rect 149866 366938 150102 367174
rect 149546 366618 149782 366854
rect 149866 366618 150102 366854
rect 149546 330938 149782 331174
rect 149866 330938 150102 331174
rect 149546 330618 149782 330854
rect 149866 330618 150102 330854
rect 149546 294938 149782 295174
rect 149866 294938 150102 295174
rect 149546 294618 149782 294854
rect 149866 294618 150102 294854
rect 149546 258938 149782 259174
rect 149866 258938 150102 259174
rect 149546 258618 149782 258854
rect 149866 258618 150102 258854
rect 149546 222938 149782 223174
rect 149866 222938 150102 223174
rect 149546 222618 149782 222854
rect 149866 222618 150102 222854
rect 149546 186938 149782 187174
rect 149866 186938 150102 187174
rect 149546 186618 149782 186854
rect 149866 186618 150102 186854
rect 149546 150938 149782 151174
rect 149866 150938 150102 151174
rect 149546 150618 149782 150854
rect 149866 150618 150102 150854
rect 149546 114938 149782 115174
rect 149866 114938 150102 115174
rect 149546 114618 149782 114854
rect 149866 114618 150102 114854
rect 149546 78938 149782 79174
rect 149866 78938 150102 79174
rect 149546 78618 149782 78854
rect 149866 78618 150102 78854
rect 149546 42938 149782 43174
rect 149866 42938 150102 43174
rect 149546 42618 149782 42854
rect 149866 42618 150102 42854
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 149546 -2502 149782 -2266
rect 149866 -2502 150102 -2266
rect 149546 -2822 149782 -2586
rect 149866 -2822 150102 -2586
rect 153266 694658 153502 694894
rect 153586 694658 153822 694894
rect 153266 694338 153502 694574
rect 153586 694338 153822 694574
rect 153266 658658 153502 658894
rect 153586 658658 153822 658894
rect 153266 658338 153502 658574
rect 153586 658338 153822 658574
rect 153266 622658 153502 622894
rect 153586 622658 153822 622894
rect 153266 622338 153502 622574
rect 153586 622338 153822 622574
rect 153266 586658 153502 586894
rect 153586 586658 153822 586894
rect 153266 586338 153502 586574
rect 153586 586338 153822 586574
rect 153266 550658 153502 550894
rect 153586 550658 153822 550894
rect 153266 550338 153502 550574
rect 153586 550338 153822 550574
rect 153266 514658 153502 514894
rect 153586 514658 153822 514894
rect 153266 514338 153502 514574
rect 153586 514338 153822 514574
rect 153266 478658 153502 478894
rect 153586 478658 153822 478894
rect 153266 478338 153502 478574
rect 153586 478338 153822 478574
rect 153266 442658 153502 442894
rect 153586 442658 153822 442894
rect 153266 442338 153502 442574
rect 153586 442338 153822 442574
rect 153266 406658 153502 406894
rect 153586 406658 153822 406894
rect 153266 406338 153502 406574
rect 153586 406338 153822 406574
rect 153266 370658 153502 370894
rect 153586 370658 153822 370894
rect 153266 370338 153502 370574
rect 153586 370338 153822 370574
rect 153266 334658 153502 334894
rect 153586 334658 153822 334894
rect 153266 334338 153502 334574
rect 153586 334338 153822 334574
rect 153266 298658 153502 298894
rect 153586 298658 153822 298894
rect 153266 298338 153502 298574
rect 153586 298338 153822 298574
rect 153266 262658 153502 262894
rect 153586 262658 153822 262894
rect 153266 262338 153502 262574
rect 153586 262338 153822 262574
rect 153266 226658 153502 226894
rect 153586 226658 153822 226894
rect 153266 226338 153502 226574
rect 153586 226338 153822 226574
rect 153266 190658 153502 190894
rect 153586 190658 153822 190894
rect 153266 190338 153502 190574
rect 153586 190338 153822 190574
rect 153266 154658 153502 154894
rect 153586 154658 153822 154894
rect 153266 154338 153502 154574
rect 153586 154338 153822 154574
rect 153266 118658 153502 118894
rect 153586 118658 153822 118894
rect 153266 118338 153502 118574
rect 153586 118338 153822 118574
rect 153266 82658 153502 82894
rect 153586 82658 153822 82894
rect 153266 82338 153502 82574
rect 153586 82338 153822 82574
rect 153266 46658 153502 46894
rect 153586 46658 153822 46894
rect 153266 46338 153502 46574
rect 153586 46338 153822 46574
rect 153266 10658 153502 10894
rect 153586 10658 153822 10894
rect 153266 10338 153502 10574
rect 153586 10338 153822 10574
rect 153266 -4422 153502 -4186
rect 153586 -4422 153822 -4186
rect 153266 -4742 153502 -4506
rect 153586 -4742 153822 -4506
rect 174986 711322 175222 711558
rect 175306 711322 175542 711558
rect 174986 711002 175222 711238
rect 175306 711002 175542 711238
rect 171266 709402 171502 709638
rect 171586 709402 171822 709638
rect 171266 709082 171502 709318
rect 171586 709082 171822 709318
rect 167546 707482 167782 707718
rect 167866 707482 168102 707718
rect 167546 707162 167782 707398
rect 167866 707162 168102 707398
rect 156986 698378 157222 698614
rect 157306 698378 157542 698614
rect 156986 698058 157222 698294
rect 157306 698058 157542 698294
rect 156986 662378 157222 662614
rect 157306 662378 157542 662614
rect 156986 662058 157222 662294
rect 157306 662058 157542 662294
rect 156986 626378 157222 626614
rect 157306 626378 157542 626614
rect 156986 626058 157222 626294
rect 157306 626058 157542 626294
rect 156986 590378 157222 590614
rect 157306 590378 157542 590614
rect 156986 590058 157222 590294
rect 157306 590058 157542 590294
rect 156986 554378 157222 554614
rect 157306 554378 157542 554614
rect 156986 554058 157222 554294
rect 157306 554058 157542 554294
rect 156986 518378 157222 518614
rect 157306 518378 157542 518614
rect 156986 518058 157222 518294
rect 157306 518058 157542 518294
rect 156986 482378 157222 482614
rect 157306 482378 157542 482614
rect 156986 482058 157222 482294
rect 157306 482058 157542 482294
rect 156986 446378 157222 446614
rect 157306 446378 157542 446614
rect 156986 446058 157222 446294
rect 157306 446058 157542 446294
rect 156986 410378 157222 410614
rect 157306 410378 157542 410614
rect 156986 410058 157222 410294
rect 157306 410058 157542 410294
rect 156986 374378 157222 374614
rect 157306 374378 157542 374614
rect 156986 374058 157222 374294
rect 157306 374058 157542 374294
rect 156986 338378 157222 338614
rect 157306 338378 157542 338614
rect 156986 338058 157222 338294
rect 157306 338058 157542 338294
rect 156986 302378 157222 302614
rect 157306 302378 157542 302614
rect 156986 302058 157222 302294
rect 157306 302058 157542 302294
rect 156986 266378 157222 266614
rect 157306 266378 157542 266614
rect 156986 266058 157222 266294
rect 157306 266058 157542 266294
rect 156986 230378 157222 230614
rect 157306 230378 157542 230614
rect 156986 230058 157222 230294
rect 157306 230058 157542 230294
rect 156986 194378 157222 194614
rect 157306 194378 157542 194614
rect 156986 194058 157222 194294
rect 157306 194058 157542 194294
rect 163826 705562 164062 705798
rect 164146 705562 164382 705798
rect 163826 705242 164062 705478
rect 164146 705242 164382 705478
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 163826 561218 164062 561454
rect 164146 561218 164382 561454
rect 163826 560898 164062 561134
rect 164146 560898 164382 561134
rect 163826 525218 164062 525454
rect 164146 525218 164382 525454
rect 163826 524898 164062 525134
rect 164146 524898 164382 525134
rect 163826 489218 164062 489454
rect 164146 489218 164382 489454
rect 163826 488898 164062 489134
rect 164146 488898 164382 489134
rect 163826 453218 164062 453454
rect 164146 453218 164382 453454
rect 163826 452898 164062 453134
rect 164146 452898 164382 453134
rect 163826 417218 164062 417454
rect 164146 417218 164382 417454
rect 163826 416898 164062 417134
rect 164146 416898 164382 417134
rect 163826 381218 164062 381454
rect 164146 381218 164382 381454
rect 163826 380898 164062 381134
rect 164146 380898 164382 381134
rect 163826 345218 164062 345454
rect 164146 345218 164382 345454
rect 163826 344898 164062 345134
rect 164146 344898 164382 345134
rect 163826 309218 164062 309454
rect 164146 309218 164382 309454
rect 163826 308898 164062 309134
rect 164146 308898 164382 309134
rect 163826 273218 164062 273454
rect 164146 273218 164382 273454
rect 163826 272898 164062 273134
rect 164146 272898 164382 273134
rect 163826 237218 164062 237454
rect 164146 237218 164382 237454
rect 163826 236898 164062 237134
rect 164146 236898 164382 237134
rect 163826 201218 164062 201454
rect 164146 201218 164382 201454
rect 163826 200898 164062 201134
rect 164146 200898 164382 201134
rect 167546 672938 167782 673174
rect 167866 672938 168102 673174
rect 167546 672618 167782 672854
rect 167866 672618 168102 672854
rect 167546 636938 167782 637174
rect 167866 636938 168102 637174
rect 167546 636618 167782 636854
rect 167866 636618 168102 636854
rect 167546 600938 167782 601174
rect 167866 600938 168102 601174
rect 167546 600618 167782 600854
rect 167866 600618 168102 600854
rect 167546 564938 167782 565174
rect 167866 564938 168102 565174
rect 167546 564618 167782 564854
rect 167866 564618 168102 564854
rect 167546 528938 167782 529174
rect 167866 528938 168102 529174
rect 167546 528618 167782 528854
rect 167866 528618 168102 528854
rect 167546 492938 167782 493174
rect 167866 492938 168102 493174
rect 167546 492618 167782 492854
rect 167866 492618 168102 492854
rect 167546 456938 167782 457174
rect 167866 456938 168102 457174
rect 167546 456618 167782 456854
rect 167866 456618 168102 456854
rect 167546 420938 167782 421174
rect 167866 420938 168102 421174
rect 167546 420618 167782 420854
rect 167866 420618 168102 420854
rect 167546 384938 167782 385174
rect 167866 384938 168102 385174
rect 167546 384618 167782 384854
rect 167866 384618 168102 384854
rect 167546 348938 167782 349174
rect 167866 348938 168102 349174
rect 167546 348618 167782 348854
rect 167866 348618 168102 348854
rect 167546 312938 167782 313174
rect 167866 312938 168102 313174
rect 167546 312618 167782 312854
rect 167866 312618 168102 312854
rect 167546 276938 167782 277174
rect 167866 276938 168102 277174
rect 167546 276618 167782 276854
rect 167866 276618 168102 276854
rect 167546 240938 167782 241174
rect 167866 240938 168102 241174
rect 167546 240618 167782 240854
rect 167866 240618 168102 240854
rect 167546 204938 167782 205174
rect 167866 204938 168102 205174
rect 167546 204618 167782 204854
rect 167866 204618 168102 204854
rect 171266 676658 171502 676894
rect 171586 676658 171822 676894
rect 171266 676338 171502 676574
rect 171586 676338 171822 676574
rect 171266 640658 171502 640894
rect 171586 640658 171822 640894
rect 171266 640338 171502 640574
rect 171586 640338 171822 640574
rect 171266 604658 171502 604894
rect 171586 604658 171822 604894
rect 171266 604338 171502 604574
rect 171586 604338 171822 604574
rect 171266 568658 171502 568894
rect 171586 568658 171822 568894
rect 171266 568338 171502 568574
rect 171586 568338 171822 568574
rect 171266 532658 171502 532894
rect 171586 532658 171822 532894
rect 171266 532338 171502 532574
rect 171586 532338 171822 532574
rect 171266 496658 171502 496894
rect 171586 496658 171822 496894
rect 171266 496338 171502 496574
rect 171586 496338 171822 496574
rect 171266 460658 171502 460894
rect 171586 460658 171822 460894
rect 171266 460338 171502 460574
rect 171586 460338 171822 460574
rect 171266 424658 171502 424894
rect 171586 424658 171822 424894
rect 171266 424338 171502 424574
rect 171586 424338 171822 424574
rect 171266 388658 171502 388894
rect 171586 388658 171822 388894
rect 171266 388338 171502 388574
rect 171586 388338 171822 388574
rect 171266 352658 171502 352894
rect 171586 352658 171822 352894
rect 171266 352338 171502 352574
rect 171586 352338 171822 352574
rect 171266 316658 171502 316894
rect 171586 316658 171822 316894
rect 171266 316338 171502 316574
rect 171586 316338 171822 316574
rect 171266 280658 171502 280894
rect 171586 280658 171822 280894
rect 171266 280338 171502 280574
rect 171586 280338 171822 280574
rect 171266 244658 171502 244894
rect 171586 244658 171822 244894
rect 171266 244338 171502 244574
rect 171586 244338 171822 244574
rect 171266 208658 171502 208894
rect 171586 208658 171822 208894
rect 171266 208338 171502 208574
rect 171586 208338 171822 208574
rect 192986 710362 193222 710598
rect 193306 710362 193542 710598
rect 192986 710042 193222 710278
rect 193306 710042 193542 710278
rect 189266 708442 189502 708678
rect 189586 708442 189822 708678
rect 189266 708122 189502 708358
rect 189586 708122 189822 708358
rect 185546 706522 185782 706758
rect 185866 706522 186102 706758
rect 185546 706202 185782 706438
rect 185866 706202 186102 706438
rect 174986 680378 175222 680614
rect 175306 680378 175542 680614
rect 174986 680058 175222 680294
rect 175306 680058 175542 680294
rect 174986 644378 175222 644614
rect 175306 644378 175542 644614
rect 174986 644058 175222 644294
rect 175306 644058 175542 644294
rect 174986 608378 175222 608614
rect 175306 608378 175542 608614
rect 174986 608058 175222 608294
rect 175306 608058 175542 608294
rect 174986 572378 175222 572614
rect 175306 572378 175542 572614
rect 174986 572058 175222 572294
rect 175306 572058 175542 572294
rect 174986 536378 175222 536614
rect 175306 536378 175542 536614
rect 174986 536058 175222 536294
rect 175306 536058 175542 536294
rect 174986 500378 175222 500614
rect 175306 500378 175542 500614
rect 174986 500058 175222 500294
rect 175306 500058 175542 500294
rect 174986 464378 175222 464614
rect 175306 464378 175542 464614
rect 174986 464058 175222 464294
rect 175306 464058 175542 464294
rect 174986 428378 175222 428614
rect 175306 428378 175542 428614
rect 174986 428058 175222 428294
rect 175306 428058 175542 428294
rect 174986 392378 175222 392614
rect 175306 392378 175542 392614
rect 174986 392058 175222 392294
rect 175306 392058 175542 392294
rect 174986 356378 175222 356614
rect 175306 356378 175542 356614
rect 174986 356058 175222 356294
rect 175306 356058 175542 356294
rect 174986 320378 175222 320614
rect 175306 320378 175542 320614
rect 174986 320058 175222 320294
rect 175306 320058 175542 320294
rect 174986 284378 175222 284614
rect 175306 284378 175542 284614
rect 174986 284058 175222 284294
rect 175306 284058 175542 284294
rect 174986 248378 175222 248614
rect 175306 248378 175542 248614
rect 174986 248058 175222 248294
rect 175306 248058 175542 248294
rect 174986 212378 175222 212614
rect 175306 212378 175542 212614
rect 174986 212058 175222 212294
rect 175306 212058 175542 212294
rect 162285 183218 162521 183454
rect 162285 182898 162521 183134
rect 164882 183218 165118 183454
rect 164882 182898 165118 183134
rect 167479 183218 167715 183454
rect 167479 182898 167715 183134
rect 174986 176378 175222 176614
rect 175306 176378 175542 176614
rect 174986 176058 175222 176294
rect 175306 176058 175542 176294
rect 163583 165218 163819 165454
rect 163583 164898 163819 165134
rect 166180 165218 166416 165454
rect 166180 164898 166416 165134
rect 156986 158378 157222 158614
rect 157306 158378 157542 158614
rect 156986 158058 157222 158294
rect 157306 158058 157542 158294
rect 162285 147218 162521 147454
rect 162285 146898 162521 147134
rect 164882 147218 165118 147454
rect 164882 146898 165118 147134
rect 167479 147218 167715 147454
rect 167479 146898 167715 147134
rect 174986 140378 175222 140614
rect 175306 140378 175542 140614
rect 174986 140058 175222 140294
rect 175306 140058 175542 140294
rect 163583 129218 163819 129454
rect 163583 128898 163819 129134
rect 166180 129218 166416 129454
rect 166180 128898 166416 129134
rect 156986 122378 157222 122614
rect 157306 122378 157542 122614
rect 156986 122058 157222 122294
rect 157306 122058 157542 122294
rect 156986 86378 157222 86614
rect 157306 86378 157542 86614
rect 156986 86058 157222 86294
rect 157306 86058 157542 86294
rect 156986 50378 157222 50614
rect 157306 50378 157542 50614
rect 156986 50058 157222 50294
rect 157306 50058 157542 50294
rect 156986 14378 157222 14614
rect 157306 14378 157542 14614
rect 156986 14058 157222 14294
rect 157306 14058 157542 14294
rect 138986 -7302 139222 -7066
rect 139306 -7302 139542 -7066
rect 138986 -7622 139222 -7386
rect 139306 -7622 139542 -7386
rect 163826 93218 164062 93454
rect 164146 93218 164382 93454
rect 163826 92898 164062 93134
rect 164146 92898 164382 93134
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -1542 164062 -1306
rect 164146 -1542 164382 -1306
rect 163826 -1862 164062 -1626
rect 164146 -1862 164382 -1626
rect 167546 96938 167782 97174
rect 167866 96938 168102 97174
rect 167546 96618 167782 96854
rect 167866 96618 168102 96854
rect 167546 60938 167782 61174
rect 167866 60938 168102 61174
rect 167546 60618 167782 60854
rect 167866 60618 168102 60854
rect 167546 24938 167782 25174
rect 167866 24938 168102 25174
rect 167546 24618 167782 24854
rect 167866 24618 168102 24854
rect 167546 -3462 167782 -3226
rect 167866 -3462 168102 -3226
rect 167546 -3782 167782 -3546
rect 167866 -3782 168102 -3546
rect 171266 100658 171502 100894
rect 171586 100658 171822 100894
rect 171266 100338 171502 100574
rect 171586 100338 171822 100574
rect 171266 64658 171502 64894
rect 171586 64658 171822 64894
rect 171266 64338 171502 64574
rect 171586 64338 171822 64574
rect 171266 28658 171502 28894
rect 171586 28658 171822 28894
rect 171266 28338 171502 28574
rect 171586 28338 171822 28574
rect 171266 -5382 171502 -5146
rect 171586 -5382 171822 -5146
rect 171266 -5702 171502 -5466
rect 171586 -5702 171822 -5466
rect 174986 104378 175222 104614
rect 175306 104378 175542 104614
rect 174986 104058 175222 104294
rect 175306 104058 175542 104294
rect 174986 68378 175222 68614
rect 175306 68378 175542 68614
rect 174986 68058 175222 68294
rect 175306 68058 175542 68294
rect 174986 32378 175222 32614
rect 175306 32378 175542 32614
rect 174986 32058 175222 32294
rect 175306 32058 175542 32294
rect 156986 -6342 157222 -6106
rect 157306 -6342 157542 -6106
rect 156986 -6662 157222 -6426
rect 157306 -6662 157542 -6426
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 181826 435218 182062 435454
rect 182146 435218 182382 435454
rect 181826 434898 182062 435134
rect 182146 434898 182382 435134
rect 181826 399218 182062 399454
rect 182146 399218 182382 399454
rect 181826 398898 182062 399134
rect 182146 398898 182382 399134
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 181826 327218 182062 327454
rect 182146 327218 182382 327454
rect 181826 326898 182062 327134
rect 182146 326898 182382 327134
rect 181826 291218 182062 291454
rect 182146 291218 182382 291454
rect 181826 290898 182062 291134
rect 182146 290898 182382 291134
rect 181826 255218 182062 255454
rect 182146 255218 182382 255454
rect 181826 254898 182062 255134
rect 182146 254898 182382 255134
rect 181826 219218 182062 219454
rect 182146 219218 182382 219454
rect 181826 218898 182062 219134
rect 182146 218898 182382 219134
rect 181826 183218 182062 183454
rect 182146 183218 182382 183454
rect 181826 182898 182062 183134
rect 182146 182898 182382 183134
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 181826 111218 182062 111454
rect 182146 111218 182382 111454
rect 181826 110898 182062 111134
rect 182146 110898 182382 111134
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 185546 690938 185782 691174
rect 185866 690938 186102 691174
rect 185546 690618 185782 690854
rect 185866 690618 186102 690854
rect 185546 654938 185782 655174
rect 185866 654938 186102 655174
rect 185546 654618 185782 654854
rect 185866 654618 186102 654854
rect 185546 618938 185782 619174
rect 185866 618938 186102 619174
rect 185546 618618 185782 618854
rect 185866 618618 186102 618854
rect 185546 582938 185782 583174
rect 185866 582938 186102 583174
rect 185546 582618 185782 582854
rect 185866 582618 186102 582854
rect 185546 546938 185782 547174
rect 185866 546938 186102 547174
rect 185546 546618 185782 546854
rect 185866 546618 186102 546854
rect 185546 510938 185782 511174
rect 185866 510938 186102 511174
rect 185546 510618 185782 510854
rect 185866 510618 186102 510854
rect 185546 474938 185782 475174
rect 185866 474938 186102 475174
rect 185546 474618 185782 474854
rect 185866 474618 186102 474854
rect 185546 438938 185782 439174
rect 185866 438938 186102 439174
rect 185546 438618 185782 438854
rect 185866 438618 186102 438854
rect 185546 402938 185782 403174
rect 185866 402938 186102 403174
rect 185546 402618 185782 402854
rect 185866 402618 186102 402854
rect 185546 366938 185782 367174
rect 185866 366938 186102 367174
rect 185546 366618 185782 366854
rect 185866 366618 186102 366854
rect 185546 330938 185782 331174
rect 185866 330938 186102 331174
rect 185546 330618 185782 330854
rect 185866 330618 186102 330854
rect 185546 294938 185782 295174
rect 185866 294938 186102 295174
rect 185546 294618 185782 294854
rect 185866 294618 186102 294854
rect 185546 258938 185782 259174
rect 185866 258938 186102 259174
rect 185546 258618 185782 258854
rect 185866 258618 186102 258854
rect 185546 222938 185782 223174
rect 185866 222938 186102 223174
rect 185546 222618 185782 222854
rect 185866 222618 186102 222854
rect 185546 186938 185782 187174
rect 185866 186938 186102 187174
rect 185546 186618 185782 186854
rect 185866 186618 186102 186854
rect 185546 150938 185782 151174
rect 185866 150938 186102 151174
rect 185546 150618 185782 150854
rect 185866 150618 186102 150854
rect 185546 114938 185782 115174
rect 185866 114938 186102 115174
rect 185546 114618 185782 114854
rect 185866 114618 186102 114854
rect 185546 78938 185782 79174
rect 185866 78938 186102 79174
rect 185546 78618 185782 78854
rect 185866 78618 186102 78854
rect 185546 42938 185782 43174
rect 185866 42938 186102 43174
rect 185546 42618 185782 42854
rect 185866 42618 186102 42854
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 185546 -2502 185782 -2266
rect 185866 -2502 186102 -2266
rect 185546 -2822 185782 -2586
rect 185866 -2822 186102 -2586
rect 189266 694658 189502 694894
rect 189586 694658 189822 694894
rect 189266 694338 189502 694574
rect 189586 694338 189822 694574
rect 189266 658658 189502 658894
rect 189586 658658 189822 658894
rect 189266 658338 189502 658574
rect 189586 658338 189822 658574
rect 189266 622658 189502 622894
rect 189586 622658 189822 622894
rect 189266 622338 189502 622574
rect 189586 622338 189822 622574
rect 189266 586658 189502 586894
rect 189586 586658 189822 586894
rect 189266 586338 189502 586574
rect 189586 586338 189822 586574
rect 189266 550658 189502 550894
rect 189586 550658 189822 550894
rect 189266 550338 189502 550574
rect 189586 550338 189822 550574
rect 189266 514658 189502 514894
rect 189586 514658 189822 514894
rect 189266 514338 189502 514574
rect 189586 514338 189822 514574
rect 189266 478658 189502 478894
rect 189586 478658 189822 478894
rect 189266 478338 189502 478574
rect 189586 478338 189822 478574
rect 189266 442658 189502 442894
rect 189586 442658 189822 442894
rect 189266 442338 189502 442574
rect 189586 442338 189822 442574
rect 189266 406658 189502 406894
rect 189586 406658 189822 406894
rect 189266 406338 189502 406574
rect 189586 406338 189822 406574
rect 189266 370658 189502 370894
rect 189586 370658 189822 370894
rect 189266 370338 189502 370574
rect 189586 370338 189822 370574
rect 189266 334658 189502 334894
rect 189586 334658 189822 334894
rect 189266 334338 189502 334574
rect 189586 334338 189822 334574
rect 189266 298658 189502 298894
rect 189586 298658 189822 298894
rect 189266 298338 189502 298574
rect 189586 298338 189822 298574
rect 189266 262658 189502 262894
rect 189586 262658 189822 262894
rect 189266 262338 189502 262574
rect 189586 262338 189822 262574
rect 189266 226658 189502 226894
rect 189586 226658 189822 226894
rect 189266 226338 189502 226574
rect 189586 226338 189822 226574
rect 189266 190658 189502 190894
rect 189586 190658 189822 190894
rect 189266 190338 189502 190574
rect 189586 190338 189822 190574
rect 189266 154658 189502 154894
rect 189586 154658 189822 154894
rect 189266 154338 189502 154574
rect 189586 154338 189822 154574
rect 189266 118658 189502 118894
rect 189586 118658 189822 118894
rect 189266 118338 189502 118574
rect 189586 118338 189822 118574
rect 189266 82658 189502 82894
rect 189586 82658 189822 82894
rect 189266 82338 189502 82574
rect 189586 82338 189822 82574
rect 189266 46658 189502 46894
rect 189586 46658 189822 46894
rect 189266 46338 189502 46574
rect 189586 46338 189822 46574
rect 189266 10658 189502 10894
rect 189586 10658 189822 10894
rect 189266 10338 189502 10574
rect 189586 10338 189822 10574
rect 189266 -4422 189502 -4186
rect 189586 -4422 189822 -4186
rect 189266 -4742 189502 -4506
rect 189586 -4742 189822 -4506
rect 210986 711322 211222 711558
rect 211306 711322 211542 711558
rect 210986 711002 211222 711238
rect 211306 711002 211542 711238
rect 207266 709402 207502 709638
rect 207586 709402 207822 709638
rect 207266 709082 207502 709318
rect 207586 709082 207822 709318
rect 203546 707482 203782 707718
rect 203866 707482 204102 707718
rect 203546 707162 203782 707398
rect 203866 707162 204102 707398
rect 192986 698378 193222 698614
rect 193306 698378 193542 698614
rect 192986 698058 193222 698294
rect 193306 698058 193542 698294
rect 192986 662378 193222 662614
rect 193306 662378 193542 662614
rect 192986 662058 193222 662294
rect 193306 662058 193542 662294
rect 192986 626378 193222 626614
rect 193306 626378 193542 626614
rect 192986 626058 193222 626294
rect 193306 626058 193542 626294
rect 192986 590378 193222 590614
rect 193306 590378 193542 590614
rect 192986 590058 193222 590294
rect 193306 590058 193542 590294
rect 192986 554378 193222 554614
rect 193306 554378 193542 554614
rect 192986 554058 193222 554294
rect 193306 554058 193542 554294
rect 192986 518378 193222 518614
rect 193306 518378 193542 518614
rect 192986 518058 193222 518294
rect 193306 518058 193542 518294
rect 192986 482378 193222 482614
rect 193306 482378 193542 482614
rect 192986 482058 193222 482294
rect 193306 482058 193542 482294
rect 192986 446378 193222 446614
rect 193306 446378 193542 446614
rect 192986 446058 193222 446294
rect 193306 446058 193542 446294
rect 192986 410378 193222 410614
rect 193306 410378 193542 410614
rect 192986 410058 193222 410294
rect 193306 410058 193542 410294
rect 192986 374378 193222 374614
rect 193306 374378 193542 374614
rect 192986 374058 193222 374294
rect 193306 374058 193542 374294
rect 192986 338378 193222 338614
rect 193306 338378 193542 338614
rect 192986 338058 193222 338294
rect 193306 338058 193542 338294
rect 192986 302378 193222 302614
rect 193306 302378 193542 302614
rect 192986 302058 193222 302294
rect 193306 302058 193542 302294
rect 199826 705562 200062 705798
rect 200146 705562 200382 705798
rect 199826 705242 200062 705478
rect 200146 705242 200382 705478
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 199826 561218 200062 561454
rect 200146 561218 200382 561454
rect 199826 560898 200062 561134
rect 200146 560898 200382 561134
rect 199826 525218 200062 525454
rect 200146 525218 200382 525454
rect 199826 524898 200062 525134
rect 200146 524898 200382 525134
rect 199826 489218 200062 489454
rect 200146 489218 200382 489454
rect 199826 488898 200062 489134
rect 200146 488898 200382 489134
rect 199826 453218 200062 453454
rect 200146 453218 200382 453454
rect 199826 452898 200062 453134
rect 200146 452898 200382 453134
rect 199826 417218 200062 417454
rect 200146 417218 200382 417454
rect 199826 416898 200062 417134
rect 200146 416898 200382 417134
rect 199826 381218 200062 381454
rect 200146 381218 200382 381454
rect 199826 380898 200062 381134
rect 200146 380898 200382 381134
rect 199826 345218 200062 345454
rect 200146 345218 200382 345454
rect 199826 344898 200062 345134
rect 200146 344898 200382 345134
rect 199826 309218 200062 309454
rect 200146 309218 200382 309454
rect 199826 308898 200062 309134
rect 200146 308898 200382 309134
rect 203546 672938 203782 673174
rect 203866 672938 204102 673174
rect 203546 672618 203782 672854
rect 203866 672618 204102 672854
rect 203546 636938 203782 637174
rect 203866 636938 204102 637174
rect 203546 636618 203782 636854
rect 203866 636618 204102 636854
rect 203546 600938 203782 601174
rect 203866 600938 204102 601174
rect 203546 600618 203782 600854
rect 203866 600618 204102 600854
rect 203546 564938 203782 565174
rect 203866 564938 204102 565174
rect 203546 564618 203782 564854
rect 203866 564618 204102 564854
rect 203546 528938 203782 529174
rect 203866 528938 204102 529174
rect 203546 528618 203782 528854
rect 203866 528618 204102 528854
rect 203546 492938 203782 493174
rect 203866 492938 204102 493174
rect 203546 492618 203782 492854
rect 203866 492618 204102 492854
rect 203546 456938 203782 457174
rect 203866 456938 204102 457174
rect 203546 456618 203782 456854
rect 203866 456618 204102 456854
rect 203546 420938 203782 421174
rect 203866 420938 204102 421174
rect 203546 420618 203782 420854
rect 203866 420618 204102 420854
rect 203546 384938 203782 385174
rect 203866 384938 204102 385174
rect 203546 384618 203782 384854
rect 203866 384618 204102 384854
rect 203546 348938 203782 349174
rect 203866 348938 204102 349174
rect 203546 348618 203782 348854
rect 203866 348618 204102 348854
rect 203546 312938 203782 313174
rect 203866 312938 204102 313174
rect 203546 312618 203782 312854
rect 203866 312618 204102 312854
rect 207266 676658 207502 676894
rect 207586 676658 207822 676894
rect 207266 676338 207502 676574
rect 207586 676338 207822 676574
rect 207266 640658 207502 640894
rect 207586 640658 207822 640894
rect 207266 640338 207502 640574
rect 207586 640338 207822 640574
rect 207266 604658 207502 604894
rect 207586 604658 207822 604894
rect 207266 604338 207502 604574
rect 207586 604338 207822 604574
rect 207266 568658 207502 568894
rect 207586 568658 207822 568894
rect 207266 568338 207502 568574
rect 207586 568338 207822 568574
rect 207266 532658 207502 532894
rect 207586 532658 207822 532894
rect 207266 532338 207502 532574
rect 207586 532338 207822 532574
rect 207266 496658 207502 496894
rect 207586 496658 207822 496894
rect 207266 496338 207502 496574
rect 207586 496338 207822 496574
rect 207266 460658 207502 460894
rect 207586 460658 207822 460894
rect 207266 460338 207502 460574
rect 207586 460338 207822 460574
rect 207266 424658 207502 424894
rect 207586 424658 207822 424894
rect 207266 424338 207502 424574
rect 207586 424338 207822 424574
rect 207266 388658 207502 388894
rect 207586 388658 207822 388894
rect 207266 388338 207502 388574
rect 207586 388338 207822 388574
rect 207266 352658 207502 352894
rect 207586 352658 207822 352894
rect 207266 352338 207502 352574
rect 207586 352338 207822 352574
rect 207266 316658 207502 316894
rect 207586 316658 207822 316894
rect 207266 316338 207502 316574
rect 207586 316338 207822 316574
rect 228986 710362 229222 710598
rect 229306 710362 229542 710598
rect 228986 710042 229222 710278
rect 229306 710042 229542 710278
rect 225266 708442 225502 708678
rect 225586 708442 225822 708678
rect 225266 708122 225502 708358
rect 225586 708122 225822 708358
rect 221546 706522 221782 706758
rect 221866 706522 222102 706758
rect 221546 706202 221782 706438
rect 221866 706202 222102 706438
rect 210986 680378 211222 680614
rect 211306 680378 211542 680614
rect 210986 680058 211222 680294
rect 211306 680058 211542 680294
rect 210986 644378 211222 644614
rect 211306 644378 211542 644614
rect 210986 644058 211222 644294
rect 211306 644058 211542 644294
rect 210986 608378 211222 608614
rect 211306 608378 211542 608614
rect 210986 608058 211222 608294
rect 211306 608058 211542 608294
rect 210986 572378 211222 572614
rect 211306 572378 211542 572614
rect 210986 572058 211222 572294
rect 211306 572058 211542 572294
rect 210986 536378 211222 536614
rect 211306 536378 211542 536614
rect 210986 536058 211222 536294
rect 211306 536058 211542 536294
rect 210986 500378 211222 500614
rect 211306 500378 211542 500614
rect 210986 500058 211222 500294
rect 211306 500058 211542 500294
rect 210986 464378 211222 464614
rect 211306 464378 211542 464614
rect 210986 464058 211222 464294
rect 211306 464058 211542 464294
rect 210986 428378 211222 428614
rect 211306 428378 211542 428614
rect 210986 428058 211222 428294
rect 211306 428058 211542 428294
rect 210986 392378 211222 392614
rect 211306 392378 211542 392614
rect 210986 392058 211222 392294
rect 211306 392058 211542 392294
rect 210986 356378 211222 356614
rect 211306 356378 211542 356614
rect 210986 356058 211222 356294
rect 211306 356058 211542 356294
rect 210986 320378 211222 320614
rect 211306 320378 211542 320614
rect 210986 320058 211222 320294
rect 211306 320058 211542 320294
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 217826 543218 218062 543454
rect 218146 543218 218382 543454
rect 217826 542898 218062 543134
rect 218146 542898 218382 543134
rect 217826 507218 218062 507454
rect 218146 507218 218382 507454
rect 217826 506898 218062 507134
rect 218146 506898 218382 507134
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 217826 435218 218062 435454
rect 218146 435218 218382 435454
rect 217826 434898 218062 435134
rect 218146 434898 218382 435134
rect 217826 399218 218062 399454
rect 218146 399218 218382 399454
rect 217826 398898 218062 399134
rect 218146 398898 218382 399134
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 217826 327218 218062 327454
rect 218146 327218 218382 327454
rect 217826 326898 218062 327134
rect 218146 326898 218382 327134
rect 221546 690938 221782 691174
rect 221866 690938 222102 691174
rect 221546 690618 221782 690854
rect 221866 690618 222102 690854
rect 221546 654938 221782 655174
rect 221866 654938 222102 655174
rect 221546 654618 221782 654854
rect 221866 654618 222102 654854
rect 221546 618938 221782 619174
rect 221866 618938 222102 619174
rect 221546 618618 221782 618854
rect 221866 618618 222102 618854
rect 221546 582938 221782 583174
rect 221866 582938 222102 583174
rect 221546 582618 221782 582854
rect 221866 582618 222102 582854
rect 221546 546938 221782 547174
rect 221866 546938 222102 547174
rect 221546 546618 221782 546854
rect 221866 546618 222102 546854
rect 221546 510938 221782 511174
rect 221866 510938 222102 511174
rect 221546 510618 221782 510854
rect 221866 510618 222102 510854
rect 221546 474938 221782 475174
rect 221866 474938 222102 475174
rect 221546 474618 221782 474854
rect 221866 474618 222102 474854
rect 221546 438938 221782 439174
rect 221866 438938 222102 439174
rect 221546 438618 221782 438854
rect 221866 438618 222102 438854
rect 221546 402938 221782 403174
rect 221866 402938 222102 403174
rect 221546 402618 221782 402854
rect 221866 402618 222102 402854
rect 221546 366938 221782 367174
rect 221866 366938 222102 367174
rect 221546 366618 221782 366854
rect 221866 366618 222102 366854
rect 221546 330938 221782 331174
rect 221866 330938 222102 331174
rect 221546 330618 221782 330854
rect 221866 330618 222102 330854
rect 225266 694658 225502 694894
rect 225586 694658 225822 694894
rect 225266 694338 225502 694574
rect 225586 694338 225822 694574
rect 225266 658658 225502 658894
rect 225586 658658 225822 658894
rect 225266 658338 225502 658574
rect 225586 658338 225822 658574
rect 225266 622658 225502 622894
rect 225586 622658 225822 622894
rect 225266 622338 225502 622574
rect 225586 622338 225822 622574
rect 225266 586658 225502 586894
rect 225586 586658 225822 586894
rect 225266 586338 225502 586574
rect 225586 586338 225822 586574
rect 225266 550658 225502 550894
rect 225586 550658 225822 550894
rect 225266 550338 225502 550574
rect 225586 550338 225822 550574
rect 225266 514658 225502 514894
rect 225586 514658 225822 514894
rect 225266 514338 225502 514574
rect 225586 514338 225822 514574
rect 225266 478658 225502 478894
rect 225586 478658 225822 478894
rect 225266 478338 225502 478574
rect 225586 478338 225822 478574
rect 225266 442658 225502 442894
rect 225586 442658 225822 442894
rect 225266 442338 225502 442574
rect 225586 442338 225822 442574
rect 225266 406658 225502 406894
rect 225586 406658 225822 406894
rect 225266 406338 225502 406574
rect 225586 406338 225822 406574
rect 225266 370658 225502 370894
rect 225586 370658 225822 370894
rect 225266 370338 225502 370574
rect 225586 370338 225822 370574
rect 225266 334658 225502 334894
rect 225586 334658 225822 334894
rect 225266 334338 225502 334574
rect 225586 334338 225822 334574
rect 246986 711322 247222 711558
rect 247306 711322 247542 711558
rect 246986 711002 247222 711238
rect 247306 711002 247542 711238
rect 243266 709402 243502 709638
rect 243586 709402 243822 709638
rect 243266 709082 243502 709318
rect 243586 709082 243822 709318
rect 239546 707482 239782 707718
rect 239866 707482 240102 707718
rect 239546 707162 239782 707398
rect 239866 707162 240102 707398
rect 228986 698378 229222 698614
rect 229306 698378 229542 698614
rect 228986 698058 229222 698294
rect 229306 698058 229542 698294
rect 228986 662378 229222 662614
rect 229306 662378 229542 662614
rect 228986 662058 229222 662294
rect 229306 662058 229542 662294
rect 228986 626378 229222 626614
rect 229306 626378 229542 626614
rect 228986 626058 229222 626294
rect 229306 626058 229542 626294
rect 228986 590378 229222 590614
rect 229306 590378 229542 590614
rect 228986 590058 229222 590294
rect 229306 590058 229542 590294
rect 228986 554378 229222 554614
rect 229306 554378 229542 554614
rect 228986 554058 229222 554294
rect 229306 554058 229542 554294
rect 228986 518378 229222 518614
rect 229306 518378 229542 518614
rect 228986 518058 229222 518294
rect 229306 518058 229542 518294
rect 228986 482378 229222 482614
rect 229306 482378 229542 482614
rect 228986 482058 229222 482294
rect 229306 482058 229542 482294
rect 228986 446378 229222 446614
rect 229306 446378 229542 446614
rect 228986 446058 229222 446294
rect 229306 446058 229542 446294
rect 228986 410378 229222 410614
rect 229306 410378 229542 410614
rect 228986 410058 229222 410294
rect 229306 410058 229542 410294
rect 228986 374378 229222 374614
rect 229306 374378 229542 374614
rect 228986 374058 229222 374294
rect 229306 374058 229542 374294
rect 228986 338378 229222 338614
rect 229306 338378 229542 338614
rect 228986 338058 229222 338294
rect 229306 338058 229542 338294
rect 228986 302378 229222 302614
rect 229306 302378 229542 302614
rect 228986 302058 229222 302294
rect 229306 302058 229542 302294
rect 235826 705562 236062 705798
rect 236146 705562 236382 705798
rect 235826 705242 236062 705478
rect 236146 705242 236382 705478
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 235826 561218 236062 561454
rect 236146 561218 236382 561454
rect 235826 560898 236062 561134
rect 236146 560898 236382 561134
rect 235826 525218 236062 525454
rect 236146 525218 236382 525454
rect 235826 524898 236062 525134
rect 236146 524898 236382 525134
rect 235826 489218 236062 489454
rect 236146 489218 236382 489454
rect 235826 488898 236062 489134
rect 236146 488898 236382 489134
rect 235826 453218 236062 453454
rect 236146 453218 236382 453454
rect 235826 452898 236062 453134
rect 236146 452898 236382 453134
rect 235826 417218 236062 417454
rect 236146 417218 236382 417454
rect 235826 416898 236062 417134
rect 236146 416898 236382 417134
rect 235826 381218 236062 381454
rect 236146 381218 236382 381454
rect 235826 380898 236062 381134
rect 236146 380898 236382 381134
rect 235826 345218 236062 345454
rect 236146 345218 236382 345454
rect 235826 344898 236062 345134
rect 236146 344898 236382 345134
rect 235826 309218 236062 309454
rect 236146 309218 236382 309454
rect 235826 308898 236062 309134
rect 236146 308898 236382 309134
rect 239546 672938 239782 673174
rect 239866 672938 240102 673174
rect 239546 672618 239782 672854
rect 239866 672618 240102 672854
rect 239546 636938 239782 637174
rect 239866 636938 240102 637174
rect 239546 636618 239782 636854
rect 239866 636618 240102 636854
rect 239546 600938 239782 601174
rect 239866 600938 240102 601174
rect 239546 600618 239782 600854
rect 239866 600618 240102 600854
rect 239546 564938 239782 565174
rect 239866 564938 240102 565174
rect 239546 564618 239782 564854
rect 239866 564618 240102 564854
rect 239546 528938 239782 529174
rect 239866 528938 240102 529174
rect 239546 528618 239782 528854
rect 239866 528618 240102 528854
rect 239546 492938 239782 493174
rect 239866 492938 240102 493174
rect 239546 492618 239782 492854
rect 239866 492618 240102 492854
rect 239546 456938 239782 457174
rect 239866 456938 240102 457174
rect 239546 456618 239782 456854
rect 239866 456618 240102 456854
rect 239546 420938 239782 421174
rect 239866 420938 240102 421174
rect 239546 420618 239782 420854
rect 239866 420618 240102 420854
rect 239546 384938 239782 385174
rect 239866 384938 240102 385174
rect 239546 384618 239782 384854
rect 239866 384618 240102 384854
rect 239546 348938 239782 349174
rect 239866 348938 240102 349174
rect 239546 348618 239782 348854
rect 239866 348618 240102 348854
rect 239546 312938 239782 313174
rect 239866 312938 240102 313174
rect 239546 312618 239782 312854
rect 239866 312618 240102 312854
rect 243266 676658 243502 676894
rect 243586 676658 243822 676894
rect 243266 676338 243502 676574
rect 243586 676338 243822 676574
rect 243266 640658 243502 640894
rect 243586 640658 243822 640894
rect 243266 640338 243502 640574
rect 243586 640338 243822 640574
rect 243266 604658 243502 604894
rect 243586 604658 243822 604894
rect 243266 604338 243502 604574
rect 243586 604338 243822 604574
rect 243266 568658 243502 568894
rect 243586 568658 243822 568894
rect 243266 568338 243502 568574
rect 243586 568338 243822 568574
rect 243266 532658 243502 532894
rect 243586 532658 243822 532894
rect 243266 532338 243502 532574
rect 243586 532338 243822 532574
rect 243266 496658 243502 496894
rect 243586 496658 243822 496894
rect 243266 496338 243502 496574
rect 243586 496338 243822 496574
rect 243266 460658 243502 460894
rect 243586 460658 243822 460894
rect 243266 460338 243502 460574
rect 243586 460338 243822 460574
rect 243266 424658 243502 424894
rect 243586 424658 243822 424894
rect 243266 424338 243502 424574
rect 243586 424338 243822 424574
rect 243266 388658 243502 388894
rect 243586 388658 243822 388894
rect 243266 388338 243502 388574
rect 243586 388338 243822 388574
rect 243266 352658 243502 352894
rect 243586 352658 243822 352894
rect 243266 352338 243502 352574
rect 243586 352338 243822 352574
rect 243266 316658 243502 316894
rect 243586 316658 243822 316894
rect 243266 316338 243502 316574
rect 243586 316338 243822 316574
rect 264986 710362 265222 710598
rect 265306 710362 265542 710598
rect 264986 710042 265222 710278
rect 265306 710042 265542 710278
rect 261266 708442 261502 708678
rect 261586 708442 261822 708678
rect 261266 708122 261502 708358
rect 261586 708122 261822 708358
rect 257546 706522 257782 706758
rect 257866 706522 258102 706758
rect 257546 706202 257782 706438
rect 257866 706202 258102 706438
rect 246986 680378 247222 680614
rect 247306 680378 247542 680614
rect 246986 680058 247222 680294
rect 247306 680058 247542 680294
rect 246986 644378 247222 644614
rect 247306 644378 247542 644614
rect 246986 644058 247222 644294
rect 247306 644058 247542 644294
rect 246986 608378 247222 608614
rect 247306 608378 247542 608614
rect 246986 608058 247222 608294
rect 247306 608058 247542 608294
rect 246986 572378 247222 572614
rect 247306 572378 247542 572614
rect 246986 572058 247222 572294
rect 247306 572058 247542 572294
rect 246986 536378 247222 536614
rect 247306 536378 247542 536614
rect 246986 536058 247222 536294
rect 247306 536058 247542 536294
rect 246986 500378 247222 500614
rect 247306 500378 247542 500614
rect 246986 500058 247222 500294
rect 247306 500058 247542 500294
rect 246986 464378 247222 464614
rect 247306 464378 247542 464614
rect 246986 464058 247222 464294
rect 247306 464058 247542 464294
rect 246986 428378 247222 428614
rect 247306 428378 247542 428614
rect 246986 428058 247222 428294
rect 247306 428058 247542 428294
rect 246986 392378 247222 392614
rect 247306 392378 247542 392614
rect 246986 392058 247222 392294
rect 247306 392058 247542 392294
rect 246986 356378 247222 356614
rect 247306 356378 247542 356614
rect 246986 356058 247222 356294
rect 247306 356058 247542 356294
rect 246986 320378 247222 320614
rect 247306 320378 247542 320614
rect 246986 320058 247222 320294
rect 247306 320058 247542 320294
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 253826 543218 254062 543454
rect 254146 543218 254382 543454
rect 253826 542898 254062 543134
rect 254146 542898 254382 543134
rect 253826 507218 254062 507454
rect 254146 507218 254382 507454
rect 253826 506898 254062 507134
rect 254146 506898 254382 507134
rect 253826 471218 254062 471454
rect 254146 471218 254382 471454
rect 253826 470898 254062 471134
rect 254146 470898 254382 471134
rect 253826 435218 254062 435454
rect 254146 435218 254382 435454
rect 253826 434898 254062 435134
rect 254146 434898 254382 435134
rect 253826 399218 254062 399454
rect 254146 399218 254382 399454
rect 253826 398898 254062 399134
rect 254146 398898 254382 399134
rect 253826 363218 254062 363454
rect 254146 363218 254382 363454
rect 253826 362898 254062 363134
rect 254146 362898 254382 363134
rect 253826 327218 254062 327454
rect 254146 327218 254382 327454
rect 253826 326898 254062 327134
rect 254146 326898 254382 327134
rect 257546 690938 257782 691174
rect 257866 690938 258102 691174
rect 257546 690618 257782 690854
rect 257866 690618 258102 690854
rect 257546 654938 257782 655174
rect 257866 654938 258102 655174
rect 257546 654618 257782 654854
rect 257866 654618 258102 654854
rect 257546 618938 257782 619174
rect 257866 618938 258102 619174
rect 257546 618618 257782 618854
rect 257866 618618 258102 618854
rect 257546 582938 257782 583174
rect 257866 582938 258102 583174
rect 257546 582618 257782 582854
rect 257866 582618 258102 582854
rect 257546 546938 257782 547174
rect 257866 546938 258102 547174
rect 257546 546618 257782 546854
rect 257866 546618 258102 546854
rect 257546 510938 257782 511174
rect 257866 510938 258102 511174
rect 257546 510618 257782 510854
rect 257866 510618 258102 510854
rect 257546 474938 257782 475174
rect 257866 474938 258102 475174
rect 257546 474618 257782 474854
rect 257866 474618 258102 474854
rect 257546 438938 257782 439174
rect 257866 438938 258102 439174
rect 257546 438618 257782 438854
rect 257866 438618 258102 438854
rect 257546 402938 257782 403174
rect 257866 402938 258102 403174
rect 257546 402618 257782 402854
rect 257866 402618 258102 402854
rect 257546 366938 257782 367174
rect 257866 366938 258102 367174
rect 257546 366618 257782 366854
rect 257866 366618 258102 366854
rect 257546 330938 257782 331174
rect 257866 330938 258102 331174
rect 257546 330618 257782 330854
rect 257866 330618 258102 330854
rect 261266 694658 261502 694894
rect 261586 694658 261822 694894
rect 261266 694338 261502 694574
rect 261586 694338 261822 694574
rect 261266 658658 261502 658894
rect 261586 658658 261822 658894
rect 261266 658338 261502 658574
rect 261586 658338 261822 658574
rect 261266 622658 261502 622894
rect 261586 622658 261822 622894
rect 261266 622338 261502 622574
rect 261586 622338 261822 622574
rect 261266 586658 261502 586894
rect 261586 586658 261822 586894
rect 261266 586338 261502 586574
rect 261586 586338 261822 586574
rect 261266 550658 261502 550894
rect 261586 550658 261822 550894
rect 261266 550338 261502 550574
rect 261586 550338 261822 550574
rect 261266 514658 261502 514894
rect 261586 514658 261822 514894
rect 261266 514338 261502 514574
rect 261586 514338 261822 514574
rect 261266 478658 261502 478894
rect 261586 478658 261822 478894
rect 261266 478338 261502 478574
rect 261586 478338 261822 478574
rect 261266 442658 261502 442894
rect 261586 442658 261822 442894
rect 261266 442338 261502 442574
rect 261586 442338 261822 442574
rect 261266 406658 261502 406894
rect 261586 406658 261822 406894
rect 261266 406338 261502 406574
rect 261586 406338 261822 406574
rect 261266 370658 261502 370894
rect 261586 370658 261822 370894
rect 261266 370338 261502 370574
rect 261586 370338 261822 370574
rect 261266 334658 261502 334894
rect 261586 334658 261822 334894
rect 261266 334338 261502 334574
rect 261586 334338 261822 334574
rect 282986 711322 283222 711558
rect 283306 711322 283542 711558
rect 282986 711002 283222 711238
rect 283306 711002 283542 711238
rect 279266 709402 279502 709638
rect 279586 709402 279822 709638
rect 279266 709082 279502 709318
rect 279586 709082 279822 709318
rect 275546 707482 275782 707718
rect 275866 707482 276102 707718
rect 275546 707162 275782 707398
rect 275866 707162 276102 707398
rect 264986 698378 265222 698614
rect 265306 698378 265542 698614
rect 264986 698058 265222 698294
rect 265306 698058 265542 698294
rect 264986 662378 265222 662614
rect 265306 662378 265542 662614
rect 264986 662058 265222 662294
rect 265306 662058 265542 662294
rect 264986 626378 265222 626614
rect 265306 626378 265542 626614
rect 264986 626058 265222 626294
rect 265306 626058 265542 626294
rect 264986 590378 265222 590614
rect 265306 590378 265542 590614
rect 264986 590058 265222 590294
rect 265306 590058 265542 590294
rect 264986 554378 265222 554614
rect 265306 554378 265542 554614
rect 264986 554058 265222 554294
rect 265306 554058 265542 554294
rect 264986 518378 265222 518614
rect 265306 518378 265542 518614
rect 264986 518058 265222 518294
rect 265306 518058 265542 518294
rect 264986 482378 265222 482614
rect 265306 482378 265542 482614
rect 264986 482058 265222 482294
rect 265306 482058 265542 482294
rect 264986 446378 265222 446614
rect 265306 446378 265542 446614
rect 264986 446058 265222 446294
rect 265306 446058 265542 446294
rect 264986 410378 265222 410614
rect 265306 410378 265542 410614
rect 264986 410058 265222 410294
rect 265306 410058 265542 410294
rect 264986 374378 265222 374614
rect 265306 374378 265542 374614
rect 264986 374058 265222 374294
rect 265306 374058 265542 374294
rect 264986 338378 265222 338614
rect 265306 338378 265542 338614
rect 264986 338058 265222 338294
rect 265306 338058 265542 338294
rect 264986 302378 265222 302614
rect 265306 302378 265542 302614
rect 264986 302058 265222 302294
rect 265306 302058 265542 302294
rect 271826 705562 272062 705798
rect 272146 705562 272382 705798
rect 271826 705242 272062 705478
rect 272146 705242 272382 705478
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 271826 561218 272062 561454
rect 272146 561218 272382 561454
rect 271826 560898 272062 561134
rect 272146 560898 272382 561134
rect 271826 525218 272062 525454
rect 272146 525218 272382 525454
rect 271826 524898 272062 525134
rect 272146 524898 272382 525134
rect 271826 489218 272062 489454
rect 272146 489218 272382 489454
rect 271826 488898 272062 489134
rect 272146 488898 272382 489134
rect 271826 453218 272062 453454
rect 272146 453218 272382 453454
rect 271826 452898 272062 453134
rect 272146 452898 272382 453134
rect 271826 417218 272062 417454
rect 272146 417218 272382 417454
rect 271826 416898 272062 417134
rect 272146 416898 272382 417134
rect 271826 381218 272062 381454
rect 272146 381218 272382 381454
rect 271826 380898 272062 381134
rect 272146 380898 272382 381134
rect 271826 345218 272062 345454
rect 272146 345218 272382 345454
rect 271826 344898 272062 345134
rect 272146 344898 272382 345134
rect 271826 309218 272062 309454
rect 272146 309218 272382 309454
rect 271826 308898 272062 309134
rect 272146 308898 272382 309134
rect 275546 672938 275782 673174
rect 275866 672938 276102 673174
rect 275546 672618 275782 672854
rect 275866 672618 276102 672854
rect 275546 636938 275782 637174
rect 275866 636938 276102 637174
rect 275546 636618 275782 636854
rect 275866 636618 276102 636854
rect 275546 600938 275782 601174
rect 275866 600938 276102 601174
rect 275546 600618 275782 600854
rect 275866 600618 276102 600854
rect 275546 564938 275782 565174
rect 275866 564938 276102 565174
rect 275546 564618 275782 564854
rect 275866 564618 276102 564854
rect 275546 528938 275782 529174
rect 275866 528938 276102 529174
rect 275546 528618 275782 528854
rect 275866 528618 276102 528854
rect 275546 492938 275782 493174
rect 275866 492938 276102 493174
rect 275546 492618 275782 492854
rect 275866 492618 276102 492854
rect 275546 456938 275782 457174
rect 275866 456938 276102 457174
rect 275546 456618 275782 456854
rect 275866 456618 276102 456854
rect 275546 420938 275782 421174
rect 275866 420938 276102 421174
rect 275546 420618 275782 420854
rect 275866 420618 276102 420854
rect 275546 384938 275782 385174
rect 275866 384938 276102 385174
rect 275546 384618 275782 384854
rect 275866 384618 276102 384854
rect 275546 348938 275782 349174
rect 275866 348938 276102 349174
rect 275546 348618 275782 348854
rect 275866 348618 276102 348854
rect 275546 312938 275782 313174
rect 275866 312938 276102 313174
rect 275546 312618 275782 312854
rect 275866 312618 276102 312854
rect 279266 676658 279502 676894
rect 279586 676658 279822 676894
rect 279266 676338 279502 676574
rect 279586 676338 279822 676574
rect 279266 640658 279502 640894
rect 279586 640658 279822 640894
rect 279266 640338 279502 640574
rect 279586 640338 279822 640574
rect 279266 604658 279502 604894
rect 279586 604658 279822 604894
rect 279266 604338 279502 604574
rect 279586 604338 279822 604574
rect 279266 568658 279502 568894
rect 279586 568658 279822 568894
rect 279266 568338 279502 568574
rect 279586 568338 279822 568574
rect 279266 532658 279502 532894
rect 279586 532658 279822 532894
rect 279266 532338 279502 532574
rect 279586 532338 279822 532574
rect 279266 496658 279502 496894
rect 279586 496658 279822 496894
rect 279266 496338 279502 496574
rect 279586 496338 279822 496574
rect 279266 460658 279502 460894
rect 279586 460658 279822 460894
rect 279266 460338 279502 460574
rect 279586 460338 279822 460574
rect 279266 424658 279502 424894
rect 279586 424658 279822 424894
rect 279266 424338 279502 424574
rect 279586 424338 279822 424574
rect 279266 388658 279502 388894
rect 279586 388658 279822 388894
rect 279266 388338 279502 388574
rect 279586 388338 279822 388574
rect 279266 352658 279502 352894
rect 279586 352658 279822 352894
rect 279266 352338 279502 352574
rect 279586 352338 279822 352574
rect 279266 316658 279502 316894
rect 279586 316658 279822 316894
rect 279266 316338 279502 316574
rect 279586 316338 279822 316574
rect 300986 710362 301222 710598
rect 301306 710362 301542 710598
rect 300986 710042 301222 710278
rect 301306 710042 301542 710278
rect 297266 708442 297502 708678
rect 297586 708442 297822 708678
rect 297266 708122 297502 708358
rect 297586 708122 297822 708358
rect 293546 706522 293782 706758
rect 293866 706522 294102 706758
rect 293546 706202 293782 706438
rect 293866 706202 294102 706438
rect 282986 680378 283222 680614
rect 283306 680378 283542 680614
rect 282986 680058 283222 680294
rect 283306 680058 283542 680294
rect 282986 644378 283222 644614
rect 283306 644378 283542 644614
rect 282986 644058 283222 644294
rect 283306 644058 283542 644294
rect 282986 608378 283222 608614
rect 283306 608378 283542 608614
rect 282986 608058 283222 608294
rect 283306 608058 283542 608294
rect 282986 572378 283222 572614
rect 283306 572378 283542 572614
rect 282986 572058 283222 572294
rect 283306 572058 283542 572294
rect 282986 536378 283222 536614
rect 283306 536378 283542 536614
rect 282986 536058 283222 536294
rect 283306 536058 283542 536294
rect 282986 500378 283222 500614
rect 283306 500378 283542 500614
rect 282986 500058 283222 500294
rect 283306 500058 283542 500294
rect 282986 464378 283222 464614
rect 283306 464378 283542 464614
rect 282986 464058 283222 464294
rect 283306 464058 283542 464294
rect 282986 428378 283222 428614
rect 283306 428378 283542 428614
rect 282986 428058 283222 428294
rect 283306 428058 283542 428294
rect 282986 392378 283222 392614
rect 283306 392378 283542 392614
rect 282986 392058 283222 392294
rect 283306 392058 283542 392294
rect 282986 356378 283222 356614
rect 283306 356378 283542 356614
rect 282986 356058 283222 356294
rect 283306 356058 283542 356294
rect 282986 320378 283222 320614
rect 283306 320378 283542 320614
rect 282986 320058 283222 320294
rect 283306 320058 283542 320294
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 289826 507218 290062 507454
rect 290146 507218 290382 507454
rect 289826 506898 290062 507134
rect 290146 506898 290382 507134
rect 289826 471218 290062 471454
rect 290146 471218 290382 471454
rect 289826 470898 290062 471134
rect 290146 470898 290382 471134
rect 289826 435218 290062 435454
rect 290146 435218 290382 435454
rect 289826 434898 290062 435134
rect 290146 434898 290382 435134
rect 289826 399218 290062 399454
rect 290146 399218 290382 399454
rect 289826 398898 290062 399134
rect 290146 398898 290382 399134
rect 289826 363218 290062 363454
rect 290146 363218 290382 363454
rect 289826 362898 290062 363134
rect 290146 362898 290382 363134
rect 289826 327218 290062 327454
rect 290146 327218 290382 327454
rect 289826 326898 290062 327134
rect 290146 326898 290382 327134
rect 293546 690938 293782 691174
rect 293866 690938 294102 691174
rect 293546 690618 293782 690854
rect 293866 690618 294102 690854
rect 293546 654938 293782 655174
rect 293866 654938 294102 655174
rect 293546 654618 293782 654854
rect 293866 654618 294102 654854
rect 293546 618938 293782 619174
rect 293866 618938 294102 619174
rect 293546 618618 293782 618854
rect 293866 618618 294102 618854
rect 293546 582938 293782 583174
rect 293866 582938 294102 583174
rect 293546 582618 293782 582854
rect 293866 582618 294102 582854
rect 293546 546938 293782 547174
rect 293866 546938 294102 547174
rect 293546 546618 293782 546854
rect 293866 546618 294102 546854
rect 293546 510938 293782 511174
rect 293866 510938 294102 511174
rect 293546 510618 293782 510854
rect 293866 510618 294102 510854
rect 293546 474938 293782 475174
rect 293866 474938 294102 475174
rect 293546 474618 293782 474854
rect 293866 474618 294102 474854
rect 293546 438938 293782 439174
rect 293866 438938 294102 439174
rect 293546 438618 293782 438854
rect 293866 438618 294102 438854
rect 293546 402938 293782 403174
rect 293866 402938 294102 403174
rect 293546 402618 293782 402854
rect 293866 402618 294102 402854
rect 293546 366938 293782 367174
rect 293866 366938 294102 367174
rect 293546 366618 293782 366854
rect 293866 366618 294102 366854
rect 293546 330938 293782 331174
rect 293866 330938 294102 331174
rect 293546 330618 293782 330854
rect 293866 330618 294102 330854
rect 297266 694658 297502 694894
rect 297586 694658 297822 694894
rect 297266 694338 297502 694574
rect 297586 694338 297822 694574
rect 297266 658658 297502 658894
rect 297586 658658 297822 658894
rect 297266 658338 297502 658574
rect 297586 658338 297822 658574
rect 297266 622658 297502 622894
rect 297586 622658 297822 622894
rect 297266 622338 297502 622574
rect 297586 622338 297822 622574
rect 297266 586658 297502 586894
rect 297586 586658 297822 586894
rect 297266 586338 297502 586574
rect 297586 586338 297822 586574
rect 297266 550658 297502 550894
rect 297586 550658 297822 550894
rect 297266 550338 297502 550574
rect 297586 550338 297822 550574
rect 297266 514658 297502 514894
rect 297586 514658 297822 514894
rect 297266 514338 297502 514574
rect 297586 514338 297822 514574
rect 297266 478658 297502 478894
rect 297586 478658 297822 478894
rect 297266 478338 297502 478574
rect 297586 478338 297822 478574
rect 297266 442658 297502 442894
rect 297586 442658 297822 442894
rect 297266 442338 297502 442574
rect 297586 442338 297822 442574
rect 297266 406658 297502 406894
rect 297586 406658 297822 406894
rect 297266 406338 297502 406574
rect 297586 406338 297822 406574
rect 297266 370658 297502 370894
rect 297586 370658 297822 370894
rect 297266 370338 297502 370574
rect 297586 370338 297822 370574
rect 297266 334658 297502 334894
rect 297586 334658 297822 334894
rect 297266 334338 297502 334574
rect 297586 334338 297822 334574
rect 318986 711322 319222 711558
rect 319306 711322 319542 711558
rect 318986 711002 319222 711238
rect 319306 711002 319542 711238
rect 315266 709402 315502 709638
rect 315586 709402 315822 709638
rect 315266 709082 315502 709318
rect 315586 709082 315822 709318
rect 311546 707482 311782 707718
rect 311866 707482 312102 707718
rect 311546 707162 311782 707398
rect 311866 707162 312102 707398
rect 300986 698378 301222 698614
rect 301306 698378 301542 698614
rect 300986 698058 301222 698294
rect 301306 698058 301542 698294
rect 300986 662378 301222 662614
rect 301306 662378 301542 662614
rect 300986 662058 301222 662294
rect 301306 662058 301542 662294
rect 300986 626378 301222 626614
rect 301306 626378 301542 626614
rect 300986 626058 301222 626294
rect 301306 626058 301542 626294
rect 300986 590378 301222 590614
rect 301306 590378 301542 590614
rect 300986 590058 301222 590294
rect 301306 590058 301542 590294
rect 300986 554378 301222 554614
rect 301306 554378 301542 554614
rect 300986 554058 301222 554294
rect 301306 554058 301542 554294
rect 300986 518378 301222 518614
rect 301306 518378 301542 518614
rect 300986 518058 301222 518294
rect 301306 518058 301542 518294
rect 300986 482378 301222 482614
rect 301306 482378 301542 482614
rect 300986 482058 301222 482294
rect 301306 482058 301542 482294
rect 300986 446378 301222 446614
rect 301306 446378 301542 446614
rect 300986 446058 301222 446294
rect 301306 446058 301542 446294
rect 300986 410378 301222 410614
rect 301306 410378 301542 410614
rect 300986 410058 301222 410294
rect 301306 410058 301542 410294
rect 300986 374378 301222 374614
rect 301306 374378 301542 374614
rect 300986 374058 301222 374294
rect 301306 374058 301542 374294
rect 300986 338378 301222 338614
rect 301306 338378 301542 338614
rect 300986 338058 301222 338294
rect 301306 338058 301542 338294
rect 300986 302378 301222 302614
rect 301306 302378 301542 302614
rect 300986 302058 301222 302294
rect 301306 302058 301542 302294
rect 307826 705562 308062 705798
rect 308146 705562 308382 705798
rect 307826 705242 308062 705478
rect 308146 705242 308382 705478
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 307826 561218 308062 561454
rect 308146 561218 308382 561454
rect 307826 560898 308062 561134
rect 308146 560898 308382 561134
rect 307826 525218 308062 525454
rect 308146 525218 308382 525454
rect 307826 524898 308062 525134
rect 308146 524898 308382 525134
rect 307826 489218 308062 489454
rect 308146 489218 308382 489454
rect 307826 488898 308062 489134
rect 308146 488898 308382 489134
rect 307826 453218 308062 453454
rect 308146 453218 308382 453454
rect 307826 452898 308062 453134
rect 308146 452898 308382 453134
rect 307826 417218 308062 417454
rect 308146 417218 308382 417454
rect 307826 416898 308062 417134
rect 308146 416898 308382 417134
rect 307826 381218 308062 381454
rect 308146 381218 308382 381454
rect 307826 380898 308062 381134
rect 308146 380898 308382 381134
rect 307826 345218 308062 345454
rect 308146 345218 308382 345454
rect 307826 344898 308062 345134
rect 308146 344898 308382 345134
rect 307826 309218 308062 309454
rect 308146 309218 308382 309454
rect 307826 308898 308062 309134
rect 308146 308898 308382 309134
rect 204250 291218 204486 291454
rect 204250 290898 204486 291134
rect 234970 291218 235206 291454
rect 234970 290898 235206 291134
rect 265690 291218 265926 291454
rect 265690 290898 265926 291134
rect 296410 291218 296646 291454
rect 296410 290898 296646 291134
rect 219610 273218 219846 273454
rect 219610 272898 219846 273134
rect 250330 273218 250566 273454
rect 250330 272898 250566 273134
rect 281050 273218 281286 273454
rect 281050 272898 281286 273134
rect 307826 273218 308062 273454
rect 308146 273218 308382 273454
rect 307826 272898 308062 273134
rect 308146 272898 308382 273134
rect 192986 266378 193222 266614
rect 193306 266378 193542 266614
rect 192986 266058 193222 266294
rect 193306 266058 193542 266294
rect 204250 255218 204486 255454
rect 204250 254898 204486 255134
rect 234970 255218 235206 255454
rect 234970 254898 235206 255134
rect 265690 255218 265926 255454
rect 265690 254898 265926 255134
rect 296410 255218 296646 255454
rect 296410 254898 296646 255134
rect 219610 237218 219846 237454
rect 219610 236898 219846 237134
rect 250330 237218 250566 237454
rect 250330 236898 250566 237134
rect 281050 237218 281286 237454
rect 281050 236898 281286 237134
rect 307826 237218 308062 237454
rect 308146 237218 308382 237454
rect 307826 236898 308062 237134
rect 308146 236898 308382 237134
rect 192986 230378 193222 230614
rect 193306 230378 193542 230614
rect 192986 230058 193222 230294
rect 193306 230058 193542 230294
rect 204250 219218 204486 219454
rect 204250 218898 204486 219134
rect 234970 219218 235206 219454
rect 234970 218898 235206 219134
rect 265690 219218 265926 219454
rect 265690 218898 265926 219134
rect 296410 219218 296646 219454
rect 296410 218898 296646 219134
rect 219610 201218 219846 201454
rect 219610 200898 219846 201134
rect 250330 201218 250566 201454
rect 250330 200898 250566 201134
rect 281050 201218 281286 201454
rect 281050 200898 281286 201134
rect 307826 201218 308062 201454
rect 308146 201218 308382 201454
rect 307826 200898 308062 201134
rect 308146 200898 308382 201134
rect 192986 194378 193222 194614
rect 193306 194378 193542 194614
rect 192986 194058 193222 194294
rect 193306 194058 193542 194294
rect 204250 183218 204486 183454
rect 204250 182898 204486 183134
rect 234970 183218 235206 183454
rect 234970 182898 235206 183134
rect 265690 183218 265926 183454
rect 265690 182898 265926 183134
rect 296410 183218 296646 183454
rect 296410 182898 296646 183134
rect 219610 165218 219846 165454
rect 219610 164898 219846 165134
rect 250330 165218 250566 165454
rect 250330 164898 250566 165134
rect 281050 165218 281286 165454
rect 281050 164898 281286 165134
rect 307826 165218 308062 165454
rect 308146 165218 308382 165454
rect 307826 164898 308062 165134
rect 308146 164898 308382 165134
rect 192986 158378 193222 158614
rect 193306 158378 193542 158614
rect 192986 158058 193222 158294
rect 193306 158058 193542 158294
rect 204250 147218 204486 147454
rect 204250 146898 204486 147134
rect 234970 147218 235206 147454
rect 234970 146898 235206 147134
rect 265690 147218 265926 147454
rect 265690 146898 265926 147134
rect 296410 147218 296646 147454
rect 296410 146898 296646 147134
rect 219610 129218 219846 129454
rect 219610 128898 219846 129134
rect 250330 129218 250566 129454
rect 250330 128898 250566 129134
rect 281050 129218 281286 129454
rect 281050 128898 281286 129134
rect 307826 129218 308062 129454
rect 308146 129218 308382 129454
rect 307826 128898 308062 129134
rect 308146 128898 308382 129134
rect 192986 122378 193222 122614
rect 193306 122378 193542 122614
rect 192986 122058 193222 122294
rect 193306 122058 193542 122294
rect 204250 111218 204486 111454
rect 204250 110898 204486 111134
rect 234970 111218 235206 111454
rect 234970 110898 235206 111134
rect 265690 111218 265926 111454
rect 265690 110898 265926 111134
rect 296410 111218 296646 111454
rect 296410 110898 296646 111134
rect 192986 86378 193222 86614
rect 193306 86378 193542 86614
rect 192986 86058 193222 86294
rect 193306 86058 193542 86294
rect 192986 50378 193222 50614
rect 193306 50378 193542 50614
rect 192986 50058 193222 50294
rect 193306 50058 193542 50294
rect 192986 14378 193222 14614
rect 193306 14378 193542 14614
rect 192986 14058 193222 14294
rect 193306 14058 193542 14294
rect 174986 -7302 175222 -7066
rect 175306 -7302 175542 -7066
rect 174986 -7622 175222 -7386
rect 175306 -7622 175542 -7386
rect 199826 93218 200062 93454
rect 200146 93218 200382 93454
rect 199826 92898 200062 93134
rect 200146 92898 200382 93134
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -1542 200062 -1306
rect 200146 -1542 200382 -1306
rect 199826 -1862 200062 -1626
rect 200146 -1862 200382 -1626
rect 203546 96938 203782 97174
rect 203866 96938 204102 97174
rect 203546 96618 203782 96854
rect 203866 96618 204102 96854
rect 203546 60938 203782 61174
rect 203866 60938 204102 61174
rect 203546 60618 203782 60854
rect 203866 60618 204102 60854
rect 203546 24938 203782 25174
rect 203866 24938 204102 25174
rect 203546 24618 203782 24854
rect 203866 24618 204102 24854
rect 203546 -3462 203782 -3226
rect 203866 -3462 204102 -3226
rect 203546 -3782 203782 -3546
rect 203866 -3782 204102 -3546
rect 207266 64658 207502 64894
rect 207586 64658 207822 64894
rect 207266 64338 207502 64574
rect 207586 64338 207822 64574
rect 207266 28658 207502 28894
rect 207586 28658 207822 28894
rect 207266 28338 207502 28574
rect 207586 28338 207822 28574
rect 207266 -5382 207502 -5146
rect 207586 -5382 207822 -5146
rect 207266 -5702 207502 -5466
rect 207586 -5702 207822 -5466
rect 210986 68378 211222 68614
rect 211306 68378 211542 68614
rect 210986 68058 211222 68294
rect 211306 68058 211542 68294
rect 210986 32378 211222 32614
rect 211306 32378 211542 32614
rect 210986 32058 211222 32294
rect 211306 32058 211542 32294
rect 192986 -6342 193222 -6106
rect 193306 -6342 193542 -6106
rect 192986 -6662 193222 -6426
rect 193306 -6662 193542 -6426
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 221546 78938 221782 79174
rect 221866 78938 222102 79174
rect 221546 78618 221782 78854
rect 221866 78618 222102 78854
rect 221546 42938 221782 43174
rect 221866 42938 222102 43174
rect 221546 42618 221782 42854
rect 221866 42618 222102 42854
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 221546 -2502 221782 -2266
rect 221866 -2502 222102 -2266
rect 221546 -2822 221782 -2586
rect 221866 -2822 222102 -2586
rect 225266 82658 225502 82894
rect 225586 82658 225822 82894
rect 225266 82338 225502 82574
rect 225586 82338 225822 82574
rect 225266 46658 225502 46894
rect 225586 46658 225822 46894
rect 225266 46338 225502 46574
rect 225586 46338 225822 46574
rect 225266 10658 225502 10894
rect 225586 10658 225822 10894
rect 225266 10338 225502 10574
rect 225586 10338 225822 10574
rect 225266 -4422 225502 -4186
rect 225586 -4422 225822 -4186
rect 225266 -4742 225502 -4506
rect 225586 -4742 225822 -4506
rect 228986 86378 229222 86614
rect 229306 86378 229542 86614
rect 228986 86058 229222 86294
rect 229306 86058 229542 86294
rect 228986 50378 229222 50614
rect 229306 50378 229542 50614
rect 228986 50058 229222 50294
rect 229306 50058 229542 50294
rect 228986 14378 229222 14614
rect 229306 14378 229542 14614
rect 228986 14058 229222 14294
rect 229306 14058 229542 14294
rect 210986 -7302 211222 -7066
rect 211306 -7302 211542 -7066
rect 210986 -7622 211222 -7386
rect 211306 -7622 211542 -7386
rect 235826 93218 236062 93454
rect 236146 93218 236382 93454
rect 235826 92898 236062 93134
rect 236146 92898 236382 93134
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -1542 236062 -1306
rect 236146 -1542 236382 -1306
rect 235826 -1862 236062 -1626
rect 236146 -1862 236382 -1626
rect 239546 96938 239782 97174
rect 239866 96938 240102 97174
rect 239546 96618 239782 96854
rect 239866 96618 240102 96854
rect 239546 60938 239782 61174
rect 239866 60938 240102 61174
rect 239546 60618 239782 60854
rect 239866 60618 240102 60854
rect 239546 24938 239782 25174
rect 239866 24938 240102 25174
rect 239546 24618 239782 24854
rect 239866 24618 240102 24854
rect 239546 -3462 239782 -3226
rect 239866 -3462 240102 -3226
rect 239546 -3782 239782 -3546
rect 239866 -3782 240102 -3546
rect 243266 64658 243502 64894
rect 243586 64658 243822 64894
rect 243266 64338 243502 64574
rect 243586 64338 243822 64574
rect 243266 28658 243502 28894
rect 243586 28658 243822 28894
rect 243266 28338 243502 28574
rect 243586 28338 243822 28574
rect 243266 -5382 243502 -5146
rect 243586 -5382 243822 -5146
rect 243266 -5702 243502 -5466
rect 243586 -5702 243822 -5466
rect 246986 68378 247222 68614
rect 247306 68378 247542 68614
rect 246986 68058 247222 68294
rect 247306 68058 247542 68294
rect 246986 32378 247222 32614
rect 247306 32378 247542 32614
rect 246986 32058 247222 32294
rect 247306 32058 247542 32294
rect 228986 -6342 229222 -6106
rect 229306 -6342 229542 -6106
rect 228986 -6662 229222 -6426
rect 229306 -6662 229542 -6426
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 257546 78938 257782 79174
rect 257866 78938 258102 79174
rect 257546 78618 257782 78854
rect 257866 78618 258102 78854
rect 257546 42938 257782 43174
rect 257866 42938 258102 43174
rect 257546 42618 257782 42854
rect 257866 42618 258102 42854
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 257546 -2502 257782 -2266
rect 257866 -2502 258102 -2266
rect 257546 -2822 257782 -2586
rect 257866 -2822 258102 -2586
rect 261266 82658 261502 82894
rect 261586 82658 261822 82894
rect 261266 82338 261502 82574
rect 261586 82338 261822 82574
rect 261266 46658 261502 46894
rect 261586 46658 261822 46894
rect 261266 46338 261502 46574
rect 261586 46338 261822 46574
rect 261266 10658 261502 10894
rect 261586 10658 261822 10894
rect 261266 10338 261502 10574
rect 261586 10338 261822 10574
rect 261266 -4422 261502 -4186
rect 261586 -4422 261822 -4186
rect 261266 -4742 261502 -4506
rect 261586 -4742 261822 -4506
rect 264986 86378 265222 86614
rect 265306 86378 265542 86614
rect 264986 86058 265222 86294
rect 265306 86058 265542 86294
rect 264986 50378 265222 50614
rect 265306 50378 265542 50614
rect 264986 50058 265222 50294
rect 265306 50058 265542 50294
rect 264986 14378 265222 14614
rect 265306 14378 265542 14614
rect 264986 14058 265222 14294
rect 265306 14058 265542 14294
rect 246986 -7302 247222 -7066
rect 247306 -7302 247542 -7066
rect 246986 -7622 247222 -7386
rect 247306 -7622 247542 -7386
rect 271826 93218 272062 93454
rect 272146 93218 272382 93454
rect 271826 92898 272062 93134
rect 272146 92898 272382 93134
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -1542 272062 -1306
rect 272146 -1542 272382 -1306
rect 271826 -1862 272062 -1626
rect 272146 -1862 272382 -1626
rect 275546 96938 275782 97174
rect 275866 96938 276102 97174
rect 275546 96618 275782 96854
rect 275866 96618 276102 96854
rect 275546 60938 275782 61174
rect 275866 60938 276102 61174
rect 275546 60618 275782 60854
rect 275866 60618 276102 60854
rect 275546 24938 275782 25174
rect 275866 24938 276102 25174
rect 275546 24618 275782 24854
rect 275866 24618 276102 24854
rect 275546 -3462 275782 -3226
rect 275866 -3462 276102 -3226
rect 275546 -3782 275782 -3546
rect 275866 -3782 276102 -3546
rect 279266 64658 279502 64894
rect 279586 64658 279822 64894
rect 279266 64338 279502 64574
rect 279586 64338 279822 64574
rect 279266 28658 279502 28894
rect 279586 28658 279822 28894
rect 279266 28338 279502 28574
rect 279586 28338 279822 28574
rect 279266 -5382 279502 -5146
rect 279586 -5382 279822 -5146
rect 279266 -5702 279502 -5466
rect 279586 -5702 279822 -5466
rect 282986 68378 283222 68614
rect 283306 68378 283542 68614
rect 282986 68058 283222 68294
rect 283306 68058 283542 68294
rect 282986 32378 283222 32614
rect 283306 32378 283542 32614
rect 282986 32058 283222 32294
rect 283306 32058 283542 32294
rect 264986 -6342 265222 -6106
rect 265306 -6342 265542 -6106
rect 264986 -6662 265222 -6426
rect 265306 -6662 265542 -6426
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 293546 78938 293782 79174
rect 293866 78938 294102 79174
rect 293546 78618 293782 78854
rect 293866 78618 294102 78854
rect 293546 42938 293782 43174
rect 293866 42938 294102 43174
rect 293546 42618 293782 42854
rect 293866 42618 294102 42854
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 293546 -2502 293782 -2266
rect 293866 -2502 294102 -2266
rect 293546 -2822 293782 -2586
rect 293866 -2822 294102 -2586
rect 297266 82658 297502 82894
rect 297586 82658 297822 82894
rect 297266 82338 297502 82574
rect 297586 82338 297822 82574
rect 297266 46658 297502 46894
rect 297586 46658 297822 46894
rect 297266 46338 297502 46574
rect 297586 46338 297822 46574
rect 297266 10658 297502 10894
rect 297586 10658 297822 10894
rect 297266 10338 297502 10574
rect 297586 10338 297822 10574
rect 297266 -4422 297502 -4186
rect 297586 -4422 297822 -4186
rect 297266 -4742 297502 -4506
rect 297586 -4742 297822 -4506
rect 300986 86378 301222 86614
rect 301306 86378 301542 86614
rect 300986 86058 301222 86294
rect 301306 86058 301542 86294
rect 300986 50378 301222 50614
rect 301306 50378 301542 50614
rect 300986 50058 301222 50294
rect 301306 50058 301542 50294
rect 300986 14378 301222 14614
rect 301306 14378 301542 14614
rect 300986 14058 301222 14294
rect 301306 14058 301542 14294
rect 282986 -7302 283222 -7066
rect 283306 -7302 283542 -7066
rect 282986 -7622 283222 -7386
rect 283306 -7622 283542 -7386
rect 307826 93218 308062 93454
rect 308146 93218 308382 93454
rect 307826 92898 308062 93134
rect 308146 92898 308382 93134
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -1542 308062 -1306
rect 308146 -1542 308382 -1306
rect 307826 -1862 308062 -1626
rect 308146 -1862 308382 -1626
rect 311546 672938 311782 673174
rect 311866 672938 312102 673174
rect 311546 672618 311782 672854
rect 311866 672618 312102 672854
rect 311546 636938 311782 637174
rect 311866 636938 312102 637174
rect 311546 636618 311782 636854
rect 311866 636618 312102 636854
rect 311546 600938 311782 601174
rect 311866 600938 312102 601174
rect 311546 600618 311782 600854
rect 311866 600618 312102 600854
rect 311546 564938 311782 565174
rect 311866 564938 312102 565174
rect 311546 564618 311782 564854
rect 311866 564618 312102 564854
rect 311546 528938 311782 529174
rect 311866 528938 312102 529174
rect 311546 528618 311782 528854
rect 311866 528618 312102 528854
rect 311546 492938 311782 493174
rect 311866 492938 312102 493174
rect 311546 492618 311782 492854
rect 311866 492618 312102 492854
rect 311546 456938 311782 457174
rect 311866 456938 312102 457174
rect 311546 456618 311782 456854
rect 311866 456618 312102 456854
rect 311546 420938 311782 421174
rect 311866 420938 312102 421174
rect 311546 420618 311782 420854
rect 311866 420618 312102 420854
rect 311546 384938 311782 385174
rect 311866 384938 312102 385174
rect 311546 384618 311782 384854
rect 311866 384618 312102 384854
rect 311546 348938 311782 349174
rect 311866 348938 312102 349174
rect 311546 348618 311782 348854
rect 311866 348618 312102 348854
rect 311546 312938 311782 313174
rect 311866 312938 312102 313174
rect 311546 312618 311782 312854
rect 311866 312618 312102 312854
rect 311546 276938 311782 277174
rect 311866 276938 312102 277174
rect 311546 276618 311782 276854
rect 311866 276618 312102 276854
rect 311546 240938 311782 241174
rect 311866 240938 312102 241174
rect 311546 240618 311782 240854
rect 311866 240618 312102 240854
rect 311546 204938 311782 205174
rect 311866 204938 312102 205174
rect 311546 204618 311782 204854
rect 311866 204618 312102 204854
rect 311546 168938 311782 169174
rect 311866 168938 312102 169174
rect 311546 168618 311782 168854
rect 311866 168618 312102 168854
rect 311546 132938 311782 133174
rect 311866 132938 312102 133174
rect 311546 132618 311782 132854
rect 311866 132618 312102 132854
rect 311546 96938 311782 97174
rect 311866 96938 312102 97174
rect 311546 96618 311782 96854
rect 311866 96618 312102 96854
rect 311546 60938 311782 61174
rect 311866 60938 312102 61174
rect 311546 60618 311782 60854
rect 311866 60618 312102 60854
rect 311546 24938 311782 25174
rect 311866 24938 312102 25174
rect 311546 24618 311782 24854
rect 311866 24618 312102 24854
rect 311546 -3462 311782 -3226
rect 311866 -3462 312102 -3226
rect 311546 -3782 311782 -3546
rect 311866 -3782 312102 -3546
rect 315266 676658 315502 676894
rect 315586 676658 315822 676894
rect 315266 676338 315502 676574
rect 315586 676338 315822 676574
rect 315266 640658 315502 640894
rect 315586 640658 315822 640894
rect 315266 640338 315502 640574
rect 315586 640338 315822 640574
rect 315266 604658 315502 604894
rect 315586 604658 315822 604894
rect 315266 604338 315502 604574
rect 315586 604338 315822 604574
rect 315266 568658 315502 568894
rect 315586 568658 315822 568894
rect 315266 568338 315502 568574
rect 315586 568338 315822 568574
rect 315266 532658 315502 532894
rect 315586 532658 315822 532894
rect 315266 532338 315502 532574
rect 315586 532338 315822 532574
rect 315266 496658 315502 496894
rect 315586 496658 315822 496894
rect 315266 496338 315502 496574
rect 315586 496338 315822 496574
rect 315266 460658 315502 460894
rect 315586 460658 315822 460894
rect 315266 460338 315502 460574
rect 315586 460338 315822 460574
rect 315266 424658 315502 424894
rect 315586 424658 315822 424894
rect 315266 424338 315502 424574
rect 315586 424338 315822 424574
rect 315266 388658 315502 388894
rect 315586 388658 315822 388894
rect 315266 388338 315502 388574
rect 315586 388338 315822 388574
rect 315266 352658 315502 352894
rect 315586 352658 315822 352894
rect 315266 352338 315502 352574
rect 315586 352338 315822 352574
rect 315266 316658 315502 316894
rect 315586 316658 315822 316894
rect 315266 316338 315502 316574
rect 315586 316338 315822 316574
rect 315266 280658 315502 280894
rect 315586 280658 315822 280894
rect 315266 280338 315502 280574
rect 315586 280338 315822 280574
rect 315266 244658 315502 244894
rect 315586 244658 315822 244894
rect 315266 244338 315502 244574
rect 315586 244338 315822 244574
rect 315266 208658 315502 208894
rect 315586 208658 315822 208894
rect 315266 208338 315502 208574
rect 315586 208338 315822 208574
rect 315266 172658 315502 172894
rect 315586 172658 315822 172894
rect 315266 172338 315502 172574
rect 315586 172338 315822 172574
rect 315266 136658 315502 136894
rect 315586 136658 315822 136894
rect 315266 136338 315502 136574
rect 315586 136338 315822 136574
rect 315266 100658 315502 100894
rect 315586 100658 315822 100894
rect 315266 100338 315502 100574
rect 315586 100338 315822 100574
rect 315266 64658 315502 64894
rect 315586 64658 315822 64894
rect 315266 64338 315502 64574
rect 315586 64338 315822 64574
rect 315266 28658 315502 28894
rect 315586 28658 315822 28894
rect 315266 28338 315502 28574
rect 315586 28338 315822 28574
rect 315266 -5382 315502 -5146
rect 315586 -5382 315822 -5146
rect 315266 -5702 315502 -5466
rect 315586 -5702 315822 -5466
rect 336986 710362 337222 710598
rect 337306 710362 337542 710598
rect 336986 710042 337222 710278
rect 337306 710042 337542 710278
rect 333266 708442 333502 708678
rect 333586 708442 333822 708678
rect 333266 708122 333502 708358
rect 333586 708122 333822 708358
rect 329546 706522 329782 706758
rect 329866 706522 330102 706758
rect 329546 706202 329782 706438
rect 329866 706202 330102 706438
rect 318986 680378 319222 680614
rect 319306 680378 319542 680614
rect 318986 680058 319222 680294
rect 319306 680058 319542 680294
rect 318986 644378 319222 644614
rect 319306 644378 319542 644614
rect 318986 644058 319222 644294
rect 319306 644058 319542 644294
rect 318986 608378 319222 608614
rect 319306 608378 319542 608614
rect 318986 608058 319222 608294
rect 319306 608058 319542 608294
rect 318986 572378 319222 572614
rect 319306 572378 319542 572614
rect 318986 572058 319222 572294
rect 319306 572058 319542 572294
rect 318986 536378 319222 536614
rect 319306 536378 319542 536614
rect 318986 536058 319222 536294
rect 319306 536058 319542 536294
rect 318986 500378 319222 500614
rect 319306 500378 319542 500614
rect 318986 500058 319222 500294
rect 319306 500058 319542 500294
rect 318986 464378 319222 464614
rect 319306 464378 319542 464614
rect 318986 464058 319222 464294
rect 319306 464058 319542 464294
rect 318986 428378 319222 428614
rect 319306 428378 319542 428614
rect 318986 428058 319222 428294
rect 319306 428058 319542 428294
rect 318986 392378 319222 392614
rect 319306 392378 319542 392614
rect 318986 392058 319222 392294
rect 319306 392058 319542 392294
rect 318986 356378 319222 356614
rect 319306 356378 319542 356614
rect 318986 356058 319222 356294
rect 319306 356058 319542 356294
rect 318986 320378 319222 320614
rect 319306 320378 319542 320614
rect 318986 320058 319222 320294
rect 319306 320058 319542 320294
rect 318986 284378 319222 284614
rect 319306 284378 319542 284614
rect 318986 284058 319222 284294
rect 319306 284058 319542 284294
rect 318986 248378 319222 248614
rect 319306 248378 319542 248614
rect 318986 248058 319222 248294
rect 319306 248058 319542 248294
rect 318986 212378 319222 212614
rect 319306 212378 319542 212614
rect 318986 212058 319222 212294
rect 319306 212058 319542 212294
rect 318986 176378 319222 176614
rect 319306 176378 319542 176614
rect 318986 176058 319222 176294
rect 319306 176058 319542 176294
rect 318986 140378 319222 140614
rect 319306 140378 319542 140614
rect 318986 140058 319222 140294
rect 319306 140058 319542 140294
rect 318986 104378 319222 104614
rect 319306 104378 319542 104614
rect 318986 104058 319222 104294
rect 319306 104058 319542 104294
rect 318986 68378 319222 68614
rect 319306 68378 319542 68614
rect 318986 68058 319222 68294
rect 319306 68058 319542 68294
rect 318986 32378 319222 32614
rect 319306 32378 319542 32614
rect 318986 32058 319222 32294
rect 319306 32058 319542 32294
rect 300986 -6342 301222 -6106
rect 301306 -6342 301542 -6106
rect 300986 -6662 301222 -6426
rect 301306 -6662 301542 -6426
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 325826 543218 326062 543454
rect 326146 543218 326382 543454
rect 325826 542898 326062 543134
rect 326146 542898 326382 543134
rect 325826 507218 326062 507454
rect 326146 507218 326382 507454
rect 325826 506898 326062 507134
rect 326146 506898 326382 507134
rect 325826 471218 326062 471454
rect 326146 471218 326382 471454
rect 325826 470898 326062 471134
rect 326146 470898 326382 471134
rect 325826 435218 326062 435454
rect 326146 435218 326382 435454
rect 325826 434898 326062 435134
rect 326146 434898 326382 435134
rect 325826 399218 326062 399454
rect 326146 399218 326382 399454
rect 325826 398898 326062 399134
rect 326146 398898 326382 399134
rect 325826 363218 326062 363454
rect 326146 363218 326382 363454
rect 325826 362898 326062 363134
rect 326146 362898 326382 363134
rect 325826 327218 326062 327454
rect 326146 327218 326382 327454
rect 325826 326898 326062 327134
rect 326146 326898 326382 327134
rect 325826 291218 326062 291454
rect 326146 291218 326382 291454
rect 325826 290898 326062 291134
rect 326146 290898 326382 291134
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 325826 219218 326062 219454
rect 326146 219218 326382 219454
rect 325826 218898 326062 219134
rect 326146 218898 326382 219134
rect 325826 183218 326062 183454
rect 326146 183218 326382 183454
rect 325826 182898 326062 183134
rect 326146 182898 326382 183134
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 325826 111218 326062 111454
rect 326146 111218 326382 111454
rect 325826 110898 326062 111134
rect 326146 110898 326382 111134
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 690938 329782 691174
rect 329866 690938 330102 691174
rect 329546 690618 329782 690854
rect 329866 690618 330102 690854
rect 329546 654938 329782 655174
rect 329866 654938 330102 655174
rect 329546 654618 329782 654854
rect 329866 654618 330102 654854
rect 329546 618938 329782 619174
rect 329866 618938 330102 619174
rect 329546 618618 329782 618854
rect 329866 618618 330102 618854
rect 329546 582938 329782 583174
rect 329866 582938 330102 583174
rect 329546 582618 329782 582854
rect 329866 582618 330102 582854
rect 329546 546938 329782 547174
rect 329866 546938 330102 547174
rect 329546 546618 329782 546854
rect 329866 546618 330102 546854
rect 329546 510938 329782 511174
rect 329866 510938 330102 511174
rect 329546 510618 329782 510854
rect 329866 510618 330102 510854
rect 329546 474938 329782 475174
rect 329866 474938 330102 475174
rect 329546 474618 329782 474854
rect 329866 474618 330102 474854
rect 329546 438938 329782 439174
rect 329866 438938 330102 439174
rect 329546 438618 329782 438854
rect 329866 438618 330102 438854
rect 329546 402938 329782 403174
rect 329866 402938 330102 403174
rect 329546 402618 329782 402854
rect 329866 402618 330102 402854
rect 329546 366938 329782 367174
rect 329866 366938 330102 367174
rect 329546 366618 329782 366854
rect 329866 366618 330102 366854
rect 329546 330938 329782 331174
rect 329866 330938 330102 331174
rect 329546 330618 329782 330854
rect 329866 330618 330102 330854
rect 329546 294938 329782 295174
rect 329866 294938 330102 295174
rect 329546 294618 329782 294854
rect 329866 294618 330102 294854
rect 329546 258938 329782 259174
rect 329866 258938 330102 259174
rect 329546 258618 329782 258854
rect 329866 258618 330102 258854
rect 329546 222938 329782 223174
rect 329866 222938 330102 223174
rect 329546 222618 329782 222854
rect 329866 222618 330102 222854
rect 329546 186938 329782 187174
rect 329866 186938 330102 187174
rect 329546 186618 329782 186854
rect 329866 186618 330102 186854
rect 329546 150938 329782 151174
rect 329866 150938 330102 151174
rect 329546 150618 329782 150854
rect 329866 150618 330102 150854
rect 329546 114938 329782 115174
rect 329866 114938 330102 115174
rect 329546 114618 329782 114854
rect 329866 114618 330102 114854
rect 329546 78938 329782 79174
rect 329866 78938 330102 79174
rect 329546 78618 329782 78854
rect 329866 78618 330102 78854
rect 329546 42938 329782 43174
rect 329866 42938 330102 43174
rect 329546 42618 329782 42854
rect 329866 42618 330102 42854
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 329546 -2502 329782 -2266
rect 329866 -2502 330102 -2266
rect 329546 -2822 329782 -2586
rect 329866 -2822 330102 -2586
rect 333266 694658 333502 694894
rect 333586 694658 333822 694894
rect 333266 694338 333502 694574
rect 333586 694338 333822 694574
rect 333266 658658 333502 658894
rect 333586 658658 333822 658894
rect 333266 658338 333502 658574
rect 333586 658338 333822 658574
rect 333266 622658 333502 622894
rect 333586 622658 333822 622894
rect 333266 622338 333502 622574
rect 333586 622338 333822 622574
rect 333266 586658 333502 586894
rect 333586 586658 333822 586894
rect 333266 586338 333502 586574
rect 333586 586338 333822 586574
rect 333266 550658 333502 550894
rect 333586 550658 333822 550894
rect 333266 550338 333502 550574
rect 333586 550338 333822 550574
rect 333266 514658 333502 514894
rect 333586 514658 333822 514894
rect 333266 514338 333502 514574
rect 333586 514338 333822 514574
rect 333266 478658 333502 478894
rect 333586 478658 333822 478894
rect 333266 478338 333502 478574
rect 333586 478338 333822 478574
rect 333266 442658 333502 442894
rect 333586 442658 333822 442894
rect 333266 442338 333502 442574
rect 333586 442338 333822 442574
rect 333266 406658 333502 406894
rect 333586 406658 333822 406894
rect 333266 406338 333502 406574
rect 333586 406338 333822 406574
rect 333266 370658 333502 370894
rect 333586 370658 333822 370894
rect 333266 370338 333502 370574
rect 333586 370338 333822 370574
rect 333266 334658 333502 334894
rect 333586 334658 333822 334894
rect 333266 334338 333502 334574
rect 333586 334338 333822 334574
rect 333266 298658 333502 298894
rect 333586 298658 333822 298894
rect 333266 298338 333502 298574
rect 333586 298338 333822 298574
rect 333266 262658 333502 262894
rect 333586 262658 333822 262894
rect 333266 262338 333502 262574
rect 333586 262338 333822 262574
rect 333266 226658 333502 226894
rect 333586 226658 333822 226894
rect 333266 226338 333502 226574
rect 333586 226338 333822 226574
rect 333266 190658 333502 190894
rect 333586 190658 333822 190894
rect 333266 190338 333502 190574
rect 333586 190338 333822 190574
rect 333266 154658 333502 154894
rect 333586 154658 333822 154894
rect 333266 154338 333502 154574
rect 333586 154338 333822 154574
rect 333266 118658 333502 118894
rect 333586 118658 333822 118894
rect 333266 118338 333502 118574
rect 333586 118338 333822 118574
rect 333266 82658 333502 82894
rect 333586 82658 333822 82894
rect 333266 82338 333502 82574
rect 333586 82338 333822 82574
rect 333266 46658 333502 46894
rect 333586 46658 333822 46894
rect 333266 46338 333502 46574
rect 333586 46338 333822 46574
rect 333266 10658 333502 10894
rect 333586 10658 333822 10894
rect 333266 10338 333502 10574
rect 333586 10338 333822 10574
rect 333266 -4422 333502 -4186
rect 333586 -4422 333822 -4186
rect 333266 -4742 333502 -4506
rect 333586 -4742 333822 -4506
rect 354986 711322 355222 711558
rect 355306 711322 355542 711558
rect 354986 711002 355222 711238
rect 355306 711002 355542 711238
rect 351266 709402 351502 709638
rect 351586 709402 351822 709638
rect 351266 709082 351502 709318
rect 351586 709082 351822 709318
rect 347546 707482 347782 707718
rect 347866 707482 348102 707718
rect 347546 707162 347782 707398
rect 347866 707162 348102 707398
rect 336986 698378 337222 698614
rect 337306 698378 337542 698614
rect 336986 698058 337222 698294
rect 337306 698058 337542 698294
rect 336986 662378 337222 662614
rect 337306 662378 337542 662614
rect 336986 662058 337222 662294
rect 337306 662058 337542 662294
rect 336986 626378 337222 626614
rect 337306 626378 337542 626614
rect 336986 626058 337222 626294
rect 337306 626058 337542 626294
rect 336986 590378 337222 590614
rect 337306 590378 337542 590614
rect 336986 590058 337222 590294
rect 337306 590058 337542 590294
rect 336986 554378 337222 554614
rect 337306 554378 337542 554614
rect 336986 554058 337222 554294
rect 337306 554058 337542 554294
rect 336986 518378 337222 518614
rect 337306 518378 337542 518614
rect 336986 518058 337222 518294
rect 337306 518058 337542 518294
rect 336986 482378 337222 482614
rect 337306 482378 337542 482614
rect 336986 482058 337222 482294
rect 337306 482058 337542 482294
rect 336986 446378 337222 446614
rect 337306 446378 337542 446614
rect 336986 446058 337222 446294
rect 337306 446058 337542 446294
rect 336986 410378 337222 410614
rect 337306 410378 337542 410614
rect 336986 410058 337222 410294
rect 337306 410058 337542 410294
rect 336986 374378 337222 374614
rect 337306 374378 337542 374614
rect 336986 374058 337222 374294
rect 337306 374058 337542 374294
rect 336986 338378 337222 338614
rect 337306 338378 337542 338614
rect 336986 338058 337222 338294
rect 337306 338058 337542 338294
rect 336986 302378 337222 302614
rect 337306 302378 337542 302614
rect 336986 302058 337222 302294
rect 337306 302058 337542 302294
rect 336986 266378 337222 266614
rect 337306 266378 337542 266614
rect 336986 266058 337222 266294
rect 337306 266058 337542 266294
rect 336986 230378 337222 230614
rect 337306 230378 337542 230614
rect 336986 230058 337222 230294
rect 337306 230058 337542 230294
rect 336986 194378 337222 194614
rect 337306 194378 337542 194614
rect 336986 194058 337222 194294
rect 337306 194058 337542 194294
rect 336986 158378 337222 158614
rect 337306 158378 337542 158614
rect 336986 158058 337222 158294
rect 337306 158058 337542 158294
rect 336986 122378 337222 122614
rect 337306 122378 337542 122614
rect 336986 122058 337222 122294
rect 337306 122058 337542 122294
rect 336986 86378 337222 86614
rect 337306 86378 337542 86614
rect 336986 86058 337222 86294
rect 337306 86058 337542 86294
rect 336986 50378 337222 50614
rect 337306 50378 337542 50614
rect 336986 50058 337222 50294
rect 337306 50058 337542 50294
rect 336986 14378 337222 14614
rect 337306 14378 337542 14614
rect 336986 14058 337222 14294
rect 337306 14058 337542 14294
rect 318986 -7302 319222 -7066
rect 319306 -7302 319542 -7066
rect 318986 -7622 319222 -7386
rect 319306 -7622 319542 -7386
rect 343826 705562 344062 705798
rect 344146 705562 344382 705798
rect 343826 705242 344062 705478
rect 344146 705242 344382 705478
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 343826 561218 344062 561454
rect 344146 561218 344382 561454
rect 343826 560898 344062 561134
rect 344146 560898 344382 561134
rect 343826 525218 344062 525454
rect 344146 525218 344382 525454
rect 343826 524898 344062 525134
rect 344146 524898 344382 525134
rect 343826 489218 344062 489454
rect 344146 489218 344382 489454
rect 343826 488898 344062 489134
rect 344146 488898 344382 489134
rect 343826 453218 344062 453454
rect 344146 453218 344382 453454
rect 343826 452898 344062 453134
rect 344146 452898 344382 453134
rect 343826 417218 344062 417454
rect 344146 417218 344382 417454
rect 343826 416898 344062 417134
rect 344146 416898 344382 417134
rect 343826 381218 344062 381454
rect 344146 381218 344382 381454
rect 343826 380898 344062 381134
rect 344146 380898 344382 381134
rect 343826 345218 344062 345454
rect 344146 345218 344382 345454
rect 343826 344898 344062 345134
rect 344146 344898 344382 345134
rect 343826 309218 344062 309454
rect 344146 309218 344382 309454
rect 343826 308898 344062 309134
rect 344146 308898 344382 309134
rect 343826 273218 344062 273454
rect 344146 273218 344382 273454
rect 343826 272898 344062 273134
rect 344146 272898 344382 273134
rect 343826 237218 344062 237454
rect 344146 237218 344382 237454
rect 343826 236898 344062 237134
rect 344146 236898 344382 237134
rect 343826 201218 344062 201454
rect 344146 201218 344382 201454
rect 343826 200898 344062 201134
rect 344146 200898 344382 201134
rect 343826 165218 344062 165454
rect 344146 165218 344382 165454
rect 343826 164898 344062 165134
rect 344146 164898 344382 165134
rect 343826 129218 344062 129454
rect 344146 129218 344382 129454
rect 343826 128898 344062 129134
rect 344146 128898 344382 129134
rect 343826 93218 344062 93454
rect 344146 93218 344382 93454
rect 343826 92898 344062 93134
rect 344146 92898 344382 93134
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -1542 344062 -1306
rect 344146 -1542 344382 -1306
rect 343826 -1862 344062 -1626
rect 344146 -1862 344382 -1626
rect 347546 672938 347782 673174
rect 347866 672938 348102 673174
rect 347546 672618 347782 672854
rect 347866 672618 348102 672854
rect 347546 636938 347782 637174
rect 347866 636938 348102 637174
rect 347546 636618 347782 636854
rect 347866 636618 348102 636854
rect 347546 600938 347782 601174
rect 347866 600938 348102 601174
rect 347546 600618 347782 600854
rect 347866 600618 348102 600854
rect 347546 564938 347782 565174
rect 347866 564938 348102 565174
rect 347546 564618 347782 564854
rect 347866 564618 348102 564854
rect 347546 528938 347782 529174
rect 347866 528938 348102 529174
rect 347546 528618 347782 528854
rect 347866 528618 348102 528854
rect 347546 492938 347782 493174
rect 347866 492938 348102 493174
rect 347546 492618 347782 492854
rect 347866 492618 348102 492854
rect 347546 456938 347782 457174
rect 347866 456938 348102 457174
rect 347546 456618 347782 456854
rect 347866 456618 348102 456854
rect 347546 420938 347782 421174
rect 347866 420938 348102 421174
rect 347546 420618 347782 420854
rect 347866 420618 348102 420854
rect 347546 384938 347782 385174
rect 347866 384938 348102 385174
rect 347546 384618 347782 384854
rect 347866 384618 348102 384854
rect 347546 348938 347782 349174
rect 347866 348938 348102 349174
rect 347546 348618 347782 348854
rect 347866 348618 348102 348854
rect 347546 312938 347782 313174
rect 347866 312938 348102 313174
rect 347546 312618 347782 312854
rect 347866 312618 348102 312854
rect 347546 276938 347782 277174
rect 347866 276938 348102 277174
rect 347546 276618 347782 276854
rect 347866 276618 348102 276854
rect 347546 240938 347782 241174
rect 347866 240938 348102 241174
rect 347546 240618 347782 240854
rect 347866 240618 348102 240854
rect 347546 204938 347782 205174
rect 347866 204938 348102 205174
rect 347546 204618 347782 204854
rect 347866 204618 348102 204854
rect 347546 168938 347782 169174
rect 347866 168938 348102 169174
rect 347546 168618 347782 168854
rect 347866 168618 348102 168854
rect 347546 132938 347782 133174
rect 347866 132938 348102 133174
rect 347546 132618 347782 132854
rect 347866 132618 348102 132854
rect 347546 96938 347782 97174
rect 347866 96938 348102 97174
rect 347546 96618 347782 96854
rect 347866 96618 348102 96854
rect 347546 60938 347782 61174
rect 347866 60938 348102 61174
rect 347546 60618 347782 60854
rect 347866 60618 348102 60854
rect 347546 24938 347782 25174
rect 347866 24938 348102 25174
rect 347546 24618 347782 24854
rect 347866 24618 348102 24854
rect 347546 -3462 347782 -3226
rect 347866 -3462 348102 -3226
rect 347546 -3782 347782 -3546
rect 347866 -3782 348102 -3546
rect 351266 676658 351502 676894
rect 351586 676658 351822 676894
rect 351266 676338 351502 676574
rect 351586 676338 351822 676574
rect 351266 640658 351502 640894
rect 351586 640658 351822 640894
rect 351266 640338 351502 640574
rect 351586 640338 351822 640574
rect 351266 604658 351502 604894
rect 351586 604658 351822 604894
rect 351266 604338 351502 604574
rect 351586 604338 351822 604574
rect 351266 568658 351502 568894
rect 351586 568658 351822 568894
rect 351266 568338 351502 568574
rect 351586 568338 351822 568574
rect 351266 532658 351502 532894
rect 351586 532658 351822 532894
rect 351266 532338 351502 532574
rect 351586 532338 351822 532574
rect 351266 496658 351502 496894
rect 351586 496658 351822 496894
rect 351266 496338 351502 496574
rect 351586 496338 351822 496574
rect 351266 460658 351502 460894
rect 351586 460658 351822 460894
rect 351266 460338 351502 460574
rect 351586 460338 351822 460574
rect 351266 424658 351502 424894
rect 351586 424658 351822 424894
rect 351266 424338 351502 424574
rect 351586 424338 351822 424574
rect 351266 388658 351502 388894
rect 351586 388658 351822 388894
rect 351266 388338 351502 388574
rect 351586 388338 351822 388574
rect 351266 352658 351502 352894
rect 351586 352658 351822 352894
rect 351266 352338 351502 352574
rect 351586 352338 351822 352574
rect 351266 316658 351502 316894
rect 351586 316658 351822 316894
rect 351266 316338 351502 316574
rect 351586 316338 351822 316574
rect 351266 280658 351502 280894
rect 351586 280658 351822 280894
rect 351266 280338 351502 280574
rect 351586 280338 351822 280574
rect 351266 244658 351502 244894
rect 351586 244658 351822 244894
rect 351266 244338 351502 244574
rect 351586 244338 351822 244574
rect 351266 208658 351502 208894
rect 351586 208658 351822 208894
rect 351266 208338 351502 208574
rect 351586 208338 351822 208574
rect 351266 172658 351502 172894
rect 351586 172658 351822 172894
rect 351266 172338 351502 172574
rect 351586 172338 351822 172574
rect 351266 136658 351502 136894
rect 351586 136658 351822 136894
rect 351266 136338 351502 136574
rect 351586 136338 351822 136574
rect 351266 100658 351502 100894
rect 351586 100658 351822 100894
rect 351266 100338 351502 100574
rect 351586 100338 351822 100574
rect 351266 64658 351502 64894
rect 351586 64658 351822 64894
rect 351266 64338 351502 64574
rect 351586 64338 351822 64574
rect 351266 28658 351502 28894
rect 351586 28658 351822 28894
rect 351266 28338 351502 28574
rect 351586 28338 351822 28574
rect 351266 -5382 351502 -5146
rect 351586 -5382 351822 -5146
rect 351266 -5702 351502 -5466
rect 351586 -5702 351822 -5466
rect 372986 710362 373222 710598
rect 373306 710362 373542 710598
rect 372986 710042 373222 710278
rect 373306 710042 373542 710278
rect 369266 708442 369502 708678
rect 369586 708442 369822 708678
rect 369266 708122 369502 708358
rect 369586 708122 369822 708358
rect 365546 706522 365782 706758
rect 365866 706522 366102 706758
rect 365546 706202 365782 706438
rect 365866 706202 366102 706438
rect 354986 680378 355222 680614
rect 355306 680378 355542 680614
rect 354986 680058 355222 680294
rect 355306 680058 355542 680294
rect 354986 644378 355222 644614
rect 355306 644378 355542 644614
rect 354986 644058 355222 644294
rect 355306 644058 355542 644294
rect 354986 608378 355222 608614
rect 355306 608378 355542 608614
rect 354986 608058 355222 608294
rect 355306 608058 355542 608294
rect 354986 572378 355222 572614
rect 355306 572378 355542 572614
rect 354986 572058 355222 572294
rect 355306 572058 355542 572294
rect 354986 536378 355222 536614
rect 355306 536378 355542 536614
rect 354986 536058 355222 536294
rect 355306 536058 355542 536294
rect 354986 500378 355222 500614
rect 355306 500378 355542 500614
rect 354986 500058 355222 500294
rect 355306 500058 355542 500294
rect 354986 464378 355222 464614
rect 355306 464378 355542 464614
rect 354986 464058 355222 464294
rect 355306 464058 355542 464294
rect 354986 428378 355222 428614
rect 355306 428378 355542 428614
rect 354986 428058 355222 428294
rect 355306 428058 355542 428294
rect 354986 392378 355222 392614
rect 355306 392378 355542 392614
rect 354986 392058 355222 392294
rect 355306 392058 355542 392294
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 361826 435218 362062 435454
rect 362146 435218 362382 435454
rect 361826 434898 362062 435134
rect 362146 434898 362382 435134
rect 361826 399218 362062 399454
rect 362146 399218 362382 399454
rect 361826 398898 362062 399134
rect 362146 398898 362382 399134
rect 365546 690938 365782 691174
rect 365866 690938 366102 691174
rect 365546 690618 365782 690854
rect 365866 690618 366102 690854
rect 365546 654938 365782 655174
rect 365866 654938 366102 655174
rect 365546 654618 365782 654854
rect 365866 654618 366102 654854
rect 365546 618938 365782 619174
rect 365866 618938 366102 619174
rect 365546 618618 365782 618854
rect 365866 618618 366102 618854
rect 365546 582938 365782 583174
rect 365866 582938 366102 583174
rect 365546 582618 365782 582854
rect 365866 582618 366102 582854
rect 365546 546938 365782 547174
rect 365866 546938 366102 547174
rect 365546 546618 365782 546854
rect 365866 546618 366102 546854
rect 365546 510938 365782 511174
rect 365866 510938 366102 511174
rect 365546 510618 365782 510854
rect 365866 510618 366102 510854
rect 365546 474938 365782 475174
rect 365866 474938 366102 475174
rect 365546 474618 365782 474854
rect 365866 474618 366102 474854
rect 365546 438938 365782 439174
rect 365866 438938 366102 439174
rect 365546 438618 365782 438854
rect 365866 438618 366102 438854
rect 365546 402938 365782 403174
rect 365866 402938 366102 403174
rect 365546 402618 365782 402854
rect 365866 402618 366102 402854
rect 369266 694658 369502 694894
rect 369586 694658 369822 694894
rect 369266 694338 369502 694574
rect 369586 694338 369822 694574
rect 369266 658658 369502 658894
rect 369586 658658 369822 658894
rect 369266 658338 369502 658574
rect 369586 658338 369822 658574
rect 369266 622658 369502 622894
rect 369586 622658 369822 622894
rect 369266 622338 369502 622574
rect 369586 622338 369822 622574
rect 369266 586658 369502 586894
rect 369586 586658 369822 586894
rect 369266 586338 369502 586574
rect 369586 586338 369822 586574
rect 369266 550658 369502 550894
rect 369586 550658 369822 550894
rect 369266 550338 369502 550574
rect 369586 550338 369822 550574
rect 369266 514658 369502 514894
rect 369586 514658 369822 514894
rect 369266 514338 369502 514574
rect 369586 514338 369822 514574
rect 369266 478658 369502 478894
rect 369586 478658 369822 478894
rect 369266 478338 369502 478574
rect 369586 478338 369822 478574
rect 369266 442658 369502 442894
rect 369586 442658 369822 442894
rect 369266 442338 369502 442574
rect 369586 442338 369822 442574
rect 369266 406658 369502 406894
rect 369586 406658 369822 406894
rect 369266 406338 369502 406574
rect 369586 406338 369822 406574
rect 390986 711322 391222 711558
rect 391306 711322 391542 711558
rect 390986 711002 391222 711238
rect 391306 711002 391542 711238
rect 387266 709402 387502 709638
rect 387586 709402 387822 709638
rect 387266 709082 387502 709318
rect 387586 709082 387822 709318
rect 383546 707482 383782 707718
rect 383866 707482 384102 707718
rect 383546 707162 383782 707398
rect 383866 707162 384102 707398
rect 372986 698378 373222 698614
rect 373306 698378 373542 698614
rect 372986 698058 373222 698294
rect 373306 698058 373542 698294
rect 372986 662378 373222 662614
rect 373306 662378 373542 662614
rect 372986 662058 373222 662294
rect 373306 662058 373542 662294
rect 372986 626378 373222 626614
rect 373306 626378 373542 626614
rect 372986 626058 373222 626294
rect 373306 626058 373542 626294
rect 372986 590378 373222 590614
rect 373306 590378 373542 590614
rect 372986 590058 373222 590294
rect 373306 590058 373542 590294
rect 372986 554378 373222 554614
rect 373306 554378 373542 554614
rect 372986 554058 373222 554294
rect 373306 554058 373542 554294
rect 372986 518378 373222 518614
rect 373306 518378 373542 518614
rect 372986 518058 373222 518294
rect 373306 518058 373542 518294
rect 372986 482378 373222 482614
rect 373306 482378 373542 482614
rect 372986 482058 373222 482294
rect 373306 482058 373542 482294
rect 372986 446378 373222 446614
rect 373306 446378 373542 446614
rect 372986 446058 373222 446294
rect 373306 446058 373542 446294
rect 372986 410378 373222 410614
rect 373306 410378 373542 410614
rect 372986 410058 373222 410294
rect 373306 410058 373542 410294
rect 372986 374378 373222 374614
rect 373306 374378 373542 374614
rect 372986 374058 373222 374294
rect 373306 374058 373542 374294
rect 362285 363218 362521 363454
rect 362285 362898 362521 363134
rect 364882 363218 365118 363454
rect 364882 362898 365118 363134
rect 367479 363218 367715 363454
rect 367479 362898 367715 363134
rect 354986 356378 355222 356614
rect 355306 356378 355542 356614
rect 354986 356058 355222 356294
rect 355306 356058 355542 356294
rect 363583 345218 363819 345454
rect 363583 344898 363819 345134
rect 366180 345218 366416 345454
rect 366180 344898 366416 345134
rect 354986 320378 355222 320614
rect 355306 320378 355542 320614
rect 354986 320058 355222 320294
rect 355306 320058 355542 320294
rect 354986 284378 355222 284614
rect 355306 284378 355542 284614
rect 354986 284058 355222 284294
rect 355306 284058 355542 284294
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 362285 291218 362521 291454
rect 362285 290898 362521 291134
rect 363583 273218 363819 273454
rect 363583 272898 363819 273134
rect 365546 330938 365782 331174
rect 365866 330938 366102 331174
rect 365546 330618 365782 330854
rect 365866 330618 366102 330854
rect 369266 334658 369502 334894
rect 369586 334658 369822 334894
rect 369266 334338 369502 334574
rect 369586 334338 369822 334574
rect 364882 291218 365118 291454
rect 364882 290898 365118 291134
rect 367479 291218 367715 291454
rect 367479 290898 367715 291134
rect 366180 273218 366416 273454
rect 366180 272898 366416 273134
rect 354986 248378 355222 248614
rect 355306 248378 355542 248614
rect 354986 248058 355222 248294
rect 355306 248058 355542 248294
rect 354986 212378 355222 212614
rect 355306 212378 355542 212614
rect 354986 212058 355222 212294
rect 355306 212058 355542 212294
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 362285 219218 362521 219454
rect 362285 218898 362521 219134
rect 363583 201218 363819 201454
rect 363583 200898 363819 201134
rect 365546 258938 365782 259174
rect 365866 258938 366102 259174
rect 365546 258618 365782 258854
rect 365866 258618 366102 258854
rect 369266 262658 369502 262894
rect 369586 262658 369822 262894
rect 369266 262338 369502 262574
rect 369586 262338 369822 262574
rect 364882 219218 365118 219454
rect 364882 218898 365118 219134
rect 367479 219218 367715 219454
rect 367479 218898 367715 219134
rect 366180 201218 366416 201454
rect 366180 200898 366416 201134
rect 372986 338378 373222 338614
rect 373306 338378 373542 338614
rect 372986 338058 373222 338294
rect 373306 338058 373542 338294
rect 372986 302378 373222 302614
rect 373306 302378 373542 302614
rect 372986 302058 373222 302294
rect 373306 302058 373542 302294
rect 372986 266378 373222 266614
rect 373306 266378 373542 266614
rect 372986 266058 373222 266294
rect 373306 266058 373542 266294
rect 372986 230378 373222 230614
rect 373306 230378 373542 230614
rect 372986 230058 373222 230294
rect 373306 230058 373542 230294
rect 354986 176378 355222 176614
rect 355306 176378 355542 176614
rect 354986 176058 355222 176294
rect 355306 176058 355542 176294
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 362285 147218 362521 147454
rect 362285 146898 362521 147134
rect 354986 140378 355222 140614
rect 355306 140378 355542 140614
rect 354986 140058 355222 140294
rect 355306 140058 355542 140294
rect 364882 147218 365118 147454
rect 364882 146898 365118 147134
rect 363583 129218 363819 129454
rect 363583 128898 363819 129134
rect 372986 194378 373222 194614
rect 373306 194378 373542 194614
rect 372986 194058 373222 194294
rect 373306 194058 373542 194294
rect 365546 186938 365782 187174
rect 365866 186938 366102 187174
rect 365546 186618 365782 186854
rect 365866 186618 366102 186854
rect 369266 190658 369502 190894
rect 369586 190658 369822 190894
rect 369266 190338 369502 190574
rect 369586 190338 369822 190574
rect 367479 147218 367715 147454
rect 367479 146898 367715 147134
rect 366180 129218 366416 129454
rect 366180 128898 366416 129134
rect 372986 158378 373222 158614
rect 373306 158378 373542 158614
rect 372986 158058 373222 158294
rect 373306 158058 373542 158294
rect 372986 122378 373222 122614
rect 373306 122378 373542 122614
rect 372986 122058 373222 122294
rect 373306 122058 373542 122294
rect 354986 104378 355222 104614
rect 355306 104378 355542 104614
rect 354986 104058 355222 104294
rect 355306 104058 355542 104294
rect 354986 68378 355222 68614
rect 355306 68378 355542 68614
rect 354986 68058 355222 68294
rect 355306 68058 355542 68294
rect 354986 32378 355222 32614
rect 355306 32378 355542 32614
rect 354986 32058 355222 32294
rect 355306 32058 355542 32294
rect 336986 -6342 337222 -6106
rect 337306 -6342 337542 -6106
rect 336986 -6662 337222 -6426
rect 337306 -6662 337542 -6426
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 365546 114938 365782 115174
rect 365866 114938 366102 115174
rect 365546 114618 365782 114854
rect 365866 114618 366102 114854
rect 365546 78938 365782 79174
rect 365866 78938 366102 79174
rect 365546 78618 365782 78854
rect 365866 78618 366102 78854
rect 365546 42938 365782 43174
rect 365866 42938 366102 43174
rect 365546 42618 365782 42854
rect 365866 42618 366102 42854
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 365546 -2502 365782 -2266
rect 365866 -2502 366102 -2266
rect 365546 -2822 365782 -2586
rect 365866 -2822 366102 -2586
rect 369266 118658 369502 118894
rect 369586 118658 369822 118894
rect 369266 118338 369502 118574
rect 369586 118338 369822 118574
rect 369266 82658 369502 82894
rect 369586 82658 369822 82894
rect 369266 82338 369502 82574
rect 369586 82338 369822 82574
rect 369266 46658 369502 46894
rect 369586 46658 369822 46894
rect 369266 46338 369502 46574
rect 369586 46338 369822 46574
rect 369266 10658 369502 10894
rect 369586 10658 369822 10894
rect 369266 10338 369502 10574
rect 369586 10338 369822 10574
rect 369266 -4422 369502 -4186
rect 369586 -4422 369822 -4186
rect 369266 -4742 369502 -4506
rect 369586 -4742 369822 -4506
rect 372986 86378 373222 86614
rect 373306 86378 373542 86614
rect 372986 86058 373222 86294
rect 373306 86058 373542 86294
rect 372986 50378 373222 50614
rect 373306 50378 373542 50614
rect 372986 50058 373222 50294
rect 373306 50058 373542 50294
rect 372986 14378 373222 14614
rect 373306 14378 373542 14614
rect 372986 14058 373222 14294
rect 373306 14058 373542 14294
rect 354986 -7302 355222 -7066
rect 355306 -7302 355542 -7066
rect 354986 -7622 355222 -7386
rect 355306 -7622 355542 -7386
rect 379826 705562 380062 705798
rect 380146 705562 380382 705798
rect 379826 705242 380062 705478
rect 380146 705242 380382 705478
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 379826 561218 380062 561454
rect 380146 561218 380382 561454
rect 379826 560898 380062 561134
rect 380146 560898 380382 561134
rect 379826 525218 380062 525454
rect 380146 525218 380382 525454
rect 379826 524898 380062 525134
rect 380146 524898 380382 525134
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 379826 453218 380062 453454
rect 380146 453218 380382 453454
rect 379826 452898 380062 453134
rect 380146 452898 380382 453134
rect 379826 417218 380062 417454
rect 380146 417218 380382 417454
rect 379826 416898 380062 417134
rect 380146 416898 380382 417134
rect 379826 381218 380062 381454
rect 380146 381218 380382 381454
rect 379826 380898 380062 381134
rect 380146 380898 380382 381134
rect 379826 345218 380062 345454
rect 380146 345218 380382 345454
rect 379826 344898 380062 345134
rect 380146 344898 380382 345134
rect 379826 309218 380062 309454
rect 380146 309218 380382 309454
rect 379826 308898 380062 309134
rect 380146 308898 380382 309134
rect 379826 273218 380062 273454
rect 380146 273218 380382 273454
rect 379826 272898 380062 273134
rect 380146 272898 380382 273134
rect 379826 237218 380062 237454
rect 380146 237218 380382 237454
rect 379826 236898 380062 237134
rect 380146 236898 380382 237134
rect 379826 201218 380062 201454
rect 380146 201218 380382 201454
rect 379826 200898 380062 201134
rect 380146 200898 380382 201134
rect 379826 165218 380062 165454
rect 380146 165218 380382 165454
rect 379826 164898 380062 165134
rect 380146 164898 380382 165134
rect 379826 129218 380062 129454
rect 380146 129218 380382 129454
rect 379826 128898 380062 129134
rect 380146 128898 380382 129134
rect 379826 93218 380062 93454
rect 380146 93218 380382 93454
rect 379826 92898 380062 93134
rect 380146 92898 380382 93134
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -1542 380062 -1306
rect 380146 -1542 380382 -1306
rect 379826 -1862 380062 -1626
rect 380146 -1862 380382 -1626
rect 383546 672938 383782 673174
rect 383866 672938 384102 673174
rect 383546 672618 383782 672854
rect 383866 672618 384102 672854
rect 383546 636938 383782 637174
rect 383866 636938 384102 637174
rect 383546 636618 383782 636854
rect 383866 636618 384102 636854
rect 383546 600938 383782 601174
rect 383866 600938 384102 601174
rect 383546 600618 383782 600854
rect 383866 600618 384102 600854
rect 383546 564938 383782 565174
rect 383866 564938 384102 565174
rect 383546 564618 383782 564854
rect 383866 564618 384102 564854
rect 383546 528938 383782 529174
rect 383866 528938 384102 529174
rect 383546 528618 383782 528854
rect 383866 528618 384102 528854
rect 383546 492938 383782 493174
rect 383866 492938 384102 493174
rect 383546 492618 383782 492854
rect 383866 492618 384102 492854
rect 383546 456938 383782 457174
rect 383866 456938 384102 457174
rect 383546 456618 383782 456854
rect 383866 456618 384102 456854
rect 383546 420938 383782 421174
rect 383866 420938 384102 421174
rect 383546 420618 383782 420854
rect 383866 420618 384102 420854
rect 383546 384938 383782 385174
rect 383866 384938 384102 385174
rect 383546 384618 383782 384854
rect 383866 384618 384102 384854
rect 383546 348938 383782 349174
rect 383866 348938 384102 349174
rect 383546 348618 383782 348854
rect 383866 348618 384102 348854
rect 383546 312938 383782 313174
rect 383866 312938 384102 313174
rect 383546 312618 383782 312854
rect 383866 312618 384102 312854
rect 383546 276938 383782 277174
rect 383866 276938 384102 277174
rect 383546 276618 383782 276854
rect 383866 276618 384102 276854
rect 383546 240938 383782 241174
rect 383866 240938 384102 241174
rect 383546 240618 383782 240854
rect 383866 240618 384102 240854
rect 383546 204938 383782 205174
rect 383866 204938 384102 205174
rect 383546 204618 383782 204854
rect 383866 204618 384102 204854
rect 383546 168938 383782 169174
rect 383866 168938 384102 169174
rect 383546 168618 383782 168854
rect 383866 168618 384102 168854
rect 383546 132938 383782 133174
rect 383866 132938 384102 133174
rect 383546 132618 383782 132854
rect 383866 132618 384102 132854
rect 383546 96938 383782 97174
rect 383866 96938 384102 97174
rect 383546 96618 383782 96854
rect 383866 96618 384102 96854
rect 383546 60938 383782 61174
rect 383866 60938 384102 61174
rect 383546 60618 383782 60854
rect 383866 60618 384102 60854
rect 383546 24938 383782 25174
rect 383866 24938 384102 25174
rect 383546 24618 383782 24854
rect 383866 24618 384102 24854
rect 383546 -3462 383782 -3226
rect 383866 -3462 384102 -3226
rect 383546 -3782 383782 -3546
rect 383866 -3782 384102 -3546
rect 387266 676658 387502 676894
rect 387586 676658 387822 676894
rect 387266 676338 387502 676574
rect 387586 676338 387822 676574
rect 387266 640658 387502 640894
rect 387586 640658 387822 640894
rect 387266 640338 387502 640574
rect 387586 640338 387822 640574
rect 387266 604658 387502 604894
rect 387586 604658 387822 604894
rect 387266 604338 387502 604574
rect 387586 604338 387822 604574
rect 387266 568658 387502 568894
rect 387586 568658 387822 568894
rect 387266 568338 387502 568574
rect 387586 568338 387822 568574
rect 387266 532658 387502 532894
rect 387586 532658 387822 532894
rect 387266 532338 387502 532574
rect 387586 532338 387822 532574
rect 387266 496658 387502 496894
rect 387586 496658 387822 496894
rect 387266 496338 387502 496574
rect 387586 496338 387822 496574
rect 387266 460658 387502 460894
rect 387586 460658 387822 460894
rect 387266 460338 387502 460574
rect 387586 460338 387822 460574
rect 387266 424658 387502 424894
rect 387586 424658 387822 424894
rect 387266 424338 387502 424574
rect 387586 424338 387822 424574
rect 387266 388658 387502 388894
rect 387586 388658 387822 388894
rect 387266 388338 387502 388574
rect 387586 388338 387822 388574
rect 387266 352658 387502 352894
rect 387586 352658 387822 352894
rect 387266 352338 387502 352574
rect 387586 352338 387822 352574
rect 387266 316658 387502 316894
rect 387586 316658 387822 316894
rect 387266 316338 387502 316574
rect 387586 316338 387822 316574
rect 387266 280658 387502 280894
rect 387586 280658 387822 280894
rect 387266 280338 387502 280574
rect 387586 280338 387822 280574
rect 387266 244658 387502 244894
rect 387586 244658 387822 244894
rect 387266 244338 387502 244574
rect 387586 244338 387822 244574
rect 387266 208658 387502 208894
rect 387586 208658 387822 208894
rect 387266 208338 387502 208574
rect 387586 208338 387822 208574
rect 387266 172658 387502 172894
rect 387586 172658 387822 172894
rect 387266 172338 387502 172574
rect 387586 172338 387822 172574
rect 387266 136658 387502 136894
rect 387586 136658 387822 136894
rect 387266 136338 387502 136574
rect 387586 136338 387822 136574
rect 387266 100658 387502 100894
rect 387586 100658 387822 100894
rect 387266 100338 387502 100574
rect 387586 100338 387822 100574
rect 387266 64658 387502 64894
rect 387586 64658 387822 64894
rect 387266 64338 387502 64574
rect 387586 64338 387822 64574
rect 387266 28658 387502 28894
rect 387586 28658 387822 28894
rect 387266 28338 387502 28574
rect 387586 28338 387822 28574
rect 387266 -5382 387502 -5146
rect 387586 -5382 387822 -5146
rect 387266 -5702 387502 -5466
rect 387586 -5702 387822 -5466
rect 408986 710362 409222 710598
rect 409306 710362 409542 710598
rect 408986 710042 409222 710278
rect 409306 710042 409542 710278
rect 405266 708442 405502 708678
rect 405586 708442 405822 708678
rect 405266 708122 405502 708358
rect 405586 708122 405822 708358
rect 401546 706522 401782 706758
rect 401866 706522 402102 706758
rect 401546 706202 401782 706438
rect 401866 706202 402102 706438
rect 390986 680378 391222 680614
rect 391306 680378 391542 680614
rect 390986 680058 391222 680294
rect 391306 680058 391542 680294
rect 390986 644378 391222 644614
rect 391306 644378 391542 644614
rect 390986 644058 391222 644294
rect 391306 644058 391542 644294
rect 390986 608378 391222 608614
rect 391306 608378 391542 608614
rect 390986 608058 391222 608294
rect 391306 608058 391542 608294
rect 390986 572378 391222 572614
rect 391306 572378 391542 572614
rect 390986 572058 391222 572294
rect 391306 572058 391542 572294
rect 390986 536378 391222 536614
rect 391306 536378 391542 536614
rect 390986 536058 391222 536294
rect 391306 536058 391542 536294
rect 390986 500378 391222 500614
rect 391306 500378 391542 500614
rect 390986 500058 391222 500294
rect 391306 500058 391542 500294
rect 390986 464378 391222 464614
rect 391306 464378 391542 464614
rect 390986 464058 391222 464294
rect 391306 464058 391542 464294
rect 390986 428378 391222 428614
rect 391306 428378 391542 428614
rect 390986 428058 391222 428294
rect 391306 428058 391542 428294
rect 390986 392378 391222 392614
rect 391306 392378 391542 392614
rect 390986 392058 391222 392294
rect 391306 392058 391542 392294
rect 390986 356378 391222 356614
rect 391306 356378 391542 356614
rect 390986 356058 391222 356294
rect 391306 356058 391542 356294
rect 390986 320378 391222 320614
rect 391306 320378 391542 320614
rect 390986 320058 391222 320294
rect 391306 320058 391542 320294
rect 390986 284378 391222 284614
rect 391306 284378 391542 284614
rect 390986 284058 391222 284294
rect 391306 284058 391542 284294
rect 390986 248378 391222 248614
rect 391306 248378 391542 248614
rect 390986 248058 391222 248294
rect 391306 248058 391542 248294
rect 390986 212378 391222 212614
rect 391306 212378 391542 212614
rect 390986 212058 391222 212294
rect 391306 212058 391542 212294
rect 390986 176378 391222 176614
rect 391306 176378 391542 176614
rect 390986 176058 391222 176294
rect 391306 176058 391542 176294
rect 390986 140378 391222 140614
rect 391306 140378 391542 140614
rect 390986 140058 391222 140294
rect 391306 140058 391542 140294
rect 390986 104378 391222 104614
rect 391306 104378 391542 104614
rect 390986 104058 391222 104294
rect 391306 104058 391542 104294
rect 390986 68378 391222 68614
rect 391306 68378 391542 68614
rect 390986 68058 391222 68294
rect 391306 68058 391542 68294
rect 390986 32378 391222 32614
rect 391306 32378 391542 32614
rect 390986 32058 391222 32294
rect 391306 32058 391542 32294
rect 372986 -6342 373222 -6106
rect 373306 -6342 373542 -6106
rect 372986 -6662 373222 -6426
rect 373306 -6662 373542 -6426
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 690938 401782 691174
rect 401866 690938 402102 691174
rect 401546 690618 401782 690854
rect 401866 690618 402102 690854
rect 401546 654938 401782 655174
rect 401866 654938 402102 655174
rect 401546 654618 401782 654854
rect 401866 654618 402102 654854
rect 401546 618938 401782 619174
rect 401866 618938 402102 619174
rect 401546 618618 401782 618854
rect 401866 618618 402102 618854
rect 401546 582938 401782 583174
rect 401866 582938 402102 583174
rect 401546 582618 401782 582854
rect 401866 582618 402102 582854
rect 401546 546938 401782 547174
rect 401866 546938 402102 547174
rect 401546 546618 401782 546854
rect 401866 546618 402102 546854
rect 401546 510938 401782 511174
rect 401866 510938 402102 511174
rect 401546 510618 401782 510854
rect 401866 510618 402102 510854
rect 401546 474938 401782 475174
rect 401866 474938 402102 475174
rect 401546 474618 401782 474854
rect 401866 474618 402102 474854
rect 401546 438938 401782 439174
rect 401866 438938 402102 439174
rect 401546 438618 401782 438854
rect 401866 438618 402102 438854
rect 401546 402938 401782 403174
rect 401866 402938 402102 403174
rect 401546 402618 401782 402854
rect 401866 402618 402102 402854
rect 401546 366938 401782 367174
rect 401866 366938 402102 367174
rect 401546 366618 401782 366854
rect 401866 366618 402102 366854
rect 401546 330938 401782 331174
rect 401866 330938 402102 331174
rect 401546 330618 401782 330854
rect 401866 330618 402102 330854
rect 401546 294938 401782 295174
rect 401866 294938 402102 295174
rect 401546 294618 401782 294854
rect 401866 294618 402102 294854
rect 401546 258938 401782 259174
rect 401866 258938 402102 259174
rect 401546 258618 401782 258854
rect 401866 258618 402102 258854
rect 401546 222938 401782 223174
rect 401866 222938 402102 223174
rect 401546 222618 401782 222854
rect 401866 222618 402102 222854
rect 401546 186938 401782 187174
rect 401866 186938 402102 187174
rect 401546 186618 401782 186854
rect 401866 186618 402102 186854
rect 401546 150938 401782 151174
rect 401866 150938 402102 151174
rect 401546 150618 401782 150854
rect 401866 150618 402102 150854
rect 401546 114938 401782 115174
rect 401866 114938 402102 115174
rect 401546 114618 401782 114854
rect 401866 114618 402102 114854
rect 401546 78938 401782 79174
rect 401866 78938 402102 79174
rect 401546 78618 401782 78854
rect 401866 78618 402102 78854
rect 401546 42938 401782 43174
rect 401866 42938 402102 43174
rect 401546 42618 401782 42854
rect 401866 42618 402102 42854
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 401546 -2502 401782 -2266
rect 401866 -2502 402102 -2266
rect 401546 -2822 401782 -2586
rect 401866 -2822 402102 -2586
rect 405266 694658 405502 694894
rect 405586 694658 405822 694894
rect 405266 694338 405502 694574
rect 405586 694338 405822 694574
rect 405266 658658 405502 658894
rect 405586 658658 405822 658894
rect 405266 658338 405502 658574
rect 405586 658338 405822 658574
rect 405266 622658 405502 622894
rect 405586 622658 405822 622894
rect 405266 622338 405502 622574
rect 405586 622338 405822 622574
rect 405266 586658 405502 586894
rect 405586 586658 405822 586894
rect 405266 586338 405502 586574
rect 405586 586338 405822 586574
rect 405266 550658 405502 550894
rect 405586 550658 405822 550894
rect 405266 550338 405502 550574
rect 405586 550338 405822 550574
rect 405266 514658 405502 514894
rect 405586 514658 405822 514894
rect 405266 514338 405502 514574
rect 405586 514338 405822 514574
rect 405266 478658 405502 478894
rect 405586 478658 405822 478894
rect 405266 478338 405502 478574
rect 405586 478338 405822 478574
rect 405266 442658 405502 442894
rect 405586 442658 405822 442894
rect 405266 442338 405502 442574
rect 405586 442338 405822 442574
rect 405266 406658 405502 406894
rect 405586 406658 405822 406894
rect 405266 406338 405502 406574
rect 405586 406338 405822 406574
rect 405266 370658 405502 370894
rect 405586 370658 405822 370894
rect 405266 370338 405502 370574
rect 405586 370338 405822 370574
rect 405266 334658 405502 334894
rect 405586 334658 405822 334894
rect 405266 334338 405502 334574
rect 405586 334338 405822 334574
rect 405266 298658 405502 298894
rect 405586 298658 405822 298894
rect 405266 298338 405502 298574
rect 405586 298338 405822 298574
rect 405266 262658 405502 262894
rect 405586 262658 405822 262894
rect 405266 262338 405502 262574
rect 405586 262338 405822 262574
rect 405266 226658 405502 226894
rect 405586 226658 405822 226894
rect 405266 226338 405502 226574
rect 405586 226338 405822 226574
rect 405266 190658 405502 190894
rect 405586 190658 405822 190894
rect 405266 190338 405502 190574
rect 405586 190338 405822 190574
rect 405266 154658 405502 154894
rect 405586 154658 405822 154894
rect 405266 154338 405502 154574
rect 405586 154338 405822 154574
rect 405266 118658 405502 118894
rect 405586 118658 405822 118894
rect 405266 118338 405502 118574
rect 405586 118338 405822 118574
rect 405266 82658 405502 82894
rect 405586 82658 405822 82894
rect 405266 82338 405502 82574
rect 405586 82338 405822 82574
rect 405266 46658 405502 46894
rect 405586 46658 405822 46894
rect 405266 46338 405502 46574
rect 405586 46338 405822 46574
rect 405266 10658 405502 10894
rect 405586 10658 405822 10894
rect 405266 10338 405502 10574
rect 405586 10338 405822 10574
rect 405266 -4422 405502 -4186
rect 405586 -4422 405822 -4186
rect 405266 -4742 405502 -4506
rect 405586 -4742 405822 -4506
rect 426986 711322 427222 711558
rect 427306 711322 427542 711558
rect 426986 711002 427222 711238
rect 427306 711002 427542 711238
rect 423266 709402 423502 709638
rect 423586 709402 423822 709638
rect 423266 709082 423502 709318
rect 423586 709082 423822 709318
rect 419546 707482 419782 707718
rect 419866 707482 420102 707718
rect 419546 707162 419782 707398
rect 419866 707162 420102 707398
rect 408986 698378 409222 698614
rect 409306 698378 409542 698614
rect 408986 698058 409222 698294
rect 409306 698058 409542 698294
rect 408986 662378 409222 662614
rect 409306 662378 409542 662614
rect 408986 662058 409222 662294
rect 409306 662058 409542 662294
rect 408986 626378 409222 626614
rect 409306 626378 409542 626614
rect 408986 626058 409222 626294
rect 409306 626058 409542 626294
rect 408986 590378 409222 590614
rect 409306 590378 409542 590614
rect 408986 590058 409222 590294
rect 409306 590058 409542 590294
rect 408986 554378 409222 554614
rect 409306 554378 409542 554614
rect 408986 554058 409222 554294
rect 409306 554058 409542 554294
rect 408986 518378 409222 518614
rect 409306 518378 409542 518614
rect 408986 518058 409222 518294
rect 409306 518058 409542 518294
rect 408986 482378 409222 482614
rect 409306 482378 409542 482614
rect 408986 482058 409222 482294
rect 409306 482058 409542 482294
rect 408986 446378 409222 446614
rect 409306 446378 409542 446614
rect 408986 446058 409222 446294
rect 409306 446058 409542 446294
rect 408986 410378 409222 410614
rect 409306 410378 409542 410614
rect 408986 410058 409222 410294
rect 409306 410058 409542 410294
rect 408986 374378 409222 374614
rect 409306 374378 409542 374614
rect 408986 374058 409222 374294
rect 409306 374058 409542 374294
rect 408986 338378 409222 338614
rect 409306 338378 409542 338614
rect 408986 338058 409222 338294
rect 409306 338058 409542 338294
rect 408986 302378 409222 302614
rect 409306 302378 409542 302614
rect 408986 302058 409222 302294
rect 409306 302058 409542 302294
rect 408986 266378 409222 266614
rect 409306 266378 409542 266614
rect 408986 266058 409222 266294
rect 409306 266058 409542 266294
rect 408986 230378 409222 230614
rect 409306 230378 409542 230614
rect 408986 230058 409222 230294
rect 409306 230058 409542 230294
rect 408986 194378 409222 194614
rect 409306 194378 409542 194614
rect 408986 194058 409222 194294
rect 409306 194058 409542 194294
rect 408986 158378 409222 158614
rect 409306 158378 409542 158614
rect 408986 158058 409222 158294
rect 409306 158058 409542 158294
rect 408986 122378 409222 122614
rect 409306 122378 409542 122614
rect 408986 122058 409222 122294
rect 409306 122058 409542 122294
rect 408986 86378 409222 86614
rect 409306 86378 409542 86614
rect 408986 86058 409222 86294
rect 409306 86058 409542 86294
rect 408986 50378 409222 50614
rect 409306 50378 409542 50614
rect 408986 50058 409222 50294
rect 409306 50058 409542 50294
rect 408986 14378 409222 14614
rect 409306 14378 409542 14614
rect 408986 14058 409222 14294
rect 409306 14058 409542 14294
rect 390986 -7302 391222 -7066
rect 391306 -7302 391542 -7066
rect 390986 -7622 391222 -7386
rect 391306 -7622 391542 -7386
rect 415826 705562 416062 705798
rect 416146 705562 416382 705798
rect 415826 705242 416062 705478
rect 416146 705242 416382 705478
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 415826 561218 416062 561454
rect 416146 561218 416382 561454
rect 415826 560898 416062 561134
rect 416146 560898 416382 561134
rect 415826 525218 416062 525454
rect 416146 525218 416382 525454
rect 415826 524898 416062 525134
rect 416146 524898 416382 525134
rect 415826 489218 416062 489454
rect 416146 489218 416382 489454
rect 415826 488898 416062 489134
rect 416146 488898 416382 489134
rect 415826 453218 416062 453454
rect 416146 453218 416382 453454
rect 415826 452898 416062 453134
rect 416146 452898 416382 453134
rect 415826 417218 416062 417454
rect 416146 417218 416382 417454
rect 415826 416898 416062 417134
rect 416146 416898 416382 417134
rect 415826 381218 416062 381454
rect 416146 381218 416382 381454
rect 415826 380898 416062 381134
rect 416146 380898 416382 381134
rect 415826 345218 416062 345454
rect 416146 345218 416382 345454
rect 415826 344898 416062 345134
rect 416146 344898 416382 345134
rect 415826 309218 416062 309454
rect 416146 309218 416382 309454
rect 415826 308898 416062 309134
rect 416146 308898 416382 309134
rect 415826 273218 416062 273454
rect 416146 273218 416382 273454
rect 415826 272898 416062 273134
rect 416146 272898 416382 273134
rect 415826 237218 416062 237454
rect 416146 237218 416382 237454
rect 415826 236898 416062 237134
rect 416146 236898 416382 237134
rect 415826 201218 416062 201454
rect 416146 201218 416382 201454
rect 415826 200898 416062 201134
rect 416146 200898 416382 201134
rect 415826 165218 416062 165454
rect 416146 165218 416382 165454
rect 415826 164898 416062 165134
rect 416146 164898 416382 165134
rect 415826 129218 416062 129454
rect 416146 129218 416382 129454
rect 415826 128898 416062 129134
rect 416146 128898 416382 129134
rect 415826 93218 416062 93454
rect 416146 93218 416382 93454
rect 415826 92898 416062 93134
rect 416146 92898 416382 93134
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -1542 416062 -1306
rect 416146 -1542 416382 -1306
rect 415826 -1862 416062 -1626
rect 416146 -1862 416382 -1626
rect 419546 672938 419782 673174
rect 419866 672938 420102 673174
rect 419546 672618 419782 672854
rect 419866 672618 420102 672854
rect 419546 636938 419782 637174
rect 419866 636938 420102 637174
rect 419546 636618 419782 636854
rect 419866 636618 420102 636854
rect 419546 600938 419782 601174
rect 419866 600938 420102 601174
rect 419546 600618 419782 600854
rect 419866 600618 420102 600854
rect 419546 564938 419782 565174
rect 419866 564938 420102 565174
rect 419546 564618 419782 564854
rect 419866 564618 420102 564854
rect 419546 528938 419782 529174
rect 419866 528938 420102 529174
rect 419546 528618 419782 528854
rect 419866 528618 420102 528854
rect 419546 492938 419782 493174
rect 419866 492938 420102 493174
rect 419546 492618 419782 492854
rect 419866 492618 420102 492854
rect 419546 456938 419782 457174
rect 419866 456938 420102 457174
rect 419546 456618 419782 456854
rect 419866 456618 420102 456854
rect 419546 420938 419782 421174
rect 419866 420938 420102 421174
rect 419546 420618 419782 420854
rect 419866 420618 420102 420854
rect 419546 384938 419782 385174
rect 419866 384938 420102 385174
rect 419546 384618 419782 384854
rect 419866 384618 420102 384854
rect 419546 348938 419782 349174
rect 419866 348938 420102 349174
rect 419546 348618 419782 348854
rect 419866 348618 420102 348854
rect 419546 312938 419782 313174
rect 419866 312938 420102 313174
rect 419546 312618 419782 312854
rect 419866 312618 420102 312854
rect 419546 276938 419782 277174
rect 419866 276938 420102 277174
rect 419546 276618 419782 276854
rect 419866 276618 420102 276854
rect 419546 240938 419782 241174
rect 419866 240938 420102 241174
rect 419546 240618 419782 240854
rect 419866 240618 420102 240854
rect 419546 204938 419782 205174
rect 419866 204938 420102 205174
rect 419546 204618 419782 204854
rect 419866 204618 420102 204854
rect 419546 168938 419782 169174
rect 419866 168938 420102 169174
rect 419546 168618 419782 168854
rect 419866 168618 420102 168854
rect 419546 132938 419782 133174
rect 419866 132938 420102 133174
rect 419546 132618 419782 132854
rect 419866 132618 420102 132854
rect 419546 96938 419782 97174
rect 419866 96938 420102 97174
rect 419546 96618 419782 96854
rect 419866 96618 420102 96854
rect 419546 60938 419782 61174
rect 419866 60938 420102 61174
rect 419546 60618 419782 60854
rect 419866 60618 420102 60854
rect 419546 24938 419782 25174
rect 419866 24938 420102 25174
rect 419546 24618 419782 24854
rect 419866 24618 420102 24854
rect 419546 -3462 419782 -3226
rect 419866 -3462 420102 -3226
rect 419546 -3782 419782 -3546
rect 419866 -3782 420102 -3546
rect 423266 676658 423502 676894
rect 423586 676658 423822 676894
rect 423266 676338 423502 676574
rect 423586 676338 423822 676574
rect 423266 640658 423502 640894
rect 423586 640658 423822 640894
rect 423266 640338 423502 640574
rect 423586 640338 423822 640574
rect 423266 604658 423502 604894
rect 423586 604658 423822 604894
rect 423266 604338 423502 604574
rect 423586 604338 423822 604574
rect 423266 568658 423502 568894
rect 423586 568658 423822 568894
rect 423266 568338 423502 568574
rect 423586 568338 423822 568574
rect 423266 532658 423502 532894
rect 423586 532658 423822 532894
rect 423266 532338 423502 532574
rect 423586 532338 423822 532574
rect 423266 496658 423502 496894
rect 423586 496658 423822 496894
rect 423266 496338 423502 496574
rect 423586 496338 423822 496574
rect 423266 460658 423502 460894
rect 423586 460658 423822 460894
rect 423266 460338 423502 460574
rect 423586 460338 423822 460574
rect 423266 424658 423502 424894
rect 423586 424658 423822 424894
rect 423266 424338 423502 424574
rect 423586 424338 423822 424574
rect 423266 388658 423502 388894
rect 423586 388658 423822 388894
rect 423266 388338 423502 388574
rect 423586 388338 423822 388574
rect 423266 352658 423502 352894
rect 423586 352658 423822 352894
rect 423266 352338 423502 352574
rect 423586 352338 423822 352574
rect 423266 316658 423502 316894
rect 423586 316658 423822 316894
rect 423266 316338 423502 316574
rect 423586 316338 423822 316574
rect 423266 280658 423502 280894
rect 423586 280658 423822 280894
rect 423266 280338 423502 280574
rect 423586 280338 423822 280574
rect 423266 244658 423502 244894
rect 423586 244658 423822 244894
rect 423266 244338 423502 244574
rect 423586 244338 423822 244574
rect 423266 208658 423502 208894
rect 423586 208658 423822 208894
rect 423266 208338 423502 208574
rect 423586 208338 423822 208574
rect 423266 172658 423502 172894
rect 423586 172658 423822 172894
rect 423266 172338 423502 172574
rect 423586 172338 423822 172574
rect 423266 136658 423502 136894
rect 423586 136658 423822 136894
rect 423266 136338 423502 136574
rect 423586 136338 423822 136574
rect 423266 100658 423502 100894
rect 423586 100658 423822 100894
rect 423266 100338 423502 100574
rect 423586 100338 423822 100574
rect 423266 64658 423502 64894
rect 423586 64658 423822 64894
rect 423266 64338 423502 64574
rect 423586 64338 423822 64574
rect 423266 28658 423502 28894
rect 423586 28658 423822 28894
rect 423266 28338 423502 28574
rect 423586 28338 423822 28574
rect 423266 -5382 423502 -5146
rect 423586 -5382 423822 -5146
rect 423266 -5702 423502 -5466
rect 423586 -5702 423822 -5466
rect 444986 710362 445222 710598
rect 445306 710362 445542 710598
rect 444986 710042 445222 710278
rect 445306 710042 445542 710278
rect 441266 708442 441502 708678
rect 441586 708442 441822 708678
rect 441266 708122 441502 708358
rect 441586 708122 441822 708358
rect 437546 706522 437782 706758
rect 437866 706522 438102 706758
rect 437546 706202 437782 706438
rect 437866 706202 438102 706438
rect 426986 680378 427222 680614
rect 427306 680378 427542 680614
rect 426986 680058 427222 680294
rect 427306 680058 427542 680294
rect 426986 644378 427222 644614
rect 427306 644378 427542 644614
rect 426986 644058 427222 644294
rect 427306 644058 427542 644294
rect 426986 608378 427222 608614
rect 427306 608378 427542 608614
rect 426986 608058 427222 608294
rect 427306 608058 427542 608294
rect 426986 572378 427222 572614
rect 427306 572378 427542 572614
rect 426986 572058 427222 572294
rect 427306 572058 427542 572294
rect 426986 536378 427222 536614
rect 427306 536378 427542 536614
rect 426986 536058 427222 536294
rect 427306 536058 427542 536294
rect 426986 500378 427222 500614
rect 427306 500378 427542 500614
rect 426986 500058 427222 500294
rect 427306 500058 427542 500294
rect 426986 464378 427222 464614
rect 427306 464378 427542 464614
rect 426986 464058 427222 464294
rect 427306 464058 427542 464294
rect 426986 428378 427222 428614
rect 427306 428378 427542 428614
rect 426986 428058 427222 428294
rect 427306 428058 427542 428294
rect 426986 392378 427222 392614
rect 427306 392378 427542 392614
rect 426986 392058 427222 392294
rect 427306 392058 427542 392294
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 433826 435218 434062 435454
rect 434146 435218 434382 435454
rect 433826 434898 434062 435134
rect 434146 434898 434382 435134
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 437546 690938 437782 691174
rect 437866 690938 438102 691174
rect 437546 690618 437782 690854
rect 437866 690618 438102 690854
rect 437546 654938 437782 655174
rect 437866 654938 438102 655174
rect 437546 654618 437782 654854
rect 437866 654618 438102 654854
rect 437546 618938 437782 619174
rect 437866 618938 438102 619174
rect 437546 618618 437782 618854
rect 437866 618618 438102 618854
rect 437546 582938 437782 583174
rect 437866 582938 438102 583174
rect 437546 582618 437782 582854
rect 437866 582618 438102 582854
rect 437546 546938 437782 547174
rect 437866 546938 438102 547174
rect 437546 546618 437782 546854
rect 437866 546618 438102 546854
rect 437546 510938 437782 511174
rect 437866 510938 438102 511174
rect 437546 510618 437782 510854
rect 437866 510618 438102 510854
rect 437546 474938 437782 475174
rect 437866 474938 438102 475174
rect 437546 474618 437782 474854
rect 437866 474618 438102 474854
rect 437546 438938 437782 439174
rect 437866 438938 438102 439174
rect 437546 438618 437782 438854
rect 437866 438618 438102 438854
rect 437546 402938 437782 403174
rect 437866 402938 438102 403174
rect 437546 402618 437782 402854
rect 437866 402618 438102 402854
rect 441266 694658 441502 694894
rect 441586 694658 441822 694894
rect 441266 694338 441502 694574
rect 441586 694338 441822 694574
rect 441266 658658 441502 658894
rect 441586 658658 441822 658894
rect 441266 658338 441502 658574
rect 441586 658338 441822 658574
rect 441266 622658 441502 622894
rect 441586 622658 441822 622894
rect 441266 622338 441502 622574
rect 441586 622338 441822 622574
rect 441266 586658 441502 586894
rect 441586 586658 441822 586894
rect 441266 586338 441502 586574
rect 441586 586338 441822 586574
rect 441266 550658 441502 550894
rect 441586 550658 441822 550894
rect 441266 550338 441502 550574
rect 441586 550338 441822 550574
rect 441266 514658 441502 514894
rect 441586 514658 441822 514894
rect 441266 514338 441502 514574
rect 441586 514338 441822 514574
rect 441266 478658 441502 478894
rect 441586 478658 441822 478894
rect 441266 478338 441502 478574
rect 441586 478338 441822 478574
rect 441266 442658 441502 442894
rect 441586 442658 441822 442894
rect 441266 442338 441502 442574
rect 441586 442338 441822 442574
rect 441266 406658 441502 406894
rect 441586 406658 441822 406894
rect 441266 406338 441502 406574
rect 441586 406338 441822 406574
rect 462986 711322 463222 711558
rect 463306 711322 463542 711558
rect 462986 711002 463222 711238
rect 463306 711002 463542 711238
rect 459266 709402 459502 709638
rect 459586 709402 459822 709638
rect 459266 709082 459502 709318
rect 459586 709082 459822 709318
rect 455546 707482 455782 707718
rect 455866 707482 456102 707718
rect 455546 707162 455782 707398
rect 455866 707162 456102 707398
rect 444986 698378 445222 698614
rect 445306 698378 445542 698614
rect 444986 698058 445222 698294
rect 445306 698058 445542 698294
rect 444986 662378 445222 662614
rect 445306 662378 445542 662614
rect 444986 662058 445222 662294
rect 445306 662058 445542 662294
rect 444986 626378 445222 626614
rect 445306 626378 445542 626614
rect 444986 626058 445222 626294
rect 445306 626058 445542 626294
rect 444986 590378 445222 590614
rect 445306 590378 445542 590614
rect 444986 590058 445222 590294
rect 445306 590058 445542 590294
rect 444986 554378 445222 554614
rect 445306 554378 445542 554614
rect 444986 554058 445222 554294
rect 445306 554058 445542 554294
rect 444986 518378 445222 518614
rect 445306 518378 445542 518614
rect 444986 518058 445222 518294
rect 445306 518058 445542 518294
rect 444986 482378 445222 482614
rect 445306 482378 445542 482614
rect 444986 482058 445222 482294
rect 445306 482058 445542 482294
rect 444986 446378 445222 446614
rect 445306 446378 445542 446614
rect 444986 446058 445222 446294
rect 445306 446058 445542 446294
rect 444986 410378 445222 410614
rect 445306 410378 445542 410614
rect 444986 410058 445222 410294
rect 445306 410058 445542 410294
rect 444986 374378 445222 374614
rect 445306 374378 445542 374614
rect 444986 374058 445222 374294
rect 445306 374058 445542 374294
rect 434285 363218 434521 363454
rect 434285 362898 434521 363134
rect 436882 363218 437118 363454
rect 436882 362898 437118 363134
rect 439479 363218 439715 363454
rect 439479 362898 439715 363134
rect 426986 356378 427222 356614
rect 427306 356378 427542 356614
rect 426986 356058 427222 356294
rect 427306 356058 427542 356294
rect 435583 345218 435819 345454
rect 435583 344898 435819 345134
rect 438180 345218 438416 345454
rect 438180 344898 438416 345134
rect 444986 338378 445222 338614
rect 445306 338378 445542 338614
rect 444986 338058 445222 338294
rect 445306 338058 445542 338294
rect 426986 320378 427222 320614
rect 427306 320378 427542 320614
rect 426986 320058 427222 320294
rect 427306 320058 427542 320294
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 437546 330938 437782 331174
rect 437866 330938 438102 331174
rect 437546 330618 437782 330854
rect 437866 330618 438102 330854
rect 441266 334658 441502 334894
rect 441586 334658 441822 334894
rect 441266 334338 441502 334574
rect 441586 334338 441822 334574
rect 444986 302378 445222 302614
rect 445306 302378 445542 302614
rect 444986 302058 445222 302294
rect 445306 302058 445542 302294
rect 434285 291218 434521 291454
rect 434285 290898 434521 291134
rect 436882 291218 437118 291454
rect 436882 290898 437118 291134
rect 439479 291218 439715 291454
rect 439479 290898 439715 291134
rect 426986 284378 427222 284614
rect 427306 284378 427542 284614
rect 426986 284058 427222 284294
rect 427306 284058 427542 284294
rect 435583 273218 435819 273454
rect 435583 272898 435819 273134
rect 438180 273218 438416 273454
rect 438180 272898 438416 273134
rect 444986 266378 445222 266614
rect 445306 266378 445542 266614
rect 444986 266058 445222 266294
rect 445306 266058 445542 266294
rect 426986 248378 427222 248614
rect 427306 248378 427542 248614
rect 426986 248058 427222 248294
rect 427306 248058 427542 248294
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 437546 258938 437782 259174
rect 437866 258938 438102 259174
rect 437546 258618 437782 258854
rect 437866 258618 438102 258854
rect 441266 262658 441502 262894
rect 441586 262658 441822 262894
rect 441266 262338 441502 262574
rect 441586 262338 441822 262574
rect 444986 230378 445222 230614
rect 445306 230378 445542 230614
rect 444986 230058 445222 230294
rect 445306 230058 445542 230294
rect 434285 219218 434521 219454
rect 434285 218898 434521 219134
rect 436882 219218 437118 219454
rect 436882 218898 437118 219134
rect 439479 219218 439715 219454
rect 439479 218898 439715 219134
rect 426986 212378 427222 212614
rect 427306 212378 427542 212614
rect 426986 212058 427222 212294
rect 427306 212058 427542 212294
rect 435583 201218 435819 201454
rect 435583 200898 435819 201134
rect 438180 201218 438416 201454
rect 438180 200898 438416 201134
rect 444986 194378 445222 194614
rect 445306 194378 445542 194614
rect 444986 194058 445222 194294
rect 445306 194058 445542 194294
rect 426986 176378 427222 176614
rect 427306 176378 427542 176614
rect 426986 176058 427222 176294
rect 427306 176058 427542 176294
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 437546 186938 437782 187174
rect 437866 186938 438102 187174
rect 437546 186618 437782 186854
rect 437866 186618 438102 186854
rect 441266 190658 441502 190894
rect 441586 190658 441822 190894
rect 441266 190338 441502 190574
rect 441586 190338 441822 190574
rect 444986 158378 445222 158614
rect 445306 158378 445542 158614
rect 444986 158058 445222 158294
rect 445306 158058 445542 158294
rect 434285 147218 434521 147454
rect 434285 146898 434521 147134
rect 436882 147218 437118 147454
rect 436882 146898 437118 147134
rect 439479 147218 439715 147454
rect 439479 146898 439715 147134
rect 426986 140378 427222 140614
rect 427306 140378 427542 140614
rect 426986 140058 427222 140294
rect 427306 140058 427542 140294
rect 435583 129218 435819 129454
rect 435583 128898 435819 129134
rect 438180 129218 438416 129454
rect 438180 128898 438416 129134
rect 444986 122378 445222 122614
rect 445306 122378 445542 122614
rect 444986 122058 445222 122294
rect 445306 122058 445542 122294
rect 426986 104378 427222 104614
rect 427306 104378 427542 104614
rect 426986 104058 427222 104294
rect 427306 104058 427542 104294
rect 426986 68378 427222 68614
rect 427306 68378 427542 68614
rect 426986 68058 427222 68294
rect 427306 68058 427542 68294
rect 426986 32378 427222 32614
rect 427306 32378 427542 32614
rect 426986 32058 427222 32294
rect 427306 32058 427542 32294
rect 408986 -6342 409222 -6106
rect 409306 -6342 409542 -6106
rect 408986 -6662 409222 -6426
rect 409306 -6662 409542 -6426
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 437546 114938 437782 115174
rect 437866 114938 438102 115174
rect 437546 114618 437782 114854
rect 437866 114618 438102 114854
rect 437546 78938 437782 79174
rect 437866 78938 438102 79174
rect 437546 78618 437782 78854
rect 437866 78618 438102 78854
rect 437546 42938 437782 43174
rect 437866 42938 438102 43174
rect 437546 42618 437782 42854
rect 437866 42618 438102 42854
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 437546 -2502 437782 -2266
rect 437866 -2502 438102 -2266
rect 437546 -2822 437782 -2586
rect 437866 -2822 438102 -2586
rect 441266 118658 441502 118894
rect 441586 118658 441822 118894
rect 441266 118338 441502 118574
rect 441586 118338 441822 118574
rect 441266 82658 441502 82894
rect 441586 82658 441822 82894
rect 441266 82338 441502 82574
rect 441586 82338 441822 82574
rect 441266 46658 441502 46894
rect 441586 46658 441822 46894
rect 441266 46338 441502 46574
rect 441586 46338 441822 46574
rect 441266 10658 441502 10894
rect 441586 10658 441822 10894
rect 441266 10338 441502 10574
rect 441586 10338 441822 10574
rect 441266 -4422 441502 -4186
rect 441586 -4422 441822 -4186
rect 441266 -4742 441502 -4506
rect 441586 -4742 441822 -4506
rect 444986 86378 445222 86614
rect 445306 86378 445542 86614
rect 444986 86058 445222 86294
rect 445306 86058 445542 86294
rect 444986 50378 445222 50614
rect 445306 50378 445542 50614
rect 444986 50058 445222 50294
rect 445306 50058 445542 50294
rect 444986 14378 445222 14614
rect 445306 14378 445542 14614
rect 444986 14058 445222 14294
rect 445306 14058 445542 14294
rect 426986 -7302 427222 -7066
rect 427306 -7302 427542 -7066
rect 426986 -7622 427222 -7386
rect 427306 -7622 427542 -7386
rect 451826 705562 452062 705798
rect 452146 705562 452382 705798
rect 451826 705242 452062 705478
rect 452146 705242 452382 705478
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 451826 453218 452062 453454
rect 452146 453218 452382 453454
rect 451826 452898 452062 453134
rect 452146 452898 452382 453134
rect 451826 417218 452062 417454
rect 452146 417218 452382 417454
rect 451826 416898 452062 417134
rect 452146 416898 452382 417134
rect 451826 381218 452062 381454
rect 452146 381218 452382 381454
rect 451826 380898 452062 381134
rect 452146 380898 452382 381134
rect 451826 345218 452062 345454
rect 452146 345218 452382 345454
rect 451826 344898 452062 345134
rect 452146 344898 452382 345134
rect 451826 309218 452062 309454
rect 452146 309218 452382 309454
rect 451826 308898 452062 309134
rect 452146 308898 452382 309134
rect 451826 273218 452062 273454
rect 452146 273218 452382 273454
rect 451826 272898 452062 273134
rect 452146 272898 452382 273134
rect 451826 237218 452062 237454
rect 452146 237218 452382 237454
rect 451826 236898 452062 237134
rect 452146 236898 452382 237134
rect 451826 201218 452062 201454
rect 452146 201218 452382 201454
rect 451826 200898 452062 201134
rect 452146 200898 452382 201134
rect 451826 165218 452062 165454
rect 452146 165218 452382 165454
rect 451826 164898 452062 165134
rect 452146 164898 452382 165134
rect 451826 129218 452062 129454
rect 452146 129218 452382 129454
rect 451826 128898 452062 129134
rect 452146 128898 452382 129134
rect 451826 93218 452062 93454
rect 452146 93218 452382 93454
rect 451826 92898 452062 93134
rect 452146 92898 452382 93134
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -1542 452062 -1306
rect 452146 -1542 452382 -1306
rect 451826 -1862 452062 -1626
rect 452146 -1862 452382 -1626
rect 455546 672938 455782 673174
rect 455866 672938 456102 673174
rect 455546 672618 455782 672854
rect 455866 672618 456102 672854
rect 455546 636938 455782 637174
rect 455866 636938 456102 637174
rect 455546 636618 455782 636854
rect 455866 636618 456102 636854
rect 455546 600938 455782 601174
rect 455866 600938 456102 601174
rect 455546 600618 455782 600854
rect 455866 600618 456102 600854
rect 455546 564938 455782 565174
rect 455866 564938 456102 565174
rect 455546 564618 455782 564854
rect 455866 564618 456102 564854
rect 455546 528938 455782 529174
rect 455866 528938 456102 529174
rect 455546 528618 455782 528854
rect 455866 528618 456102 528854
rect 455546 492938 455782 493174
rect 455866 492938 456102 493174
rect 455546 492618 455782 492854
rect 455866 492618 456102 492854
rect 455546 456938 455782 457174
rect 455866 456938 456102 457174
rect 455546 456618 455782 456854
rect 455866 456618 456102 456854
rect 455546 420938 455782 421174
rect 455866 420938 456102 421174
rect 455546 420618 455782 420854
rect 455866 420618 456102 420854
rect 455546 384938 455782 385174
rect 455866 384938 456102 385174
rect 455546 384618 455782 384854
rect 455866 384618 456102 384854
rect 455546 348938 455782 349174
rect 455866 348938 456102 349174
rect 455546 348618 455782 348854
rect 455866 348618 456102 348854
rect 455546 312938 455782 313174
rect 455866 312938 456102 313174
rect 455546 312618 455782 312854
rect 455866 312618 456102 312854
rect 455546 276938 455782 277174
rect 455866 276938 456102 277174
rect 455546 276618 455782 276854
rect 455866 276618 456102 276854
rect 455546 240938 455782 241174
rect 455866 240938 456102 241174
rect 455546 240618 455782 240854
rect 455866 240618 456102 240854
rect 455546 204938 455782 205174
rect 455866 204938 456102 205174
rect 455546 204618 455782 204854
rect 455866 204618 456102 204854
rect 455546 168938 455782 169174
rect 455866 168938 456102 169174
rect 455546 168618 455782 168854
rect 455866 168618 456102 168854
rect 455546 132938 455782 133174
rect 455866 132938 456102 133174
rect 455546 132618 455782 132854
rect 455866 132618 456102 132854
rect 455546 96938 455782 97174
rect 455866 96938 456102 97174
rect 455546 96618 455782 96854
rect 455866 96618 456102 96854
rect 455546 60938 455782 61174
rect 455866 60938 456102 61174
rect 455546 60618 455782 60854
rect 455866 60618 456102 60854
rect 455546 24938 455782 25174
rect 455866 24938 456102 25174
rect 455546 24618 455782 24854
rect 455866 24618 456102 24854
rect 455546 -3462 455782 -3226
rect 455866 -3462 456102 -3226
rect 455546 -3782 455782 -3546
rect 455866 -3782 456102 -3546
rect 459266 676658 459502 676894
rect 459586 676658 459822 676894
rect 459266 676338 459502 676574
rect 459586 676338 459822 676574
rect 459266 640658 459502 640894
rect 459586 640658 459822 640894
rect 459266 640338 459502 640574
rect 459586 640338 459822 640574
rect 459266 604658 459502 604894
rect 459586 604658 459822 604894
rect 459266 604338 459502 604574
rect 459586 604338 459822 604574
rect 459266 568658 459502 568894
rect 459586 568658 459822 568894
rect 459266 568338 459502 568574
rect 459586 568338 459822 568574
rect 459266 532658 459502 532894
rect 459586 532658 459822 532894
rect 459266 532338 459502 532574
rect 459586 532338 459822 532574
rect 459266 496658 459502 496894
rect 459586 496658 459822 496894
rect 459266 496338 459502 496574
rect 459586 496338 459822 496574
rect 459266 460658 459502 460894
rect 459586 460658 459822 460894
rect 459266 460338 459502 460574
rect 459586 460338 459822 460574
rect 459266 424658 459502 424894
rect 459586 424658 459822 424894
rect 459266 424338 459502 424574
rect 459586 424338 459822 424574
rect 459266 388658 459502 388894
rect 459586 388658 459822 388894
rect 459266 388338 459502 388574
rect 459586 388338 459822 388574
rect 459266 352658 459502 352894
rect 459586 352658 459822 352894
rect 459266 352338 459502 352574
rect 459586 352338 459822 352574
rect 459266 316658 459502 316894
rect 459586 316658 459822 316894
rect 459266 316338 459502 316574
rect 459586 316338 459822 316574
rect 459266 280658 459502 280894
rect 459586 280658 459822 280894
rect 459266 280338 459502 280574
rect 459586 280338 459822 280574
rect 459266 244658 459502 244894
rect 459586 244658 459822 244894
rect 459266 244338 459502 244574
rect 459586 244338 459822 244574
rect 459266 208658 459502 208894
rect 459586 208658 459822 208894
rect 459266 208338 459502 208574
rect 459586 208338 459822 208574
rect 459266 172658 459502 172894
rect 459586 172658 459822 172894
rect 459266 172338 459502 172574
rect 459586 172338 459822 172574
rect 459266 136658 459502 136894
rect 459586 136658 459822 136894
rect 459266 136338 459502 136574
rect 459586 136338 459822 136574
rect 459266 100658 459502 100894
rect 459586 100658 459822 100894
rect 459266 100338 459502 100574
rect 459586 100338 459822 100574
rect 459266 64658 459502 64894
rect 459586 64658 459822 64894
rect 459266 64338 459502 64574
rect 459586 64338 459822 64574
rect 459266 28658 459502 28894
rect 459586 28658 459822 28894
rect 459266 28338 459502 28574
rect 459586 28338 459822 28574
rect 459266 -5382 459502 -5146
rect 459586 -5382 459822 -5146
rect 459266 -5702 459502 -5466
rect 459586 -5702 459822 -5466
rect 480986 710362 481222 710598
rect 481306 710362 481542 710598
rect 480986 710042 481222 710278
rect 481306 710042 481542 710278
rect 477266 708442 477502 708678
rect 477586 708442 477822 708678
rect 477266 708122 477502 708358
rect 477586 708122 477822 708358
rect 473546 706522 473782 706758
rect 473866 706522 474102 706758
rect 473546 706202 473782 706438
rect 473866 706202 474102 706438
rect 462986 680378 463222 680614
rect 463306 680378 463542 680614
rect 462986 680058 463222 680294
rect 463306 680058 463542 680294
rect 462986 644378 463222 644614
rect 463306 644378 463542 644614
rect 462986 644058 463222 644294
rect 463306 644058 463542 644294
rect 462986 608378 463222 608614
rect 463306 608378 463542 608614
rect 462986 608058 463222 608294
rect 463306 608058 463542 608294
rect 462986 572378 463222 572614
rect 463306 572378 463542 572614
rect 462986 572058 463222 572294
rect 463306 572058 463542 572294
rect 462986 536378 463222 536614
rect 463306 536378 463542 536614
rect 462986 536058 463222 536294
rect 463306 536058 463542 536294
rect 462986 500378 463222 500614
rect 463306 500378 463542 500614
rect 462986 500058 463222 500294
rect 463306 500058 463542 500294
rect 462986 464378 463222 464614
rect 463306 464378 463542 464614
rect 462986 464058 463222 464294
rect 463306 464058 463542 464294
rect 462986 428378 463222 428614
rect 463306 428378 463542 428614
rect 462986 428058 463222 428294
rect 463306 428058 463542 428294
rect 462986 392378 463222 392614
rect 463306 392378 463542 392614
rect 462986 392058 463222 392294
rect 463306 392058 463542 392294
rect 462986 356378 463222 356614
rect 463306 356378 463542 356614
rect 462986 356058 463222 356294
rect 463306 356058 463542 356294
rect 462986 320378 463222 320614
rect 463306 320378 463542 320614
rect 462986 320058 463222 320294
rect 463306 320058 463542 320294
rect 462986 284378 463222 284614
rect 463306 284378 463542 284614
rect 462986 284058 463222 284294
rect 463306 284058 463542 284294
rect 462986 248378 463222 248614
rect 463306 248378 463542 248614
rect 462986 248058 463222 248294
rect 463306 248058 463542 248294
rect 462986 212378 463222 212614
rect 463306 212378 463542 212614
rect 462986 212058 463222 212294
rect 463306 212058 463542 212294
rect 462986 176378 463222 176614
rect 463306 176378 463542 176614
rect 462986 176058 463222 176294
rect 463306 176058 463542 176294
rect 462986 140378 463222 140614
rect 463306 140378 463542 140614
rect 462986 140058 463222 140294
rect 463306 140058 463542 140294
rect 462986 104378 463222 104614
rect 463306 104378 463542 104614
rect 462986 104058 463222 104294
rect 463306 104058 463542 104294
rect 462986 68378 463222 68614
rect 463306 68378 463542 68614
rect 462986 68058 463222 68294
rect 463306 68058 463542 68294
rect 462986 32378 463222 32614
rect 463306 32378 463542 32614
rect 462986 32058 463222 32294
rect 463306 32058 463542 32294
rect 444986 -6342 445222 -6106
rect 445306 -6342 445542 -6106
rect 444986 -6662 445222 -6426
rect 445306 -6662 445542 -6426
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 690938 473782 691174
rect 473866 690938 474102 691174
rect 473546 690618 473782 690854
rect 473866 690618 474102 690854
rect 473546 654938 473782 655174
rect 473866 654938 474102 655174
rect 473546 654618 473782 654854
rect 473866 654618 474102 654854
rect 473546 618938 473782 619174
rect 473866 618938 474102 619174
rect 473546 618618 473782 618854
rect 473866 618618 474102 618854
rect 473546 582938 473782 583174
rect 473866 582938 474102 583174
rect 473546 582618 473782 582854
rect 473866 582618 474102 582854
rect 473546 546938 473782 547174
rect 473866 546938 474102 547174
rect 473546 546618 473782 546854
rect 473866 546618 474102 546854
rect 473546 510938 473782 511174
rect 473866 510938 474102 511174
rect 473546 510618 473782 510854
rect 473866 510618 474102 510854
rect 473546 474938 473782 475174
rect 473866 474938 474102 475174
rect 473546 474618 473782 474854
rect 473866 474618 474102 474854
rect 473546 438938 473782 439174
rect 473866 438938 474102 439174
rect 473546 438618 473782 438854
rect 473866 438618 474102 438854
rect 473546 402938 473782 403174
rect 473866 402938 474102 403174
rect 473546 402618 473782 402854
rect 473866 402618 474102 402854
rect 473546 366938 473782 367174
rect 473866 366938 474102 367174
rect 473546 366618 473782 366854
rect 473866 366618 474102 366854
rect 473546 330938 473782 331174
rect 473866 330938 474102 331174
rect 473546 330618 473782 330854
rect 473866 330618 474102 330854
rect 473546 294938 473782 295174
rect 473866 294938 474102 295174
rect 473546 294618 473782 294854
rect 473866 294618 474102 294854
rect 473546 258938 473782 259174
rect 473866 258938 474102 259174
rect 473546 258618 473782 258854
rect 473866 258618 474102 258854
rect 473546 222938 473782 223174
rect 473866 222938 474102 223174
rect 473546 222618 473782 222854
rect 473866 222618 474102 222854
rect 473546 186938 473782 187174
rect 473866 186938 474102 187174
rect 473546 186618 473782 186854
rect 473866 186618 474102 186854
rect 473546 150938 473782 151174
rect 473866 150938 474102 151174
rect 473546 150618 473782 150854
rect 473866 150618 474102 150854
rect 473546 114938 473782 115174
rect 473866 114938 474102 115174
rect 473546 114618 473782 114854
rect 473866 114618 474102 114854
rect 473546 78938 473782 79174
rect 473866 78938 474102 79174
rect 473546 78618 473782 78854
rect 473866 78618 474102 78854
rect 473546 42938 473782 43174
rect 473866 42938 474102 43174
rect 473546 42618 473782 42854
rect 473866 42618 474102 42854
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -2502 473782 -2266
rect 473866 -2502 474102 -2266
rect 473546 -2822 473782 -2586
rect 473866 -2822 474102 -2586
rect 477266 694658 477502 694894
rect 477586 694658 477822 694894
rect 477266 694338 477502 694574
rect 477586 694338 477822 694574
rect 477266 658658 477502 658894
rect 477586 658658 477822 658894
rect 477266 658338 477502 658574
rect 477586 658338 477822 658574
rect 477266 622658 477502 622894
rect 477586 622658 477822 622894
rect 477266 622338 477502 622574
rect 477586 622338 477822 622574
rect 477266 586658 477502 586894
rect 477586 586658 477822 586894
rect 477266 586338 477502 586574
rect 477586 586338 477822 586574
rect 477266 550658 477502 550894
rect 477586 550658 477822 550894
rect 477266 550338 477502 550574
rect 477586 550338 477822 550574
rect 477266 514658 477502 514894
rect 477586 514658 477822 514894
rect 477266 514338 477502 514574
rect 477586 514338 477822 514574
rect 477266 478658 477502 478894
rect 477586 478658 477822 478894
rect 477266 478338 477502 478574
rect 477586 478338 477822 478574
rect 477266 442658 477502 442894
rect 477586 442658 477822 442894
rect 477266 442338 477502 442574
rect 477586 442338 477822 442574
rect 477266 406658 477502 406894
rect 477586 406658 477822 406894
rect 477266 406338 477502 406574
rect 477586 406338 477822 406574
rect 477266 370658 477502 370894
rect 477586 370658 477822 370894
rect 477266 370338 477502 370574
rect 477586 370338 477822 370574
rect 477266 334658 477502 334894
rect 477586 334658 477822 334894
rect 477266 334338 477502 334574
rect 477586 334338 477822 334574
rect 477266 298658 477502 298894
rect 477586 298658 477822 298894
rect 477266 298338 477502 298574
rect 477586 298338 477822 298574
rect 477266 262658 477502 262894
rect 477586 262658 477822 262894
rect 477266 262338 477502 262574
rect 477586 262338 477822 262574
rect 477266 226658 477502 226894
rect 477586 226658 477822 226894
rect 477266 226338 477502 226574
rect 477586 226338 477822 226574
rect 477266 190658 477502 190894
rect 477586 190658 477822 190894
rect 477266 190338 477502 190574
rect 477586 190338 477822 190574
rect 477266 154658 477502 154894
rect 477586 154658 477822 154894
rect 477266 154338 477502 154574
rect 477586 154338 477822 154574
rect 477266 118658 477502 118894
rect 477586 118658 477822 118894
rect 477266 118338 477502 118574
rect 477586 118338 477822 118574
rect 477266 82658 477502 82894
rect 477586 82658 477822 82894
rect 477266 82338 477502 82574
rect 477586 82338 477822 82574
rect 477266 46658 477502 46894
rect 477586 46658 477822 46894
rect 477266 46338 477502 46574
rect 477586 46338 477822 46574
rect 477266 10658 477502 10894
rect 477586 10658 477822 10894
rect 477266 10338 477502 10574
rect 477586 10338 477822 10574
rect 477266 -4422 477502 -4186
rect 477586 -4422 477822 -4186
rect 477266 -4742 477502 -4506
rect 477586 -4742 477822 -4506
rect 498986 711322 499222 711558
rect 499306 711322 499542 711558
rect 498986 711002 499222 711238
rect 499306 711002 499542 711238
rect 495266 709402 495502 709638
rect 495586 709402 495822 709638
rect 495266 709082 495502 709318
rect 495586 709082 495822 709318
rect 491546 707482 491782 707718
rect 491866 707482 492102 707718
rect 491546 707162 491782 707398
rect 491866 707162 492102 707398
rect 480986 698378 481222 698614
rect 481306 698378 481542 698614
rect 480986 698058 481222 698294
rect 481306 698058 481542 698294
rect 480986 662378 481222 662614
rect 481306 662378 481542 662614
rect 480986 662058 481222 662294
rect 481306 662058 481542 662294
rect 480986 626378 481222 626614
rect 481306 626378 481542 626614
rect 480986 626058 481222 626294
rect 481306 626058 481542 626294
rect 480986 590378 481222 590614
rect 481306 590378 481542 590614
rect 480986 590058 481222 590294
rect 481306 590058 481542 590294
rect 480986 554378 481222 554614
rect 481306 554378 481542 554614
rect 480986 554058 481222 554294
rect 481306 554058 481542 554294
rect 480986 518378 481222 518614
rect 481306 518378 481542 518614
rect 480986 518058 481222 518294
rect 481306 518058 481542 518294
rect 480986 482378 481222 482614
rect 481306 482378 481542 482614
rect 480986 482058 481222 482294
rect 481306 482058 481542 482294
rect 480986 446378 481222 446614
rect 481306 446378 481542 446614
rect 480986 446058 481222 446294
rect 481306 446058 481542 446294
rect 480986 410378 481222 410614
rect 481306 410378 481542 410614
rect 480986 410058 481222 410294
rect 481306 410058 481542 410294
rect 480986 374378 481222 374614
rect 481306 374378 481542 374614
rect 480986 374058 481222 374294
rect 481306 374058 481542 374294
rect 480986 338378 481222 338614
rect 481306 338378 481542 338614
rect 480986 338058 481222 338294
rect 481306 338058 481542 338294
rect 480986 302378 481222 302614
rect 481306 302378 481542 302614
rect 480986 302058 481222 302294
rect 481306 302058 481542 302294
rect 480986 266378 481222 266614
rect 481306 266378 481542 266614
rect 480986 266058 481222 266294
rect 481306 266058 481542 266294
rect 480986 230378 481222 230614
rect 481306 230378 481542 230614
rect 480986 230058 481222 230294
rect 481306 230058 481542 230294
rect 480986 194378 481222 194614
rect 481306 194378 481542 194614
rect 480986 194058 481222 194294
rect 481306 194058 481542 194294
rect 480986 158378 481222 158614
rect 481306 158378 481542 158614
rect 480986 158058 481222 158294
rect 481306 158058 481542 158294
rect 480986 122378 481222 122614
rect 481306 122378 481542 122614
rect 480986 122058 481222 122294
rect 481306 122058 481542 122294
rect 480986 86378 481222 86614
rect 481306 86378 481542 86614
rect 480986 86058 481222 86294
rect 481306 86058 481542 86294
rect 480986 50378 481222 50614
rect 481306 50378 481542 50614
rect 480986 50058 481222 50294
rect 481306 50058 481542 50294
rect 480986 14378 481222 14614
rect 481306 14378 481542 14614
rect 480986 14058 481222 14294
rect 481306 14058 481542 14294
rect 462986 -7302 463222 -7066
rect 463306 -7302 463542 -7066
rect 462986 -7622 463222 -7386
rect 463306 -7622 463542 -7386
rect 487826 705562 488062 705798
rect 488146 705562 488382 705798
rect 487826 705242 488062 705478
rect 488146 705242 488382 705478
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 487826 453218 488062 453454
rect 488146 453218 488382 453454
rect 487826 452898 488062 453134
rect 488146 452898 488382 453134
rect 487826 417218 488062 417454
rect 488146 417218 488382 417454
rect 487826 416898 488062 417134
rect 488146 416898 488382 417134
rect 487826 381218 488062 381454
rect 488146 381218 488382 381454
rect 487826 380898 488062 381134
rect 488146 380898 488382 381134
rect 487826 345218 488062 345454
rect 488146 345218 488382 345454
rect 487826 344898 488062 345134
rect 488146 344898 488382 345134
rect 487826 309218 488062 309454
rect 488146 309218 488382 309454
rect 487826 308898 488062 309134
rect 488146 308898 488382 309134
rect 487826 273218 488062 273454
rect 488146 273218 488382 273454
rect 487826 272898 488062 273134
rect 488146 272898 488382 273134
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 487826 129218 488062 129454
rect 488146 129218 488382 129454
rect 487826 128898 488062 129134
rect 488146 128898 488382 129134
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -1542 488062 -1306
rect 488146 -1542 488382 -1306
rect 487826 -1862 488062 -1626
rect 488146 -1862 488382 -1626
rect 491546 672938 491782 673174
rect 491866 672938 492102 673174
rect 491546 672618 491782 672854
rect 491866 672618 492102 672854
rect 491546 636938 491782 637174
rect 491866 636938 492102 637174
rect 491546 636618 491782 636854
rect 491866 636618 492102 636854
rect 491546 600938 491782 601174
rect 491866 600938 492102 601174
rect 491546 600618 491782 600854
rect 491866 600618 492102 600854
rect 491546 564938 491782 565174
rect 491866 564938 492102 565174
rect 491546 564618 491782 564854
rect 491866 564618 492102 564854
rect 491546 528938 491782 529174
rect 491866 528938 492102 529174
rect 491546 528618 491782 528854
rect 491866 528618 492102 528854
rect 491546 492938 491782 493174
rect 491866 492938 492102 493174
rect 491546 492618 491782 492854
rect 491866 492618 492102 492854
rect 491546 456938 491782 457174
rect 491866 456938 492102 457174
rect 491546 456618 491782 456854
rect 491866 456618 492102 456854
rect 491546 420938 491782 421174
rect 491866 420938 492102 421174
rect 491546 420618 491782 420854
rect 491866 420618 492102 420854
rect 491546 384938 491782 385174
rect 491866 384938 492102 385174
rect 491546 384618 491782 384854
rect 491866 384618 492102 384854
rect 491546 348938 491782 349174
rect 491866 348938 492102 349174
rect 491546 348618 491782 348854
rect 491866 348618 492102 348854
rect 491546 312938 491782 313174
rect 491866 312938 492102 313174
rect 491546 312618 491782 312854
rect 491866 312618 492102 312854
rect 491546 276938 491782 277174
rect 491866 276938 492102 277174
rect 491546 276618 491782 276854
rect 491866 276618 492102 276854
rect 491546 240938 491782 241174
rect 491866 240938 492102 241174
rect 491546 240618 491782 240854
rect 491866 240618 492102 240854
rect 491546 204938 491782 205174
rect 491866 204938 492102 205174
rect 491546 204618 491782 204854
rect 491866 204618 492102 204854
rect 491546 168938 491782 169174
rect 491866 168938 492102 169174
rect 491546 168618 491782 168854
rect 491866 168618 492102 168854
rect 491546 132938 491782 133174
rect 491866 132938 492102 133174
rect 491546 132618 491782 132854
rect 491866 132618 492102 132854
rect 491546 96938 491782 97174
rect 491866 96938 492102 97174
rect 491546 96618 491782 96854
rect 491866 96618 492102 96854
rect 491546 60938 491782 61174
rect 491866 60938 492102 61174
rect 491546 60618 491782 60854
rect 491866 60618 492102 60854
rect 491546 24938 491782 25174
rect 491866 24938 492102 25174
rect 491546 24618 491782 24854
rect 491866 24618 492102 24854
rect 491546 -3462 491782 -3226
rect 491866 -3462 492102 -3226
rect 491546 -3782 491782 -3546
rect 491866 -3782 492102 -3546
rect 495266 676658 495502 676894
rect 495586 676658 495822 676894
rect 495266 676338 495502 676574
rect 495586 676338 495822 676574
rect 495266 640658 495502 640894
rect 495586 640658 495822 640894
rect 495266 640338 495502 640574
rect 495586 640338 495822 640574
rect 495266 604658 495502 604894
rect 495586 604658 495822 604894
rect 495266 604338 495502 604574
rect 495586 604338 495822 604574
rect 495266 568658 495502 568894
rect 495586 568658 495822 568894
rect 495266 568338 495502 568574
rect 495586 568338 495822 568574
rect 495266 532658 495502 532894
rect 495586 532658 495822 532894
rect 495266 532338 495502 532574
rect 495586 532338 495822 532574
rect 495266 496658 495502 496894
rect 495586 496658 495822 496894
rect 495266 496338 495502 496574
rect 495586 496338 495822 496574
rect 495266 460658 495502 460894
rect 495586 460658 495822 460894
rect 495266 460338 495502 460574
rect 495586 460338 495822 460574
rect 495266 424658 495502 424894
rect 495586 424658 495822 424894
rect 495266 424338 495502 424574
rect 495586 424338 495822 424574
rect 495266 388658 495502 388894
rect 495586 388658 495822 388894
rect 495266 388338 495502 388574
rect 495586 388338 495822 388574
rect 495266 352658 495502 352894
rect 495586 352658 495822 352894
rect 495266 352338 495502 352574
rect 495586 352338 495822 352574
rect 495266 316658 495502 316894
rect 495586 316658 495822 316894
rect 495266 316338 495502 316574
rect 495586 316338 495822 316574
rect 495266 280658 495502 280894
rect 495586 280658 495822 280894
rect 495266 280338 495502 280574
rect 495586 280338 495822 280574
rect 495266 244658 495502 244894
rect 495586 244658 495822 244894
rect 495266 244338 495502 244574
rect 495586 244338 495822 244574
rect 495266 208658 495502 208894
rect 495586 208658 495822 208894
rect 495266 208338 495502 208574
rect 495586 208338 495822 208574
rect 495266 172658 495502 172894
rect 495586 172658 495822 172894
rect 495266 172338 495502 172574
rect 495586 172338 495822 172574
rect 495266 136658 495502 136894
rect 495586 136658 495822 136894
rect 495266 136338 495502 136574
rect 495586 136338 495822 136574
rect 495266 100658 495502 100894
rect 495586 100658 495822 100894
rect 495266 100338 495502 100574
rect 495586 100338 495822 100574
rect 495266 64658 495502 64894
rect 495586 64658 495822 64894
rect 495266 64338 495502 64574
rect 495586 64338 495822 64574
rect 495266 28658 495502 28894
rect 495586 28658 495822 28894
rect 495266 28338 495502 28574
rect 495586 28338 495822 28574
rect 495266 -5382 495502 -5146
rect 495586 -5382 495822 -5146
rect 495266 -5702 495502 -5466
rect 495586 -5702 495822 -5466
rect 516986 710362 517222 710598
rect 517306 710362 517542 710598
rect 516986 710042 517222 710278
rect 517306 710042 517542 710278
rect 513266 708442 513502 708678
rect 513586 708442 513822 708678
rect 513266 708122 513502 708358
rect 513586 708122 513822 708358
rect 509546 706522 509782 706758
rect 509866 706522 510102 706758
rect 509546 706202 509782 706438
rect 509866 706202 510102 706438
rect 498986 680378 499222 680614
rect 499306 680378 499542 680614
rect 498986 680058 499222 680294
rect 499306 680058 499542 680294
rect 498986 644378 499222 644614
rect 499306 644378 499542 644614
rect 498986 644058 499222 644294
rect 499306 644058 499542 644294
rect 498986 608378 499222 608614
rect 499306 608378 499542 608614
rect 498986 608058 499222 608294
rect 499306 608058 499542 608294
rect 498986 572378 499222 572614
rect 499306 572378 499542 572614
rect 498986 572058 499222 572294
rect 499306 572058 499542 572294
rect 498986 536378 499222 536614
rect 499306 536378 499542 536614
rect 498986 536058 499222 536294
rect 499306 536058 499542 536294
rect 498986 500378 499222 500614
rect 499306 500378 499542 500614
rect 498986 500058 499222 500294
rect 499306 500058 499542 500294
rect 498986 464378 499222 464614
rect 499306 464378 499542 464614
rect 498986 464058 499222 464294
rect 499306 464058 499542 464294
rect 498986 428378 499222 428614
rect 499306 428378 499542 428614
rect 498986 428058 499222 428294
rect 499306 428058 499542 428294
rect 498986 392378 499222 392614
rect 499306 392378 499542 392614
rect 498986 392058 499222 392294
rect 499306 392058 499542 392294
rect 498986 356378 499222 356614
rect 499306 356378 499542 356614
rect 498986 356058 499222 356294
rect 499306 356058 499542 356294
rect 498986 320378 499222 320614
rect 499306 320378 499542 320614
rect 498986 320058 499222 320294
rect 499306 320058 499542 320294
rect 498986 284378 499222 284614
rect 499306 284378 499542 284614
rect 498986 284058 499222 284294
rect 499306 284058 499542 284294
rect 498986 248378 499222 248614
rect 499306 248378 499542 248614
rect 498986 248058 499222 248294
rect 499306 248058 499542 248294
rect 498986 212378 499222 212614
rect 499306 212378 499542 212614
rect 498986 212058 499222 212294
rect 499306 212058 499542 212294
rect 498986 176378 499222 176614
rect 499306 176378 499542 176614
rect 498986 176058 499222 176294
rect 499306 176058 499542 176294
rect 498986 140378 499222 140614
rect 499306 140378 499542 140614
rect 498986 140058 499222 140294
rect 499306 140058 499542 140294
rect 498986 104378 499222 104614
rect 499306 104378 499542 104614
rect 498986 104058 499222 104294
rect 499306 104058 499542 104294
rect 498986 68378 499222 68614
rect 499306 68378 499542 68614
rect 498986 68058 499222 68294
rect 499306 68058 499542 68294
rect 498986 32378 499222 32614
rect 499306 32378 499542 32614
rect 498986 32058 499222 32294
rect 499306 32058 499542 32294
rect 480986 -6342 481222 -6106
rect 481306 -6342 481542 -6106
rect 480986 -6662 481222 -6426
rect 481306 -6662 481542 -6426
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 690938 509782 691174
rect 509866 690938 510102 691174
rect 509546 690618 509782 690854
rect 509866 690618 510102 690854
rect 509546 654938 509782 655174
rect 509866 654938 510102 655174
rect 509546 654618 509782 654854
rect 509866 654618 510102 654854
rect 509546 618938 509782 619174
rect 509866 618938 510102 619174
rect 509546 618618 509782 618854
rect 509866 618618 510102 618854
rect 509546 582938 509782 583174
rect 509866 582938 510102 583174
rect 509546 582618 509782 582854
rect 509866 582618 510102 582854
rect 509546 546938 509782 547174
rect 509866 546938 510102 547174
rect 509546 546618 509782 546854
rect 509866 546618 510102 546854
rect 509546 510938 509782 511174
rect 509866 510938 510102 511174
rect 509546 510618 509782 510854
rect 509866 510618 510102 510854
rect 509546 474938 509782 475174
rect 509866 474938 510102 475174
rect 509546 474618 509782 474854
rect 509866 474618 510102 474854
rect 509546 438938 509782 439174
rect 509866 438938 510102 439174
rect 509546 438618 509782 438854
rect 509866 438618 510102 438854
rect 509546 402938 509782 403174
rect 509866 402938 510102 403174
rect 509546 402618 509782 402854
rect 509866 402618 510102 402854
rect 509546 366938 509782 367174
rect 509866 366938 510102 367174
rect 509546 366618 509782 366854
rect 509866 366618 510102 366854
rect 509546 330938 509782 331174
rect 509866 330938 510102 331174
rect 509546 330618 509782 330854
rect 509866 330618 510102 330854
rect 509546 294938 509782 295174
rect 509866 294938 510102 295174
rect 509546 294618 509782 294854
rect 509866 294618 510102 294854
rect 509546 258938 509782 259174
rect 509866 258938 510102 259174
rect 509546 258618 509782 258854
rect 509866 258618 510102 258854
rect 509546 222938 509782 223174
rect 509866 222938 510102 223174
rect 509546 222618 509782 222854
rect 509866 222618 510102 222854
rect 509546 186938 509782 187174
rect 509866 186938 510102 187174
rect 509546 186618 509782 186854
rect 509866 186618 510102 186854
rect 509546 150938 509782 151174
rect 509866 150938 510102 151174
rect 509546 150618 509782 150854
rect 509866 150618 510102 150854
rect 509546 114938 509782 115174
rect 509866 114938 510102 115174
rect 509546 114618 509782 114854
rect 509866 114618 510102 114854
rect 509546 78938 509782 79174
rect 509866 78938 510102 79174
rect 509546 78618 509782 78854
rect 509866 78618 510102 78854
rect 509546 42938 509782 43174
rect 509866 42938 510102 43174
rect 509546 42618 509782 42854
rect 509866 42618 510102 42854
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -2502 509782 -2266
rect 509866 -2502 510102 -2266
rect 509546 -2822 509782 -2586
rect 509866 -2822 510102 -2586
rect 513266 694658 513502 694894
rect 513586 694658 513822 694894
rect 513266 694338 513502 694574
rect 513586 694338 513822 694574
rect 513266 658658 513502 658894
rect 513586 658658 513822 658894
rect 513266 658338 513502 658574
rect 513586 658338 513822 658574
rect 513266 622658 513502 622894
rect 513586 622658 513822 622894
rect 513266 622338 513502 622574
rect 513586 622338 513822 622574
rect 513266 586658 513502 586894
rect 513586 586658 513822 586894
rect 513266 586338 513502 586574
rect 513586 586338 513822 586574
rect 513266 550658 513502 550894
rect 513586 550658 513822 550894
rect 513266 550338 513502 550574
rect 513586 550338 513822 550574
rect 513266 514658 513502 514894
rect 513586 514658 513822 514894
rect 513266 514338 513502 514574
rect 513586 514338 513822 514574
rect 513266 478658 513502 478894
rect 513586 478658 513822 478894
rect 513266 478338 513502 478574
rect 513586 478338 513822 478574
rect 513266 442658 513502 442894
rect 513586 442658 513822 442894
rect 513266 442338 513502 442574
rect 513586 442338 513822 442574
rect 513266 406658 513502 406894
rect 513586 406658 513822 406894
rect 513266 406338 513502 406574
rect 513586 406338 513822 406574
rect 513266 370658 513502 370894
rect 513586 370658 513822 370894
rect 513266 370338 513502 370574
rect 513586 370338 513822 370574
rect 513266 334658 513502 334894
rect 513586 334658 513822 334894
rect 513266 334338 513502 334574
rect 513586 334338 513822 334574
rect 513266 298658 513502 298894
rect 513586 298658 513822 298894
rect 513266 298338 513502 298574
rect 513586 298338 513822 298574
rect 513266 262658 513502 262894
rect 513586 262658 513822 262894
rect 513266 262338 513502 262574
rect 513586 262338 513822 262574
rect 513266 226658 513502 226894
rect 513586 226658 513822 226894
rect 513266 226338 513502 226574
rect 513586 226338 513822 226574
rect 513266 190658 513502 190894
rect 513586 190658 513822 190894
rect 513266 190338 513502 190574
rect 513586 190338 513822 190574
rect 513266 154658 513502 154894
rect 513586 154658 513822 154894
rect 513266 154338 513502 154574
rect 513586 154338 513822 154574
rect 513266 118658 513502 118894
rect 513586 118658 513822 118894
rect 513266 118338 513502 118574
rect 513586 118338 513822 118574
rect 513266 82658 513502 82894
rect 513586 82658 513822 82894
rect 513266 82338 513502 82574
rect 513586 82338 513822 82574
rect 513266 46658 513502 46894
rect 513586 46658 513822 46894
rect 513266 46338 513502 46574
rect 513586 46338 513822 46574
rect 513266 10658 513502 10894
rect 513586 10658 513822 10894
rect 513266 10338 513502 10574
rect 513586 10338 513822 10574
rect 513266 -4422 513502 -4186
rect 513586 -4422 513822 -4186
rect 513266 -4742 513502 -4506
rect 513586 -4742 513822 -4506
rect 534986 711322 535222 711558
rect 535306 711322 535542 711558
rect 534986 711002 535222 711238
rect 535306 711002 535542 711238
rect 531266 709402 531502 709638
rect 531586 709402 531822 709638
rect 531266 709082 531502 709318
rect 531586 709082 531822 709318
rect 527546 707482 527782 707718
rect 527866 707482 528102 707718
rect 527546 707162 527782 707398
rect 527866 707162 528102 707398
rect 516986 698378 517222 698614
rect 517306 698378 517542 698614
rect 516986 698058 517222 698294
rect 517306 698058 517542 698294
rect 516986 662378 517222 662614
rect 517306 662378 517542 662614
rect 516986 662058 517222 662294
rect 517306 662058 517542 662294
rect 516986 626378 517222 626614
rect 517306 626378 517542 626614
rect 516986 626058 517222 626294
rect 517306 626058 517542 626294
rect 516986 590378 517222 590614
rect 517306 590378 517542 590614
rect 516986 590058 517222 590294
rect 517306 590058 517542 590294
rect 516986 554378 517222 554614
rect 517306 554378 517542 554614
rect 516986 554058 517222 554294
rect 517306 554058 517542 554294
rect 516986 518378 517222 518614
rect 517306 518378 517542 518614
rect 516986 518058 517222 518294
rect 517306 518058 517542 518294
rect 516986 482378 517222 482614
rect 517306 482378 517542 482614
rect 516986 482058 517222 482294
rect 517306 482058 517542 482294
rect 516986 446378 517222 446614
rect 517306 446378 517542 446614
rect 516986 446058 517222 446294
rect 517306 446058 517542 446294
rect 516986 410378 517222 410614
rect 517306 410378 517542 410614
rect 516986 410058 517222 410294
rect 517306 410058 517542 410294
rect 516986 374378 517222 374614
rect 517306 374378 517542 374614
rect 516986 374058 517222 374294
rect 517306 374058 517542 374294
rect 516986 338378 517222 338614
rect 517306 338378 517542 338614
rect 516986 338058 517222 338294
rect 517306 338058 517542 338294
rect 516986 302378 517222 302614
rect 517306 302378 517542 302614
rect 516986 302058 517222 302294
rect 517306 302058 517542 302294
rect 516986 266378 517222 266614
rect 517306 266378 517542 266614
rect 516986 266058 517222 266294
rect 517306 266058 517542 266294
rect 516986 230378 517222 230614
rect 517306 230378 517542 230614
rect 516986 230058 517222 230294
rect 517306 230058 517542 230294
rect 516986 194378 517222 194614
rect 517306 194378 517542 194614
rect 516986 194058 517222 194294
rect 517306 194058 517542 194294
rect 516986 158378 517222 158614
rect 517306 158378 517542 158614
rect 516986 158058 517222 158294
rect 517306 158058 517542 158294
rect 516986 122378 517222 122614
rect 517306 122378 517542 122614
rect 516986 122058 517222 122294
rect 517306 122058 517542 122294
rect 516986 86378 517222 86614
rect 517306 86378 517542 86614
rect 516986 86058 517222 86294
rect 517306 86058 517542 86294
rect 516986 50378 517222 50614
rect 517306 50378 517542 50614
rect 516986 50058 517222 50294
rect 517306 50058 517542 50294
rect 516986 14378 517222 14614
rect 517306 14378 517542 14614
rect 516986 14058 517222 14294
rect 517306 14058 517542 14294
rect 498986 -7302 499222 -7066
rect 499306 -7302 499542 -7066
rect 498986 -7622 499222 -7386
rect 499306 -7622 499542 -7386
rect 523826 705562 524062 705798
rect 524146 705562 524382 705798
rect 523826 705242 524062 705478
rect 524146 705242 524382 705478
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -1542 524062 -1306
rect 524146 -1542 524382 -1306
rect 523826 -1862 524062 -1626
rect 524146 -1862 524382 -1626
rect 527546 672938 527782 673174
rect 527866 672938 528102 673174
rect 527546 672618 527782 672854
rect 527866 672618 528102 672854
rect 527546 636938 527782 637174
rect 527866 636938 528102 637174
rect 527546 636618 527782 636854
rect 527866 636618 528102 636854
rect 527546 600938 527782 601174
rect 527866 600938 528102 601174
rect 527546 600618 527782 600854
rect 527866 600618 528102 600854
rect 527546 564938 527782 565174
rect 527866 564938 528102 565174
rect 527546 564618 527782 564854
rect 527866 564618 528102 564854
rect 527546 528938 527782 529174
rect 527866 528938 528102 529174
rect 527546 528618 527782 528854
rect 527866 528618 528102 528854
rect 527546 492938 527782 493174
rect 527866 492938 528102 493174
rect 527546 492618 527782 492854
rect 527866 492618 528102 492854
rect 527546 456938 527782 457174
rect 527866 456938 528102 457174
rect 527546 456618 527782 456854
rect 527866 456618 528102 456854
rect 527546 420938 527782 421174
rect 527866 420938 528102 421174
rect 527546 420618 527782 420854
rect 527866 420618 528102 420854
rect 527546 384938 527782 385174
rect 527866 384938 528102 385174
rect 527546 384618 527782 384854
rect 527866 384618 528102 384854
rect 527546 348938 527782 349174
rect 527866 348938 528102 349174
rect 527546 348618 527782 348854
rect 527866 348618 528102 348854
rect 527546 312938 527782 313174
rect 527866 312938 528102 313174
rect 527546 312618 527782 312854
rect 527866 312618 528102 312854
rect 527546 276938 527782 277174
rect 527866 276938 528102 277174
rect 527546 276618 527782 276854
rect 527866 276618 528102 276854
rect 527546 240938 527782 241174
rect 527866 240938 528102 241174
rect 527546 240618 527782 240854
rect 527866 240618 528102 240854
rect 527546 204938 527782 205174
rect 527866 204938 528102 205174
rect 527546 204618 527782 204854
rect 527866 204618 528102 204854
rect 527546 168938 527782 169174
rect 527866 168938 528102 169174
rect 527546 168618 527782 168854
rect 527866 168618 528102 168854
rect 527546 132938 527782 133174
rect 527866 132938 528102 133174
rect 527546 132618 527782 132854
rect 527866 132618 528102 132854
rect 527546 96938 527782 97174
rect 527866 96938 528102 97174
rect 527546 96618 527782 96854
rect 527866 96618 528102 96854
rect 527546 60938 527782 61174
rect 527866 60938 528102 61174
rect 527546 60618 527782 60854
rect 527866 60618 528102 60854
rect 527546 24938 527782 25174
rect 527866 24938 528102 25174
rect 527546 24618 527782 24854
rect 527866 24618 528102 24854
rect 527546 -3462 527782 -3226
rect 527866 -3462 528102 -3226
rect 527546 -3782 527782 -3546
rect 527866 -3782 528102 -3546
rect 531266 676658 531502 676894
rect 531586 676658 531822 676894
rect 531266 676338 531502 676574
rect 531586 676338 531822 676574
rect 531266 640658 531502 640894
rect 531586 640658 531822 640894
rect 531266 640338 531502 640574
rect 531586 640338 531822 640574
rect 531266 604658 531502 604894
rect 531586 604658 531822 604894
rect 531266 604338 531502 604574
rect 531586 604338 531822 604574
rect 531266 568658 531502 568894
rect 531586 568658 531822 568894
rect 531266 568338 531502 568574
rect 531586 568338 531822 568574
rect 531266 532658 531502 532894
rect 531586 532658 531822 532894
rect 531266 532338 531502 532574
rect 531586 532338 531822 532574
rect 531266 496658 531502 496894
rect 531586 496658 531822 496894
rect 531266 496338 531502 496574
rect 531586 496338 531822 496574
rect 531266 460658 531502 460894
rect 531586 460658 531822 460894
rect 531266 460338 531502 460574
rect 531586 460338 531822 460574
rect 531266 424658 531502 424894
rect 531586 424658 531822 424894
rect 531266 424338 531502 424574
rect 531586 424338 531822 424574
rect 531266 388658 531502 388894
rect 531586 388658 531822 388894
rect 531266 388338 531502 388574
rect 531586 388338 531822 388574
rect 531266 352658 531502 352894
rect 531586 352658 531822 352894
rect 531266 352338 531502 352574
rect 531586 352338 531822 352574
rect 531266 316658 531502 316894
rect 531586 316658 531822 316894
rect 531266 316338 531502 316574
rect 531586 316338 531822 316574
rect 531266 280658 531502 280894
rect 531586 280658 531822 280894
rect 531266 280338 531502 280574
rect 531586 280338 531822 280574
rect 531266 244658 531502 244894
rect 531586 244658 531822 244894
rect 531266 244338 531502 244574
rect 531586 244338 531822 244574
rect 531266 208658 531502 208894
rect 531586 208658 531822 208894
rect 531266 208338 531502 208574
rect 531586 208338 531822 208574
rect 531266 172658 531502 172894
rect 531586 172658 531822 172894
rect 531266 172338 531502 172574
rect 531586 172338 531822 172574
rect 531266 136658 531502 136894
rect 531586 136658 531822 136894
rect 531266 136338 531502 136574
rect 531586 136338 531822 136574
rect 531266 100658 531502 100894
rect 531586 100658 531822 100894
rect 531266 100338 531502 100574
rect 531586 100338 531822 100574
rect 531266 64658 531502 64894
rect 531586 64658 531822 64894
rect 531266 64338 531502 64574
rect 531586 64338 531822 64574
rect 531266 28658 531502 28894
rect 531586 28658 531822 28894
rect 531266 28338 531502 28574
rect 531586 28338 531822 28574
rect 531266 -5382 531502 -5146
rect 531586 -5382 531822 -5146
rect 531266 -5702 531502 -5466
rect 531586 -5702 531822 -5466
rect 552986 710362 553222 710598
rect 553306 710362 553542 710598
rect 552986 710042 553222 710278
rect 553306 710042 553542 710278
rect 549266 708442 549502 708678
rect 549586 708442 549822 708678
rect 549266 708122 549502 708358
rect 549586 708122 549822 708358
rect 545546 706522 545782 706758
rect 545866 706522 546102 706758
rect 545546 706202 545782 706438
rect 545866 706202 546102 706438
rect 534986 680378 535222 680614
rect 535306 680378 535542 680614
rect 534986 680058 535222 680294
rect 535306 680058 535542 680294
rect 534986 644378 535222 644614
rect 535306 644378 535542 644614
rect 534986 644058 535222 644294
rect 535306 644058 535542 644294
rect 534986 608378 535222 608614
rect 535306 608378 535542 608614
rect 534986 608058 535222 608294
rect 535306 608058 535542 608294
rect 534986 572378 535222 572614
rect 535306 572378 535542 572614
rect 534986 572058 535222 572294
rect 535306 572058 535542 572294
rect 534986 536378 535222 536614
rect 535306 536378 535542 536614
rect 534986 536058 535222 536294
rect 535306 536058 535542 536294
rect 534986 500378 535222 500614
rect 535306 500378 535542 500614
rect 534986 500058 535222 500294
rect 535306 500058 535542 500294
rect 534986 464378 535222 464614
rect 535306 464378 535542 464614
rect 534986 464058 535222 464294
rect 535306 464058 535542 464294
rect 534986 428378 535222 428614
rect 535306 428378 535542 428614
rect 534986 428058 535222 428294
rect 535306 428058 535542 428294
rect 534986 392378 535222 392614
rect 535306 392378 535542 392614
rect 534986 392058 535222 392294
rect 535306 392058 535542 392294
rect 534986 356378 535222 356614
rect 535306 356378 535542 356614
rect 534986 356058 535222 356294
rect 535306 356058 535542 356294
rect 534986 320378 535222 320614
rect 535306 320378 535542 320614
rect 534986 320058 535222 320294
rect 535306 320058 535542 320294
rect 534986 284378 535222 284614
rect 535306 284378 535542 284614
rect 534986 284058 535222 284294
rect 535306 284058 535542 284294
rect 534986 248378 535222 248614
rect 535306 248378 535542 248614
rect 534986 248058 535222 248294
rect 535306 248058 535542 248294
rect 534986 212378 535222 212614
rect 535306 212378 535542 212614
rect 534986 212058 535222 212294
rect 535306 212058 535542 212294
rect 534986 176378 535222 176614
rect 535306 176378 535542 176614
rect 534986 176058 535222 176294
rect 535306 176058 535542 176294
rect 534986 140378 535222 140614
rect 535306 140378 535542 140614
rect 534986 140058 535222 140294
rect 535306 140058 535542 140294
rect 534986 104378 535222 104614
rect 535306 104378 535542 104614
rect 534986 104058 535222 104294
rect 535306 104058 535542 104294
rect 534986 68378 535222 68614
rect 535306 68378 535542 68614
rect 534986 68058 535222 68294
rect 535306 68058 535542 68294
rect 534986 32378 535222 32614
rect 535306 32378 535542 32614
rect 534986 32058 535222 32294
rect 535306 32058 535542 32294
rect 516986 -6342 517222 -6106
rect 517306 -6342 517542 -6106
rect 516986 -6662 517222 -6426
rect 517306 -6662 517542 -6426
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 690938 545782 691174
rect 545866 690938 546102 691174
rect 545546 690618 545782 690854
rect 545866 690618 546102 690854
rect 545546 654938 545782 655174
rect 545866 654938 546102 655174
rect 545546 654618 545782 654854
rect 545866 654618 546102 654854
rect 545546 618938 545782 619174
rect 545866 618938 546102 619174
rect 545546 618618 545782 618854
rect 545866 618618 546102 618854
rect 545546 582938 545782 583174
rect 545866 582938 546102 583174
rect 545546 582618 545782 582854
rect 545866 582618 546102 582854
rect 545546 546938 545782 547174
rect 545866 546938 546102 547174
rect 545546 546618 545782 546854
rect 545866 546618 546102 546854
rect 545546 510938 545782 511174
rect 545866 510938 546102 511174
rect 545546 510618 545782 510854
rect 545866 510618 546102 510854
rect 545546 474938 545782 475174
rect 545866 474938 546102 475174
rect 545546 474618 545782 474854
rect 545866 474618 546102 474854
rect 545546 438938 545782 439174
rect 545866 438938 546102 439174
rect 545546 438618 545782 438854
rect 545866 438618 546102 438854
rect 545546 402938 545782 403174
rect 545866 402938 546102 403174
rect 545546 402618 545782 402854
rect 545866 402618 546102 402854
rect 545546 366938 545782 367174
rect 545866 366938 546102 367174
rect 545546 366618 545782 366854
rect 545866 366618 546102 366854
rect 545546 330938 545782 331174
rect 545866 330938 546102 331174
rect 545546 330618 545782 330854
rect 545866 330618 546102 330854
rect 545546 294938 545782 295174
rect 545866 294938 546102 295174
rect 545546 294618 545782 294854
rect 545866 294618 546102 294854
rect 545546 258938 545782 259174
rect 545866 258938 546102 259174
rect 545546 258618 545782 258854
rect 545866 258618 546102 258854
rect 545546 222938 545782 223174
rect 545866 222938 546102 223174
rect 545546 222618 545782 222854
rect 545866 222618 546102 222854
rect 545546 186938 545782 187174
rect 545866 186938 546102 187174
rect 545546 186618 545782 186854
rect 545866 186618 546102 186854
rect 545546 150938 545782 151174
rect 545866 150938 546102 151174
rect 545546 150618 545782 150854
rect 545866 150618 546102 150854
rect 545546 114938 545782 115174
rect 545866 114938 546102 115174
rect 545546 114618 545782 114854
rect 545866 114618 546102 114854
rect 545546 78938 545782 79174
rect 545866 78938 546102 79174
rect 545546 78618 545782 78854
rect 545866 78618 546102 78854
rect 545546 42938 545782 43174
rect 545866 42938 546102 43174
rect 545546 42618 545782 42854
rect 545866 42618 546102 42854
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -2502 545782 -2266
rect 545866 -2502 546102 -2266
rect 545546 -2822 545782 -2586
rect 545866 -2822 546102 -2586
rect 549266 694658 549502 694894
rect 549586 694658 549822 694894
rect 549266 694338 549502 694574
rect 549586 694338 549822 694574
rect 549266 658658 549502 658894
rect 549586 658658 549822 658894
rect 549266 658338 549502 658574
rect 549586 658338 549822 658574
rect 549266 622658 549502 622894
rect 549586 622658 549822 622894
rect 549266 622338 549502 622574
rect 549586 622338 549822 622574
rect 549266 586658 549502 586894
rect 549586 586658 549822 586894
rect 549266 586338 549502 586574
rect 549586 586338 549822 586574
rect 549266 550658 549502 550894
rect 549586 550658 549822 550894
rect 549266 550338 549502 550574
rect 549586 550338 549822 550574
rect 549266 514658 549502 514894
rect 549586 514658 549822 514894
rect 549266 514338 549502 514574
rect 549586 514338 549822 514574
rect 549266 478658 549502 478894
rect 549586 478658 549822 478894
rect 549266 478338 549502 478574
rect 549586 478338 549822 478574
rect 549266 442658 549502 442894
rect 549586 442658 549822 442894
rect 549266 442338 549502 442574
rect 549586 442338 549822 442574
rect 549266 406658 549502 406894
rect 549586 406658 549822 406894
rect 549266 406338 549502 406574
rect 549586 406338 549822 406574
rect 549266 370658 549502 370894
rect 549586 370658 549822 370894
rect 549266 370338 549502 370574
rect 549586 370338 549822 370574
rect 549266 334658 549502 334894
rect 549586 334658 549822 334894
rect 549266 334338 549502 334574
rect 549586 334338 549822 334574
rect 549266 298658 549502 298894
rect 549586 298658 549822 298894
rect 549266 298338 549502 298574
rect 549586 298338 549822 298574
rect 549266 262658 549502 262894
rect 549586 262658 549822 262894
rect 549266 262338 549502 262574
rect 549586 262338 549822 262574
rect 549266 226658 549502 226894
rect 549586 226658 549822 226894
rect 549266 226338 549502 226574
rect 549586 226338 549822 226574
rect 549266 190658 549502 190894
rect 549586 190658 549822 190894
rect 549266 190338 549502 190574
rect 549586 190338 549822 190574
rect 549266 154658 549502 154894
rect 549586 154658 549822 154894
rect 549266 154338 549502 154574
rect 549586 154338 549822 154574
rect 549266 118658 549502 118894
rect 549586 118658 549822 118894
rect 549266 118338 549502 118574
rect 549586 118338 549822 118574
rect 549266 82658 549502 82894
rect 549586 82658 549822 82894
rect 549266 82338 549502 82574
rect 549586 82338 549822 82574
rect 549266 46658 549502 46894
rect 549586 46658 549822 46894
rect 549266 46338 549502 46574
rect 549586 46338 549822 46574
rect 549266 10658 549502 10894
rect 549586 10658 549822 10894
rect 549266 10338 549502 10574
rect 549586 10338 549822 10574
rect 549266 -4422 549502 -4186
rect 549586 -4422 549822 -4186
rect 549266 -4742 549502 -4506
rect 549586 -4742 549822 -4506
rect 570986 711322 571222 711558
rect 571306 711322 571542 711558
rect 570986 711002 571222 711238
rect 571306 711002 571542 711238
rect 567266 709402 567502 709638
rect 567586 709402 567822 709638
rect 567266 709082 567502 709318
rect 567586 709082 567822 709318
rect 563546 707482 563782 707718
rect 563866 707482 564102 707718
rect 563546 707162 563782 707398
rect 563866 707162 564102 707398
rect 552986 698378 553222 698614
rect 553306 698378 553542 698614
rect 552986 698058 553222 698294
rect 553306 698058 553542 698294
rect 552986 662378 553222 662614
rect 553306 662378 553542 662614
rect 552986 662058 553222 662294
rect 553306 662058 553542 662294
rect 552986 626378 553222 626614
rect 553306 626378 553542 626614
rect 552986 626058 553222 626294
rect 553306 626058 553542 626294
rect 552986 590378 553222 590614
rect 553306 590378 553542 590614
rect 552986 590058 553222 590294
rect 553306 590058 553542 590294
rect 552986 554378 553222 554614
rect 553306 554378 553542 554614
rect 552986 554058 553222 554294
rect 553306 554058 553542 554294
rect 552986 518378 553222 518614
rect 553306 518378 553542 518614
rect 552986 518058 553222 518294
rect 553306 518058 553542 518294
rect 552986 482378 553222 482614
rect 553306 482378 553542 482614
rect 552986 482058 553222 482294
rect 553306 482058 553542 482294
rect 552986 446378 553222 446614
rect 553306 446378 553542 446614
rect 552986 446058 553222 446294
rect 553306 446058 553542 446294
rect 552986 410378 553222 410614
rect 553306 410378 553542 410614
rect 552986 410058 553222 410294
rect 553306 410058 553542 410294
rect 552986 374378 553222 374614
rect 553306 374378 553542 374614
rect 552986 374058 553222 374294
rect 553306 374058 553542 374294
rect 552986 338378 553222 338614
rect 553306 338378 553542 338614
rect 552986 338058 553222 338294
rect 553306 338058 553542 338294
rect 552986 302378 553222 302614
rect 553306 302378 553542 302614
rect 552986 302058 553222 302294
rect 553306 302058 553542 302294
rect 552986 266378 553222 266614
rect 553306 266378 553542 266614
rect 552986 266058 553222 266294
rect 553306 266058 553542 266294
rect 552986 230378 553222 230614
rect 553306 230378 553542 230614
rect 552986 230058 553222 230294
rect 553306 230058 553542 230294
rect 552986 194378 553222 194614
rect 553306 194378 553542 194614
rect 552986 194058 553222 194294
rect 553306 194058 553542 194294
rect 552986 158378 553222 158614
rect 553306 158378 553542 158614
rect 552986 158058 553222 158294
rect 553306 158058 553542 158294
rect 552986 122378 553222 122614
rect 553306 122378 553542 122614
rect 552986 122058 553222 122294
rect 553306 122058 553542 122294
rect 552986 86378 553222 86614
rect 553306 86378 553542 86614
rect 552986 86058 553222 86294
rect 553306 86058 553542 86294
rect 552986 50378 553222 50614
rect 553306 50378 553542 50614
rect 552986 50058 553222 50294
rect 553306 50058 553542 50294
rect 552986 14378 553222 14614
rect 553306 14378 553542 14614
rect 552986 14058 553222 14294
rect 553306 14058 553542 14294
rect 534986 -7302 535222 -7066
rect 535306 -7302 535542 -7066
rect 534986 -7622 535222 -7386
rect 535306 -7622 535542 -7386
rect 559826 705562 560062 705798
rect 560146 705562 560382 705798
rect 559826 705242 560062 705478
rect 560146 705242 560382 705478
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -1542 560062 -1306
rect 560146 -1542 560382 -1306
rect 559826 -1862 560062 -1626
rect 560146 -1862 560382 -1626
rect 563546 672938 563782 673174
rect 563866 672938 564102 673174
rect 563546 672618 563782 672854
rect 563866 672618 564102 672854
rect 563546 636938 563782 637174
rect 563866 636938 564102 637174
rect 563546 636618 563782 636854
rect 563866 636618 564102 636854
rect 563546 600938 563782 601174
rect 563866 600938 564102 601174
rect 563546 600618 563782 600854
rect 563866 600618 564102 600854
rect 563546 564938 563782 565174
rect 563866 564938 564102 565174
rect 563546 564618 563782 564854
rect 563866 564618 564102 564854
rect 563546 528938 563782 529174
rect 563866 528938 564102 529174
rect 563546 528618 563782 528854
rect 563866 528618 564102 528854
rect 563546 492938 563782 493174
rect 563866 492938 564102 493174
rect 563546 492618 563782 492854
rect 563866 492618 564102 492854
rect 563546 456938 563782 457174
rect 563866 456938 564102 457174
rect 563546 456618 563782 456854
rect 563866 456618 564102 456854
rect 563546 420938 563782 421174
rect 563866 420938 564102 421174
rect 563546 420618 563782 420854
rect 563866 420618 564102 420854
rect 563546 384938 563782 385174
rect 563866 384938 564102 385174
rect 563546 384618 563782 384854
rect 563866 384618 564102 384854
rect 563546 348938 563782 349174
rect 563866 348938 564102 349174
rect 563546 348618 563782 348854
rect 563866 348618 564102 348854
rect 563546 312938 563782 313174
rect 563866 312938 564102 313174
rect 563546 312618 563782 312854
rect 563866 312618 564102 312854
rect 563546 276938 563782 277174
rect 563866 276938 564102 277174
rect 563546 276618 563782 276854
rect 563866 276618 564102 276854
rect 563546 240938 563782 241174
rect 563866 240938 564102 241174
rect 563546 240618 563782 240854
rect 563866 240618 564102 240854
rect 563546 204938 563782 205174
rect 563866 204938 564102 205174
rect 563546 204618 563782 204854
rect 563866 204618 564102 204854
rect 563546 168938 563782 169174
rect 563866 168938 564102 169174
rect 563546 168618 563782 168854
rect 563866 168618 564102 168854
rect 563546 132938 563782 133174
rect 563866 132938 564102 133174
rect 563546 132618 563782 132854
rect 563866 132618 564102 132854
rect 563546 96938 563782 97174
rect 563866 96938 564102 97174
rect 563546 96618 563782 96854
rect 563866 96618 564102 96854
rect 563546 60938 563782 61174
rect 563866 60938 564102 61174
rect 563546 60618 563782 60854
rect 563866 60618 564102 60854
rect 563546 24938 563782 25174
rect 563866 24938 564102 25174
rect 563546 24618 563782 24854
rect 563866 24618 564102 24854
rect 563546 -3462 563782 -3226
rect 563866 -3462 564102 -3226
rect 563546 -3782 563782 -3546
rect 563866 -3782 564102 -3546
rect 567266 676658 567502 676894
rect 567586 676658 567822 676894
rect 567266 676338 567502 676574
rect 567586 676338 567822 676574
rect 567266 640658 567502 640894
rect 567586 640658 567822 640894
rect 567266 640338 567502 640574
rect 567586 640338 567822 640574
rect 567266 604658 567502 604894
rect 567586 604658 567822 604894
rect 567266 604338 567502 604574
rect 567586 604338 567822 604574
rect 567266 568658 567502 568894
rect 567586 568658 567822 568894
rect 567266 568338 567502 568574
rect 567586 568338 567822 568574
rect 567266 532658 567502 532894
rect 567586 532658 567822 532894
rect 567266 532338 567502 532574
rect 567586 532338 567822 532574
rect 567266 496658 567502 496894
rect 567586 496658 567822 496894
rect 567266 496338 567502 496574
rect 567586 496338 567822 496574
rect 567266 460658 567502 460894
rect 567586 460658 567822 460894
rect 567266 460338 567502 460574
rect 567586 460338 567822 460574
rect 567266 424658 567502 424894
rect 567586 424658 567822 424894
rect 567266 424338 567502 424574
rect 567586 424338 567822 424574
rect 567266 388658 567502 388894
rect 567586 388658 567822 388894
rect 567266 388338 567502 388574
rect 567586 388338 567822 388574
rect 567266 352658 567502 352894
rect 567586 352658 567822 352894
rect 567266 352338 567502 352574
rect 567586 352338 567822 352574
rect 567266 316658 567502 316894
rect 567586 316658 567822 316894
rect 567266 316338 567502 316574
rect 567586 316338 567822 316574
rect 567266 280658 567502 280894
rect 567586 280658 567822 280894
rect 567266 280338 567502 280574
rect 567586 280338 567822 280574
rect 567266 244658 567502 244894
rect 567586 244658 567822 244894
rect 567266 244338 567502 244574
rect 567586 244338 567822 244574
rect 567266 208658 567502 208894
rect 567586 208658 567822 208894
rect 567266 208338 567502 208574
rect 567586 208338 567822 208574
rect 567266 172658 567502 172894
rect 567586 172658 567822 172894
rect 567266 172338 567502 172574
rect 567586 172338 567822 172574
rect 567266 136658 567502 136894
rect 567586 136658 567822 136894
rect 567266 136338 567502 136574
rect 567586 136338 567822 136574
rect 567266 100658 567502 100894
rect 567586 100658 567822 100894
rect 567266 100338 567502 100574
rect 567586 100338 567822 100574
rect 567266 64658 567502 64894
rect 567586 64658 567822 64894
rect 567266 64338 567502 64574
rect 567586 64338 567822 64574
rect 567266 28658 567502 28894
rect 567586 28658 567822 28894
rect 567266 28338 567502 28574
rect 567586 28338 567822 28574
rect 567266 -5382 567502 -5146
rect 567586 -5382 567822 -5146
rect 567266 -5702 567502 -5466
rect 567586 -5702 567822 -5466
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 581546 706522 581782 706758
rect 581866 706522 582102 706758
rect 581546 706202 581782 706438
rect 581866 706202 582102 706438
rect 570986 680378 571222 680614
rect 571306 680378 571542 680614
rect 570986 680058 571222 680294
rect 571306 680058 571542 680294
rect 570986 644378 571222 644614
rect 571306 644378 571542 644614
rect 570986 644058 571222 644294
rect 571306 644058 571542 644294
rect 570986 608378 571222 608614
rect 571306 608378 571542 608614
rect 570986 608058 571222 608294
rect 571306 608058 571542 608294
rect 570986 572378 571222 572614
rect 571306 572378 571542 572614
rect 570986 572058 571222 572294
rect 571306 572058 571542 572294
rect 570986 536378 571222 536614
rect 571306 536378 571542 536614
rect 570986 536058 571222 536294
rect 571306 536058 571542 536294
rect 570986 500378 571222 500614
rect 571306 500378 571542 500614
rect 570986 500058 571222 500294
rect 571306 500058 571542 500294
rect 570986 464378 571222 464614
rect 571306 464378 571542 464614
rect 570986 464058 571222 464294
rect 571306 464058 571542 464294
rect 570986 428378 571222 428614
rect 571306 428378 571542 428614
rect 570986 428058 571222 428294
rect 571306 428058 571542 428294
rect 570986 392378 571222 392614
rect 571306 392378 571542 392614
rect 570986 392058 571222 392294
rect 571306 392058 571542 392294
rect 570986 356378 571222 356614
rect 571306 356378 571542 356614
rect 570986 356058 571222 356294
rect 571306 356058 571542 356294
rect 570986 320378 571222 320614
rect 571306 320378 571542 320614
rect 570986 320058 571222 320294
rect 571306 320058 571542 320294
rect 570986 284378 571222 284614
rect 571306 284378 571542 284614
rect 570986 284058 571222 284294
rect 571306 284058 571542 284294
rect 570986 248378 571222 248614
rect 571306 248378 571542 248614
rect 570986 248058 571222 248294
rect 571306 248058 571542 248294
rect 570986 212378 571222 212614
rect 571306 212378 571542 212614
rect 570986 212058 571222 212294
rect 571306 212058 571542 212294
rect 570986 176378 571222 176614
rect 571306 176378 571542 176614
rect 570986 176058 571222 176294
rect 571306 176058 571542 176294
rect 570986 140378 571222 140614
rect 571306 140378 571542 140614
rect 570986 140058 571222 140294
rect 571306 140058 571542 140294
rect 570986 104378 571222 104614
rect 571306 104378 571542 104614
rect 570986 104058 571222 104294
rect 571306 104058 571542 104294
rect 570986 68378 571222 68614
rect 571306 68378 571542 68614
rect 570986 68058 571222 68294
rect 571306 68058 571542 68294
rect 570986 32378 571222 32614
rect 571306 32378 571542 32614
rect 570986 32058 571222 32294
rect 571306 32058 571542 32294
rect 552986 -6342 553222 -6106
rect 553306 -6342 553542 -6106
rect 552986 -6662 553222 -6426
rect 553306 -6662 553542 -6426
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 669218 586538 669454
rect 586622 669218 586858 669454
rect 586302 668898 586538 669134
rect 586622 668898 586858 669134
rect 586302 633218 586538 633454
rect 586622 633218 586858 633454
rect 586302 632898 586538 633134
rect 586622 632898 586858 633134
rect 586302 597218 586538 597454
rect 586622 597218 586858 597454
rect 586302 596898 586538 597134
rect 586622 596898 586858 597134
rect 586302 561218 586538 561454
rect 586622 561218 586858 561454
rect 586302 560898 586538 561134
rect 586622 560898 586858 561134
rect 586302 525218 586538 525454
rect 586622 525218 586858 525454
rect 586302 524898 586538 525134
rect 586622 524898 586858 525134
rect 586302 489218 586538 489454
rect 586622 489218 586858 489454
rect 586302 488898 586538 489134
rect 586622 488898 586858 489134
rect 586302 453218 586538 453454
rect 586622 453218 586858 453454
rect 586302 452898 586538 453134
rect 586622 452898 586858 453134
rect 586302 417218 586538 417454
rect 586622 417218 586858 417454
rect 586302 416898 586538 417134
rect 586622 416898 586858 417134
rect 586302 381218 586538 381454
rect 586622 381218 586858 381454
rect 586302 380898 586538 381134
rect 586622 380898 586858 381134
rect 586302 345218 586538 345454
rect 586622 345218 586858 345454
rect 586302 344898 586538 345134
rect 586622 344898 586858 345134
rect 586302 309218 586538 309454
rect 586622 309218 586858 309454
rect 586302 308898 586538 309134
rect 586622 308898 586858 309134
rect 586302 273218 586538 273454
rect 586622 273218 586858 273454
rect 586302 272898 586538 273134
rect 586622 272898 586858 273134
rect 586302 237218 586538 237454
rect 586622 237218 586858 237454
rect 586302 236898 586538 237134
rect 586622 236898 586858 237134
rect 586302 201218 586538 201454
rect 586622 201218 586858 201454
rect 586302 200898 586538 201134
rect 586622 200898 586858 201134
rect 586302 165218 586538 165454
rect 586622 165218 586858 165454
rect 586302 164898 586538 165134
rect 586622 164898 586858 165134
rect 586302 129218 586538 129454
rect 586622 129218 586858 129454
rect 586302 128898 586538 129134
rect 586622 128898 586858 129134
rect 586302 93218 586538 93454
rect 586622 93218 586858 93454
rect 586302 92898 586538 93134
rect 586622 92898 586858 93134
rect 586302 57218 586538 57454
rect 586622 57218 586858 57454
rect 586302 56898 586538 57134
rect 586622 56898 586858 57134
rect 586302 21218 586538 21454
rect 586622 21218 586858 21454
rect 586302 20898 586538 21134
rect 586622 20898 586858 21134
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 690938 587498 691174
rect 587582 690938 587818 691174
rect 587262 690618 587498 690854
rect 587582 690618 587818 690854
rect 587262 654938 587498 655174
rect 587582 654938 587818 655174
rect 587262 654618 587498 654854
rect 587582 654618 587818 654854
rect 587262 618938 587498 619174
rect 587582 618938 587818 619174
rect 587262 618618 587498 618854
rect 587582 618618 587818 618854
rect 587262 582938 587498 583174
rect 587582 582938 587818 583174
rect 587262 582618 587498 582854
rect 587582 582618 587818 582854
rect 587262 546938 587498 547174
rect 587582 546938 587818 547174
rect 587262 546618 587498 546854
rect 587582 546618 587818 546854
rect 587262 510938 587498 511174
rect 587582 510938 587818 511174
rect 587262 510618 587498 510854
rect 587582 510618 587818 510854
rect 587262 474938 587498 475174
rect 587582 474938 587818 475174
rect 587262 474618 587498 474854
rect 587582 474618 587818 474854
rect 587262 438938 587498 439174
rect 587582 438938 587818 439174
rect 587262 438618 587498 438854
rect 587582 438618 587818 438854
rect 587262 402938 587498 403174
rect 587582 402938 587818 403174
rect 587262 402618 587498 402854
rect 587582 402618 587818 402854
rect 587262 366938 587498 367174
rect 587582 366938 587818 367174
rect 587262 366618 587498 366854
rect 587582 366618 587818 366854
rect 587262 330938 587498 331174
rect 587582 330938 587818 331174
rect 587262 330618 587498 330854
rect 587582 330618 587818 330854
rect 587262 294938 587498 295174
rect 587582 294938 587818 295174
rect 587262 294618 587498 294854
rect 587582 294618 587818 294854
rect 587262 258938 587498 259174
rect 587582 258938 587818 259174
rect 587262 258618 587498 258854
rect 587582 258618 587818 258854
rect 587262 222938 587498 223174
rect 587582 222938 587818 223174
rect 587262 222618 587498 222854
rect 587582 222618 587818 222854
rect 587262 186938 587498 187174
rect 587582 186938 587818 187174
rect 587262 186618 587498 186854
rect 587582 186618 587818 186854
rect 587262 150938 587498 151174
rect 587582 150938 587818 151174
rect 587262 150618 587498 150854
rect 587582 150618 587818 150854
rect 587262 114938 587498 115174
rect 587582 114938 587818 115174
rect 587262 114618 587498 114854
rect 587582 114618 587818 114854
rect 587262 78938 587498 79174
rect 587582 78938 587818 79174
rect 587262 78618 587498 78854
rect 587582 78618 587818 78854
rect 587262 42938 587498 43174
rect 587582 42938 587818 43174
rect 587262 42618 587498 42854
rect 587582 42618 587818 42854
rect 587262 6938 587498 7174
rect 587582 6938 587818 7174
rect 587262 6618 587498 6854
rect 587582 6618 587818 6854
rect 581546 -2502 581782 -2266
rect 581866 -2502 582102 -2266
rect 581546 -2822 581782 -2586
rect 581866 -2822 582102 -2586
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 672938 588458 673174
rect 588542 672938 588778 673174
rect 588222 672618 588458 672854
rect 588542 672618 588778 672854
rect 588222 636938 588458 637174
rect 588542 636938 588778 637174
rect 588222 636618 588458 636854
rect 588542 636618 588778 636854
rect 588222 600938 588458 601174
rect 588542 600938 588778 601174
rect 588222 600618 588458 600854
rect 588542 600618 588778 600854
rect 588222 564938 588458 565174
rect 588542 564938 588778 565174
rect 588222 564618 588458 564854
rect 588542 564618 588778 564854
rect 588222 528938 588458 529174
rect 588542 528938 588778 529174
rect 588222 528618 588458 528854
rect 588542 528618 588778 528854
rect 588222 492938 588458 493174
rect 588542 492938 588778 493174
rect 588222 492618 588458 492854
rect 588542 492618 588778 492854
rect 588222 456938 588458 457174
rect 588542 456938 588778 457174
rect 588222 456618 588458 456854
rect 588542 456618 588778 456854
rect 588222 420938 588458 421174
rect 588542 420938 588778 421174
rect 588222 420618 588458 420854
rect 588542 420618 588778 420854
rect 588222 384938 588458 385174
rect 588542 384938 588778 385174
rect 588222 384618 588458 384854
rect 588542 384618 588778 384854
rect 588222 348938 588458 349174
rect 588542 348938 588778 349174
rect 588222 348618 588458 348854
rect 588542 348618 588778 348854
rect 588222 312938 588458 313174
rect 588542 312938 588778 313174
rect 588222 312618 588458 312854
rect 588542 312618 588778 312854
rect 588222 276938 588458 277174
rect 588542 276938 588778 277174
rect 588222 276618 588458 276854
rect 588542 276618 588778 276854
rect 588222 240938 588458 241174
rect 588542 240938 588778 241174
rect 588222 240618 588458 240854
rect 588542 240618 588778 240854
rect 588222 204938 588458 205174
rect 588542 204938 588778 205174
rect 588222 204618 588458 204854
rect 588542 204618 588778 204854
rect 588222 168938 588458 169174
rect 588542 168938 588778 169174
rect 588222 168618 588458 168854
rect 588542 168618 588778 168854
rect 588222 132938 588458 133174
rect 588542 132938 588778 133174
rect 588222 132618 588458 132854
rect 588542 132618 588778 132854
rect 588222 96938 588458 97174
rect 588542 96938 588778 97174
rect 588222 96618 588458 96854
rect 588542 96618 588778 96854
rect 588222 60938 588458 61174
rect 588542 60938 588778 61174
rect 588222 60618 588458 60854
rect 588542 60618 588778 60854
rect 588222 24938 588458 25174
rect 588542 24938 588778 25174
rect 588222 24618 588458 24854
rect 588542 24618 588778 24854
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 694658 589418 694894
rect 589502 694658 589738 694894
rect 589182 694338 589418 694574
rect 589502 694338 589738 694574
rect 589182 658658 589418 658894
rect 589502 658658 589738 658894
rect 589182 658338 589418 658574
rect 589502 658338 589738 658574
rect 589182 622658 589418 622894
rect 589502 622658 589738 622894
rect 589182 622338 589418 622574
rect 589502 622338 589738 622574
rect 589182 586658 589418 586894
rect 589502 586658 589738 586894
rect 589182 586338 589418 586574
rect 589502 586338 589738 586574
rect 589182 550658 589418 550894
rect 589502 550658 589738 550894
rect 589182 550338 589418 550574
rect 589502 550338 589738 550574
rect 589182 514658 589418 514894
rect 589502 514658 589738 514894
rect 589182 514338 589418 514574
rect 589502 514338 589738 514574
rect 589182 478658 589418 478894
rect 589502 478658 589738 478894
rect 589182 478338 589418 478574
rect 589502 478338 589738 478574
rect 589182 442658 589418 442894
rect 589502 442658 589738 442894
rect 589182 442338 589418 442574
rect 589502 442338 589738 442574
rect 589182 406658 589418 406894
rect 589502 406658 589738 406894
rect 589182 406338 589418 406574
rect 589502 406338 589738 406574
rect 589182 370658 589418 370894
rect 589502 370658 589738 370894
rect 589182 370338 589418 370574
rect 589502 370338 589738 370574
rect 589182 334658 589418 334894
rect 589502 334658 589738 334894
rect 589182 334338 589418 334574
rect 589502 334338 589738 334574
rect 589182 298658 589418 298894
rect 589502 298658 589738 298894
rect 589182 298338 589418 298574
rect 589502 298338 589738 298574
rect 589182 262658 589418 262894
rect 589502 262658 589738 262894
rect 589182 262338 589418 262574
rect 589502 262338 589738 262574
rect 589182 226658 589418 226894
rect 589502 226658 589738 226894
rect 589182 226338 589418 226574
rect 589502 226338 589738 226574
rect 589182 190658 589418 190894
rect 589502 190658 589738 190894
rect 589182 190338 589418 190574
rect 589502 190338 589738 190574
rect 589182 154658 589418 154894
rect 589502 154658 589738 154894
rect 589182 154338 589418 154574
rect 589502 154338 589738 154574
rect 589182 118658 589418 118894
rect 589502 118658 589738 118894
rect 589182 118338 589418 118574
rect 589502 118338 589738 118574
rect 589182 82658 589418 82894
rect 589502 82658 589738 82894
rect 589182 82338 589418 82574
rect 589502 82338 589738 82574
rect 589182 46658 589418 46894
rect 589502 46658 589738 46894
rect 589182 46338 589418 46574
rect 589502 46338 589738 46574
rect 589182 10658 589418 10894
rect 589502 10658 589738 10894
rect 589182 10338 589418 10574
rect 589502 10338 589738 10574
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 676658 590378 676894
rect 590462 676658 590698 676894
rect 590142 676338 590378 676574
rect 590462 676338 590698 676574
rect 590142 640658 590378 640894
rect 590462 640658 590698 640894
rect 590142 640338 590378 640574
rect 590462 640338 590698 640574
rect 590142 604658 590378 604894
rect 590462 604658 590698 604894
rect 590142 604338 590378 604574
rect 590462 604338 590698 604574
rect 590142 568658 590378 568894
rect 590462 568658 590698 568894
rect 590142 568338 590378 568574
rect 590462 568338 590698 568574
rect 590142 532658 590378 532894
rect 590462 532658 590698 532894
rect 590142 532338 590378 532574
rect 590462 532338 590698 532574
rect 590142 496658 590378 496894
rect 590462 496658 590698 496894
rect 590142 496338 590378 496574
rect 590462 496338 590698 496574
rect 590142 460658 590378 460894
rect 590462 460658 590698 460894
rect 590142 460338 590378 460574
rect 590462 460338 590698 460574
rect 590142 424658 590378 424894
rect 590462 424658 590698 424894
rect 590142 424338 590378 424574
rect 590462 424338 590698 424574
rect 590142 388658 590378 388894
rect 590462 388658 590698 388894
rect 590142 388338 590378 388574
rect 590462 388338 590698 388574
rect 590142 352658 590378 352894
rect 590462 352658 590698 352894
rect 590142 352338 590378 352574
rect 590462 352338 590698 352574
rect 590142 316658 590378 316894
rect 590462 316658 590698 316894
rect 590142 316338 590378 316574
rect 590462 316338 590698 316574
rect 590142 280658 590378 280894
rect 590462 280658 590698 280894
rect 590142 280338 590378 280574
rect 590462 280338 590698 280574
rect 590142 244658 590378 244894
rect 590462 244658 590698 244894
rect 590142 244338 590378 244574
rect 590462 244338 590698 244574
rect 590142 208658 590378 208894
rect 590462 208658 590698 208894
rect 590142 208338 590378 208574
rect 590462 208338 590698 208574
rect 590142 172658 590378 172894
rect 590462 172658 590698 172894
rect 590142 172338 590378 172574
rect 590462 172338 590698 172574
rect 590142 136658 590378 136894
rect 590462 136658 590698 136894
rect 590142 136338 590378 136574
rect 590462 136338 590698 136574
rect 590142 100658 590378 100894
rect 590462 100658 590698 100894
rect 590142 100338 590378 100574
rect 590462 100338 590698 100574
rect 590142 64658 590378 64894
rect 590462 64658 590698 64894
rect 590142 64338 590378 64574
rect 590462 64338 590698 64574
rect 590142 28658 590378 28894
rect 590462 28658 590698 28894
rect 590142 28338 590378 28574
rect 590462 28338 590698 28574
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 698378 591338 698614
rect 591422 698378 591658 698614
rect 591102 698058 591338 698294
rect 591422 698058 591658 698294
rect 591102 662378 591338 662614
rect 591422 662378 591658 662614
rect 591102 662058 591338 662294
rect 591422 662058 591658 662294
rect 591102 626378 591338 626614
rect 591422 626378 591658 626614
rect 591102 626058 591338 626294
rect 591422 626058 591658 626294
rect 591102 590378 591338 590614
rect 591422 590378 591658 590614
rect 591102 590058 591338 590294
rect 591422 590058 591658 590294
rect 591102 554378 591338 554614
rect 591422 554378 591658 554614
rect 591102 554058 591338 554294
rect 591422 554058 591658 554294
rect 591102 518378 591338 518614
rect 591422 518378 591658 518614
rect 591102 518058 591338 518294
rect 591422 518058 591658 518294
rect 591102 482378 591338 482614
rect 591422 482378 591658 482614
rect 591102 482058 591338 482294
rect 591422 482058 591658 482294
rect 591102 446378 591338 446614
rect 591422 446378 591658 446614
rect 591102 446058 591338 446294
rect 591422 446058 591658 446294
rect 591102 410378 591338 410614
rect 591422 410378 591658 410614
rect 591102 410058 591338 410294
rect 591422 410058 591658 410294
rect 591102 374378 591338 374614
rect 591422 374378 591658 374614
rect 591102 374058 591338 374294
rect 591422 374058 591658 374294
rect 591102 338378 591338 338614
rect 591422 338378 591658 338614
rect 591102 338058 591338 338294
rect 591422 338058 591658 338294
rect 591102 302378 591338 302614
rect 591422 302378 591658 302614
rect 591102 302058 591338 302294
rect 591422 302058 591658 302294
rect 591102 266378 591338 266614
rect 591422 266378 591658 266614
rect 591102 266058 591338 266294
rect 591422 266058 591658 266294
rect 591102 230378 591338 230614
rect 591422 230378 591658 230614
rect 591102 230058 591338 230294
rect 591422 230058 591658 230294
rect 591102 194378 591338 194614
rect 591422 194378 591658 194614
rect 591102 194058 591338 194294
rect 591422 194058 591658 194294
rect 591102 158378 591338 158614
rect 591422 158378 591658 158614
rect 591102 158058 591338 158294
rect 591422 158058 591658 158294
rect 591102 122378 591338 122614
rect 591422 122378 591658 122614
rect 591102 122058 591338 122294
rect 591422 122058 591658 122294
rect 591102 86378 591338 86614
rect 591422 86378 591658 86614
rect 591102 86058 591338 86294
rect 591422 86058 591658 86294
rect 591102 50378 591338 50614
rect 591422 50378 591658 50614
rect 591102 50058 591338 50294
rect 591422 50058 591658 50294
rect 591102 14378 591338 14614
rect 591422 14378 591658 14614
rect 591102 14058 591338 14294
rect 591422 14058 591658 14294
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 680378 592298 680614
rect 592382 680378 592618 680614
rect 592062 680058 592298 680294
rect 592382 680058 592618 680294
rect 592062 644378 592298 644614
rect 592382 644378 592618 644614
rect 592062 644058 592298 644294
rect 592382 644058 592618 644294
rect 592062 608378 592298 608614
rect 592382 608378 592618 608614
rect 592062 608058 592298 608294
rect 592382 608058 592618 608294
rect 592062 572378 592298 572614
rect 592382 572378 592618 572614
rect 592062 572058 592298 572294
rect 592382 572058 592618 572294
rect 592062 536378 592298 536614
rect 592382 536378 592618 536614
rect 592062 536058 592298 536294
rect 592382 536058 592618 536294
rect 592062 500378 592298 500614
rect 592382 500378 592618 500614
rect 592062 500058 592298 500294
rect 592382 500058 592618 500294
rect 592062 464378 592298 464614
rect 592382 464378 592618 464614
rect 592062 464058 592298 464294
rect 592382 464058 592618 464294
rect 592062 428378 592298 428614
rect 592382 428378 592618 428614
rect 592062 428058 592298 428294
rect 592382 428058 592618 428294
rect 592062 392378 592298 392614
rect 592382 392378 592618 392614
rect 592062 392058 592298 392294
rect 592382 392058 592618 392294
rect 592062 356378 592298 356614
rect 592382 356378 592618 356614
rect 592062 356058 592298 356294
rect 592382 356058 592618 356294
rect 592062 320378 592298 320614
rect 592382 320378 592618 320614
rect 592062 320058 592298 320294
rect 592382 320058 592618 320294
rect 592062 284378 592298 284614
rect 592382 284378 592618 284614
rect 592062 284058 592298 284294
rect 592382 284058 592618 284294
rect 592062 248378 592298 248614
rect 592382 248378 592618 248614
rect 592062 248058 592298 248294
rect 592382 248058 592618 248294
rect 592062 212378 592298 212614
rect 592382 212378 592618 212614
rect 592062 212058 592298 212294
rect 592382 212058 592618 212294
rect 592062 176378 592298 176614
rect 592382 176378 592618 176614
rect 592062 176058 592298 176294
rect 592382 176058 592618 176294
rect 592062 140378 592298 140614
rect 592382 140378 592618 140614
rect 592062 140058 592298 140294
rect 592382 140058 592618 140294
rect 592062 104378 592298 104614
rect 592382 104378 592618 104614
rect 592062 104058 592298 104294
rect 592382 104058 592618 104294
rect 592062 68378 592298 68614
rect 592382 68378 592618 68614
rect 592062 68058 592298 68294
rect 592382 68058 592618 68294
rect 592062 32378 592298 32614
rect 592382 32378 592618 32614
rect 592062 32058 592298 32294
rect 592382 32058 592618 32294
rect 570986 -7302 571222 -7066
rect 571306 -7302 571542 -7066
rect 570986 -7622 571222 -7386
rect 571306 -7622 571542 -7386
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 592650 698294
rect -8726 698026 592650 698058
rect -6806 694894 590730 694926
rect -6806 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 590730 694894
rect -6806 694574 590730 694658
rect -6806 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 590730 694574
rect -6806 694306 590730 694338
rect -4886 691174 588810 691206
rect -4886 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 588810 691174
rect -4886 690854 588810 690938
rect -4886 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 588810 690854
rect -4886 690586 588810 690618
rect -2966 687454 586890 687486
rect -2966 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 586890 687454
rect -2966 687134 586890 687218
rect -2966 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 586890 687134
rect -2966 686866 586890 686898
rect -8726 680614 592650 680646
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect -8726 680294 592650 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect -8726 680026 592650 680058
rect -6806 676894 590730 676926
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect -6806 676574 590730 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect -6806 676306 590730 676338
rect -4886 673174 588810 673206
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect -4886 672854 588810 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect -4886 672586 588810 672618
rect -2966 669454 586890 669486
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect -2966 669134 586890 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect -2966 668866 586890 668898
rect -8726 662614 592650 662646
rect -8726 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 592650 662294
rect -8726 662026 592650 662058
rect -6806 658894 590730 658926
rect -6806 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 590730 658894
rect -6806 658574 590730 658658
rect -6806 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 590730 658574
rect -6806 658306 590730 658338
rect -4886 655174 588810 655206
rect -4886 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 588810 655174
rect -4886 654854 588810 654938
rect -4886 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 588810 654854
rect -4886 654586 588810 654618
rect -2966 651454 586890 651486
rect -2966 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 586890 651454
rect -2966 651134 586890 651218
rect -2966 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 586890 651134
rect -2966 650866 586890 650898
rect -8726 644614 592650 644646
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect -8726 644294 592650 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect -8726 644026 592650 644058
rect -6806 640894 590730 640926
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect -6806 640574 590730 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect -6806 640306 590730 640338
rect -4886 637174 588810 637206
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect -4886 636854 588810 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect -4886 636586 588810 636618
rect -2966 633454 586890 633486
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect -2966 633134 586890 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect -2966 632866 586890 632898
rect -8726 626614 592650 626646
rect -8726 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 592650 626294
rect -8726 626026 592650 626058
rect -6806 622894 590730 622926
rect -6806 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 590730 622894
rect -6806 622574 590730 622658
rect -6806 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 590730 622574
rect -6806 622306 590730 622338
rect -4886 619174 588810 619206
rect -4886 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 588810 619174
rect -4886 618854 588810 618938
rect -4886 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 588810 618854
rect -4886 618586 588810 618618
rect -2966 615454 586890 615486
rect -2966 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 586890 615454
rect -2966 615134 586890 615218
rect -2966 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 586890 615134
rect -2966 614866 586890 614898
rect -8726 608614 592650 608646
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect -8726 608294 592650 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect -8726 608026 592650 608058
rect -6806 604894 590730 604926
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect -6806 604574 590730 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect -6806 604306 590730 604338
rect -4886 601174 588810 601206
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect -4886 600854 588810 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect -4886 600586 588810 600618
rect -2966 597454 586890 597486
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect -2966 597134 586890 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect -2966 596866 586890 596898
rect -8726 590614 592650 590646
rect -8726 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 592650 590294
rect -8726 590026 592650 590058
rect -6806 586894 590730 586926
rect -6806 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 590730 586894
rect -6806 586574 590730 586658
rect -6806 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 590730 586574
rect -6806 586306 590730 586338
rect -4886 583174 588810 583206
rect -4886 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 77546 583174
rect 77782 582938 77866 583174
rect 78102 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 588810 583174
rect -4886 582854 588810 582938
rect -4886 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 77546 582854
rect 77782 582618 77866 582854
rect 78102 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 588810 582854
rect -4886 582586 588810 582618
rect -2966 579454 586890 579486
rect -2966 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 586890 579454
rect -2966 579134 586890 579218
rect -2966 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 586890 579134
rect -2966 578866 586890 578898
rect -8726 572614 592650 572646
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect -8726 572294 592650 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect -8726 572026 592650 572058
rect -6806 568894 590730 568926
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect -6806 568574 590730 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect -6806 568306 590730 568338
rect -4886 565174 588810 565206
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 95546 565174
rect 95782 564938 95866 565174
rect 96102 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect -4886 564854 588810 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 95546 564854
rect 95782 564618 95866 564854
rect 96102 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect -4886 564586 588810 564618
rect -2966 561454 586890 561486
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect -2966 561134 586890 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect -2966 560866 586890 560898
rect -8726 554614 592650 554646
rect -8726 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 84986 554614
rect 85222 554378 85306 554614
rect 85542 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 84986 554294
rect 85222 554058 85306 554294
rect 85542 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 592650 554294
rect -8726 554026 592650 554058
rect -6806 550894 590730 550926
rect -6806 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 81266 550894
rect 81502 550658 81586 550894
rect 81822 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 590730 550894
rect -6806 550574 590730 550658
rect -6806 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 81266 550574
rect 81502 550338 81586 550574
rect 81822 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 590730 550574
rect -6806 550306 590730 550338
rect -4886 547174 588810 547206
rect -4886 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 77546 547174
rect 77782 546938 77866 547174
rect 78102 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 588810 547174
rect -4886 546854 588810 546938
rect -4886 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 77546 546854
rect 77782 546618 77866 546854
rect 78102 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 588810 546854
rect -4886 546586 588810 546618
rect -2966 543454 586890 543486
rect -2966 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 586890 543454
rect -2966 543134 586890 543218
rect -2966 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 586890 543134
rect -2966 542866 586890 542898
rect -8726 536614 592650 536646
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 174986 536614
rect 175222 536378 175306 536614
rect 175542 536378 210986 536614
rect 211222 536378 211306 536614
rect 211542 536378 246986 536614
rect 247222 536378 247306 536614
rect 247542 536378 282986 536614
rect 283222 536378 283306 536614
rect 283542 536378 318986 536614
rect 319222 536378 319306 536614
rect 319542 536378 354986 536614
rect 355222 536378 355306 536614
rect 355542 536378 390986 536614
rect 391222 536378 391306 536614
rect 391542 536378 426986 536614
rect 427222 536378 427306 536614
rect 427542 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect -8726 536294 592650 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 174986 536294
rect 175222 536058 175306 536294
rect 175542 536058 210986 536294
rect 211222 536058 211306 536294
rect 211542 536058 246986 536294
rect 247222 536058 247306 536294
rect 247542 536058 282986 536294
rect 283222 536058 283306 536294
rect 283542 536058 318986 536294
rect 319222 536058 319306 536294
rect 319542 536058 354986 536294
rect 355222 536058 355306 536294
rect 355542 536058 390986 536294
rect 391222 536058 391306 536294
rect 391542 536058 426986 536294
rect 427222 536058 427306 536294
rect 427542 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect -8726 536026 592650 536058
rect -6806 532894 590730 532926
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 171266 532894
rect 171502 532658 171586 532894
rect 171822 532658 207266 532894
rect 207502 532658 207586 532894
rect 207822 532658 243266 532894
rect 243502 532658 243586 532894
rect 243822 532658 279266 532894
rect 279502 532658 279586 532894
rect 279822 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 351266 532894
rect 351502 532658 351586 532894
rect 351822 532658 387266 532894
rect 387502 532658 387586 532894
rect 387822 532658 423266 532894
rect 423502 532658 423586 532894
rect 423822 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect -6806 532574 590730 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 171266 532574
rect 171502 532338 171586 532574
rect 171822 532338 207266 532574
rect 207502 532338 207586 532574
rect 207822 532338 243266 532574
rect 243502 532338 243586 532574
rect 243822 532338 279266 532574
rect 279502 532338 279586 532574
rect 279822 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 351266 532574
rect 351502 532338 351586 532574
rect 351822 532338 387266 532574
rect 387502 532338 387586 532574
rect 387822 532338 423266 532574
rect 423502 532338 423586 532574
rect 423822 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect -6806 532306 590730 532338
rect -4886 529174 588810 529206
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 167546 529174
rect 167782 528938 167866 529174
rect 168102 528938 203546 529174
rect 203782 528938 203866 529174
rect 204102 528938 239546 529174
rect 239782 528938 239866 529174
rect 240102 528938 275546 529174
rect 275782 528938 275866 529174
rect 276102 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 347546 529174
rect 347782 528938 347866 529174
rect 348102 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 419546 529174
rect 419782 528938 419866 529174
rect 420102 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect -4886 528854 588810 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 167546 528854
rect 167782 528618 167866 528854
rect 168102 528618 203546 528854
rect 203782 528618 203866 528854
rect 204102 528618 239546 528854
rect 239782 528618 239866 528854
rect 240102 528618 275546 528854
rect 275782 528618 275866 528854
rect 276102 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 347546 528854
rect 347782 528618 347866 528854
rect 348102 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 419546 528854
rect 419782 528618 419866 528854
rect 420102 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect -4886 528586 588810 528618
rect -2966 525454 586890 525486
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect -2966 525134 586890 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect -2966 524866 586890 524898
rect -8726 518614 592650 518646
rect -8726 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 592650 518294
rect -8726 518026 592650 518058
rect -6806 514894 590730 514926
rect -6806 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 590730 514894
rect -6806 514574 590730 514658
rect -6806 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 590730 514574
rect -6806 514306 590730 514338
rect -4886 511174 588810 511206
rect -4886 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 588810 511174
rect -4886 510854 588810 510938
rect -4886 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 588810 510854
rect -4886 510586 588810 510618
rect -2966 507454 586890 507486
rect -2966 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 586890 507454
rect -2966 507134 586890 507218
rect -2966 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 586890 507134
rect -2966 506866 586890 506898
rect -8726 500614 592650 500646
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 138986 500614
rect 139222 500378 139306 500614
rect 139542 500378 174986 500614
rect 175222 500378 175306 500614
rect 175542 500378 210986 500614
rect 211222 500378 211306 500614
rect 211542 500378 246986 500614
rect 247222 500378 247306 500614
rect 247542 500378 282986 500614
rect 283222 500378 283306 500614
rect 283542 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect -8726 500294 592650 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 138986 500294
rect 139222 500058 139306 500294
rect 139542 500058 174986 500294
rect 175222 500058 175306 500294
rect 175542 500058 210986 500294
rect 211222 500058 211306 500294
rect 211542 500058 246986 500294
rect 247222 500058 247306 500294
rect 247542 500058 282986 500294
rect 283222 500058 283306 500294
rect 283542 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect -8726 500026 592650 500058
rect -6806 496894 590730 496926
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 171266 496894
rect 171502 496658 171586 496894
rect 171822 496658 207266 496894
rect 207502 496658 207586 496894
rect 207822 496658 243266 496894
rect 243502 496658 243586 496894
rect 243822 496658 279266 496894
rect 279502 496658 279586 496894
rect 279822 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect -6806 496574 590730 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 171266 496574
rect 171502 496338 171586 496574
rect 171822 496338 207266 496574
rect 207502 496338 207586 496574
rect 207822 496338 243266 496574
rect 243502 496338 243586 496574
rect 243822 496338 279266 496574
rect 279502 496338 279586 496574
rect 279822 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect -6806 496306 590730 496338
rect -4886 493174 588810 493206
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 167546 493174
rect 167782 492938 167866 493174
rect 168102 492938 203546 493174
rect 203782 492938 203866 493174
rect 204102 492938 239546 493174
rect 239782 492938 239866 493174
rect 240102 492938 275546 493174
rect 275782 492938 275866 493174
rect 276102 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect -4886 492854 588810 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 167546 492854
rect 167782 492618 167866 492854
rect 168102 492618 203546 492854
rect 203782 492618 203866 492854
rect 204102 492618 239546 492854
rect 239782 492618 239866 492854
rect 240102 492618 275546 492854
rect 275782 492618 275866 492854
rect 276102 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect -4886 492586 588810 492618
rect -2966 489454 586890 489486
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect -2966 489134 586890 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect -2966 488866 586890 488898
rect -8726 482614 592650 482646
rect -8726 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 592650 482294
rect -8726 482026 592650 482058
rect -6806 478894 590730 478926
rect -6806 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 590730 478894
rect -6806 478574 590730 478658
rect -6806 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 590730 478574
rect -6806 478306 590730 478338
rect -4886 475174 588810 475206
rect -4886 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 588810 475174
rect -4886 474854 588810 474938
rect -4886 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 588810 474854
rect -4886 474586 588810 474618
rect -2966 471454 586890 471486
rect -2966 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 586890 471454
rect -2966 471134 586890 471218
rect -2966 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 586890 471134
rect -2966 470866 586890 470898
rect -8726 464614 592650 464646
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 102986 464614
rect 103222 464378 103306 464614
rect 103542 464378 138986 464614
rect 139222 464378 139306 464614
rect 139542 464378 174986 464614
rect 175222 464378 175306 464614
rect 175542 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 246986 464614
rect 247222 464378 247306 464614
rect 247542 464378 282986 464614
rect 283222 464378 283306 464614
rect 283542 464378 318986 464614
rect 319222 464378 319306 464614
rect 319542 464378 354986 464614
rect 355222 464378 355306 464614
rect 355542 464378 390986 464614
rect 391222 464378 391306 464614
rect 391542 464378 426986 464614
rect 427222 464378 427306 464614
rect 427542 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect -8726 464294 592650 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 102986 464294
rect 103222 464058 103306 464294
rect 103542 464058 138986 464294
rect 139222 464058 139306 464294
rect 139542 464058 174986 464294
rect 175222 464058 175306 464294
rect 175542 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 246986 464294
rect 247222 464058 247306 464294
rect 247542 464058 282986 464294
rect 283222 464058 283306 464294
rect 283542 464058 318986 464294
rect 319222 464058 319306 464294
rect 319542 464058 354986 464294
rect 355222 464058 355306 464294
rect 355542 464058 390986 464294
rect 391222 464058 391306 464294
rect 391542 464058 426986 464294
rect 427222 464058 427306 464294
rect 427542 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect -8726 464026 592650 464058
rect -6806 460894 590730 460926
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 99266 460894
rect 99502 460658 99586 460894
rect 99822 460658 135266 460894
rect 135502 460658 135586 460894
rect 135822 460658 171266 460894
rect 171502 460658 171586 460894
rect 171822 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 243266 460894
rect 243502 460658 243586 460894
rect 243822 460658 279266 460894
rect 279502 460658 279586 460894
rect 279822 460658 315266 460894
rect 315502 460658 315586 460894
rect 315822 460658 351266 460894
rect 351502 460658 351586 460894
rect 351822 460658 387266 460894
rect 387502 460658 387586 460894
rect 387822 460658 423266 460894
rect 423502 460658 423586 460894
rect 423822 460658 459266 460894
rect 459502 460658 459586 460894
rect 459822 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect -6806 460574 590730 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 99266 460574
rect 99502 460338 99586 460574
rect 99822 460338 135266 460574
rect 135502 460338 135586 460574
rect 135822 460338 171266 460574
rect 171502 460338 171586 460574
rect 171822 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 243266 460574
rect 243502 460338 243586 460574
rect 243822 460338 279266 460574
rect 279502 460338 279586 460574
rect 279822 460338 315266 460574
rect 315502 460338 315586 460574
rect 315822 460338 351266 460574
rect 351502 460338 351586 460574
rect 351822 460338 387266 460574
rect 387502 460338 387586 460574
rect 387822 460338 423266 460574
rect 423502 460338 423586 460574
rect 423822 460338 459266 460574
rect 459502 460338 459586 460574
rect 459822 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect -6806 460306 590730 460338
rect -4886 457174 588810 457206
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 95546 457174
rect 95782 456938 95866 457174
rect 96102 456938 131546 457174
rect 131782 456938 131866 457174
rect 132102 456938 167546 457174
rect 167782 456938 167866 457174
rect 168102 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 239546 457174
rect 239782 456938 239866 457174
rect 240102 456938 275546 457174
rect 275782 456938 275866 457174
rect 276102 456938 311546 457174
rect 311782 456938 311866 457174
rect 312102 456938 347546 457174
rect 347782 456938 347866 457174
rect 348102 456938 383546 457174
rect 383782 456938 383866 457174
rect 384102 456938 419546 457174
rect 419782 456938 419866 457174
rect 420102 456938 455546 457174
rect 455782 456938 455866 457174
rect 456102 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect -4886 456854 588810 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 95546 456854
rect 95782 456618 95866 456854
rect 96102 456618 131546 456854
rect 131782 456618 131866 456854
rect 132102 456618 167546 456854
rect 167782 456618 167866 456854
rect 168102 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 239546 456854
rect 239782 456618 239866 456854
rect 240102 456618 275546 456854
rect 275782 456618 275866 456854
rect 276102 456618 311546 456854
rect 311782 456618 311866 456854
rect 312102 456618 347546 456854
rect 347782 456618 347866 456854
rect 348102 456618 383546 456854
rect 383782 456618 383866 456854
rect 384102 456618 419546 456854
rect 419782 456618 419866 456854
rect 420102 456618 455546 456854
rect 455782 456618 455866 456854
rect 456102 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect -4886 456586 588810 456618
rect -2966 453454 586890 453486
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect -2966 453134 586890 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect -2966 452866 586890 452898
rect -8726 446614 592650 446646
rect -8726 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 84986 446614
rect 85222 446378 85306 446614
rect 85542 446378 120986 446614
rect 121222 446378 121306 446614
rect 121542 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 192986 446614
rect 193222 446378 193306 446614
rect 193542 446378 228986 446614
rect 229222 446378 229306 446614
rect 229542 446378 264986 446614
rect 265222 446378 265306 446614
rect 265542 446378 300986 446614
rect 301222 446378 301306 446614
rect 301542 446378 336986 446614
rect 337222 446378 337306 446614
rect 337542 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 84986 446294
rect 85222 446058 85306 446294
rect 85542 446058 120986 446294
rect 121222 446058 121306 446294
rect 121542 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 192986 446294
rect 193222 446058 193306 446294
rect 193542 446058 228986 446294
rect 229222 446058 229306 446294
rect 229542 446058 264986 446294
rect 265222 446058 265306 446294
rect 265542 446058 300986 446294
rect 301222 446058 301306 446294
rect 301542 446058 336986 446294
rect 337222 446058 337306 446294
rect 337542 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 592650 446294
rect -8726 446026 592650 446058
rect -6806 442894 590730 442926
rect -6806 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 81266 442894
rect 81502 442658 81586 442894
rect 81822 442658 117266 442894
rect 117502 442658 117586 442894
rect 117822 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 225266 442894
rect 225502 442658 225586 442894
rect 225822 442658 261266 442894
rect 261502 442658 261586 442894
rect 261822 442658 297266 442894
rect 297502 442658 297586 442894
rect 297822 442658 333266 442894
rect 333502 442658 333586 442894
rect 333822 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 441266 442894
rect 441502 442658 441586 442894
rect 441822 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 590730 442894
rect -6806 442574 590730 442658
rect -6806 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 81266 442574
rect 81502 442338 81586 442574
rect 81822 442338 117266 442574
rect 117502 442338 117586 442574
rect 117822 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 225266 442574
rect 225502 442338 225586 442574
rect 225822 442338 261266 442574
rect 261502 442338 261586 442574
rect 261822 442338 297266 442574
rect 297502 442338 297586 442574
rect 297822 442338 333266 442574
rect 333502 442338 333586 442574
rect 333822 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 441266 442574
rect 441502 442338 441586 442574
rect 441822 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 590730 442574
rect -6806 442306 590730 442338
rect -4886 439174 588810 439206
rect -4886 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 77546 439174
rect 77782 438938 77866 439174
rect 78102 438938 113546 439174
rect 113782 438938 113866 439174
rect 114102 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 221546 439174
rect 221782 438938 221866 439174
rect 222102 438938 257546 439174
rect 257782 438938 257866 439174
rect 258102 438938 293546 439174
rect 293782 438938 293866 439174
rect 294102 438938 329546 439174
rect 329782 438938 329866 439174
rect 330102 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 588810 439174
rect -4886 438854 588810 438938
rect -4886 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 77546 438854
rect 77782 438618 77866 438854
rect 78102 438618 113546 438854
rect 113782 438618 113866 438854
rect 114102 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 221546 438854
rect 221782 438618 221866 438854
rect 222102 438618 257546 438854
rect 257782 438618 257866 438854
rect 258102 438618 293546 438854
rect 293782 438618 293866 438854
rect 294102 438618 329546 438854
rect 329782 438618 329866 438854
rect 330102 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 588810 438854
rect -4886 438586 588810 438618
rect -2966 435454 586890 435486
rect -2966 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 586890 435454
rect -2966 435134 586890 435218
rect -2966 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 586890 435134
rect -2966 434866 586890 434898
rect -8726 428614 592650 428646
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 66986 428614
rect 67222 428378 67306 428614
rect 67542 428378 102986 428614
rect 103222 428378 103306 428614
rect 103542 428378 138986 428614
rect 139222 428378 139306 428614
rect 139542 428378 174986 428614
rect 175222 428378 175306 428614
rect 175542 428378 210986 428614
rect 211222 428378 211306 428614
rect 211542 428378 246986 428614
rect 247222 428378 247306 428614
rect 247542 428378 282986 428614
rect 283222 428378 283306 428614
rect 283542 428378 318986 428614
rect 319222 428378 319306 428614
rect 319542 428378 354986 428614
rect 355222 428378 355306 428614
rect 355542 428378 390986 428614
rect 391222 428378 391306 428614
rect 391542 428378 426986 428614
rect 427222 428378 427306 428614
rect 427542 428378 462986 428614
rect 463222 428378 463306 428614
rect 463542 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect -8726 428294 592650 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 66986 428294
rect 67222 428058 67306 428294
rect 67542 428058 102986 428294
rect 103222 428058 103306 428294
rect 103542 428058 138986 428294
rect 139222 428058 139306 428294
rect 139542 428058 174986 428294
rect 175222 428058 175306 428294
rect 175542 428058 210986 428294
rect 211222 428058 211306 428294
rect 211542 428058 246986 428294
rect 247222 428058 247306 428294
rect 247542 428058 282986 428294
rect 283222 428058 283306 428294
rect 283542 428058 318986 428294
rect 319222 428058 319306 428294
rect 319542 428058 354986 428294
rect 355222 428058 355306 428294
rect 355542 428058 390986 428294
rect 391222 428058 391306 428294
rect 391542 428058 426986 428294
rect 427222 428058 427306 428294
rect 427542 428058 462986 428294
rect 463222 428058 463306 428294
rect 463542 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect -8726 428026 592650 428058
rect -6806 424894 590730 424926
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 99266 424894
rect 99502 424658 99586 424894
rect 99822 424658 135266 424894
rect 135502 424658 135586 424894
rect 135822 424658 171266 424894
rect 171502 424658 171586 424894
rect 171822 424658 207266 424894
rect 207502 424658 207586 424894
rect 207822 424658 243266 424894
rect 243502 424658 243586 424894
rect 243822 424658 279266 424894
rect 279502 424658 279586 424894
rect 279822 424658 315266 424894
rect 315502 424658 315586 424894
rect 315822 424658 351266 424894
rect 351502 424658 351586 424894
rect 351822 424658 387266 424894
rect 387502 424658 387586 424894
rect 387822 424658 423266 424894
rect 423502 424658 423586 424894
rect 423822 424658 459266 424894
rect 459502 424658 459586 424894
rect 459822 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect -6806 424574 590730 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 99266 424574
rect 99502 424338 99586 424574
rect 99822 424338 135266 424574
rect 135502 424338 135586 424574
rect 135822 424338 171266 424574
rect 171502 424338 171586 424574
rect 171822 424338 207266 424574
rect 207502 424338 207586 424574
rect 207822 424338 243266 424574
rect 243502 424338 243586 424574
rect 243822 424338 279266 424574
rect 279502 424338 279586 424574
rect 279822 424338 315266 424574
rect 315502 424338 315586 424574
rect 315822 424338 351266 424574
rect 351502 424338 351586 424574
rect 351822 424338 387266 424574
rect 387502 424338 387586 424574
rect 387822 424338 423266 424574
rect 423502 424338 423586 424574
rect 423822 424338 459266 424574
rect 459502 424338 459586 424574
rect 459822 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect -6806 424306 590730 424338
rect -4886 421174 588810 421206
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 95546 421174
rect 95782 420938 95866 421174
rect 96102 420938 131546 421174
rect 131782 420938 131866 421174
rect 132102 420938 167546 421174
rect 167782 420938 167866 421174
rect 168102 420938 203546 421174
rect 203782 420938 203866 421174
rect 204102 420938 239546 421174
rect 239782 420938 239866 421174
rect 240102 420938 275546 421174
rect 275782 420938 275866 421174
rect 276102 420938 311546 421174
rect 311782 420938 311866 421174
rect 312102 420938 347546 421174
rect 347782 420938 347866 421174
rect 348102 420938 383546 421174
rect 383782 420938 383866 421174
rect 384102 420938 419546 421174
rect 419782 420938 419866 421174
rect 420102 420938 455546 421174
rect 455782 420938 455866 421174
rect 456102 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect -4886 420854 588810 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 95546 420854
rect 95782 420618 95866 420854
rect 96102 420618 131546 420854
rect 131782 420618 131866 420854
rect 132102 420618 167546 420854
rect 167782 420618 167866 420854
rect 168102 420618 203546 420854
rect 203782 420618 203866 420854
rect 204102 420618 239546 420854
rect 239782 420618 239866 420854
rect 240102 420618 275546 420854
rect 275782 420618 275866 420854
rect 276102 420618 311546 420854
rect 311782 420618 311866 420854
rect 312102 420618 347546 420854
rect 347782 420618 347866 420854
rect 348102 420618 383546 420854
rect 383782 420618 383866 420854
rect 384102 420618 419546 420854
rect 419782 420618 419866 420854
rect 420102 420618 455546 420854
rect 455782 420618 455866 420854
rect 456102 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect -4886 420586 588810 420618
rect -2966 417454 586890 417486
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect -2966 417134 586890 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect -2966 416866 586890 416898
rect -8726 410614 592650 410646
rect -8726 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 84986 410614
rect 85222 410378 85306 410614
rect 85542 410378 120986 410614
rect 121222 410378 121306 410614
rect 121542 410378 156986 410614
rect 157222 410378 157306 410614
rect 157542 410378 192986 410614
rect 193222 410378 193306 410614
rect 193542 410378 228986 410614
rect 229222 410378 229306 410614
rect 229542 410378 264986 410614
rect 265222 410378 265306 410614
rect 265542 410378 300986 410614
rect 301222 410378 301306 410614
rect 301542 410378 336986 410614
rect 337222 410378 337306 410614
rect 337542 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 84986 410294
rect 85222 410058 85306 410294
rect 85542 410058 120986 410294
rect 121222 410058 121306 410294
rect 121542 410058 156986 410294
rect 157222 410058 157306 410294
rect 157542 410058 192986 410294
rect 193222 410058 193306 410294
rect 193542 410058 228986 410294
rect 229222 410058 229306 410294
rect 229542 410058 264986 410294
rect 265222 410058 265306 410294
rect 265542 410058 300986 410294
rect 301222 410058 301306 410294
rect 301542 410058 336986 410294
rect 337222 410058 337306 410294
rect 337542 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 592650 410294
rect -8726 410026 592650 410058
rect -6806 406894 590730 406926
rect -6806 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 81266 406894
rect 81502 406658 81586 406894
rect 81822 406658 117266 406894
rect 117502 406658 117586 406894
rect 117822 406658 153266 406894
rect 153502 406658 153586 406894
rect 153822 406658 189266 406894
rect 189502 406658 189586 406894
rect 189822 406658 225266 406894
rect 225502 406658 225586 406894
rect 225822 406658 261266 406894
rect 261502 406658 261586 406894
rect 261822 406658 297266 406894
rect 297502 406658 297586 406894
rect 297822 406658 333266 406894
rect 333502 406658 333586 406894
rect 333822 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 590730 406894
rect -6806 406574 590730 406658
rect -6806 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 81266 406574
rect 81502 406338 81586 406574
rect 81822 406338 117266 406574
rect 117502 406338 117586 406574
rect 117822 406338 153266 406574
rect 153502 406338 153586 406574
rect 153822 406338 189266 406574
rect 189502 406338 189586 406574
rect 189822 406338 225266 406574
rect 225502 406338 225586 406574
rect 225822 406338 261266 406574
rect 261502 406338 261586 406574
rect 261822 406338 297266 406574
rect 297502 406338 297586 406574
rect 297822 406338 333266 406574
rect 333502 406338 333586 406574
rect 333822 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 590730 406574
rect -6806 406306 590730 406338
rect -4886 403174 588810 403206
rect -4886 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 77546 403174
rect 77782 402938 77866 403174
rect 78102 402938 113546 403174
rect 113782 402938 113866 403174
rect 114102 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 185546 403174
rect 185782 402938 185866 403174
rect 186102 402938 221546 403174
rect 221782 402938 221866 403174
rect 222102 402938 257546 403174
rect 257782 402938 257866 403174
rect 258102 402938 293546 403174
rect 293782 402938 293866 403174
rect 294102 402938 329546 403174
rect 329782 402938 329866 403174
rect 330102 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 588810 403174
rect -4886 402854 588810 402938
rect -4886 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 77546 402854
rect 77782 402618 77866 402854
rect 78102 402618 113546 402854
rect 113782 402618 113866 402854
rect 114102 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 185546 402854
rect 185782 402618 185866 402854
rect 186102 402618 221546 402854
rect 221782 402618 221866 402854
rect 222102 402618 257546 402854
rect 257782 402618 257866 402854
rect 258102 402618 293546 402854
rect 293782 402618 293866 402854
rect 294102 402618 329546 402854
rect 329782 402618 329866 402854
rect 330102 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 588810 402854
rect -4886 402586 588810 402618
rect -2966 399454 586890 399486
rect -2966 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 586890 399454
rect -2966 399134 586890 399218
rect -2966 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 586890 399134
rect -2966 398866 586890 398898
rect -8726 392614 592650 392646
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 66986 392614
rect 67222 392378 67306 392614
rect 67542 392378 102986 392614
rect 103222 392378 103306 392614
rect 103542 392378 138986 392614
rect 139222 392378 139306 392614
rect 139542 392378 174986 392614
rect 175222 392378 175306 392614
rect 175542 392378 210986 392614
rect 211222 392378 211306 392614
rect 211542 392378 246986 392614
rect 247222 392378 247306 392614
rect 247542 392378 282986 392614
rect 283222 392378 283306 392614
rect 283542 392378 318986 392614
rect 319222 392378 319306 392614
rect 319542 392378 354986 392614
rect 355222 392378 355306 392614
rect 355542 392378 390986 392614
rect 391222 392378 391306 392614
rect 391542 392378 426986 392614
rect 427222 392378 427306 392614
rect 427542 392378 462986 392614
rect 463222 392378 463306 392614
rect 463542 392378 498986 392614
rect 499222 392378 499306 392614
rect 499542 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect -8726 392294 592650 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 66986 392294
rect 67222 392058 67306 392294
rect 67542 392058 102986 392294
rect 103222 392058 103306 392294
rect 103542 392058 138986 392294
rect 139222 392058 139306 392294
rect 139542 392058 174986 392294
rect 175222 392058 175306 392294
rect 175542 392058 210986 392294
rect 211222 392058 211306 392294
rect 211542 392058 246986 392294
rect 247222 392058 247306 392294
rect 247542 392058 282986 392294
rect 283222 392058 283306 392294
rect 283542 392058 318986 392294
rect 319222 392058 319306 392294
rect 319542 392058 354986 392294
rect 355222 392058 355306 392294
rect 355542 392058 390986 392294
rect 391222 392058 391306 392294
rect 391542 392058 426986 392294
rect 427222 392058 427306 392294
rect 427542 392058 462986 392294
rect 463222 392058 463306 392294
rect 463542 392058 498986 392294
rect 499222 392058 499306 392294
rect 499542 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect -8726 392026 592650 392058
rect -6806 388894 590730 388926
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 99266 388894
rect 99502 388658 99586 388894
rect 99822 388658 135266 388894
rect 135502 388658 135586 388894
rect 135822 388658 171266 388894
rect 171502 388658 171586 388894
rect 171822 388658 207266 388894
rect 207502 388658 207586 388894
rect 207822 388658 243266 388894
rect 243502 388658 243586 388894
rect 243822 388658 279266 388894
rect 279502 388658 279586 388894
rect 279822 388658 315266 388894
rect 315502 388658 315586 388894
rect 315822 388658 351266 388894
rect 351502 388658 351586 388894
rect 351822 388658 387266 388894
rect 387502 388658 387586 388894
rect 387822 388658 423266 388894
rect 423502 388658 423586 388894
rect 423822 388658 459266 388894
rect 459502 388658 459586 388894
rect 459822 388658 495266 388894
rect 495502 388658 495586 388894
rect 495822 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect -6806 388574 590730 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 99266 388574
rect 99502 388338 99586 388574
rect 99822 388338 135266 388574
rect 135502 388338 135586 388574
rect 135822 388338 171266 388574
rect 171502 388338 171586 388574
rect 171822 388338 207266 388574
rect 207502 388338 207586 388574
rect 207822 388338 243266 388574
rect 243502 388338 243586 388574
rect 243822 388338 279266 388574
rect 279502 388338 279586 388574
rect 279822 388338 315266 388574
rect 315502 388338 315586 388574
rect 315822 388338 351266 388574
rect 351502 388338 351586 388574
rect 351822 388338 387266 388574
rect 387502 388338 387586 388574
rect 387822 388338 423266 388574
rect 423502 388338 423586 388574
rect 423822 388338 459266 388574
rect 459502 388338 459586 388574
rect 459822 388338 495266 388574
rect 495502 388338 495586 388574
rect 495822 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect -6806 388306 590730 388338
rect -4886 385174 588810 385206
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 59546 385174
rect 59782 384938 59866 385174
rect 60102 384938 95546 385174
rect 95782 384938 95866 385174
rect 96102 384938 131546 385174
rect 131782 384938 131866 385174
rect 132102 384938 167546 385174
rect 167782 384938 167866 385174
rect 168102 384938 203546 385174
rect 203782 384938 203866 385174
rect 204102 384938 239546 385174
rect 239782 384938 239866 385174
rect 240102 384938 275546 385174
rect 275782 384938 275866 385174
rect 276102 384938 311546 385174
rect 311782 384938 311866 385174
rect 312102 384938 347546 385174
rect 347782 384938 347866 385174
rect 348102 384938 383546 385174
rect 383782 384938 383866 385174
rect 384102 384938 419546 385174
rect 419782 384938 419866 385174
rect 420102 384938 455546 385174
rect 455782 384938 455866 385174
rect 456102 384938 491546 385174
rect 491782 384938 491866 385174
rect 492102 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect -4886 384854 588810 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 59546 384854
rect 59782 384618 59866 384854
rect 60102 384618 95546 384854
rect 95782 384618 95866 384854
rect 96102 384618 131546 384854
rect 131782 384618 131866 384854
rect 132102 384618 167546 384854
rect 167782 384618 167866 384854
rect 168102 384618 203546 384854
rect 203782 384618 203866 384854
rect 204102 384618 239546 384854
rect 239782 384618 239866 384854
rect 240102 384618 275546 384854
rect 275782 384618 275866 384854
rect 276102 384618 311546 384854
rect 311782 384618 311866 384854
rect 312102 384618 347546 384854
rect 347782 384618 347866 384854
rect 348102 384618 383546 384854
rect 383782 384618 383866 384854
rect 384102 384618 419546 384854
rect 419782 384618 419866 384854
rect 420102 384618 455546 384854
rect 455782 384618 455866 384854
rect 456102 384618 491546 384854
rect 491782 384618 491866 384854
rect 492102 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect -4886 384586 588810 384618
rect -2966 381454 586890 381486
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect -2966 381134 586890 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect -2966 380866 586890 380898
rect -8726 374614 592650 374646
rect -8726 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 264986 374614
rect 265222 374378 265306 374614
rect 265542 374378 300986 374614
rect 301222 374378 301306 374614
rect 301542 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 264986 374294
rect 265222 374058 265306 374294
rect 265542 374058 300986 374294
rect 301222 374058 301306 374294
rect 301542 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 592650 374294
rect -8726 374026 592650 374058
rect -6806 370894 590730 370926
rect -6806 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 261266 370894
rect 261502 370658 261586 370894
rect 261822 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 590730 370894
rect -6806 370574 590730 370658
rect -6806 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 261266 370574
rect 261502 370338 261586 370574
rect 261822 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 590730 370574
rect -6806 370306 590730 370338
rect -4886 367174 588810 367206
rect -4886 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 257546 367174
rect 257782 366938 257866 367174
rect 258102 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 588810 367174
rect -4886 366854 588810 366938
rect -4886 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 257546 366854
rect 257782 366618 257866 366854
rect 258102 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 588810 366854
rect -4886 366586 588810 366618
rect -2966 363454 586890 363486
rect -2966 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 362285 363454
rect 362521 363218 364882 363454
rect 365118 363218 367479 363454
rect 367715 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 434285 363454
rect 434521 363218 436882 363454
rect 437118 363218 439479 363454
rect 439715 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 586890 363454
rect -2966 363134 586890 363218
rect -2966 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 362285 363134
rect 362521 362898 364882 363134
rect 365118 362898 367479 363134
rect 367715 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 434285 363134
rect 434521 362898 436882 363134
rect 437118 362898 439479 363134
rect 439715 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 586890 363134
rect -2966 362866 586890 362898
rect -8726 356614 592650 356646
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 102986 356614
rect 103222 356378 103306 356614
rect 103542 356378 138986 356614
rect 139222 356378 139306 356614
rect 139542 356378 174986 356614
rect 175222 356378 175306 356614
rect 175542 356378 210986 356614
rect 211222 356378 211306 356614
rect 211542 356378 246986 356614
rect 247222 356378 247306 356614
rect 247542 356378 282986 356614
rect 283222 356378 283306 356614
rect 283542 356378 318986 356614
rect 319222 356378 319306 356614
rect 319542 356378 354986 356614
rect 355222 356378 355306 356614
rect 355542 356378 390986 356614
rect 391222 356378 391306 356614
rect 391542 356378 426986 356614
rect 427222 356378 427306 356614
rect 427542 356378 462986 356614
rect 463222 356378 463306 356614
rect 463542 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect -8726 356294 592650 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 102986 356294
rect 103222 356058 103306 356294
rect 103542 356058 138986 356294
rect 139222 356058 139306 356294
rect 139542 356058 174986 356294
rect 175222 356058 175306 356294
rect 175542 356058 210986 356294
rect 211222 356058 211306 356294
rect 211542 356058 246986 356294
rect 247222 356058 247306 356294
rect 247542 356058 282986 356294
rect 283222 356058 283306 356294
rect 283542 356058 318986 356294
rect 319222 356058 319306 356294
rect 319542 356058 354986 356294
rect 355222 356058 355306 356294
rect 355542 356058 390986 356294
rect 391222 356058 391306 356294
rect 391542 356058 426986 356294
rect 427222 356058 427306 356294
rect 427542 356058 462986 356294
rect 463222 356058 463306 356294
rect 463542 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect -8726 356026 592650 356058
rect -6806 352894 590730 352926
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 63266 352894
rect 63502 352658 63586 352894
rect 63822 352658 99266 352894
rect 99502 352658 99586 352894
rect 99822 352658 135266 352894
rect 135502 352658 135586 352894
rect 135822 352658 171266 352894
rect 171502 352658 171586 352894
rect 171822 352658 207266 352894
rect 207502 352658 207586 352894
rect 207822 352658 243266 352894
rect 243502 352658 243586 352894
rect 243822 352658 279266 352894
rect 279502 352658 279586 352894
rect 279822 352658 315266 352894
rect 315502 352658 315586 352894
rect 315822 352658 351266 352894
rect 351502 352658 351586 352894
rect 351822 352658 387266 352894
rect 387502 352658 387586 352894
rect 387822 352658 423266 352894
rect 423502 352658 423586 352894
rect 423822 352658 459266 352894
rect 459502 352658 459586 352894
rect 459822 352658 495266 352894
rect 495502 352658 495586 352894
rect 495822 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect -6806 352574 590730 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 63266 352574
rect 63502 352338 63586 352574
rect 63822 352338 99266 352574
rect 99502 352338 99586 352574
rect 99822 352338 135266 352574
rect 135502 352338 135586 352574
rect 135822 352338 171266 352574
rect 171502 352338 171586 352574
rect 171822 352338 207266 352574
rect 207502 352338 207586 352574
rect 207822 352338 243266 352574
rect 243502 352338 243586 352574
rect 243822 352338 279266 352574
rect 279502 352338 279586 352574
rect 279822 352338 315266 352574
rect 315502 352338 315586 352574
rect 315822 352338 351266 352574
rect 351502 352338 351586 352574
rect 351822 352338 387266 352574
rect 387502 352338 387586 352574
rect 387822 352338 423266 352574
rect 423502 352338 423586 352574
rect 423822 352338 459266 352574
rect 459502 352338 459586 352574
rect 459822 352338 495266 352574
rect 495502 352338 495586 352574
rect 495822 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect -6806 352306 590730 352338
rect -4886 349174 588810 349206
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 59546 349174
rect 59782 348938 59866 349174
rect 60102 348938 95546 349174
rect 95782 348938 95866 349174
rect 96102 348938 131546 349174
rect 131782 348938 131866 349174
rect 132102 348938 167546 349174
rect 167782 348938 167866 349174
rect 168102 348938 203546 349174
rect 203782 348938 203866 349174
rect 204102 348938 239546 349174
rect 239782 348938 239866 349174
rect 240102 348938 275546 349174
rect 275782 348938 275866 349174
rect 276102 348938 311546 349174
rect 311782 348938 311866 349174
rect 312102 348938 347546 349174
rect 347782 348938 347866 349174
rect 348102 348938 383546 349174
rect 383782 348938 383866 349174
rect 384102 348938 419546 349174
rect 419782 348938 419866 349174
rect 420102 348938 455546 349174
rect 455782 348938 455866 349174
rect 456102 348938 491546 349174
rect 491782 348938 491866 349174
rect 492102 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect -4886 348854 588810 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 59546 348854
rect 59782 348618 59866 348854
rect 60102 348618 95546 348854
rect 95782 348618 95866 348854
rect 96102 348618 131546 348854
rect 131782 348618 131866 348854
rect 132102 348618 167546 348854
rect 167782 348618 167866 348854
rect 168102 348618 203546 348854
rect 203782 348618 203866 348854
rect 204102 348618 239546 348854
rect 239782 348618 239866 348854
rect 240102 348618 275546 348854
rect 275782 348618 275866 348854
rect 276102 348618 311546 348854
rect 311782 348618 311866 348854
rect 312102 348618 347546 348854
rect 347782 348618 347866 348854
rect 348102 348618 383546 348854
rect 383782 348618 383866 348854
rect 384102 348618 419546 348854
rect 419782 348618 419866 348854
rect 420102 348618 455546 348854
rect 455782 348618 455866 348854
rect 456102 348618 491546 348854
rect 491782 348618 491866 348854
rect 492102 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect -4886 348586 588810 348618
rect -2966 345454 586890 345486
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 363583 345454
rect 363819 345218 366180 345454
rect 366416 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 435583 345454
rect 435819 345218 438180 345454
rect 438416 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect -2966 345134 586890 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 363583 345134
rect 363819 344898 366180 345134
rect 366416 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 435583 345134
rect 435819 344898 438180 345134
rect 438416 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect -2966 344866 586890 344898
rect -8726 338614 592650 338646
rect -8726 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 84986 338614
rect 85222 338378 85306 338614
rect 85542 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 192986 338614
rect 193222 338378 193306 338614
rect 193542 338378 228986 338614
rect 229222 338378 229306 338614
rect 229542 338378 264986 338614
rect 265222 338378 265306 338614
rect 265542 338378 300986 338614
rect 301222 338378 301306 338614
rect 301542 338378 336986 338614
rect 337222 338378 337306 338614
rect 337542 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 84986 338294
rect 85222 338058 85306 338294
rect 85542 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 192986 338294
rect 193222 338058 193306 338294
rect 193542 338058 228986 338294
rect 229222 338058 229306 338294
rect 229542 338058 264986 338294
rect 265222 338058 265306 338294
rect 265542 338058 300986 338294
rect 301222 338058 301306 338294
rect 301542 338058 336986 338294
rect 337222 338058 337306 338294
rect 337542 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 592650 338294
rect -8726 338026 592650 338058
rect -6806 334894 590730 334926
rect -6806 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 189266 334894
rect 189502 334658 189586 334894
rect 189822 334658 225266 334894
rect 225502 334658 225586 334894
rect 225822 334658 261266 334894
rect 261502 334658 261586 334894
rect 261822 334658 297266 334894
rect 297502 334658 297586 334894
rect 297822 334658 333266 334894
rect 333502 334658 333586 334894
rect 333822 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 590730 334894
rect -6806 334574 590730 334658
rect -6806 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 189266 334574
rect 189502 334338 189586 334574
rect 189822 334338 225266 334574
rect 225502 334338 225586 334574
rect 225822 334338 261266 334574
rect 261502 334338 261586 334574
rect 261822 334338 297266 334574
rect 297502 334338 297586 334574
rect 297822 334338 333266 334574
rect 333502 334338 333586 334574
rect 333822 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 590730 334574
rect -6806 334306 590730 334338
rect -4886 331174 588810 331206
rect -4886 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 113546 331174
rect 113782 330938 113866 331174
rect 114102 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 221546 331174
rect 221782 330938 221866 331174
rect 222102 330938 257546 331174
rect 257782 330938 257866 331174
rect 258102 330938 293546 331174
rect 293782 330938 293866 331174
rect 294102 330938 329546 331174
rect 329782 330938 329866 331174
rect 330102 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 588810 331174
rect -4886 330854 588810 330938
rect -4886 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 113546 330854
rect 113782 330618 113866 330854
rect 114102 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 221546 330854
rect 221782 330618 221866 330854
rect 222102 330618 257546 330854
rect 257782 330618 257866 330854
rect 258102 330618 293546 330854
rect 293782 330618 293866 330854
rect 294102 330618 329546 330854
rect 329782 330618 329866 330854
rect 330102 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 588810 330854
rect -4886 330586 588810 330618
rect -2966 327454 586890 327486
rect -2966 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 586890 327454
rect -2966 327134 586890 327218
rect -2966 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 586890 327134
rect -2966 326866 586890 326898
rect -8726 320614 592650 320646
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 66986 320614
rect 67222 320378 67306 320614
rect 67542 320378 102986 320614
rect 103222 320378 103306 320614
rect 103542 320378 138986 320614
rect 139222 320378 139306 320614
rect 139542 320378 174986 320614
rect 175222 320378 175306 320614
rect 175542 320378 210986 320614
rect 211222 320378 211306 320614
rect 211542 320378 246986 320614
rect 247222 320378 247306 320614
rect 247542 320378 282986 320614
rect 283222 320378 283306 320614
rect 283542 320378 318986 320614
rect 319222 320378 319306 320614
rect 319542 320378 354986 320614
rect 355222 320378 355306 320614
rect 355542 320378 390986 320614
rect 391222 320378 391306 320614
rect 391542 320378 426986 320614
rect 427222 320378 427306 320614
rect 427542 320378 462986 320614
rect 463222 320378 463306 320614
rect 463542 320378 498986 320614
rect 499222 320378 499306 320614
rect 499542 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect -8726 320294 592650 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 66986 320294
rect 67222 320058 67306 320294
rect 67542 320058 102986 320294
rect 103222 320058 103306 320294
rect 103542 320058 138986 320294
rect 139222 320058 139306 320294
rect 139542 320058 174986 320294
rect 175222 320058 175306 320294
rect 175542 320058 210986 320294
rect 211222 320058 211306 320294
rect 211542 320058 246986 320294
rect 247222 320058 247306 320294
rect 247542 320058 282986 320294
rect 283222 320058 283306 320294
rect 283542 320058 318986 320294
rect 319222 320058 319306 320294
rect 319542 320058 354986 320294
rect 355222 320058 355306 320294
rect 355542 320058 390986 320294
rect 391222 320058 391306 320294
rect 391542 320058 426986 320294
rect 427222 320058 427306 320294
rect 427542 320058 462986 320294
rect 463222 320058 463306 320294
rect 463542 320058 498986 320294
rect 499222 320058 499306 320294
rect 499542 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect -8726 320026 592650 320058
rect -6806 316894 590730 316926
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 63266 316894
rect 63502 316658 63586 316894
rect 63822 316658 99266 316894
rect 99502 316658 99586 316894
rect 99822 316658 135266 316894
rect 135502 316658 135586 316894
rect 135822 316658 171266 316894
rect 171502 316658 171586 316894
rect 171822 316658 207266 316894
rect 207502 316658 207586 316894
rect 207822 316658 243266 316894
rect 243502 316658 243586 316894
rect 243822 316658 279266 316894
rect 279502 316658 279586 316894
rect 279822 316658 315266 316894
rect 315502 316658 315586 316894
rect 315822 316658 351266 316894
rect 351502 316658 351586 316894
rect 351822 316658 387266 316894
rect 387502 316658 387586 316894
rect 387822 316658 423266 316894
rect 423502 316658 423586 316894
rect 423822 316658 459266 316894
rect 459502 316658 459586 316894
rect 459822 316658 495266 316894
rect 495502 316658 495586 316894
rect 495822 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect -6806 316574 590730 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 63266 316574
rect 63502 316338 63586 316574
rect 63822 316338 99266 316574
rect 99502 316338 99586 316574
rect 99822 316338 135266 316574
rect 135502 316338 135586 316574
rect 135822 316338 171266 316574
rect 171502 316338 171586 316574
rect 171822 316338 207266 316574
rect 207502 316338 207586 316574
rect 207822 316338 243266 316574
rect 243502 316338 243586 316574
rect 243822 316338 279266 316574
rect 279502 316338 279586 316574
rect 279822 316338 315266 316574
rect 315502 316338 315586 316574
rect 315822 316338 351266 316574
rect 351502 316338 351586 316574
rect 351822 316338 387266 316574
rect 387502 316338 387586 316574
rect 387822 316338 423266 316574
rect 423502 316338 423586 316574
rect 423822 316338 459266 316574
rect 459502 316338 459586 316574
rect 459822 316338 495266 316574
rect 495502 316338 495586 316574
rect 495822 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect -6806 316306 590730 316338
rect -4886 313174 588810 313206
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 59546 313174
rect 59782 312938 59866 313174
rect 60102 312938 95546 313174
rect 95782 312938 95866 313174
rect 96102 312938 131546 313174
rect 131782 312938 131866 313174
rect 132102 312938 167546 313174
rect 167782 312938 167866 313174
rect 168102 312938 203546 313174
rect 203782 312938 203866 313174
rect 204102 312938 239546 313174
rect 239782 312938 239866 313174
rect 240102 312938 275546 313174
rect 275782 312938 275866 313174
rect 276102 312938 311546 313174
rect 311782 312938 311866 313174
rect 312102 312938 347546 313174
rect 347782 312938 347866 313174
rect 348102 312938 383546 313174
rect 383782 312938 383866 313174
rect 384102 312938 419546 313174
rect 419782 312938 419866 313174
rect 420102 312938 455546 313174
rect 455782 312938 455866 313174
rect 456102 312938 491546 313174
rect 491782 312938 491866 313174
rect 492102 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect -4886 312854 588810 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 59546 312854
rect 59782 312618 59866 312854
rect 60102 312618 95546 312854
rect 95782 312618 95866 312854
rect 96102 312618 131546 312854
rect 131782 312618 131866 312854
rect 132102 312618 167546 312854
rect 167782 312618 167866 312854
rect 168102 312618 203546 312854
rect 203782 312618 203866 312854
rect 204102 312618 239546 312854
rect 239782 312618 239866 312854
rect 240102 312618 275546 312854
rect 275782 312618 275866 312854
rect 276102 312618 311546 312854
rect 311782 312618 311866 312854
rect 312102 312618 347546 312854
rect 347782 312618 347866 312854
rect 348102 312618 383546 312854
rect 383782 312618 383866 312854
rect 384102 312618 419546 312854
rect 419782 312618 419866 312854
rect 420102 312618 455546 312854
rect 455782 312618 455866 312854
rect 456102 312618 491546 312854
rect 491782 312618 491866 312854
rect 492102 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect -4886 312586 588810 312618
rect -2966 309454 586890 309486
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect -2966 309134 586890 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect -2966 308866 586890 308898
rect -8726 302614 592650 302646
rect -8726 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 84986 302614
rect 85222 302378 85306 302614
rect 85542 302378 120986 302614
rect 121222 302378 121306 302614
rect 121542 302378 156986 302614
rect 157222 302378 157306 302614
rect 157542 302378 192986 302614
rect 193222 302378 193306 302614
rect 193542 302378 228986 302614
rect 229222 302378 229306 302614
rect 229542 302378 264986 302614
rect 265222 302378 265306 302614
rect 265542 302378 300986 302614
rect 301222 302378 301306 302614
rect 301542 302378 336986 302614
rect 337222 302378 337306 302614
rect 337542 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 84986 302294
rect 85222 302058 85306 302294
rect 85542 302058 120986 302294
rect 121222 302058 121306 302294
rect 121542 302058 156986 302294
rect 157222 302058 157306 302294
rect 157542 302058 192986 302294
rect 193222 302058 193306 302294
rect 193542 302058 228986 302294
rect 229222 302058 229306 302294
rect 229542 302058 264986 302294
rect 265222 302058 265306 302294
rect 265542 302058 300986 302294
rect 301222 302058 301306 302294
rect 301542 302058 336986 302294
rect 337222 302058 337306 302294
rect 337542 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 592650 302294
rect -8726 302026 592650 302058
rect -6806 298894 590730 298926
rect -6806 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 81266 298894
rect 81502 298658 81586 298894
rect 81822 298658 117266 298894
rect 117502 298658 117586 298894
rect 117822 298658 153266 298894
rect 153502 298658 153586 298894
rect 153822 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 333266 298894
rect 333502 298658 333586 298894
rect 333822 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 590730 298894
rect -6806 298574 590730 298658
rect -6806 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 81266 298574
rect 81502 298338 81586 298574
rect 81822 298338 117266 298574
rect 117502 298338 117586 298574
rect 117822 298338 153266 298574
rect 153502 298338 153586 298574
rect 153822 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 333266 298574
rect 333502 298338 333586 298574
rect 333822 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 590730 298574
rect -6806 298306 590730 298338
rect -4886 295174 588810 295206
rect -4886 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 77546 295174
rect 77782 294938 77866 295174
rect 78102 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 149546 295174
rect 149782 294938 149866 295174
rect 150102 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 329546 295174
rect 329782 294938 329866 295174
rect 330102 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 588810 295174
rect -4886 294854 588810 294938
rect -4886 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 77546 294854
rect 77782 294618 77866 294854
rect 78102 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 149546 294854
rect 149782 294618 149866 294854
rect 150102 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 329546 294854
rect 329782 294618 329866 294854
rect 330102 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 588810 294854
rect -4886 294586 588810 294618
rect -2966 291454 586890 291486
rect -2966 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 204250 291454
rect 204486 291218 234970 291454
rect 235206 291218 265690 291454
rect 265926 291218 296410 291454
rect 296646 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 362285 291454
rect 362521 291218 364882 291454
rect 365118 291218 367479 291454
rect 367715 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 434285 291454
rect 434521 291218 436882 291454
rect 437118 291218 439479 291454
rect 439715 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 586890 291454
rect -2966 291134 586890 291218
rect -2966 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 204250 291134
rect 204486 290898 234970 291134
rect 235206 290898 265690 291134
rect 265926 290898 296410 291134
rect 296646 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 362285 291134
rect 362521 290898 364882 291134
rect 365118 290898 367479 291134
rect 367715 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 434285 291134
rect 434521 290898 436882 291134
rect 437118 290898 439479 291134
rect 439715 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 586890 291134
rect -2966 290866 586890 290898
rect -8726 284614 592650 284646
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 66986 284614
rect 67222 284378 67306 284614
rect 67542 284378 102986 284614
rect 103222 284378 103306 284614
rect 103542 284378 138986 284614
rect 139222 284378 139306 284614
rect 139542 284378 174986 284614
rect 175222 284378 175306 284614
rect 175542 284378 318986 284614
rect 319222 284378 319306 284614
rect 319542 284378 354986 284614
rect 355222 284378 355306 284614
rect 355542 284378 390986 284614
rect 391222 284378 391306 284614
rect 391542 284378 426986 284614
rect 427222 284378 427306 284614
rect 427542 284378 462986 284614
rect 463222 284378 463306 284614
rect 463542 284378 498986 284614
rect 499222 284378 499306 284614
rect 499542 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect -8726 284294 592650 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 66986 284294
rect 67222 284058 67306 284294
rect 67542 284058 102986 284294
rect 103222 284058 103306 284294
rect 103542 284058 138986 284294
rect 139222 284058 139306 284294
rect 139542 284058 174986 284294
rect 175222 284058 175306 284294
rect 175542 284058 318986 284294
rect 319222 284058 319306 284294
rect 319542 284058 354986 284294
rect 355222 284058 355306 284294
rect 355542 284058 390986 284294
rect 391222 284058 391306 284294
rect 391542 284058 426986 284294
rect 427222 284058 427306 284294
rect 427542 284058 462986 284294
rect 463222 284058 463306 284294
rect 463542 284058 498986 284294
rect 499222 284058 499306 284294
rect 499542 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect -8726 284026 592650 284058
rect -6806 280894 590730 280926
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 63266 280894
rect 63502 280658 63586 280894
rect 63822 280658 99266 280894
rect 99502 280658 99586 280894
rect 99822 280658 135266 280894
rect 135502 280658 135586 280894
rect 135822 280658 171266 280894
rect 171502 280658 171586 280894
rect 171822 280658 315266 280894
rect 315502 280658 315586 280894
rect 315822 280658 351266 280894
rect 351502 280658 351586 280894
rect 351822 280658 387266 280894
rect 387502 280658 387586 280894
rect 387822 280658 423266 280894
rect 423502 280658 423586 280894
rect 423822 280658 459266 280894
rect 459502 280658 459586 280894
rect 459822 280658 495266 280894
rect 495502 280658 495586 280894
rect 495822 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect -6806 280574 590730 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 63266 280574
rect 63502 280338 63586 280574
rect 63822 280338 99266 280574
rect 99502 280338 99586 280574
rect 99822 280338 135266 280574
rect 135502 280338 135586 280574
rect 135822 280338 171266 280574
rect 171502 280338 171586 280574
rect 171822 280338 315266 280574
rect 315502 280338 315586 280574
rect 315822 280338 351266 280574
rect 351502 280338 351586 280574
rect 351822 280338 387266 280574
rect 387502 280338 387586 280574
rect 387822 280338 423266 280574
rect 423502 280338 423586 280574
rect 423822 280338 459266 280574
rect 459502 280338 459586 280574
rect 459822 280338 495266 280574
rect 495502 280338 495586 280574
rect 495822 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect -6806 280306 590730 280338
rect -4886 277174 588810 277206
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 59546 277174
rect 59782 276938 59866 277174
rect 60102 276938 95546 277174
rect 95782 276938 95866 277174
rect 96102 276938 131546 277174
rect 131782 276938 131866 277174
rect 132102 276938 167546 277174
rect 167782 276938 167866 277174
rect 168102 276938 311546 277174
rect 311782 276938 311866 277174
rect 312102 276938 347546 277174
rect 347782 276938 347866 277174
rect 348102 276938 383546 277174
rect 383782 276938 383866 277174
rect 384102 276938 419546 277174
rect 419782 276938 419866 277174
rect 420102 276938 455546 277174
rect 455782 276938 455866 277174
rect 456102 276938 491546 277174
rect 491782 276938 491866 277174
rect 492102 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect -4886 276854 588810 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 59546 276854
rect 59782 276618 59866 276854
rect 60102 276618 95546 276854
rect 95782 276618 95866 276854
rect 96102 276618 131546 276854
rect 131782 276618 131866 276854
rect 132102 276618 167546 276854
rect 167782 276618 167866 276854
rect 168102 276618 311546 276854
rect 311782 276618 311866 276854
rect 312102 276618 347546 276854
rect 347782 276618 347866 276854
rect 348102 276618 383546 276854
rect 383782 276618 383866 276854
rect 384102 276618 419546 276854
rect 419782 276618 419866 276854
rect 420102 276618 455546 276854
rect 455782 276618 455866 276854
rect 456102 276618 491546 276854
rect 491782 276618 491866 276854
rect 492102 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect -4886 276586 588810 276618
rect -2966 273454 586890 273486
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 219610 273454
rect 219846 273218 250330 273454
rect 250566 273218 281050 273454
rect 281286 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 363583 273454
rect 363819 273218 366180 273454
rect 366416 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 435583 273454
rect 435819 273218 438180 273454
rect 438416 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect -2966 273134 586890 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 219610 273134
rect 219846 272898 250330 273134
rect 250566 272898 281050 273134
rect 281286 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 363583 273134
rect 363819 272898 366180 273134
rect 366416 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 435583 273134
rect 435819 272898 438180 273134
rect 438416 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect -2966 272866 586890 272898
rect -8726 266614 592650 266646
rect -8726 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 84986 266614
rect 85222 266378 85306 266614
rect 85542 266378 120986 266614
rect 121222 266378 121306 266614
rect 121542 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 192986 266614
rect 193222 266378 193306 266614
rect 193542 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 84986 266294
rect 85222 266058 85306 266294
rect 85542 266058 120986 266294
rect 121222 266058 121306 266294
rect 121542 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 192986 266294
rect 193222 266058 193306 266294
rect 193542 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 592650 266294
rect -8726 266026 592650 266058
rect -6806 262894 590730 262926
rect -6806 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 81266 262894
rect 81502 262658 81586 262894
rect 81822 262658 117266 262894
rect 117502 262658 117586 262894
rect 117822 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 590730 262894
rect -6806 262574 590730 262658
rect -6806 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 81266 262574
rect 81502 262338 81586 262574
rect 81822 262338 117266 262574
rect 117502 262338 117586 262574
rect 117822 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 590730 262574
rect -6806 262306 590730 262338
rect -4886 259174 588810 259206
rect -4886 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 77546 259174
rect 77782 258938 77866 259174
rect 78102 258938 113546 259174
rect 113782 258938 113866 259174
rect 114102 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 588810 259174
rect -4886 258854 588810 258938
rect -4886 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 77546 258854
rect 77782 258618 77866 258854
rect 78102 258618 113546 258854
rect 113782 258618 113866 258854
rect 114102 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 588810 258854
rect -4886 258586 588810 258618
rect -2966 255454 586890 255486
rect -2966 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 204250 255454
rect 204486 255218 234970 255454
rect 235206 255218 265690 255454
rect 265926 255218 296410 255454
rect 296646 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 586890 255454
rect -2966 255134 586890 255218
rect -2966 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 204250 255134
rect 204486 254898 234970 255134
rect 235206 254898 265690 255134
rect 265926 254898 296410 255134
rect 296646 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 586890 255134
rect -2966 254866 586890 254898
rect -8726 248614 592650 248646
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 66986 248614
rect 67222 248378 67306 248614
rect 67542 248378 102986 248614
rect 103222 248378 103306 248614
rect 103542 248378 138986 248614
rect 139222 248378 139306 248614
rect 139542 248378 174986 248614
rect 175222 248378 175306 248614
rect 175542 248378 318986 248614
rect 319222 248378 319306 248614
rect 319542 248378 354986 248614
rect 355222 248378 355306 248614
rect 355542 248378 390986 248614
rect 391222 248378 391306 248614
rect 391542 248378 426986 248614
rect 427222 248378 427306 248614
rect 427542 248378 462986 248614
rect 463222 248378 463306 248614
rect 463542 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect -8726 248294 592650 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 66986 248294
rect 67222 248058 67306 248294
rect 67542 248058 102986 248294
rect 103222 248058 103306 248294
rect 103542 248058 138986 248294
rect 139222 248058 139306 248294
rect 139542 248058 174986 248294
rect 175222 248058 175306 248294
rect 175542 248058 318986 248294
rect 319222 248058 319306 248294
rect 319542 248058 354986 248294
rect 355222 248058 355306 248294
rect 355542 248058 390986 248294
rect 391222 248058 391306 248294
rect 391542 248058 426986 248294
rect 427222 248058 427306 248294
rect 427542 248058 462986 248294
rect 463222 248058 463306 248294
rect 463542 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect -8726 248026 592650 248058
rect -6806 244894 590730 244926
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 99266 244894
rect 99502 244658 99586 244894
rect 99822 244658 135266 244894
rect 135502 244658 135586 244894
rect 135822 244658 171266 244894
rect 171502 244658 171586 244894
rect 171822 244658 315266 244894
rect 315502 244658 315586 244894
rect 315822 244658 351266 244894
rect 351502 244658 351586 244894
rect 351822 244658 387266 244894
rect 387502 244658 387586 244894
rect 387822 244658 423266 244894
rect 423502 244658 423586 244894
rect 423822 244658 459266 244894
rect 459502 244658 459586 244894
rect 459822 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect -6806 244574 590730 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 99266 244574
rect 99502 244338 99586 244574
rect 99822 244338 135266 244574
rect 135502 244338 135586 244574
rect 135822 244338 171266 244574
rect 171502 244338 171586 244574
rect 171822 244338 315266 244574
rect 315502 244338 315586 244574
rect 315822 244338 351266 244574
rect 351502 244338 351586 244574
rect 351822 244338 387266 244574
rect 387502 244338 387586 244574
rect 387822 244338 423266 244574
rect 423502 244338 423586 244574
rect 423822 244338 459266 244574
rect 459502 244338 459586 244574
rect 459822 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect -6806 244306 590730 244338
rect -4886 241174 588810 241206
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 95546 241174
rect 95782 240938 95866 241174
rect 96102 240938 131546 241174
rect 131782 240938 131866 241174
rect 132102 240938 167546 241174
rect 167782 240938 167866 241174
rect 168102 240938 311546 241174
rect 311782 240938 311866 241174
rect 312102 240938 347546 241174
rect 347782 240938 347866 241174
rect 348102 240938 383546 241174
rect 383782 240938 383866 241174
rect 384102 240938 419546 241174
rect 419782 240938 419866 241174
rect 420102 240938 455546 241174
rect 455782 240938 455866 241174
rect 456102 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect -4886 240854 588810 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 95546 240854
rect 95782 240618 95866 240854
rect 96102 240618 131546 240854
rect 131782 240618 131866 240854
rect 132102 240618 167546 240854
rect 167782 240618 167866 240854
rect 168102 240618 311546 240854
rect 311782 240618 311866 240854
rect 312102 240618 347546 240854
rect 347782 240618 347866 240854
rect 348102 240618 383546 240854
rect 383782 240618 383866 240854
rect 384102 240618 419546 240854
rect 419782 240618 419866 240854
rect 420102 240618 455546 240854
rect 455782 240618 455866 240854
rect 456102 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect -4886 240586 588810 240618
rect -2966 237454 586890 237486
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 219610 237454
rect 219846 237218 250330 237454
rect 250566 237218 281050 237454
rect 281286 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect -2966 237134 586890 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 219610 237134
rect 219846 236898 250330 237134
rect 250566 236898 281050 237134
rect 281286 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect -2966 236866 586890 236898
rect -8726 230614 592650 230646
rect -8726 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 156986 230614
rect 157222 230378 157306 230614
rect 157542 230378 192986 230614
rect 193222 230378 193306 230614
rect 193542 230378 336986 230614
rect 337222 230378 337306 230614
rect 337542 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 156986 230294
rect 157222 230058 157306 230294
rect 157542 230058 192986 230294
rect 193222 230058 193306 230294
rect 193542 230058 336986 230294
rect 337222 230058 337306 230294
rect 337542 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 592650 230294
rect -8726 230026 592650 230058
rect -6806 226894 590730 226926
rect -6806 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 81266 226894
rect 81502 226658 81586 226894
rect 81822 226658 117266 226894
rect 117502 226658 117586 226894
rect 117822 226658 153266 226894
rect 153502 226658 153586 226894
rect 153822 226658 189266 226894
rect 189502 226658 189586 226894
rect 189822 226658 333266 226894
rect 333502 226658 333586 226894
rect 333822 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 590730 226894
rect -6806 226574 590730 226658
rect -6806 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 81266 226574
rect 81502 226338 81586 226574
rect 81822 226338 117266 226574
rect 117502 226338 117586 226574
rect 117822 226338 153266 226574
rect 153502 226338 153586 226574
rect 153822 226338 189266 226574
rect 189502 226338 189586 226574
rect 189822 226338 333266 226574
rect 333502 226338 333586 226574
rect 333822 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 590730 226574
rect -6806 226306 590730 226338
rect -4886 223174 588810 223206
rect -4886 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 113546 223174
rect 113782 222938 113866 223174
rect 114102 222938 149546 223174
rect 149782 222938 149866 223174
rect 150102 222938 185546 223174
rect 185782 222938 185866 223174
rect 186102 222938 329546 223174
rect 329782 222938 329866 223174
rect 330102 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 588810 223174
rect -4886 222854 588810 222938
rect -4886 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 113546 222854
rect 113782 222618 113866 222854
rect 114102 222618 149546 222854
rect 149782 222618 149866 222854
rect 150102 222618 185546 222854
rect 185782 222618 185866 222854
rect 186102 222618 329546 222854
rect 329782 222618 329866 222854
rect 330102 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 588810 222854
rect -4886 222586 588810 222618
rect -2966 219454 586890 219486
rect -2966 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 204250 219454
rect 204486 219218 234970 219454
rect 235206 219218 265690 219454
rect 265926 219218 296410 219454
rect 296646 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 362285 219454
rect 362521 219218 364882 219454
rect 365118 219218 367479 219454
rect 367715 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 434285 219454
rect 434521 219218 436882 219454
rect 437118 219218 439479 219454
rect 439715 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 586890 219454
rect -2966 219134 586890 219218
rect -2966 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 204250 219134
rect 204486 218898 234970 219134
rect 235206 218898 265690 219134
rect 265926 218898 296410 219134
rect 296646 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 362285 219134
rect 362521 218898 364882 219134
rect 365118 218898 367479 219134
rect 367715 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 434285 219134
rect 434521 218898 436882 219134
rect 437118 218898 439479 219134
rect 439715 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 586890 219134
rect -2966 218866 586890 218898
rect -8726 212614 592650 212646
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 66986 212614
rect 67222 212378 67306 212614
rect 67542 212378 102986 212614
rect 103222 212378 103306 212614
rect 103542 212378 138986 212614
rect 139222 212378 139306 212614
rect 139542 212378 174986 212614
rect 175222 212378 175306 212614
rect 175542 212378 318986 212614
rect 319222 212378 319306 212614
rect 319542 212378 354986 212614
rect 355222 212378 355306 212614
rect 355542 212378 390986 212614
rect 391222 212378 391306 212614
rect 391542 212378 426986 212614
rect 427222 212378 427306 212614
rect 427542 212378 462986 212614
rect 463222 212378 463306 212614
rect 463542 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect -8726 212294 592650 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 66986 212294
rect 67222 212058 67306 212294
rect 67542 212058 102986 212294
rect 103222 212058 103306 212294
rect 103542 212058 138986 212294
rect 139222 212058 139306 212294
rect 139542 212058 174986 212294
rect 175222 212058 175306 212294
rect 175542 212058 318986 212294
rect 319222 212058 319306 212294
rect 319542 212058 354986 212294
rect 355222 212058 355306 212294
rect 355542 212058 390986 212294
rect 391222 212058 391306 212294
rect 391542 212058 426986 212294
rect 427222 212058 427306 212294
rect 427542 212058 462986 212294
rect 463222 212058 463306 212294
rect 463542 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect -8726 212026 592650 212058
rect -6806 208894 590730 208926
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 63266 208894
rect 63502 208658 63586 208894
rect 63822 208658 99266 208894
rect 99502 208658 99586 208894
rect 99822 208658 135266 208894
rect 135502 208658 135586 208894
rect 135822 208658 171266 208894
rect 171502 208658 171586 208894
rect 171822 208658 315266 208894
rect 315502 208658 315586 208894
rect 315822 208658 351266 208894
rect 351502 208658 351586 208894
rect 351822 208658 387266 208894
rect 387502 208658 387586 208894
rect 387822 208658 423266 208894
rect 423502 208658 423586 208894
rect 423822 208658 459266 208894
rect 459502 208658 459586 208894
rect 459822 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect -6806 208574 590730 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 63266 208574
rect 63502 208338 63586 208574
rect 63822 208338 99266 208574
rect 99502 208338 99586 208574
rect 99822 208338 135266 208574
rect 135502 208338 135586 208574
rect 135822 208338 171266 208574
rect 171502 208338 171586 208574
rect 171822 208338 315266 208574
rect 315502 208338 315586 208574
rect 315822 208338 351266 208574
rect 351502 208338 351586 208574
rect 351822 208338 387266 208574
rect 387502 208338 387586 208574
rect 387822 208338 423266 208574
rect 423502 208338 423586 208574
rect 423822 208338 459266 208574
rect 459502 208338 459586 208574
rect 459822 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect -6806 208306 590730 208338
rect -4886 205174 588810 205206
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 59546 205174
rect 59782 204938 59866 205174
rect 60102 204938 95546 205174
rect 95782 204938 95866 205174
rect 96102 204938 131546 205174
rect 131782 204938 131866 205174
rect 132102 204938 167546 205174
rect 167782 204938 167866 205174
rect 168102 204938 311546 205174
rect 311782 204938 311866 205174
rect 312102 204938 347546 205174
rect 347782 204938 347866 205174
rect 348102 204938 383546 205174
rect 383782 204938 383866 205174
rect 384102 204938 419546 205174
rect 419782 204938 419866 205174
rect 420102 204938 455546 205174
rect 455782 204938 455866 205174
rect 456102 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect -4886 204854 588810 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 59546 204854
rect 59782 204618 59866 204854
rect 60102 204618 95546 204854
rect 95782 204618 95866 204854
rect 96102 204618 131546 204854
rect 131782 204618 131866 204854
rect 132102 204618 167546 204854
rect 167782 204618 167866 204854
rect 168102 204618 311546 204854
rect 311782 204618 311866 204854
rect 312102 204618 347546 204854
rect 347782 204618 347866 204854
rect 348102 204618 383546 204854
rect 383782 204618 383866 204854
rect 384102 204618 419546 204854
rect 419782 204618 419866 204854
rect 420102 204618 455546 204854
rect 455782 204618 455866 204854
rect 456102 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect -4886 204586 588810 204618
rect -2966 201454 586890 201486
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 219610 201454
rect 219846 201218 250330 201454
rect 250566 201218 281050 201454
rect 281286 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 363583 201454
rect 363819 201218 366180 201454
rect 366416 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 435583 201454
rect 435819 201218 438180 201454
rect 438416 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect -2966 201134 586890 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 219610 201134
rect 219846 200898 250330 201134
rect 250566 200898 281050 201134
rect 281286 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 363583 201134
rect 363819 200898 366180 201134
rect 366416 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 435583 201134
rect 435819 200898 438180 201134
rect 438416 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect -2966 200866 586890 200898
rect -8726 194614 592650 194646
rect -8726 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 120986 194614
rect 121222 194378 121306 194614
rect 121542 194378 156986 194614
rect 157222 194378 157306 194614
rect 157542 194378 192986 194614
rect 193222 194378 193306 194614
rect 193542 194378 336986 194614
rect 337222 194378 337306 194614
rect 337542 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 120986 194294
rect 121222 194058 121306 194294
rect 121542 194058 156986 194294
rect 157222 194058 157306 194294
rect 157542 194058 192986 194294
rect 193222 194058 193306 194294
rect 193542 194058 336986 194294
rect 337222 194058 337306 194294
rect 337542 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 592650 194294
rect -8726 194026 592650 194058
rect -6806 190894 590730 190926
rect -6806 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 117266 190894
rect 117502 190658 117586 190894
rect 117822 190658 153266 190894
rect 153502 190658 153586 190894
rect 153822 190658 189266 190894
rect 189502 190658 189586 190894
rect 189822 190658 333266 190894
rect 333502 190658 333586 190894
rect 333822 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 590730 190894
rect -6806 190574 590730 190658
rect -6806 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 117266 190574
rect 117502 190338 117586 190574
rect 117822 190338 153266 190574
rect 153502 190338 153586 190574
rect 153822 190338 189266 190574
rect 189502 190338 189586 190574
rect 189822 190338 333266 190574
rect 333502 190338 333586 190574
rect 333822 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 590730 190574
rect -6806 190306 590730 190338
rect -4886 187174 588810 187206
rect -4886 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 149546 187174
rect 149782 186938 149866 187174
rect 150102 186938 185546 187174
rect 185782 186938 185866 187174
rect 186102 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 588810 187174
rect -4886 186854 588810 186938
rect -4886 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 149546 186854
rect 149782 186618 149866 186854
rect 150102 186618 185546 186854
rect 185782 186618 185866 186854
rect 186102 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 588810 186854
rect -4886 186586 588810 186618
rect -2966 183454 586890 183486
rect -2966 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 162285 183454
rect 162521 183218 164882 183454
rect 165118 183218 167479 183454
rect 167715 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 204250 183454
rect 204486 183218 234970 183454
rect 235206 183218 265690 183454
rect 265926 183218 296410 183454
rect 296646 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 586890 183454
rect -2966 183134 586890 183218
rect -2966 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 162285 183134
rect 162521 182898 164882 183134
rect 165118 182898 167479 183134
rect 167715 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 204250 183134
rect 204486 182898 234970 183134
rect 235206 182898 265690 183134
rect 265926 182898 296410 183134
rect 296646 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 586890 183134
rect -2966 182866 586890 182898
rect -8726 176614 592650 176646
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 66986 176614
rect 67222 176378 67306 176614
rect 67542 176378 102986 176614
rect 103222 176378 103306 176614
rect 103542 176378 138986 176614
rect 139222 176378 139306 176614
rect 139542 176378 174986 176614
rect 175222 176378 175306 176614
rect 175542 176378 318986 176614
rect 319222 176378 319306 176614
rect 319542 176378 354986 176614
rect 355222 176378 355306 176614
rect 355542 176378 390986 176614
rect 391222 176378 391306 176614
rect 391542 176378 426986 176614
rect 427222 176378 427306 176614
rect 427542 176378 462986 176614
rect 463222 176378 463306 176614
rect 463542 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect -8726 176294 592650 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 66986 176294
rect 67222 176058 67306 176294
rect 67542 176058 102986 176294
rect 103222 176058 103306 176294
rect 103542 176058 138986 176294
rect 139222 176058 139306 176294
rect 139542 176058 174986 176294
rect 175222 176058 175306 176294
rect 175542 176058 318986 176294
rect 319222 176058 319306 176294
rect 319542 176058 354986 176294
rect 355222 176058 355306 176294
rect 355542 176058 390986 176294
rect 391222 176058 391306 176294
rect 391542 176058 426986 176294
rect 427222 176058 427306 176294
rect 427542 176058 462986 176294
rect 463222 176058 463306 176294
rect 463542 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect -8726 176026 592650 176058
rect -6806 172894 590730 172926
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 63266 172894
rect 63502 172658 63586 172894
rect 63822 172658 99266 172894
rect 99502 172658 99586 172894
rect 99822 172658 135266 172894
rect 135502 172658 135586 172894
rect 135822 172658 315266 172894
rect 315502 172658 315586 172894
rect 315822 172658 351266 172894
rect 351502 172658 351586 172894
rect 351822 172658 387266 172894
rect 387502 172658 387586 172894
rect 387822 172658 423266 172894
rect 423502 172658 423586 172894
rect 423822 172658 459266 172894
rect 459502 172658 459586 172894
rect 459822 172658 495266 172894
rect 495502 172658 495586 172894
rect 495822 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect -6806 172574 590730 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 63266 172574
rect 63502 172338 63586 172574
rect 63822 172338 99266 172574
rect 99502 172338 99586 172574
rect 99822 172338 135266 172574
rect 135502 172338 135586 172574
rect 135822 172338 315266 172574
rect 315502 172338 315586 172574
rect 315822 172338 351266 172574
rect 351502 172338 351586 172574
rect 351822 172338 387266 172574
rect 387502 172338 387586 172574
rect 387822 172338 423266 172574
rect 423502 172338 423586 172574
rect 423822 172338 459266 172574
rect 459502 172338 459586 172574
rect 459822 172338 495266 172574
rect 495502 172338 495586 172574
rect 495822 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect -6806 172306 590730 172338
rect -4886 169174 588810 169206
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 59546 169174
rect 59782 168938 59866 169174
rect 60102 168938 95546 169174
rect 95782 168938 95866 169174
rect 96102 168938 131546 169174
rect 131782 168938 131866 169174
rect 132102 168938 311546 169174
rect 311782 168938 311866 169174
rect 312102 168938 347546 169174
rect 347782 168938 347866 169174
rect 348102 168938 383546 169174
rect 383782 168938 383866 169174
rect 384102 168938 419546 169174
rect 419782 168938 419866 169174
rect 420102 168938 455546 169174
rect 455782 168938 455866 169174
rect 456102 168938 491546 169174
rect 491782 168938 491866 169174
rect 492102 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect -4886 168854 588810 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 59546 168854
rect 59782 168618 59866 168854
rect 60102 168618 95546 168854
rect 95782 168618 95866 168854
rect 96102 168618 131546 168854
rect 131782 168618 131866 168854
rect 132102 168618 311546 168854
rect 311782 168618 311866 168854
rect 312102 168618 347546 168854
rect 347782 168618 347866 168854
rect 348102 168618 383546 168854
rect 383782 168618 383866 168854
rect 384102 168618 419546 168854
rect 419782 168618 419866 168854
rect 420102 168618 455546 168854
rect 455782 168618 455866 168854
rect 456102 168618 491546 168854
rect 491782 168618 491866 168854
rect 492102 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect -4886 168586 588810 168618
rect -2966 165454 586890 165486
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 163583 165454
rect 163819 165218 166180 165454
rect 166416 165218 219610 165454
rect 219846 165218 250330 165454
rect 250566 165218 281050 165454
rect 281286 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect -2966 165134 586890 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 163583 165134
rect 163819 164898 166180 165134
rect 166416 164898 219610 165134
rect 219846 164898 250330 165134
rect 250566 164898 281050 165134
rect 281286 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect -2966 164866 586890 164898
rect -8726 158614 592650 158646
rect -8726 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 84986 158614
rect 85222 158378 85306 158614
rect 85542 158378 120986 158614
rect 121222 158378 121306 158614
rect 121542 158378 156986 158614
rect 157222 158378 157306 158614
rect 157542 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 84986 158294
rect 85222 158058 85306 158294
rect 85542 158058 120986 158294
rect 121222 158058 121306 158294
rect 121542 158058 156986 158294
rect 157222 158058 157306 158294
rect 157542 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 592650 158294
rect -8726 158026 592650 158058
rect -6806 154894 590730 154926
rect -6806 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 81266 154894
rect 81502 154658 81586 154894
rect 81822 154658 117266 154894
rect 117502 154658 117586 154894
rect 117822 154658 153266 154894
rect 153502 154658 153586 154894
rect 153822 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 590730 154894
rect -6806 154574 590730 154658
rect -6806 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 81266 154574
rect 81502 154338 81586 154574
rect 81822 154338 117266 154574
rect 117502 154338 117586 154574
rect 117822 154338 153266 154574
rect 153502 154338 153586 154574
rect 153822 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 590730 154574
rect -6806 154306 590730 154338
rect -4886 151174 588810 151206
rect -4886 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 77546 151174
rect 77782 150938 77866 151174
rect 78102 150938 113546 151174
rect 113782 150938 113866 151174
rect 114102 150938 149546 151174
rect 149782 150938 149866 151174
rect 150102 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 588810 151174
rect -4886 150854 588810 150938
rect -4886 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 77546 150854
rect 77782 150618 77866 150854
rect 78102 150618 113546 150854
rect 113782 150618 113866 150854
rect 114102 150618 149546 150854
rect 149782 150618 149866 150854
rect 150102 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 588810 150854
rect -4886 150586 588810 150618
rect -2966 147454 586890 147486
rect -2966 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 162285 147454
rect 162521 147218 164882 147454
rect 165118 147218 167479 147454
rect 167715 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 204250 147454
rect 204486 147218 234970 147454
rect 235206 147218 265690 147454
rect 265926 147218 296410 147454
rect 296646 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 362285 147454
rect 362521 147218 364882 147454
rect 365118 147218 367479 147454
rect 367715 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 434285 147454
rect 434521 147218 436882 147454
rect 437118 147218 439479 147454
rect 439715 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 586890 147454
rect -2966 147134 586890 147218
rect -2966 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 162285 147134
rect 162521 146898 164882 147134
rect 165118 146898 167479 147134
rect 167715 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 204250 147134
rect 204486 146898 234970 147134
rect 235206 146898 265690 147134
rect 265926 146898 296410 147134
rect 296646 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 362285 147134
rect 362521 146898 364882 147134
rect 365118 146898 367479 147134
rect 367715 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 434285 147134
rect 434521 146898 436882 147134
rect 437118 146898 439479 147134
rect 439715 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 586890 147134
rect -2966 146866 586890 146898
rect -8726 140614 592650 140646
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 66986 140614
rect 67222 140378 67306 140614
rect 67542 140378 102986 140614
rect 103222 140378 103306 140614
rect 103542 140378 138986 140614
rect 139222 140378 139306 140614
rect 139542 140378 174986 140614
rect 175222 140378 175306 140614
rect 175542 140378 318986 140614
rect 319222 140378 319306 140614
rect 319542 140378 354986 140614
rect 355222 140378 355306 140614
rect 355542 140378 390986 140614
rect 391222 140378 391306 140614
rect 391542 140378 426986 140614
rect 427222 140378 427306 140614
rect 427542 140378 462986 140614
rect 463222 140378 463306 140614
rect 463542 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect -8726 140294 592650 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 66986 140294
rect 67222 140058 67306 140294
rect 67542 140058 102986 140294
rect 103222 140058 103306 140294
rect 103542 140058 138986 140294
rect 139222 140058 139306 140294
rect 139542 140058 174986 140294
rect 175222 140058 175306 140294
rect 175542 140058 318986 140294
rect 319222 140058 319306 140294
rect 319542 140058 354986 140294
rect 355222 140058 355306 140294
rect 355542 140058 390986 140294
rect 391222 140058 391306 140294
rect 391542 140058 426986 140294
rect 427222 140058 427306 140294
rect 427542 140058 462986 140294
rect 463222 140058 463306 140294
rect 463542 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect -8726 140026 592650 140058
rect -6806 136894 590730 136926
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 63266 136894
rect 63502 136658 63586 136894
rect 63822 136658 99266 136894
rect 99502 136658 99586 136894
rect 99822 136658 135266 136894
rect 135502 136658 135586 136894
rect 135822 136658 315266 136894
rect 315502 136658 315586 136894
rect 315822 136658 351266 136894
rect 351502 136658 351586 136894
rect 351822 136658 387266 136894
rect 387502 136658 387586 136894
rect 387822 136658 423266 136894
rect 423502 136658 423586 136894
rect 423822 136658 459266 136894
rect 459502 136658 459586 136894
rect 459822 136658 495266 136894
rect 495502 136658 495586 136894
rect 495822 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect -6806 136574 590730 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 63266 136574
rect 63502 136338 63586 136574
rect 63822 136338 99266 136574
rect 99502 136338 99586 136574
rect 99822 136338 135266 136574
rect 135502 136338 135586 136574
rect 135822 136338 315266 136574
rect 315502 136338 315586 136574
rect 315822 136338 351266 136574
rect 351502 136338 351586 136574
rect 351822 136338 387266 136574
rect 387502 136338 387586 136574
rect 387822 136338 423266 136574
rect 423502 136338 423586 136574
rect 423822 136338 459266 136574
rect 459502 136338 459586 136574
rect 459822 136338 495266 136574
rect 495502 136338 495586 136574
rect 495822 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect -6806 136306 590730 136338
rect -4886 133174 588810 133206
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 59546 133174
rect 59782 132938 59866 133174
rect 60102 132938 95546 133174
rect 95782 132938 95866 133174
rect 96102 132938 131546 133174
rect 131782 132938 131866 133174
rect 132102 132938 311546 133174
rect 311782 132938 311866 133174
rect 312102 132938 347546 133174
rect 347782 132938 347866 133174
rect 348102 132938 383546 133174
rect 383782 132938 383866 133174
rect 384102 132938 419546 133174
rect 419782 132938 419866 133174
rect 420102 132938 455546 133174
rect 455782 132938 455866 133174
rect 456102 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect -4886 132854 588810 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 59546 132854
rect 59782 132618 59866 132854
rect 60102 132618 95546 132854
rect 95782 132618 95866 132854
rect 96102 132618 131546 132854
rect 131782 132618 131866 132854
rect 132102 132618 311546 132854
rect 311782 132618 311866 132854
rect 312102 132618 347546 132854
rect 347782 132618 347866 132854
rect 348102 132618 383546 132854
rect 383782 132618 383866 132854
rect 384102 132618 419546 132854
rect 419782 132618 419866 132854
rect 420102 132618 455546 132854
rect 455782 132618 455866 132854
rect 456102 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect -4886 132586 588810 132618
rect -2966 129454 586890 129486
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 127826 129454
rect 128062 129218 128146 129454
rect 128382 129218 163583 129454
rect 163819 129218 166180 129454
rect 166416 129218 219610 129454
rect 219846 129218 250330 129454
rect 250566 129218 281050 129454
rect 281286 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 363583 129454
rect 363819 129218 366180 129454
rect 366416 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 435583 129454
rect 435819 129218 438180 129454
rect 438416 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect -2966 129134 586890 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 127826 129134
rect 128062 128898 128146 129134
rect 128382 128898 163583 129134
rect 163819 128898 166180 129134
rect 166416 128898 219610 129134
rect 219846 128898 250330 129134
rect 250566 128898 281050 129134
rect 281286 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 363583 129134
rect 363819 128898 366180 129134
rect 366416 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 435583 129134
rect 435819 128898 438180 129134
rect 438416 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect -2966 128866 586890 128898
rect -8726 122614 592650 122646
rect -8726 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 84986 122614
rect 85222 122378 85306 122614
rect 85542 122378 120986 122614
rect 121222 122378 121306 122614
rect 121542 122378 156986 122614
rect 157222 122378 157306 122614
rect 157542 122378 192986 122614
rect 193222 122378 193306 122614
rect 193542 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 84986 122294
rect 85222 122058 85306 122294
rect 85542 122058 120986 122294
rect 121222 122058 121306 122294
rect 121542 122058 156986 122294
rect 157222 122058 157306 122294
rect 157542 122058 192986 122294
rect 193222 122058 193306 122294
rect 193542 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 592650 122294
rect -8726 122026 592650 122058
rect -6806 118894 590730 118926
rect -6806 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 81266 118894
rect 81502 118658 81586 118894
rect 81822 118658 117266 118894
rect 117502 118658 117586 118894
rect 117822 118658 153266 118894
rect 153502 118658 153586 118894
rect 153822 118658 189266 118894
rect 189502 118658 189586 118894
rect 189822 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 590730 118894
rect -6806 118574 590730 118658
rect -6806 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 81266 118574
rect 81502 118338 81586 118574
rect 81822 118338 117266 118574
rect 117502 118338 117586 118574
rect 117822 118338 153266 118574
rect 153502 118338 153586 118574
rect 153822 118338 189266 118574
rect 189502 118338 189586 118574
rect 189822 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 590730 118574
rect -6806 118306 590730 118338
rect -4886 115174 588810 115206
rect -4886 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 77546 115174
rect 77782 114938 77866 115174
rect 78102 114938 113546 115174
rect 113782 114938 113866 115174
rect 114102 114938 149546 115174
rect 149782 114938 149866 115174
rect 150102 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 588810 115174
rect -4886 114854 588810 114938
rect -4886 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 77546 114854
rect 77782 114618 77866 114854
rect 78102 114618 113546 114854
rect 113782 114618 113866 114854
rect 114102 114618 149546 114854
rect 149782 114618 149866 114854
rect 150102 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 588810 114854
rect -4886 114586 588810 114618
rect -2966 111454 586890 111486
rect -2966 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 204250 111454
rect 204486 111218 234970 111454
rect 235206 111218 265690 111454
rect 265926 111218 296410 111454
rect 296646 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 586890 111454
rect -2966 111134 586890 111218
rect -2966 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 204250 111134
rect 204486 110898 234970 111134
rect 235206 110898 265690 111134
rect 265926 110898 296410 111134
rect 296646 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 586890 111134
rect -2966 110866 586890 110898
rect -8726 104614 592650 104646
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 66986 104614
rect 67222 104378 67306 104614
rect 67542 104378 102986 104614
rect 103222 104378 103306 104614
rect 103542 104378 138986 104614
rect 139222 104378 139306 104614
rect 139542 104378 174986 104614
rect 175222 104378 175306 104614
rect 175542 104378 318986 104614
rect 319222 104378 319306 104614
rect 319542 104378 354986 104614
rect 355222 104378 355306 104614
rect 355542 104378 390986 104614
rect 391222 104378 391306 104614
rect 391542 104378 426986 104614
rect 427222 104378 427306 104614
rect 427542 104378 462986 104614
rect 463222 104378 463306 104614
rect 463542 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect -8726 104294 592650 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 66986 104294
rect 67222 104058 67306 104294
rect 67542 104058 102986 104294
rect 103222 104058 103306 104294
rect 103542 104058 138986 104294
rect 139222 104058 139306 104294
rect 139542 104058 174986 104294
rect 175222 104058 175306 104294
rect 175542 104058 318986 104294
rect 319222 104058 319306 104294
rect 319542 104058 354986 104294
rect 355222 104058 355306 104294
rect 355542 104058 390986 104294
rect 391222 104058 391306 104294
rect 391542 104058 426986 104294
rect 427222 104058 427306 104294
rect 427542 104058 462986 104294
rect 463222 104058 463306 104294
rect 463542 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect -8726 104026 592650 104058
rect -6806 100894 590730 100926
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 63266 100894
rect 63502 100658 63586 100894
rect 63822 100658 99266 100894
rect 99502 100658 99586 100894
rect 99822 100658 135266 100894
rect 135502 100658 135586 100894
rect 135822 100658 171266 100894
rect 171502 100658 171586 100894
rect 171822 100658 315266 100894
rect 315502 100658 315586 100894
rect 315822 100658 351266 100894
rect 351502 100658 351586 100894
rect 351822 100658 387266 100894
rect 387502 100658 387586 100894
rect 387822 100658 423266 100894
rect 423502 100658 423586 100894
rect 423822 100658 459266 100894
rect 459502 100658 459586 100894
rect 459822 100658 495266 100894
rect 495502 100658 495586 100894
rect 495822 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect -6806 100574 590730 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 63266 100574
rect 63502 100338 63586 100574
rect 63822 100338 99266 100574
rect 99502 100338 99586 100574
rect 99822 100338 135266 100574
rect 135502 100338 135586 100574
rect 135822 100338 171266 100574
rect 171502 100338 171586 100574
rect 171822 100338 315266 100574
rect 315502 100338 315586 100574
rect 315822 100338 351266 100574
rect 351502 100338 351586 100574
rect 351822 100338 387266 100574
rect 387502 100338 387586 100574
rect 387822 100338 423266 100574
rect 423502 100338 423586 100574
rect 423822 100338 459266 100574
rect 459502 100338 459586 100574
rect 459822 100338 495266 100574
rect 495502 100338 495586 100574
rect 495822 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect -6806 100306 590730 100338
rect -4886 97174 588810 97206
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 59546 97174
rect 59782 96938 59866 97174
rect 60102 96938 95546 97174
rect 95782 96938 95866 97174
rect 96102 96938 131546 97174
rect 131782 96938 131866 97174
rect 132102 96938 167546 97174
rect 167782 96938 167866 97174
rect 168102 96938 203546 97174
rect 203782 96938 203866 97174
rect 204102 96938 239546 97174
rect 239782 96938 239866 97174
rect 240102 96938 275546 97174
rect 275782 96938 275866 97174
rect 276102 96938 311546 97174
rect 311782 96938 311866 97174
rect 312102 96938 347546 97174
rect 347782 96938 347866 97174
rect 348102 96938 383546 97174
rect 383782 96938 383866 97174
rect 384102 96938 419546 97174
rect 419782 96938 419866 97174
rect 420102 96938 455546 97174
rect 455782 96938 455866 97174
rect 456102 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect -4886 96854 588810 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 59546 96854
rect 59782 96618 59866 96854
rect 60102 96618 95546 96854
rect 95782 96618 95866 96854
rect 96102 96618 131546 96854
rect 131782 96618 131866 96854
rect 132102 96618 167546 96854
rect 167782 96618 167866 96854
rect 168102 96618 203546 96854
rect 203782 96618 203866 96854
rect 204102 96618 239546 96854
rect 239782 96618 239866 96854
rect 240102 96618 275546 96854
rect 275782 96618 275866 96854
rect 276102 96618 311546 96854
rect 311782 96618 311866 96854
rect 312102 96618 347546 96854
rect 347782 96618 347866 96854
rect 348102 96618 383546 96854
rect 383782 96618 383866 96854
rect 384102 96618 419546 96854
rect 419782 96618 419866 96854
rect 420102 96618 455546 96854
rect 455782 96618 455866 96854
rect 456102 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect -4886 96586 588810 96618
rect -2966 93454 586890 93486
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 127826 93454
rect 128062 93218 128146 93454
rect 128382 93218 163826 93454
rect 164062 93218 164146 93454
rect 164382 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect -2966 93134 586890 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 127826 93134
rect 128062 92898 128146 93134
rect 128382 92898 163826 93134
rect 164062 92898 164146 93134
rect 164382 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect -2966 92866 586890 92898
rect -8726 86614 592650 86646
rect -8726 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 120986 86614
rect 121222 86378 121306 86614
rect 121542 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 192986 86614
rect 193222 86378 193306 86614
rect 193542 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 120986 86294
rect 121222 86058 121306 86294
rect 121542 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 192986 86294
rect 193222 86058 193306 86294
rect 193542 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 592650 86294
rect -8726 86026 592650 86058
rect -6806 82894 590730 82926
rect -6806 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 117266 82894
rect 117502 82658 117586 82894
rect 117822 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 189266 82894
rect 189502 82658 189586 82894
rect 189822 82658 225266 82894
rect 225502 82658 225586 82894
rect 225822 82658 261266 82894
rect 261502 82658 261586 82894
rect 261822 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 590730 82894
rect -6806 82574 590730 82658
rect -6806 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 117266 82574
rect 117502 82338 117586 82574
rect 117822 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 189266 82574
rect 189502 82338 189586 82574
rect 189822 82338 225266 82574
rect 225502 82338 225586 82574
rect 225822 82338 261266 82574
rect 261502 82338 261586 82574
rect 261822 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 590730 82574
rect -6806 82306 590730 82338
rect -4886 79174 588810 79206
rect -4886 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 588810 79174
rect -4886 78854 588810 78938
rect -4886 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 588810 78854
rect -4886 78586 588810 78618
rect -2966 75454 586890 75486
rect -2966 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 586890 75454
rect -2966 75134 586890 75218
rect -2966 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 586890 75134
rect -2966 74866 586890 74898
rect -8726 68614 592650 68646
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 66986 68614
rect 67222 68378 67306 68614
rect 67542 68378 102986 68614
rect 103222 68378 103306 68614
rect 103542 68378 138986 68614
rect 139222 68378 139306 68614
rect 139542 68378 174986 68614
rect 175222 68378 175306 68614
rect 175542 68378 210986 68614
rect 211222 68378 211306 68614
rect 211542 68378 246986 68614
rect 247222 68378 247306 68614
rect 247542 68378 282986 68614
rect 283222 68378 283306 68614
rect 283542 68378 318986 68614
rect 319222 68378 319306 68614
rect 319542 68378 354986 68614
rect 355222 68378 355306 68614
rect 355542 68378 390986 68614
rect 391222 68378 391306 68614
rect 391542 68378 426986 68614
rect 427222 68378 427306 68614
rect 427542 68378 462986 68614
rect 463222 68378 463306 68614
rect 463542 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect -8726 68294 592650 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 66986 68294
rect 67222 68058 67306 68294
rect 67542 68058 102986 68294
rect 103222 68058 103306 68294
rect 103542 68058 138986 68294
rect 139222 68058 139306 68294
rect 139542 68058 174986 68294
rect 175222 68058 175306 68294
rect 175542 68058 210986 68294
rect 211222 68058 211306 68294
rect 211542 68058 246986 68294
rect 247222 68058 247306 68294
rect 247542 68058 282986 68294
rect 283222 68058 283306 68294
rect 283542 68058 318986 68294
rect 319222 68058 319306 68294
rect 319542 68058 354986 68294
rect 355222 68058 355306 68294
rect 355542 68058 390986 68294
rect 391222 68058 391306 68294
rect 391542 68058 426986 68294
rect 427222 68058 427306 68294
rect 427542 68058 462986 68294
rect 463222 68058 463306 68294
rect 463542 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect -8726 68026 592650 68058
rect -6806 64894 590730 64926
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 63266 64894
rect 63502 64658 63586 64894
rect 63822 64658 99266 64894
rect 99502 64658 99586 64894
rect 99822 64658 135266 64894
rect 135502 64658 135586 64894
rect 135822 64658 171266 64894
rect 171502 64658 171586 64894
rect 171822 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 243266 64894
rect 243502 64658 243586 64894
rect 243822 64658 279266 64894
rect 279502 64658 279586 64894
rect 279822 64658 315266 64894
rect 315502 64658 315586 64894
rect 315822 64658 351266 64894
rect 351502 64658 351586 64894
rect 351822 64658 387266 64894
rect 387502 64658 387586 64894
rect 387822 64658 423266 64894
rect 423502 64658 423586 64894
rect 423822 64658 459266 64894
rect 459502 64658 459586 64894
rect 459822 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect -6806 64574 590730 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 63266 64574
rect 63502 64338 63586 64574
rect 63822 64338 99266 64574
rect 99502 64338 99586 64574
rect 99822 64338 135266 64574
rect 135502 64338 135586 64574
rect 135822 64338 171266 64574
rect 171502 64338 171586 64574
rect 171822 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 243266 64574
rect 243502 64338 243586 64574
rect 243822 64338 279266 64574
rect 279502 64338 279586 64574
rect 279822 64338 315266 64574
rect 315502 64338 315586 64574
rect 315822 64338 351266 64574
rect 351502 64338 351586 64574
rect 351822 64338 387266 64574
rect 387502 64338 387586 64574
rect 387822 64338 423266 64574
rect 423502 64338 423586 64574
rect 423822 64338 459266 64574
rect 459502 64338 459586 64574
rect 459822 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect -6806 64306 590730 64338
rect -4886 61174 588810 61206
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 59546 61174
rect 59782 60938 59866 61174
rect 60102 60938 95546 61174
rect 95782 60938 95866 61174
rect 96102 60938 131546 61174
rect 131782 60938 131866 61174
rect 132102 60938 167546 61174
rect 167782 60938 167866 61174
rect 168102 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 239546 61174
rect 239782 60938 239866 61174
rect 240102 60938 275546 61174
rect 275782 60938 275866 61174
rect 276102 60938 311546 61174
rect 311782 60938 311866 61174
rect 312102 60938 347546 61174
rect 347782 60938 347866 61174
rect 348102 60938 383546 61174
rect 383782 60938 383866 61174
rect 384102 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect -4886 60854 588810 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 59546 60854
rect 59782 60618 59866 60854
rect 60102 60618 95546 60854
rect 95782 60618 95866 60854
rect 96102 60618 131546 60854
rect 131782 60618 131866 60854
rect 132102 60618 167546 60854
rect 167782 60618 167866 60854
rect 168102 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 239546 60854
rect 239782 60618 239866 60854
rect 240102 60618 275546 60854
rect 275782 60618 275866 60854
rect 276102 60618 311546 60854
rect 311782 60618 311866 60854
rect 312102 60618 347546 60854
rect 347782 60618 347866 60854
rect 348102 60618 383546 60854
rect 383782 60618 383866 60854
rect 384102 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect -4886 60586 588810 60618
rect -2966 57454 586890 57486
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect -2966 57134 586890 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect -2966 56866 586890 56898
rect -8726 50614 592650 50646
rect -8726 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 592650 50294
rect -8726 50026 592650 50058
rect -6806 46894 590730 46926
rect -6806 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 590730 46894
rect -6806 46574 590730 46658
rect -6806 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 590730 46574
rect -6806 46306 590730 46338
rect -4886 43174 588810 43206
rect -4886 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 588810 43174
rect -4886 42854 588810 42938
rect -4886 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 588810 42854
rect -4886 42586 588810 42618
rect -2966 39454 586890 39486
rect -2966 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 586890 39454
rect -2966 39134 586890 39218
rect -2966 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 586890 39134
rect -2966 38866 586890 38898
rect -8726 32614 592650 32646
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect -8726 32294 592650 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect -8726 32026 592650 32058
rect -6806 28894 590730 28926
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect -6806 28574 590730 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect -6806 28306 590730 28338
rect -4886 25174 588810 25206
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect -4886 24854 588810 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect -4886 24586 588810 24618
rect -2966 21454 586890 21486
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect -2966 21134 586890 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect -2966 20866 586890 20898
rect -8726 14614 592650 14646
rect -8726 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 592650 14294
rect -8726 14026 592650 14058
rect -6806 10894 590730 10926
rect -6806 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 590730 10894
rect -6806 10574 590730 10658
rect -6806 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 590730 10574
rect -6806 10306 590730 10338
rect -4886 7174 588810 7206
rect -4886 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 588810 7174
rect -4886 6854 588810 6938
rect -4886 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 588810 6854
rect -4886 6586 588810 6618
rect -2966 3454 586890 3486
rect -2966 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 586890 3454
rect -2966 3134 586890 3218
rect -2966 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 586890 3134
rect -2966 2866 586890 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use digitalcore_macro  digitalcore
timestamp 1641029093
transform 1 0 200000 0 1 100000
box 0 0 100000 200000
use collapsering_macro  ring0
timestamp 1641029093
transform 1 0 160000 0 1 124000
box 934 0 10000 29776
use ringosc_macro  ring1
timestamp 1641029093
transform 1 0 160000 0 1 160000
box 934 0 10000 29504
use collapsering_macro  ring2
timestamp 1641029093
transform 1 0 360000 0 1 124000
box 934 0 10000 29776
use collapsering_macro  ring3
timestamp 1641029093
transform 1 0 360000 0 1 196000
box 934 0 10000 29776
use collapsering_macro  ring4
timestamp 1641029093
transform 1 0 360000 0 1 268000
box 934 0 10000 29776
use collapsering_macro  ring5
timestamp 1641029093
transform 1 0 360000 0 1 340000
box 934 0 10000 29776
use ringosc_macro  ring6
timestamp 1641029093
transform 1 0 432000 0 1 124000
box 934 0 10000 29504
use ringosc_macro  ring7
timestamp 1641029093
transform 1 0 432000 0 1 196000
box 934 0 10000 29504
use ringosc_macro  ring8
timestamp 1641029093
transform 1 0 432000 0 1 268000
box 934 0 10000 29504
use ringosc_macro  ring9
timestamp 1641029093
transform 1 0 432000 0 1 340000
box 934 0 10000 29504
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 38866 586890 39486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 74866 586890 75486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 110866 586890 111486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 146866 586890 147486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 182866 586890 183486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 218866 586890 219486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 254866 586890 255486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 290866 586890 291486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 326866 586890 327486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 362866 586890 363486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 398866 586890 399486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 434866 586890 435486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 470866 586890 471486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 506866 586890 507486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 542866 586890 543486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 578866 586890 579486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 614866 586890 615486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 650866 586890 651486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 686866 586890 687486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 -1894 218414 98000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 -1894 254414 98000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 -1894 290414 98000 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 -1894 362414 122000 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 -1894 434414 122000 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 156000 362414 194000 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 156000 434414 194000 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 228000 362414 266000 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 228000 434414 266000 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 300000 362414 338000 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 300000 434414 338000 6 vccd1
port 531 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 1794 -1894 2414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 -1894 38414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 -1894 74414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 -1894 110414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 -1894 146414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 -1894 182414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 302000 218414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 302000 254414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 302000 290414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 -1894 326414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 372000 362414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 -1894 398414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 372000 434414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 -1894 470414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 -1894 506414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 -1894 542414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 577794 -1894 578414 705830 6 vccd1
port 531 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 532 nsew power input
rlabel metal5 s -4886 6586 588810 7206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 42586 588810 43206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 78586 588810 79206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 114586 588810 115206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 150586 588810 151206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 186586 588810 187206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 222586 588810 223206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 258586 588810 259206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 294586 588810 295206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 330586 588810 331206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 366586 588810 367206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 402586 588810 403206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 438586 588810 439206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 474586 588810 475206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 510586 588810 511206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 546586 588810 547206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 582586 588810 583206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 618586 588810 619206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 654586 588810 655206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 690586 588810 691206 6 vccd2
port 532 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 -3814 222134 98000 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 -3814 258134 98000 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 -3814 294134 98000 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 -3814 366134 122000 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 -3814 438134 122000 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 156000 366134 194000 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 156000 438134 194000 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 228000 366134 266000 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 228000 438134 266000 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 300000 366134 338000 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 300000 438134 338000 6 vccd2
port 532 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 532 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 5514 -3814 6134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 41514 -3814 42134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 -3814 78134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 -3814 114134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 -3814 150134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 -3814 186134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 302000 222134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 302000 258134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 302000 294134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 -3814 330134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 372000 366134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 -3814 402134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 372000 438134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 -3814 474134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 -3814 510134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 545514 -3814 546134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 581514 -3814 582134 707750 6 vccd2
port 532 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 533 nsew power input
rlabel metal5 s -6806 10306 590730 10926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 46306 590730 46926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 82306 590730 82926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 118306 590730 118926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 154306 590730 154926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 190306 590730 190926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 226306 590730 226926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 262306 590730 262926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 298306 590730 298926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 334306 590730 334926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 370306 590730 370926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 406306 590730 406926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 442306 590730 442926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 478306 590730 478926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 514306 590730 514926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 550306 590730 550926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 586306 590730 586926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 622306 590730 622926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 658306 590730 658926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 694306 590730 694926 6 vdda1
port 533 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 -5734 225854 98000 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 -5734 261854 98000 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 -5734 297854 98000 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 -5734 369854 122000 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 -5734 441854 122000 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 156000 369854 194000 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 156000 441854 194000 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 228000 369854 266000 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 228000 441854 266000 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 300000 369854 338000 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 300000 441854 338000 6 vdda1
port 533 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 533 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 9234 -5734 9854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 45234 -5734 45854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 -5734 81854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 -5734 117854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 -5734 153854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 -5734 189854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 302000 225854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 302000 261854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 302000 297854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 -5734 333854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 372000 369854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 -5734 405854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 372000 441854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 -5734 477854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 -5734 513854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 549234 -5734 549854 709670 6 vdda1
port 533 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 534 nsew power input
rlabel metal5 s -8726 14026 592650 14646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 50026 592650 50646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 86026 592650 86646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 122026 592650 122646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 158026 592650 158646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 194026 592650 194646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 230026 592650 230646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 266026 592650 266646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 302026 592650 302646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 338026 592650 338646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 374026 592650 374646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 410026 592650 410646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 446026 592650 446646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 482026 592650 482646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 518026 592650 518646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 554026 592650 554646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 590026 592650 590646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 626026 592650 626646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 662026 592650 662646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 698026 592650 698646 6 vdda2
port 534 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 -7654 229574 98000 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 -7654 265574 98000 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 -7654 301574 98000 6 vdda2
port 534 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 534 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 12954 -7654 13574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 -7654 49574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 -7654 85574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 -7654 121574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 -7654 157574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 -7654 193574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 302000 229574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 302000 265574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 302000 301574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 -7654 337574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 -7654 373574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 -7654 409574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 -7654 445574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 -7654 481574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 -7654 517574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 552954 -7654 553574 711590 6 vdda2
port 534 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 28306 590730 28926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 64306 590730 64926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 100306 590730 100926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 136306 590730 136926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 172306 590730 172926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 208306 590730 208926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 244306 590730 244926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 280306 590730 280926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 316306 590730 316926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 352306 590730 352926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 388306 590730 388926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 424306 590730 424926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 460306 590730 460926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 496306 590730 496926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 532306 590730 532926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 568306 590730 568926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 604306 590730 604926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 640306 590730 640926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 676306 590730 676926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 -5734 207854 98000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 -5734 243854 98000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 -5734 279854 98000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 -5734 171854 122000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 156000 171854 158000 6 vssa1
port 535 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 535 nsew ground input
rlabel metal4 s 27234 -5734 27854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 -5734 63854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 -5734 99854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 -5734 135854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 192000 171854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 302000 207854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 302000 243854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 302000 279854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 -5734 315854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 -5734 351854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 -5734 387854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 -5734 423854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 -5734 459854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 -5734 495854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 -5734 531854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 567234 -5734 567854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 32026 592650 32646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 68026 592650 68646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 104026 592650 104646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 140026 592650 140646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 176026 592650 176646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 212026 592650 212646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 248026 592650 248646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 284026 592650 284646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 320026 592650 320646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 356026 592650 356646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 392026 592650 392646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 428026 592650 428646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 464026 592650 464646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 500026 592650 500646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 536026 592650 536646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 572026 592650 572646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 608026 592650 608646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 644026 592650 644646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 680026 592650 680646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 -7654 211574 98000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 -7654 247574 98000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 -7654 283574 98000 6 vssa2
port 536 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 536 nsew ground input
rlabel metal4 s 30954 -7654 31574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 -7654 67574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 -7654 103574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 -7654 139574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 -7654 175574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 302000 211574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 302000 247574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 302000 283574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 -7654 319574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 -7654 355574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 -7654 391574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 -7654 427574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 -7654 463574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 -7654 499574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 -7654 535574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 570954 -7654 571574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 20866 586890 21486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 56866 586890 57486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 92866 586890 93486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 128866 586890 129486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 164866 586890 165486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 200866 586890 201486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 236866 586890 237486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 272866 586890 273486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 308866 586890 309486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 344866 586890 345486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 380866 586890 381486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 416866 586890 417486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 452866 586890 453486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 488866 586890 489486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 524866 586890 525486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 560866 586890 561486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 596866 586890 597486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 632866 586890 633486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 668866 586890 669486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 -1894 200414 98000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 -1894 236414 98000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 -1894 272414 98000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 -1894 164414 122000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 156000 164414 158000 6 vssd1
port 537 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 537 nsew ground input
rlabel metal4 s 19794 -1894 20414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 -1894 56414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 -1894 92414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 -1894 128414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 192000 164414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 302000 200414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 302000 236414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 302000 272414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 -1894 308414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 -1894 344414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 -1894 380414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 -1894 416414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 -1894 452414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 -1894 488414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 -1894 524414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 559794 -1894 560414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 24586 588810 25206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 60586 588810 61206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 96586 588810 97206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 132586 588810 133206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 168586 588810 169206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 204586 588810 205206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 240586 588810 241206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 276586 588810 277206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 312586 588810 313206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 348586 588810 349206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 384586 588810 385206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 420586 588810 421206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 456586 588810 457206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 492586 588810 493206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 528586 588810 529206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 564586 588810 565206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 600586 588810 601206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 636586 588810 637206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 672586 588810 673206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 -3814 204134 98000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 -3814 240134 98000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 -3814 276134 98000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 -3814 168134 122000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 156000 168134 158000 6 vssd2
port 538 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 538 nsew ground input
rlabel metal4 s 23514 -3814 24134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 -3814 60134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 -3814 96134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 -3814 132134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 192000 168134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 302000 204134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 302000 240134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 302000 276134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 -3814 312134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 -3814 348134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 -3814 384134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 -3814 420134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 -3814 456134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 -3814 492134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 -3814 528134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 563514 -3814 564134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 539 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 540 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 541 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 542 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 543 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 544 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 545 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 546 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 547 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 548 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 549 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 550 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 551 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 552 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 553 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 554 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 555 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 556 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 557 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 558 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 559 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 560 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 561 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 562 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 563 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 564 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 565 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 566 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 567 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 568 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 569 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 570 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 571 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 572 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 573 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 574 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 575 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 576 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 577 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 578 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 579 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 580 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 581 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 582 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 583 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 584 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 585 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 586 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 587 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 588 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 589 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 590 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 591 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 592 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 593 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 594 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 595 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 596 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 597 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 598 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 599 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 600 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 601 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 602 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 603 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 604 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 605 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 606 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 607 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 608 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 609 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 610 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 611 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 612 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 613 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 614 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 615 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 616 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 617 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 618 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 619 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 620 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 621 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 622 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 623 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 624 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 625 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 626 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 627 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 628 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 629 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 630 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 631 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 632 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 633 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 634 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 635 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 636 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 637 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 638 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 639 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 640 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 641 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 642 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 643 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
